magic
tech scmos
timestamp 1617651948
<< polysilicon >>
rect -1302 -988 -1300 -986
rect -1294 -988 -1292 -986
rect -1284 -988 -1282 -986
rect -1058 -988 -1056 -986
rect -1050 -988 -1048 -986
rect -1040 -988 -1038 -986
rect -749 -988 -747 -986
rect -741 -988 -739 -986
rect -731 -988 -729 -986
rect -441 -988 -439 -986
rect -433 -988 -431 -986
rect -423 -988 -421 -986
rect -134 -988 -132 -986
rect -126 -988 -124 -986
rect -116 -988 -114 -986
rect 175 -988 177 -986
rect 183 -988 185 -986
rect 193 -988 195 -986
rect 483 -988 485 -986
rect 491 -988 493 -986
rect 501 -988 503 -986
rect 791 -988 793 -986
rect 799 -988 801 -986
rect 809 -988 811 -986
rect -1302 -1064 -1300 -996
rect -1294 -1020 -1292 -996
rect -1294 -1064 -1292 -1024
rect -1284 -1064 -1282 -996
rect -1058 -1064 -1056 -996
rect -1050 -1020 -1048 -996
rect -1050 -1064 -1048 -1024
rect -1040 -1064 -1038 -996
rect -749 -1064 -747 -996
rect -741 -1020 -739 -996
rect -741 -1064 -739 -1024
rect -731 -1064 -729 -996
rect -441 -1064 -439 -996
rect -433 -1020 -431 -996
rect -433 -1064 -431 -1024
rect -423 -1064 -421 -996
rect -134 -1064 -132 -996
rect -126 -1020 -124 -996
rect -126 -1064 -124 -1024
rect -116 -1064 -114 -996
rect 175 -1064 177 -996
rect 183 -1020 185 -996
rect 183 -1064 185 -1024
rect 193 -1064 195 -996
rect 483 -1064 485 -996
rect 491 -1020 493 -996
rect 491 -1064 493 -1024
rect 501 -1064 503 -996
rect 791 -1064 793 -996
rect 799 -1020 801 -996
rect 799 -1064 801 -1024
rect 809 -1064 811 -996
rect -1302 -1070 -1300 -1068
rect -1294 -1070 -1292 -1068
rect -1284 -1070 -1282 -1068
rect -1058 -1070 -1056 -1068
rect -1050 -1070 -1048 -1068
rect -1040 -1070 -1038 -1068
rect -749 -1070 -747 -1068
rect -741 -1070 -739 -1068
rect -731 -1070 -729 -1068
rect -441 -1070 -439 -1068
rect -433 -1070 -431 -1068
rect -423 -1070 -421 -1068
rect -134 -1070 -132 -1068
rect -126 -1070 -124 -1068
rect -116 -1070 -114 -1068
rect 175 -1070 177 -1068
rect 183 -1070 185 -1068
rect 193 -1070 195 -1068
rect 483 -1070 485 -1068
rect 491 -1070 493 -1068
rect 501 -1070 503 -1068
rect 791 -1070 793 -1068
rect 799 -1070 801 -1068
rect 809 -1070 811 -1068
rect -1304 -1138 -1302 -1136
rect -1296 -1138 -1294 -1136
rect -1286 -1138 -1284 -1136
rect -1057 -1138 -1055 -1136
rect -1049 -1138 -1047 -1136
rect -1039 -1138 -1037 -1136
rect -749 -1138 -747 -1136
rect -741 -1138 -739 -1136
rect -731 -1138 -729 -1136
rect -441 -1138 -439 -1136
rect -433 -1138 -431 -1136
rect -423 -1138 -421 -1136
rect -133 -1138 -131 -1136
rect -125 -1138 -123 -1136
rect -115 -1138 -113 -1136
rect 175 -1138 177 -1136
rect 183 -1138 185 -1136
rect 193 -1138 195 -1136
rect 483 -1138 485 -1136
rect 491 -1138 493 -1136
rect 501 -1138 503 -1136
rect 791 -1138 793 -1136
rect 799 -1138 801 -1136
rect 809 -1138 811 -1136
rect -1304 -1214 -1302 -1146
rect -1296 -1170 -1294 -1146
rect -1296 -1214 -1294 -1174
rect -1286 -1214 -1284 -1146
rect -1057 -1214 -1055 -1146
rect -1049 -1170 -1047 -1146
rect -1049 -1214 -1047 -1174
rect -1039 -1214 -1037 -1146
rect -749 -1214 -747 -1146
rect -741 -1170 -739 -1146
rect -741 -1214 -739 -1174
rect -731 -1214 -729 -1146
rect -441 -1214 -439 -1146
rect -433 -1170 -431 -1146
rect -433 -1214 -431 -1174
rect -423 -1214 -421 -1146
rect -133 -1214 -131 -1146
rect -125 -1170 -123 -1146
rect -125 -1214 -123 -1174
rect -115 -1214 -113 -1146
rect 175 -1214 177 -1146
rect 183 -1170 185 -1146
rect 183 -1214 185 -1174
rect 193 -1214 195 -1146
rect 483 -1214 485 -1146
rect 491 -1170 493 -1146
rect 491 -1214 493 -1174
rect 501 -1214 503 -1146
rect 791 -1214 793 -1146
rect 799 -1170 801 -1146
rect 799 -1214 801 -1174
rect 809 -1214 811 -1146
rect -1304 -1220 -1302 -1218
rect -1296 -1220 -1294 -1218
rect -1286 -1220 -1284 -1218
rect -1057 -1220 -1055 -1218
rect -1049 -1220 -1047 -1218
rect -1039 -1220 -1037 -1218
rect -749 -1220 -747 -1218
rect -741 -1220 -739 -1218
rect -731 -1220 -729 -1218
rect -441 -1220 -439 -1218
rect -433 -1220 -431 -1218
rect -423 -1220 -421 -1218
rect -133 -1220 -131 -1218
rect -125 -1220 -123 -1218
rect -115 -1220 -113 -1218
rect 175 -1220 177 -1218
rect 183 -1220 185 -1218
rect 193 -1220 195 -1218
rect 483 -1220 485 -1218
rect 491 -1220 493 -1218
rect 501 -1220 503 -1218
rect 791 -1220 793 -1218
rect 799 -1220 801 -1218
rect 809 -1220 811 -1218
rect -1225 -1302 -1223 -1300
rect -1215 -1302 -1213 -1300
rect -1199 -1302 -1197 -1300
rect -1189 -1302 -1187 -1300
rect -1181 -1302 -1179 -1300
rect -1171 -1302 -1169 -1300
rect -1155 -1302 -1153 -1300
rect -1147 -1302 -1145 -1300
rect -1137 -1302 -1135 -1300
rect -1057 -1302 -1055 -1300
rect -1047 -1302 -1045 -1300
rect -1031 -1302 -1029 -1300
rect -1021 -1302 -1019 -1300
rect -1005 -1302 -1003 -1300
rect -995 -1302 -993 -1300
rect -987 -1302 -985 -1300
rect -977 -1302 -975 -1300
rect -961 -1302 -959 -1300
rect -953 -1302 -951 -1300
rect -943 -1302 -941 -1300
rect -927 -1302 -925 -1300
rect -917 -1302 -915 -1300
rect -909 -1302 -907 -1300
rect -899 -1302 -897 -1300
rect -883 -1302 -881 -1300
rect -875 -1302 -873 -1300
rect -859 -1302 -857 -1300
rect -843 -1302 -841 -1300
rect -835 -1302 -833 -1300
rect -825 -1302 -823 -1300
rect -749 -1302 -747 -1300
rect -739 -1302 -737 -1300
rect -723 -1302 -721 -1300
rect -713 -1302 -711 -1300
rect -697 -1302 -695 -1300
rect -687 -1302 -685 -1300
rect -679 -1302 -677 -1300
rect -669 -1302 -667 -1300
rect -653 -1302 -651 -1300
rect -645 -1302 -643 -1300
rect -635 -1302 -633 -1300
rect -619 -1302 -617 -1300
rect -609 -1302 -607 -1300
rect -601 -1302 -599 -1300
rect -591 -1302 -589 -1300
rect -575 -1302 -573 -1300
rect -567 -1302 -565 -1300
rect -551 -1302 -549 -1300
rect -535 -1302 -533 -1300
rect -527 -1302 -525 -1300
rect -517 -1302 -515 -1300
rect -441 -1302 -439 -1300
rect -431 -1302 -429 -1300
rect -415 -1302 -413 -1300
rect -405 -1302 -403 -1300
rect -389 -1302 -387 -1300
rect -379 -1302 -377 -1300
rect -371 -1302 -369 -1300
rect -361 -1302 -359 -1300
rect -345 -1302 -343 -1300
rect -337 -1302 -335 -1300
rect -327 -1302 -325 -1300
rect -311 -1302 -309 -1300
rect -301 -1302 -299 -1300
rect -293 -1302 -291 -1300
rect -283 -1302 -281 -1300
rect -267 -1302 -265 -1300
rect -259 -1302 -257 -1300
rect -243 -1302 -241 -1300
rect -227 -1302 -225 -1300
rect -219 -1302 -217 -1300
rect -209 -1302 -207 -1300
rect -133 -1302 -131 -1300
rect -123 -1302 -121 -1300
rect -107 -1302 -105 -1300
rect -97 -1302 -95 -1300
rect -81 -1302 -79 -1300
rect -71 -1302 -69 -1300
rect -63 -1302 -61 -1300
rect -53 -1302 -51 -1300
rect -37 -1302 -35 -1300
rect -29 -1302 -27 -1300
rect -19 -1302 -17 -1300
rect -3 -1302 -1 -1300
rect 7 -1302 9 -1300
rect 15 -1302 17 -1300
rect 25 -1302 27 -1300
rect 41 -1302 43 -1300
rect 49 -1302 51 -1300
rect 65 -1302 67 -1300
rect 81 -1302 83 -1300
rect 89 -1302 91 -1300
rect 99 -1302 101 -1300
rect 175 -1302 177 -1300
rect 185 -1302 187 -1300
rect 201 -1302 203 -1300
rect 211 -1302 213 -1300
rect 227 -1302 229 -1300
rect 237 -1302 239 -1300
rect 245 -1302 247 -1300
rect 255 -1302 257 -1300
rect 271 -1302 273 -1300
rect 279 -1302 281 -1300
rect 289 -1302 291 -1300
rect 305 -1302 307 -1300
rect 315 -1302 317 -1300
rect 323 -1302 325 -1300
rect 333 -1302 335 -1300
rect 349 -1302 351 -1300
rect 357 -1302 359 -1300
rect 373 -1302 375 -1300
rect 389 -1302 391 -1300
rect 397 -1302 399 -1300
rect 407 -1302 409 -1300
rect 483 -1302 485 -1300
rect 493 -1302 495 -1300
rect 509 -1302 511 -1300
rect 519 -1302 521 -1300
rect 535 -1302 537 -1300
rect 545 -1302 547 -1300
rect 553 -1302 555 -1300
rect 563 -1302 565 -1300
rect 579 -1302 581 -1300
rect 587 -1302 589 -1300
rect 597 -1302 599 -1300
rect 613 -1302 615 -1300
rect 623 -1302 625 -1300
rect 631 -1302 633 -1300
rect 641 -1302 643 -1300
rect 657 -1302 659 -1300
rect 665 -1302 667 -1300
rect 681 -1302 683 -1300
rect 697 -1302 699 -1300
rect 705 -1302 707 -1300
rect 715 -1302 717 -1300
rect 789 -1302 791 -1300
rect 799 -1302 801 -1300
rect 815 -1302 817 -1300
rect 825 -1302 827 -1300
rect 833 -1302 835 -1300
rect 843 -1302 845 -1300
rect 859 -1302 861 -1300
rect 867 -1302 869 -1300
rect 877 -1302 879 -1300
rect -1225 -1378 -1223 -1310
rect -1215 -1378 -1213 -1310
rect -1199 -1378 -1197 -1310
rect -1189 -1378 -1187 -1310
rect -1181 -1378 -1179 -1310
rect -1171 -1378 -1169 -1310
rect -1155 -1378 -1153 -1310
rect -1147 -1378 -1145 -1310
rect -1137 -1378 -1135 -1310
rect -1057 -1378 -1055 -1310
rect -1047 -1378 -1045 -1310
rect -1031 -1378 -1029 -1310
rect -1021 -1378 -1019 -1310
rect -1005 -1378 -1003 -1310
rect -995 -1378 -993 -1310
rect -987 -1378 -985 -1310
rect -977 -1378 -975 -1310
rect -961 -1378 -959 -1310
rect -953 -1378 -951 -1310
rect -943 -1378 -941 -1310
rect -927 -1378 -925 -1310
rect -917 -1378 -915 -1310
rect -909 -1378 -907 -1310
rect -899 -1378 -897 -1310
rect -883 -1378 -881 -1310
rect -875 -1378 -873 -1310
rect -859 -1378 -857 -1310
rect -843 -1378 -841 -1310
rect -835 -1378 -833 -1310
rect -825 -1378 -823 -1310
rect -749 -1378 -747 -1310
rect -739 -1378 -737 -1310
rect -723 -1378 -721 -1310
rect -713 -1378 -711 -1310
rect -697 -1378 -695 -1310
rect -687 -1378 -685 -1310
rect -679 -1378 -677 -1310
rect -669 -1378 -667 -1310
rect -653 -1378 -651 -1310
rect -645 -1378 -643 -1310
rect -635 -1378 -633 -1310
rect -619 -1378 -617 -1310
rect -609 -1378 -607 -1310
rect -601 -1378 -599 -1310
rect -591 -1378 -589 -1310
rect -575 -1378 -573 -1310
rect -567 -1378 -565 -1310
rect -551 -1378 -549 -1310
rect -535 -1378 -533 -1310
rect -527 -1378 -525 -1310
rect -517 -1378 -515 -1310
rect -441 -1378 -439 -1310
rect -431 -1378 -429 -1310
rect -415 -1378 -413 -1310
rect -405 -1378 -403 -1310
rect -389 -1378 -387 -1310
rect -379 -1378 -377 -1310
rect -371 -1378 -369 -1310
rect -361 -1378 -359 -1310
rect -345 -1378 -343 -1310
rect -337 -1378 -335 -1310
rect -327 -1378 -325 -1310
rect -311 -1378 -309 -1310
rect -301 -1378 -299 -1310
rect -293 -1378 -291 -1310
rect -283 -1378 -281 -1310
rect -267 -1378 -265 -1310
rect -259 -1378 -257 -1310
rect -243 -1378 -241 -1310
rect -227 -1378 -225 -1310
rect -219 -1378 -217 -1310
rect -209 -1378 -207 -1310
rect -133 -1378 -131 -1310
rect -123 -1378 -121 -1310
rect -107 -1378 -105 -1310
rect -97 -1378 -95 -1310
rect -81 -1378 -79 -1310
rect -71 -1378 -69 -1310
rect -63 -1378 -61 -1310
rect -53 -1378 -51 -1310
rect -37 -1378 -35 -1310
rect -29 -1378 -27 -1310
rect -19 -1378 -17 -1310
rect -3 -1378 -1 -1310
rect 7 -1378 9 -1310
rect 15 -1378 17 -1310
rect 25 -1378 27 -1310
rect 41 -1378 43 -1310
rect 49 -1378 51 -1310
rect 65 -1378 67 -1310
rect 81 -1378 83 -1310
rect 89 -1378 91 -1310
rect 99 -1378 101 -1310
rect 175 -1378 177 -1310
rect 185 -1378 187 -1310
rect 201 -1378 203 -1310
rect 211 -1378 213 -1310
rect 227 -1378 229 -1310
rect 237 -1378 239 -1310
rect 245 -1378 247 -1310
rect 255 -1378 257 -1310
rect 271 -1378 273 -1310
rect 279 -1378 281 -1310
rect 289 -1378 291 -1310
rect 305 -1378 307 -1310
rect 315 -1378 317 -1310
rect 323 -1378 325 -1310
rect 333 -1378 335 -1310
rect 349 -1378 351 -1310
rect 357 -1378 359 -1310
rect 373 -1378 375 -1310
rect 389 -1378 391 -1310
rect 397 -1378 399 -1310
rect 407 -1378 409 -1310
rect 483 -1378 485 -1310
rect 493 -1378 495 -1310
rect 509 -1378 511 -1310
rect 519 -1378 521 -1310
rect 535 -1378 537 -1310
rect 545 -1378 547 -1310
rect 553 -1378 555 -1310
rect 563 -1378 565 -1310
rect 579 -1378 581 -1310
rect 587 -1378 589 -1310
rect 597 -1378 599 -1310
rect 613 -1378 615 -1310
rect 623 -1378 625 -1310
rect 631 -1378 633 -1310
rect 641 -1378 643 -1310
rect 657 -1378 659 -1310
rect 665 -1378 667 -1310
rect 681 -1378 683 -1310
rect 697 -1378 699 -1310
rect 705 -1378 707 -1310
rect 715 -1378 717 -1310
rect 789 -1378 791 -1310
rect 799 -1378 801 -1310
rect 815 -1378 817 -1310
rect 825 -1378 827 -1310
rect 833 -1378 835 -1310
rect 843 -1378 845 -1310
rect 859 -1378 861 -1310
rect 867 -1378 869 -1310
rect 877 -1378 879 -1310
rect -1225 -1384 -1223 -1382
rect -1215 -1384 -1213 -1382
rect -1199 -1384 -1197 -1382
rect -1189 -1384 -1187 -1382
rect -1181 -1384 -1179 -1382
rect -1171 -1384 -1169 -1382
rect -1155 -1384 -1153 -1382
rect -1147 -1384 -1145 -1382
rect -1137 -1384 -1135 -1382
rect -1057 -1384 -1055 -1382
rect -1047 -1384 -1045 -1382
rect -1031 -1384 -1029 -1382
rect -1021 -1384 -1019 -1382
rect -1005 -1384 -1003 -1382
rect -995 -1384 -993 -1382
rect -987 -1384 -985 -1382
rect -977 -1384 -975 -1382
rect -961 -1384 -959 -1382
rect -953 -1384 -951 -1382
rect -943 -1384 -941 -1382
rect -927 -1384 -925 -1382
rect -917 -1384 -915 -1382
rect -909 -1384 -907 -1382
rect -899 -1384 -897 -1382
rect -883 -1384 -881 -1382
rect -875 -1384 -873 -1382
rect -859 -1384 -857 -1382
rect -843 -1384 -841 -1382
rect -835 -1384 -833 -1382
rect -825 -1384 -823 -1382
rect -749 -1384 -747 -1382
rect -739 -1384 -737 -1382
rect -723 -1384 -721 -1382
rect -713 -1384 -711 -1382
rect -697 -1384 -695 -1382
rect -687 -1384 -685 -1382
rect -679 -1384 -677 -1382
rect -669 -1384 -667 -1382
rect -653 -1384 -651 -1382
rect -645 -1384 -643 -1382
rect -635 -1384 -633 -1382
rect -619 -1384 -617 -1382
rect -609 -1384 -607 -1382
rect -601 -1384 -599 -1382
rect -591 -1384 -589 -1382
rect -575 -1384 -573 -1382
rect -567 -1384 -565 -1382
rect -551 -1384 -549 -1382
rect -535 -1384 -533 -1382
rect -527 -1384 -525 -1382
rect -517 -1384 -515 -1382
rect -441 -1384 -439 -1382
rect -431 -1384 -429 -1382
rect -415 -1384 -413 -1382
rect -405 -1384 -403 -1382
rect -389 -1384 -387 -1382
rect -379 -1384 -377 -1382
rect -371 -1384 -369 -1382
rect -361 -1384 -359 -1382
rect -345 -1384 -343 -1382
rect -337 -1384 -335 -1382
rect -327 -1384 -325 -1382
rect -311 -1384 -309 -1382
rect -301 -1384 -299 -1382
rect -293 -1384 -291 -1382
rect -283 -1384 -281 -1382
rect -267 -1384 -265 -1382
rect -259 -1384 -257 -1382
rect -243 -1384 -241 -1382
rect -227 -1384 -225 -1382
rect -219 -1384 -217 -1382
rect -209 -1384 -207 -1382
rect -133 -1384 -131 -1382
rect -123 -1384 -121 -1382
rect -107 -1384 -105 -1382
rect -97 -1384 -95 -1382
rect -81 -1384 -79 -1382
rect -71 -1384 -69 -1382
rect -63 -1384 -61 -1382
rect -53 -1384 -51 -1382
rect -37 -1384 -35 -1382
rect -29 -1384 -27 -1382
rect -19 -1384 -17 -1382
rect -3 -1384 -1 -1382
rect 7 -1384 9 -1382
rect 15 -1384 17 -1382
rect 25 -1384 27 -1382
rect 41 -1384 43 -1382
rect 49 -1384 51 -1382
rect 65 -1384 67 -1382
rect 81 -1384 83 -1382
rect 89 -1384 91 -1382
rect 99 -1384 101 -1382
rect 175 -1384 177 -1382
rect 185 -1384 187 -1382
rect 201 -1384 203 -1382
rect 211 -1384 213 -1382
rect 227 -1384 229 -1382
rect 237 -1384 239 -1382
rect 245 -1384 247 -1382
rect 255 -1384 257 -1382
rect 271 -1384 273 -1382
rect 279 -1384 281 -1382
rect 289 -1384 291 -1382
rect 305 -1384 307 -1382
rect 315 -1384 317 -1382
rect 323 -1384 325 -1382
rect 333 -1384 335 -1382
rect 349 -1384 351 -1382
rect 357 -1384 359 -1382
rect 373 -1384 375 -1382
rect 389 -1384 391 -1382
rect 397 -1384 399 -1382
rect 407 -1384 409 -1382
rect 483 -1384 485 -1382
rect 493 -1384 495 -1382
rect 509 -1384 511 -1382
rect 519 -1384 521 -1382
rect 535 -1384 537 -1382
rect 545 -1384 547 -1382
rect 553 -1384 555 -1382
rect 563 -1384 565 -1382
rect 579 -1384 581 -1382
rect 587 -1384 589 -1382
rect 597 -1384 599 -1382
rect 613 -1384 615 -1382
rect 623 -1384 625 -1382
rect 631 -1384 633 -1382
rect 641 -1384 643 -1382
rect 657 -1384 659 -1382
rect 665 -1384 667 -1382
rect 681 -1384 683 -1382
rect 697 -1384 699 -1382
rect 705 -1384 707 -1382
rect 715 -1384 717 -1382
rect 789 -1384 791 -1382
rect 799 -1384 801 -1382
rect 815 -1384 817 -1382
rect 825 -1384 827 -1382
rect 833 -1384 835 -1382
rect 843 -1384 845 -1382
rect 859 -1384 861 -1382
rect 867 -1384 869 -1382
rect 877 -1384 879 -1382
rect -1304 -1459 -1302 -1457
rect -1296 -1459 -1294 -1457
rect -1286 -1459 -1284 -1457
rect -1057 -1459 -1055 -1457
rect -1049 -1459 -1047 -1457
rect -1039 -1459 -1037 -1457
rect -749 -1459 -747 -1457
rect -741 -1459 -739 -1457
rect -731 -1459 -729 -1457
rect -441 -1459 -439 -1457
rect -433 -1459 -431 -1457
rect -423 -1459 -421 -1457
rect -133 -1459 -131 -1457
rect -125 -1459 -123 -1457
rect -115 -1459 -113 -1457
rect 175 -1459 177 -1457
rect 183 -1459 185 -1457
rect 193 -1459 195 -1457
rect 483 -1459 485 -1457
rect 491 -1459 493 -1457
rect 501 -1459 503 -1457
rect 791 -1459 793 -1457
rect 799 -1459 801 -1457
rect 809 -1459 811 -1457
rect -1304 -1535 -1302 -1467
rect -1296 -1491 -1294 -1467
rect -1296 -1535 -1294 -1495
rect -1286 -1535 -1284 -1467
rect -1057 -1535 -1055 -1467
rect -1049 -1491 -1047 -1467
rect -1049 -1535 -1047 -1495
rect -1039 -1535 -1037 -1467
rect -749 -1535 -747 -1467
rect -741 -1491 -739 -1467
rect -741 -1535 -739 -1495
rect -731 -1535 -729 -1467
rect -441 -1535 -439 -1467
rect -433 -1491 -431 -1467
rect -433 -1535 -431 -1495
rect -423 -1535 -421 -1467
rect -133 -1535 -131 -1467
rect -125 -1491 -123 -1467
rect -125 -1535 -123 -1495
rect -115 -1535 -113 -1467
rect 175 -1535 177 -1467
rect 183 -1491 185 -1467
rect 183 -1535 185 -1495
rect 193 -1535 195 -1467
rect 483 -1535 485 -1467
rect 491 -1491 493 -1467
rect 491 -1535 493 -1495
rect 501 -1535 503 -1467
rect 791 -1535 793 -1467
rect 799 -1491 801 -1467
rect 799 -1535 801 -1495
rect 809 -1535 811 -1467
rect -1304 -1541 -1302 -1539
rect -1296 -1541 -1294 -1539
rect -1286 -1541 -1284 -1539
rect -1057 -1541 -1055 -1539
rect -1049 -1541 -1047 -1539
rect -1039 -1541 -1037 -1539
rect -749 -1541 -747 -1539
rect -741 -1541 -739 -1539
rect -731 -1541 -729 -1539
rect -441 -1541 -439 -1539
rect -433 -1541 -431 -1539
rect -423 -1541 -421 -1539
rect -133 -1541 -131 -1539
rect -125 -1541 -123 -1539
rect -115 -1541 -113 -1539
rect 175 -1541 177 -1539
rect 183 -1541 185 -1539
rect 193 -1541 195 -1539
rect 483 -1541 485 -1539
rect 491 -1541 493 -1539
rect 501 -1541 503 -1539
rect 791 -1541 793 -1539
rect 799 -1541 801 -1539
rect 809 -1541 811 -1539
rect -1229 -1618 -1227 -1616
rect -1219 -1618 -1217 -1616
rect -1203 -1618 -1201 -1616
rect -1193 -1618 -1191 -1616
rect -1185 -1618 -1183 -1616
rect -1175 -1618 -1173 -1616
rect -1159 -1618 -1157 -1616
rect -1151 -1618 -1149 -1616
rect -1141 -1618 -1139 -1616
rect -1057 -1618 -1055 -1616
rect -1047 -1618 -1045 -1616
rect -1031 -1618 -1029 -1616
rect -1021 -1618 -1019 -1616
rect -1005 -1618 -1003 -1616
rect -995 -1618 -993 -1616
rect -987 -1618 -985 -1616
rect -977 -1618 -975 -1616
rect -961 -1618 -959 -1616
rect -953 -1618 -951 -1616
rect -943 -1618 -941 -1616
rect -927 -1618 -925 -1616
rect -917 -1618 -915 -1616
rect -909 -1618 -907 -1616
rect -899 -1618 -897 -1616
rect -883 -1618 -881 -1616
rect -875 -1618 -873 -1616
rect -859 -1618 -857 -1616
rect -843 -1618 -841 -1616
rect -835 -1618 -833 -1616
rect -825 -1618 -823 -1616
rect -749 -1618 -747 -1616
rect -739 -1618 -737 -1616
rect -723 -1618 -721 -1616
rect -713 -1618 -711 -1616
rect -697 -1618 -695 -1616
rect -687 -1618 -685 -1616
rect -679 -1618 -677 -1616
rect -669 -1618 -667 -1616
rect -653 -1618 -651 -1616
rect -645 -1618 -643 -1616
rect -635 -1618 -633 -1616
rect -619 -1618 -617 -1616
rect -609 -1618 -607 -1616
rect -601 -1618 -599 -1616
rect -591 -1618 -589 -1616
rect -575 -1618 -573 -1616
rect -567 -1618 -565 -1616
rect -551 -1618 -549 -1616
rect -535 -1618 -533 -1616
rect -527 -1618 -525 -1616
rect -517 -1618 -515 -1616
rect -441 -1618 -439 -1616
rect -431 -1618 -429 -1616
rect -415 -1618 -413 -1616
rect -405 -1618 -403 -1616
rect -389 -1618 -387 -1616
rect -379 -1618 -377 -1616
rect -371 -1618 -369 -1616
rect -361 -1618 -359 -1616
rect -345 -1618 -343 -1616
rect -337 -1618 -335 -1616
rect -327 -1618 -325 -1616
rect -311 -1618 -309 -1616
rect -301 -1618 -299 -1616
rect -293 -1618 -291 -1616
rect -283 -1618 -281 -1616
rect -267 -1618 -265 -1616
rect -259 -1618 -257 -1616
rect -243 -1618 -241 -1616
rect -227 -1618 -225 -1616
rect -219 -1618 -217 -1616
rect -209 -1618 -207 -1616
rect -133 -1618 -131 -1616
rect -123 -1618 -121 -1616
rect -107 -1618 -105 -1616
rect -97 -1618 -95 -1616
rect -81 -1618 -79 -1616
rect -71 -1618 -69 -1616
rect -63 -1618 -61 -1616
rect -53 -1618 -51 -1616
rect -37 -1618 -35 -1616
rect -29 -1618 -27 -1616
rect -19 -1618 -17 -1616
rect -3 -1618 -1 -1616
rect 7 -1618 9 -1616
rect 15 -1618 17 -1616
rect 25 -1618 27 -1616
rect 41 -1618 43 -1616
rect 49 -1618 51 -1616
rect 65 -1618 67 -1616
rect 81 -1618 83 -1616
rect 89 -1618 91 -1616
rect 99 -1618 101 -1616
rect 175 -1618 177 -1616
rect 185 -1618 187 -1616
rect 201 -1618 203 -1616
rect 211 -1618 213 -1616
rect 227 -1618 229 -1616
rect 237 -1618 239 -1616
rect 245 -1618 247 -1616
rect 255 -1618 257 -1616
rect 271 -1618 273 -1616
rect 279 -1618 281 -1616
rect 289 -1618 291 -1616
rect 305 -1618 307 -1616
rect 315 -1618 317 -1616
rect 323 -1618 325 -1616
rect 333 -1618 335 -1616
rect 349 -1618 351 -1616
rect 357 -1618 359 -1616
rect 373 -1618 375 -1616
rect 389 -1618 391 -1616
rect 397 -1618 399 -1616
rect 407 -1618 409 -1616
rect 483 -1618 485 -1616
rect 493 -1618 495 -1616
rect 509 -1618 511 -1616
rect 519 -1618 521 -1616
rect 535 -1618 537 -1616
rect 545 -1618 547 -1616
rect 553 -1618 555 -1616
rect 563 -1618 565 -1616
rect 579 -1618 581 -1616
rect 587 -1618 589 -1616
rect 597 -1618 599 -1616
rect 613 -1618 615 -1616
rect 623 -1618 625 -1616
rect 631 -1618 633 -1616
rect 641 -1618 643 -1616
rect 657 -1618 659 -1616
rect 665 -1618 667 -1616
rect 681 -1618 683 -1616
rect 697 -1618 699 -1616
rect 705 -1618 707 -1616
rect 715 -1618 717 -1616
rect 791 -1618 793 -1616
rect 801 -1618 803 -1616
rect 817 -1618 819 -1616
rect 827 -1618 829 -1616
rect 843 -1618 845 -1616
rect 853 -1618 855 -1616
rect 861 -1618 863 -1616
rect 871 -1618 873 -1616
rect 887 -1618 889 -1616
rect 895 -1618 897 -1616
rect 905 -1618 907 -1616
rect 921 -1618 923 -1616
rect 931 -1618 933 -1616
rect 939 -1618 941 -1616
rect 949 -1618 951 -1616
rect 965 -1618 967 -1616
rect 973 -1618 975 -1616
rect 989 -1618 991 -1616
rect 1005 -1618 1007 -1616
rect 1013 -1618 1015 -1616
rect 1023 -1618 1025 -1616
rect -1229 -1694 -1227 -1626
rect -1219 -1694 -1217 -1626
rect -1203 -1694 -1201 -1626
rect -1193 -1694 -1191 -1626
rect -1185 -1694 -1183 -1626
rect -1175 -1694 -1173 -1626
rect -1159 -1694 -1157 -1626
rect -1151 -1694 -1149 -1626
rect -1141 -1694 -1139 -1626
rect -1057 -1694 -1055 -1626
rect -1047 -1694 -1045 -1626
rect -1031 -1694 -1029 -1626
rect -1021 -1694 -1019 -1626
rect -1005 -1694 -1003 -1626
rect -995 -1694 -993 -1626
rect -987 -1694 -985 -1626
rect -977 -1694 -975 -1626
rect -961 -1694 -959 -1626
rect -953 -1694 -951 -1626
rect -943 -1694 -941 -1626
rect -927 -1694 -925 -1626
rect -917 -1694 -915 -1626
rect -909 -1694 -907 -1626
rect -899 -1694 -897 -1626
rect -883 -1694 -881 -1626
rect -875 -1694 -873 -1626
rect -859 -1694 -857 -1626
rect -843 -1694 -841 -1626
rect -835 -1694 -833 -1626
rect -825 -1694 -823 -1626
rect -749 -1694 -747 -1626
rect -739 -1694 -737 -1626
rect -723 -1694 -721 -1626
rect -713 -1694 -711 -1626
rect -697 -1694 -695 -1626
rect -687 -1694 -685 -1626
rect -679 -1694 -677 -1626
rect -669 -1694 -667 -1626
rect -653 -1694 -651 -1626
rect -645 -1694 -643 -1626
rect -635 -1694 -633 -1626
rect -619 -1694 -617 -1626
rect -609 -1694 -607 -1626
rect -601 -1694 -599 -1626
rect -591 -1694 -589 -1626
rect -575 -1694 -573 -1626
rect -567 -1694 -565 -1626
rect -551 -1694 -549 -1626
rect -535 -1694 -533 -1626
rect -527 -1694 -525 -1626
rect -517 -1694 -515 -1626
rect -441 -1694 -439 -1626
rect -431 -1694 -429 -1626
rect -415 -1694 -413 -1626
rect -405 -1694 -403 -1626
rect -389 -1694 -387 -1626
rect -379 -1694 -377 -1626
rect -371 -1694 -369 -1626
rect -361 -1694 -359 -1626
rect -345 -1694 -343 -1626
rect -337 -1694 -335 -1626
rect -327 -1694 -325 -1626
rect -311 -1694 -309 -1626
rect -301 -1694 -299 -1626
rect -293 -1694 -291 -1626
rect -283 -1694 -281 -1626
rect -267 -1694 -265 -1626
rect -259 -1694 -257 -1626
rect -243 -1694 -241 -1626
rect -227 -1694 -225 -1626
rect -219 -1694 -217 -1626
rect -209 -1694 -207 -1626
rect -133 -1694 -131 -1626
rect -123 -1694 -121 -1626
rect -107 -1694 -105 -1626
rect -97 -1694 -95 -1626
rect -81 -1694 -79 -1626
rect -71 -1694 -69 -1626
rect -63 -1694 -61 -1626
rect -53 -1694 -51 -1626
rect -37 -1694 -35 -1626
rect -29 -1694 -27 -1626
rect -19 -1694 -17 -1626
rect -3 -1694 -1 -1626
rect 7 -1694 9 -1626
rect 15 -1694 17 -1626
rect 25 -1694 27 -1626
rect 41 -1694 43 -1626
rect 49 -1694 51 -1626
rect 65 -1694 67 -1626
rect 81 -1694 83 -1626
rect 89 -1694 91 -1626
rect 99 -1694 101 -1626
rect 175 -1694 177 -1626
rect 185 -1694 187 -1626
rect 201 -1694 203 -1626
rect 211 -1694 213 -1626
rect 227 -1694 229 -1626
rect 237 -1694 239 -1626
rect 245 -1694 247 -1626
rect 255 -1694 257 -1626
rect 271 -1694 273 -1626
rect 279 -1694 281 -1626
rect 289 -1694 291 -1626
rect 305 -1694 307 -1626
rect 315 -1694 317 -1626
rect 323 -1694 325 -1626
rect 333 -1694 335 -1626
rect 349 -1694 351 -1626
rect 357 -1694 359 -1626
rect 373 -1694 375 -1626
rect 389 -1694 391 -1626
rect 397 -1694 399 -1626
rect 407 -1694 409 -1626
rect 483 -1694 485 -1626
rect 493 -1694 495 -1626
rect 509 -1694 511 -1626
rect 519 -1694 521 -1626
rect 535 -1694 537 -1626
rect 545 -1694 547 -1626
rect 553 -1694 555 -1626
rect 563 -1694 565 -1626
rect 579 -1694 581 -1626
rect 587 -1694 589 -1626
rect 597 -1694 599 -1626
rect 613 -1694 615 -1626
rect 623 -1694 625 -1626
rect 631 -1694 633 -1626
rect 641 -1694 643 -1626
rect 657 -1694 659 -1626
rect 665 -1694 667 -1626
rect 681 -1694 683 -1626
rect 697 -1694 699 -1626
rect 705 -1694 707 -1626
rect 715 -1694 717 -1626
rect 791 -1694 793 -1626
rect 801 -1694 803 -1626
rect 817 -1694 819 -1626
rect 827 -1694 829 -1626
rect 843 -1694 845 -1626
rect 853 -1694 855 -1626
rect 861 -1694 863 -1626
rect 871 -1694 873 -1626
rect 887 -1694 889 -1626
rect 895 -1694 897 -1626
rect 905 -1694 907 -1626
rect 921 -1694 923 -1626
rect 931 -1694 933 -1626
rect 939 -1694 941 -1626
rect 949 -1694 951 -1626
rect 965 -1694 967 -1626
rect 973 -1694 975 -1626
rect 989 -1694 991 -1626
rect 1005 -1694 1007 -1626
rect 1013 -1694 1015 -1626
rect 1023 -1694 1025 -1626
rect -1229 -1700 -1227 -1698
rect -1219 -1700 -1217 -1698
rect -1203 -1700 -1201 -1698
rect -1193 -1700 -1191 -1698
rect -1185 -1700 -1183 -1698
rect -1175 -1700 -1173 -1698
rect -1159 -1700 -1157 -1698
rect -1151 -1700 -1149 -1698
rect -1141 -1700 -1139 -1698
rect -1057 -1700 -1055 -1698
rect -1047 -1700 -1045 -1698
rect -1031 -1700 -1029 -1698
rect -1021 -1700 -1019 -1698
rect -1005 -1700 -1003 -1698
rect -995 -1700 -993 -1698
rect -987 -1700 -985 -1698
rect -977 -1700 -975 -1698
rect -961 -1700 -959 -1698
rect -953 -1700 -951 -1698
rect -943 -1700 -941 -1698
rect -927 -1700 -925 -1698
rect -917 -1700 -915 -1698
rect -909 -1700 -907 -1698
rect -899 -1700 -897 -1698
rect -883 -1700 -881 -1698
rect -875 -1700 -873 -1698
rect -859 -1700 -857 -1698
rect -843 -1700 -841 -1698
rect -835 -1700 -833 -1698
rect -825 -1700 -823 -1698
rect -749 -1700 -747 -1698
rect -739 -1700 -737 -1698
rect -723 -1700 -721 -1698
rect -713 -1700 -711 -1698
rect -697 -1700 -695 -1698
rect -687 -1700 -685 -1698
rect -679 -1700 -677 -1698
rect -669 -1700 -667 -1698
rect -653 -1700 -651 -1698
rect -645 -1700 -643 -1698
rect -635 -1700 -633 -1698
rect -619 -1700 -617 -1698
rect -609 -1700 -607 -1698
rect -601 -1700 -599 -1698
rect -591 -1700 -589 -1698
rect -575 -1700 -573 -1698
rect -567 -1700 -565 -1698
rect -551 -1700 -549 -1698
rect -535 -1700 -533 -1698
rect -527 -1700 -525 -1698
rect -517 -1700 -515 -1698
rect -441 -1700 -439 -1698
rect -431 -1700 -429 -1698
rect -415 -1700 -413 -1698
rect -405 -1700 -403 -1698
rect -389 -1700 -387 -1698
rect -379 -1700 -377 -1698
rect -371 -1700 -369 -1698
rect -361 -1700 -359 -1698
rect -345 -1700 -343 -1698
rect -337 -1700 -335 -1698
rect -327 -1700 -325 -1698
rect -311 -1700 -309 -1698
rect -301 -1700 -299 -1698
rect -293 -1700 -291 -1698
rect -283 -1700 -281 -1698
rect -267 -1700 -265 -1698
rect -259 -1700 -257 -1698
rect -243 -1700 -241 -1698
rect -227 -1700 -225 -1698
rect -219 -1700 -217 -1698
rect -209 -1700 -207 -1698
rect -133 -1700 -131 -1698
rect -123 -1700 -121 -1698
rect -107 -1700 -105 -1698
rect -97 -1700 -95 -1698
rect -81 -1700 -79 -1698
rect -71 -1700 -69 -1698
rect -63 -1700 -61 -1698
rect -53 -1700 -51 -1698
rect -37 -1700 -35 -1698
rect -29 -1700 -27 -1698
rect -19 -1700 -17 -1698
rect -3 -1700 -1 -1698
rect 7 -1700 9 -1698
rect 15 -1700 17 -1698
rect 25 -1700 27 -1698
rect 41 -1700 43 -1698
rect 49 -1700 51 -1698
rect 65 -1700 67 -1698
rect 81 -1700 83 -1698
rect 89 -1700 91 -1698
rect 99 -1700 101 -1698
rect 175 -1700 177 -1698
rect 185 -1700 187 -1698
rect 201 -1700 203 -1698
rect 211 -1700 213 -1698
rect 227 -1700 229 -1698
rect 237 -1700 239 -1698
rect 245 -1700 247 -1698
rect 255 -1700 257 -1698
rect 271 -1700 273 -1698
rect 279 -1700 281 -1698
rect 289 -1700 291 -1698
rect 305 -1700 307 -1698
rect 315 -1700 317 -1698
rect 323 -1700 325 -1698
rect 333 -1700 335 -1698
rect 349 -1700 351 -1698
rect 357 -1700 359 -1698
rect 373 -1700 375 -1698
rect 389 -1700 391 -1698
rect 397 -1700 399 -1698
rect 407 -1700 409 -1698
rect 483 -1700 485 -1698
rect 493 -1700 495 -1698
rect 509 -1700 511 -1698
rect 519 -1700 521 -1698
rect 535 -1700 537 -1698
rect 545 -1700 547 -1698
rect 553 -1700 555 -1698
rect 563 -1700 565 -1698
rect 579 -1700 581 -1698
rect 587 -1700 589 -1698
rect 597 -1700 599 -1698
rect 613 -1700 615 -1698
rect 623 -1700 625 -1698
rect 631 -1700 633 -1698
rect 641 -1700 643 -1698
rect 657 -1700 659 -1698
rect 665 -1700 667 -1698
rect 681 -1700 683 -1698
rect 697 -1700 699 -1698
rect 705 -1700 707 -1698
rect 715 -1700 717 -1698
rect 791 -1700 793 -1698
rect 801 -1700 803 -1698
rect 817 -1700 819 -1698
rect 827 -1700 829 -1698
rect 843 -1700 845 -1698
rect 853 -1700 855 -1698
rect 861 -1700 863 -1698
rect 871 -1700 873 -1698
rect 887 -1700 889 -1698
rect 895 -1700 897 -1698
rect 905 -1700 907 -1698
rect 921 -1700 923 -1698
rect 931 -1700 933 -1698
rect 939 -1700 941 -1698
rect 949 -1700 951 -1698
rect 965 -1700 967 -1698
rect 973 -1700 975 -1698
rect 989 -1700 991 -1698
rect 1005 -1700 1007 -1698
rect 1013 -1700 1015 -1698
rect 1023 -1700 1025 -1698
rect -1304 -1750 -1302 -1748
rect -1296 -1750 -1294 -1748
rect -1286 -1750 -1284 -1748
rect -1057 -1750 -1055 -1748
rect -1049 -1750 -1047 -1748
rect -1039 -1750 -1037 -1748
rect -749 -1750 -747 -1748
rect -741 -1750 -739 -1748
rect -731 -1750 -729 -1748
rect -441 -1750 -439 -1748
rect -433 -1750 -431 -1748
rect -423 -1750 -421 -1748
rect -133 -1750 -131 -1748
rect -125 -1750 -123 -1748
rect -115 -1750 -113 -1748
rect 175 -1750 177 -1748
rect 183 -1750 185 -1748
rect 193 -1750 195 -1748
rect 483 -1750 485 -1748
rect 491 -1750 493 -1748
rect 501 -1750 503 -1748
rect 791 -1750 793 -1748
rect 799 -1750 801 -1748
rect 809 -1750 811 -1748
rect -1304 -1826 -1302 -1758
rect -1296 -1782 -1294 -1758
rect -1296 -1826 -1294 -1786
rect -1286 -1826 -1284 -1758
rect -1057 -1826 -1055 -1758
rect -1049 -1782 -1047 -1758
rect -1049 -1826 -1047 -1786
rect -1039 -1826 -1037 -1758
rect -749 -1826 -747 -1758
rect -741 -1782 -739 -1758
rect -741 -1826 -739 -1786
rect -731 -1826 -729 -1758
rect -441 -1826 -439 -1758
rect -433 -1782 -431 -1758
rect -433 -1826 -431 -1786
rect -423 -1826 -421 -1758
rect -133 -1826 -131 -1758
rect -125 -1782 -123 -1758
rect -125 -1826 -123 -1786
rect -115 -1826 -113 -1758
rect 175 -1826 177 -1758
rect 183 -1782 185 -1758
rect 183 -1826 185 -1786
rect 193 -1826 195 -1758
rect 483 -1826 485 -1758
rect 491 -1782 493 -1758
rect 491 -1826 493 -1786
rect 501 -1826 503 -1758
rect 791 -1826 793 -1758
rect 799 -1782 801 -1758
rect 799 -1826 801 -1786
rect 809 -1826 811 -1758
rect -1304 -1832 -1302 -1830
rect -1296 -1832 -1294 -1830
rect -1286 -1832 -1284 -1830
rect -1057 -1832 -1055 -1830
rect -1049 -1832 -1047 -1830
rect -1039 -1832 -1037 -1830
rect -749 -1832 -747 -1830
rect -741 -1832 -739 -1830
rect -731 -1832 -729 -1830
rect -441 -1832 -439 -1830
rect -433 -1832 -431 -1830
rect -423 -1832 -421 -1830
rect -133 -1832 -131 -1830
rect -125 -1832 -123 -1830
rect -115 -1832 -113 -1830
rect 175 -1832 177 -1830
rect 183 -1832 185 -1830
rect 193 -1832 195 -1830
rect 483 -1832 485 -1830
rect 491 -1832 493 -1830
rect 501 -1832 503 -1830
rect 791 -1832 793 -1830
rect 799 -1832 801 -1830
rect 809 -1832 811 -1830
rect -1229 -1909 -1227 -1907
rect -1219 -1909 -1217 -1907
rect -1203 -1909 -1201 -1907
rect -1193 -1909 -1191 -1907
rect -1185 -1909 -1183 -1907
rect -1175 -1909 -1173 -1907
rect -1159 -1909 -1157 -1907
rect -1151 -1909 -1149 -1907
rect -1141 -1909 -1139 -1907
rect -1057 -1909 -1055 -1907
rect -1047 -1909 -1045 -1907
rect -1031 -1909 -1029 -1907
rect -1021 -1909 -1019 -1907
rect -1005 -1909 -1003 -1907
rect -995 -1909 -993 -1907
rect -987 -1909 -985 -1907
rect -977 -1909 -975 -1907
rect -961 -1909 -959 -1907
rect -953 -1909 -951 -1907
rect -943 -1909 -941 -1907
rect -927 -1909 -925 -1907
rect -917 -1909 -915 -1907
rect -909 -1909 -907 -1907
rect -899 -1909 -897 -1907
rect -883 -1909 -881 -1907
rect -875 -1909 -873 -1907
rect -859 -1909 -857 -1907
rect -843 -1909 -841 -1907
rect -835 -1909 -833 -1907
rect -825 -1909 -823 -1907
rect -749 -1909 -747 -1907
rect -739 -1909 -737 -1907
rect -723 -1909 -721 -1907
rect -713 -1909 -711 -1907
rect -697 -1909 -695 -1907
rect -687 -1909 -685 -1907
rect -679 -1909 -677 -1907
rect -669 -1909 -667 -1907
rect -653 -1909 -651 -1907
rect -645 -1909 -643 -1907
rect -635 -1909 -633 -1907
rect -619 -1909 -617 -1907
rect -609 -1909 -607 -1907
rect -601 -1909 -599 -1907
rect -591 -1909 -589 -1907
rect -575 -1909 -573 -1907
rect -567 -1909 -565 -1907
rect -551 -1909 -549 -1907
rect -535 -1909 -533 -1907
rect -527 -1909 -525 -1907
rect -517 -1909 -515 -1907
rect -441 -1909 -439 -1907
rect -431 -1909 -429 -1907
rect -415 -1909 -413 -1907
rect -405 -1909 -403 -1907
rect -389 -1909 -387 -1907
rect -379 -1909 -377 -1907
rect -371 -1909 -369 -1907
rect -361 -1909 -359 -1907
rect -345 -1909 -343 -1907
rect -337 -1909 -335 -1907
rect -327 -1909 -325 -1907
rect -311 -1909 -309 -1907
rect -301 -1909 -299 -1907
rect -293 -1909 -291 -1907
rect -283 -1909 -281 -1907
rect -267 -1909 -265 -1907
rect -259 -1909 -257 -1907
rect -243 -1909 -241 -1907
rect -227 -1909 -225 -1907
rect -219 -1909 -217 -1907
rect -209 -1909 -207 -1907
rect -133 -1909 -131 -1907
rect -123 -1909 -121 -1907
rect -107 -1909 -105 -1907
rect -97 -1909 -95 -1907
rect -81 -1909 -79 -1907
rect -71 -1909 -69 -1907
rect -63 -1909 -61 -1907
rect -53 -1909 -51 -1907
rect -37 -1909 -35 -1907
rect -29 -1909 -27 -1907
rect -19 -1909 -17 -1907
rect -3 -1909 -1 -1907
rect 7 -1909 9 -1907
rect 15 -1909 17 -1907
rect 25 -1909 27 -1907
rect 41 -1909 43 -1907
rect 49 -1909 51 -1907
rect 65 -1909 67 -1907
rect 81 -1909 83 -1907
rect 89 -1909 91 -1907
rect 99 -1909 101 -1907
rect 175 -1909 177 -1907
rect 185 -1909 187 -1907
rect 201 -1909 203 -1907
rect 211 -1909 213 -1907
rect 227 -1909 229 -1907
rect 237 -1909 239 -1907
rect 245 -1909 247 -1907
rect 255 -1909 257 -1907
rect 271 -1909 273 -1907
rect 279 -1909 281 -1907
rect 289 -1909 291 -1907
rect 305 -1909 307 -1907
rect 315 -1909 317 -1907
rect 323 -1909 325 -1907
rect 333 -1909 335 -1907
rect 349 -1909 351 -1907
rect 357 -1909 359 -1907
rect 373 -1909 375 -1907
rect 389 -1909 391 -1907
rect 397 -1909 399 -1907
rect 407 -1909 409 -1907
rect 483 -1909 485 -1907
rect 493 -1909 495 -1907
rect 509 -1909 511 -1907
rect 519 -1909 521 -1907
rect 535 -1909 537 -1907
rect 545 -1909 547 -1907
rect 553 -1909 555 -1907
rect 563 -1909 565 -1907
rect 579 -1909 581 -1907
rect 587 -1909 589 -1907
rect 597 -1909 599 -1907
rect 613 -1909 615 -1907
rect 623 -1909 625 -1907
rect 631 -1909 633 -1907
rect 641 -1909 643 -1907
rect 657 -1909 659 -1907
rect 665 -1909 667 -1907
rect 681 -1909 683 -1907
rect 697 -1909 699 -1907
rect 705 -1909 707 -1907
rect 715 -1909 717 -1907
rect 791 -1909 793 -1907
rect 801 -1909 803 -1907
rect 817 -1909 819 -1907
rect 827 -1909 829 -1907
rect 843 -1909 845 -1907
rect 853 -1909 855 -1907
rect 861 -1909 863 -1907
rect 871 -1909 873 -1907
rect 887 -1909 889 -1907
rect 895 -1909 897 -1907
rect 905 -1909 907 -1907
rect 921 -1909 923 -1907
rect 931 -1909 933 -1907
rect 939 -1909 941 -1907
rect 949 -1909 951 -1907
rect 965 -1909 967 -1907
rect 973 -1909 975 -1907
rect 989 -1909 991 -1907
rect 1005 -1909 1007 -1907
rect 1013 -1909 1015 -1907
rect 1023 -1909 1025 -1907
rect -1229 -1985 -1227 -1917
rect -1219 -1985 -1217 -1917
rect -1203 -1985 -1201 -1917
rect -1193 -1985 -1191 -1917
rect -1185 -1985 -1183 -1917
rect -1175 -1985 -1173 -1917
rect -1159 -1985 -1157 -1917
rect -1151 -1985 -1149 -1917
rect -1141 -1985 -1139 -1917
rect -1057 -1985 -1055 -1917
rect -1047 -1985 -1045 -1917
rect -1031 -1985 -1029 -1917
rect -1021 -1985 -1019 -1917
rect -1005 -1985 -1003 -1917
rect -995 -1985 -993 -1917
rect -987 -1985 -985 -1917
rect -977 -1985 -975 -1917
rect -961 -1985 -959 -1917
rect -953 -1985 -951 -1917
rect -943 -1985 -941 -1917
rect -927 -1985 -925 -1917
rect -917 -1985 -915 -1917
rect -909 -1985 -907 -1917
rect -899 -1985 -897 -1917
rect -883 -1985 -881 -1917
rect -875 -1985 -873 -1917
rect -859 -1985 -857 -1917
rect -843 -1985 -841 -1917
rect -835 -1985 -833 -1917
rect -825 -1985 -823 -1917
rect -749 -1985 -747 -1917
rect -739 -1985 -737 -1917
rect -723 -1985 -721 -1917
rect -713 -1985 -711 -1917
rect -697 -1985 -695 -1917
rect -687 -1985 -685 -1917
rect -679 -1985 -677 -1917
rect -669 -1985 -667 -1917
rect -653 -1985 -651 -1917
rect -645 -1985 -643 -1917
rect -635 -1985 -633 -1917
rect -619 -1985 -617 -1917
rect -609 -1985 -607 -1917
rect -601 -1985 -599 -1917
rect -591 -1985 -589 -1917
rect -575 -1985 -573 -1917
rect -567 -1985 -565 -1917
rect -551 -1985 -549 -1917
rect -535 -1985 -533 -1917
rect -527 -1985 -525 -1917
rect -517 -1985 -515 -1917
rect -441 -1985 -439 -1917
rect -431 -1985 -429 -1917
rect -415 -1985 -413 -1917
rect -405 -1985 -403 -1917
rect -389 -1985 -387 -1917
rect -379 -1985 -377 -1917
rect -371 -1985 -369 -1917
rect -361 -1985 -359 -1917
rect -345 -1985 -343 -1917
rect -337 -1985 -335 -1917
rect -327 -1985 -325 -1917
rect -311 -1985 -309 -1917
rect -301 -1985 -299 -1917
rect -293 -1985 -291 -1917
rect -283 -1985 -281 -1917
rect -267 -1985 -265 -1917
rect -259 -1985 -257 -1917
rect -243 -1985 -241 -1917
rect -227 -1985 -225 -1917
rect -219 -1985 -217 -1917
rect -209 -1985 -207 -1917
rect -133 -1985 -131 -1917
rect -123 -1985 -121 -1917
rect -107 -1985 -105 -1917
rect -97 -1985 -95 -1917
rect -81 -1985 -79 -1917
rect -71 -1985 -69 -1917
rect -63 -1985 -61 -1917
rect -53 -1985 -51 -1917
rect -37 -1985 -35 -1917
rect -29 -1985 -27 -1917
rect -19 -1985 -17 -1917
rect -3 -1985 -1 -1917
rect 7 -1985 9 -1917
rect 15 -1985 17 -1917
rect 25 -1985 27 -1917
rect 41 -1985 43 -1917
rect 49 -1985 51 -1917
rect 65 -1985 67 -1917
rect 81 -1985 83 -1917
rect 89 -1985 91 -1917
rect 99 -1985 101 -1917
rect 175 -1985 177 -1917
rect 185 -1985 187 -1917
rect 201 -1985 203 -1917
rect 211 -1985 213 -1917
rect 227 -1985 229 -1917
rect 237 -1985 239 -1917
rect 245 -1985 247 -1917
rect 255 -1985 257 -1917
rect 271 -1985 273 -1917
rect 279 -1985 281 -1917
rect 289 -1985 291 -1917
rect 305 -1985 307 -1917
rect 315 -1985 317 -1917
rect 323 -1985 325 -1917
rect 333 -1985 335 -1917
rect 349 -1985 351 -1917
rect 357 -1985 359 -1917
rect 373 -1985 375 -1917
rect 389 -1985 391 -1917
rect 397 -1985 399 -1917
rect 407 -1985 409 -1917
rect 483 -1985 485 -1917
rect 493 -1985 495 -1917
rect 509 -1985 511 -1917
rect 519 -1985 521 -1917
rect 535 -1985 537 -1917
rect 545 -1985 547 -1917
rect 553 -1985 555 -1917
rect 563 -1985 565 -1917
rect 579 -1985 581 -1917
rect 587 -1985 589 -1917
rect 597 -1985 599 -1917
rect 613 -1985 615 -1917
rect 623 -1985 625 -1917
rect 631 -1985 633 -1917
rect 641 -1985 643 -1917
rect 657 -1985 659 -1917
rect 665 -1985 667 -1917
rect 681 -1985 683 -1917
rect 697 -1985 699 -1917
rect 705 -1985 707 -1917
rect 715 -1985 717 -1917
rect 791 -1985 793 -1917
rect 801 -1985 803 -1917
rect 817 -1985 819 -1917
rect 827 -1985 829 -1917
rect 843 -1985 845 -1917
rect 853 -1985 855 -1917
rect 861 -1985 863 -1917
rect 871 -1985 873 -1917
rect 887 -1985 889 -1917
rect 895 -1985 897 -1917
rect 905 -1985 907 -1917
rect 921 -1985 923 -1917
rect 931 -1985 933 -1917
rect 939 -1985 941 -1917
rect 949 -1985 951 -1917
rect 965 -1985 967 -1917
rect 973 -1985 975 -1917
rect 989 -1985 991 -1917
rect 1005 -1985 1007 -1917
rect 1013 -1985 1015 -1917
rect 1023 -1985 1025 -1917
rect -1229 -1991 -1227 -1989
rect -1219 -1991 -1217 -1989
rect -1203 -1991 -1201 -1989
rect -1193 -1991 -1191 -1989
rect -1185 -1991 -1183 -1989
rect -1175 -1991 -1173 -1989
rect -1159 -1991 -1157 -1989
rect -1151 -1991 -1149 -1989
rect -1141 -1991 -1139 -1989
rect -1057 -1991 -1055 -1989
rect -1047 -1991 -1045 -1989
rect -1031 -1991 -1029 -1989
rect -1021 -1991 -1019 -1989
rect -1005 -1991 -1003 -1989
rect -995 -1991 -993 -1989
rect -987 -1991 -985 -1989
rect -977 -1991 -975 -1989
rect -961 -1991 -959 -1989
rect -953 -1991 -951 -1989
rect -943 -1991 -941 -1989
rect -927 -1991 -925 -1989
rect -917 -1991 -915 -1989
rect -909 -1991 -907 -1989
rect -899 -1991 -897 -1989
rect -883 -1991 -881 -1989
rect -875 -1991 -873 -1989
rect -859 -1991 -857 -1989
rect -843 -1991 -841 -1989
rect -835 -1991 -833 -1989
rect -825 -1991 -823 -1989
rect -749 -1991 -747 -1989
rect -739 -1991 -737 -1989
rect -723 -1991 -721 -1989
rect -713 -1991 -711 -1989
rect -697 -1991 -695 -1989
rect -687 -1991 -685 -1989
rect -679 -1991 -677 -1989
rect -669 -1991 -667 -1989
rect -653 -1991 -651 -1989
rect -645 -1991 -643 -1989
rect -635 -1991 -633 -1989
rect -619 -1991 -617 -1989
rect -609 -1991 -607 -1989
rect -601 -1991 -599 -1989
rect -591 -1991 -589 -1989
rect -575 -1991 -573 -1989
rect -567 -1991 -565 -1989
rect -551 -1991 -549 -1989
rect -535 -1991 -533 -1989
rect -527 -1991 -525 -1989
rect -517 -1991 -515 -1989
rect -441 -1991 -439 -1989
rect -431 -1991 -429 -1989
rect -415 -1991 -413 -1989
rect -405 -1991 -403 -1989
rect -389 -1991 -387 -1989
rect -379 -1991 -377 -1989
rect -371 -1991 -369 -1989
rect -361 -1991 -359 -1989
rect -345 -1991 -343 -1989
rect -337 -1991 -335 -1989
rect -327 -1991 -325 -1989
rect -311 -1991 -309 -1989
rect -301 -1991 -299 -1989
rect -293 -1991 -291 -1989
rect -283 -1991 -281 -1989
rect -267 -1991 -265 -1989
rect -259 -1991 -257 -1989
rect -243 -1991 -241 -1989
rect -227 -1991 -225 -1989
rect -219 -1991 -217 -1989
rect -209 -1991 -207 -1989
rect -133 -1991 -131 -1989
rect -123 -1991 -121 -1989
rect -107 -1991 -105 -1989
rect -97 -1991 -95 -1989
rect -81 -1991 -79 -1989
rect -71 -1991 -69 -1989
rect -63 -1991 -61 -1989
rect -53 -1991 -51 -1989
rect -37 -1991 -35 -1989
rect -29 -1991 -27 -1989
rect -19 -1991 -17 -1989
rect -3 -1991 -1 -1989
rect 7 -1991 9 -1989
rect 15 -1991 17 -1989
rect 25 -1991 27 -1989
rect 41 -1991 43 -1989
rect 49 -1991 51 -1989
rect 65 -1991 67 -1989
rect 81 -1991 83 -1989
rect 89 -1991 91 -1989
rect 99 -1991 101 -1989
rect 175 -1991 177 -1989
rect 185 -1991 187 -1989
rect 201 -1991 203 -1989
rect 211 -1991 213 -1989
rect 227 -1991 229 -1989
rect 237 -1991 239 -1989
rect 245 -1991 247 -1989
rect 255 -1991 257 -1989
rect 271 -1991 273 -1989
rect 279 -1991 281 -1989
rect 289 -1991 291 -1989
rect 305 -1991 307 -1989
rect 315 -1991 317 -1989
rect 323 -1991 325 -1989
rect 333 -1991 335 -1989
rect 349 -1991 351 -1989
rect 357 -1991 359 -1989
rect 373 -1991 375 -1989
rect 389 -1991 391 -1989
rect 397 -1991 399 -1989
rect 407 -1991 409 -1989
rect 483 -1991 485 -1989
rect 493 -1991 495 -1989
rect 509 -1991 511 -1989
rect 519 -1991 521 -1989
rect 535 -1991 537 -1989
rect 545 -1991 547 -1989
rect 553 -1991 555 -1989
rect 563 -1991 565 -1989
rect 579 -1991 581 -1989
rect 587 -1991 589 -1989
rect 597 -1991 599 -1989
rect 613 -1991 615 -1989
rect 623 -1991 625 -1989
rect 631 -1991 633 -1989
rect 641 -1991 643 -1989
rect 657 -1991 659 -1989
rect 665 -1991 667 -1989
rect 681 -1991 683 -1989
rect 697 -1991 699 -1989
rect 705 -1991 707 -1989
rect 715 -1991 717 -1989
rect 791 -1991 793 -1989
rect 801 -1991 803 -1989
rect 817 -1991 819 -1989
rect 827 -1991 829 -1989
rect 843 -1991 845 -1989
rect 853 -1991 855 -1989
rect 861 -1991 863 -1989
rect 871 -1991 873 -1989
rect 887 -1991 889 -1989
rect 895 -1991 897 -1989
rect 905 -1991 907 -1989
rect 921 -1991 923 -1989
rect 931 -1991 933 -1989
rect 939 -1991 941 -1989
rect 949 -1991 951 -1989
rect 965 -1991 967 -1989
rect 973 -1991 975 -1989
rect 989 -1991 991 -1989
rect 1005 -1991 1007 -1989
rect 1013 -1991 1015 -1989
rect 1023 -1991 1025 -1989
rect -1304 -2072 -1302 -2070
rect -1296 -2072 -1294 -2070
rect -1286 -2072 -1284 -2070
rect -1057 -2072 -1055 -2070
rect -1049 -2072 -1047 -2070
rect -1039 -2072 -1037 -2070
rect -749 -2072 -747 -2070
rect -741 -2072 -739 -2070
rect -731 -2072 -729 -2070
rect -441 -2072 -439 -2070
rect -433 -2072 -431 -2070
rect -423 -2072 -421 -2070
rect -133 -2072 -131 -2070
rect -125 -2072 -123 -2070
rect -115 -2072 -113 -2070
rect 175 -2072 177 -2070
rect 183 -2072 185 -2070
rect 193 -2072 195 -2070
rect 483 -2072 485 -2070
rect 491 -2072 493 -2070
rect 501 -2072 503 -2070
rect 791 -2072 793 -2070
rect 799 -2072 801 -2070
rect 809 -2072 811 -2070
rect -1304 -2148 -1302 -2080
rect -1296 -2104 -1294 -2080
rect -1296 -2148 -1294 -2108
rect -1286 -2148 -1284 -2080
rect -1057 -2148 -1055 -2080
rect -1049 -2104 -1047 -2080
rect -1049 -2148 -1047 -2108
rect -1039 -2148 -1037 -2080
rect -749 -2148 -747 -2080
rect -741 -2104 -739 -2080
rect -741 -2148 -739 -2108
rect -731 -2148 -729 -2080
rect -441 -2148 -439 -2080
rect -433 -2104 -431 -2080
rect -433 -2148 -431 -2108
rect -423 -2148 -421 -2080
rect -133 -2148 -131 -2080
rect -125 -2104 -123 -2080
rect -125 -2148 -123 -2108
rect -115 -2148 -113 -2080
rect 175 -2148 177 -2080
rect 183 -2104 185 -2080
rect 183 -2148 185 -2108
rect 193 -2148 195 -2080
rect 483 -2148 485 -2080
rect 491 -2104 493 -2080
rect 491 -2148 493 -2108
rect 501 -2148 503 -2080
rect 791 -2148 793 -2080
rect 799 -2104 801 -2080
rect 799 -2148 801 -2108
rect 809 -2148 811 -2080
rect -1304 -2154 -1302 -2152
rect -1296 -2154 -1294 -2152
rect -1286 -2154 -1284 -2152
rect -1057 -2154 -1055 -2152
rect -1049 -2154 -1047 -2152
rect -1039 -2154 -1037 -2152
rect -749 -2154 -747 -2152
rect -741 -2154 -739 -2152
rect -731 -2154 -729 -2152
rect -441 -2154 -439 -2152
rect -433 -2154 -431 -2152
rect -423 -2154 -421 -2152
rect -133 -2154 -131 -2152
rect -125 -2154 -123 -2152
rect -115 -2154 -113 -2152
rect 175 -2154 177 -2152
rect 183 -2154 185 -2152
rect 193 -2154 195 -2152
rect 483 -2154 485 -2152
rect 491 -2154 493 -2152
rect 501 -2154 503 -2152
rect 791 -2154 793 -2152
rect 799 -2154 801 -2152
rect 809 -2154 811 -2152
rect -1229 -2231 -1227 -2229
rect -1219 -2231 -1217 -2229
rect -1203 -2231 -1201 -2229
rect -1193 -2231 -1191 -2229
rect -1185 -2231 -1183 -2229
rect -1175 -2231 -1173 -2229
rect -1159 -2231 -1157 -2229
rect -1151 -2231 -1149 -2229
rect -1141 -2231 -1139 -2229
rect -1057 -2231 -1055 -2229
rect -1047 -2231 -1045 -2229
rect -1031 -2231 -1029 -2229
rect -1021 -2231 -1019 -2229
rect -1005 -2231 -1003 -2229
rect -995 -2231 -993 -2229
rect -987 -2231 -985 -2229
rect -977 -2231 -975 -2229
rect -961 -2231 -959 -2229
rect -953 -2231 -951 -2229
rect -943 -2231 -941 -2229
rect -927 -2231 -925 -2229
rect -917 -2231 -915 -2229
rect -909 -2231 -907 -2229
rect -899 -2231 -897 -2229
rect -883 -2231 -881 -2229
rect -875 -2231 -873 -2229
rect -859 -2231 -857 -2229
rect -843 -2231 -841 -2229
rect -835 -2231 -833 -2229
rect -825 -2231 -823 -2229
rect -749 -2231 -747 -2229
rect -739 -2231 -737 -2229
rect -723 -2231 -721 -2229
rect -713 -2231 -711 -2229
rect -697 -2231 -695 -2229
rect -687 -2231 -685 -2229
rect -679 -2231 -677 -2229
rect -669 -2231 -667 -2229
rect -653 -2231 -651 -2229
rect -645 -2231 -643 -2229
rect -635 -2231 -633 -2229
rect -619 -2231 -617 -2229
rect -609 -2231 -607 -2229
rect -601 -2231 -599 -2229
rect -591 -2231 -589 -2229
rect -575 -2231 -573 -2229
rect -567 -2231 -565 -2229
rect -551 -2231 -549 -2229
rect -535 -2231 -533 -2229
rect -527 -2231 -525 -2229
rect -517 -2231 -515 -2229
rect -441 -2231 -439 -2229
rect -431 -2231 -429 -2229
rect -415 -2231 -413 -2229
rect -405 -2231 -403 -2229
rect -389 -2231 -387 -2229
rect -379 -2231 -377 -2229
rect -371 -2231 -369 -2229
rect -361 -2231 -359 -2229
rect -345 -2231 -343 -2229
rect -337 -2231 -335 -2229
rect -327 -2231 -325 -2229
rect -311 -2231 -309 -2229
rect -301 -2231 -299 -2229
rect -293 -2231 -291 -2229
rect -283 -2231 -281 -2229
rect -267 -2231 -265 -2229
rect -259 -2231 -257 -2229
rect -243 -2231 -241 -2229
rect -227 -2231 -225 -2229
rect -219 -2231 -217 -2229
rect -209 -2231 -207 -2229
rect -133 -2231 -131 -2229
rect -123 -2231 -121 -2229
rect -107 -2231 -105 -2229
rect -97 -2231 -95 -2229
rect -81 -2231 -79 -2229
rect -71 -2231 -69 -2229
rect -63 -2231 -61 -2229
rect -53 -2231 -51 -2229
rect -37 -2231 -35 -2229
rect -29 -2231 -27 -2229
rect -19 -2231 -17 -2229
rect -3 -2231 -1 -2229
rect 7 -2231 9 -2229
rect 15 -2231 17 -2229
rect 25 -2231 27 -2229
rect 41 -2231 43 -2229
rect 49 -2231 51 -2229
rect 65 -2231 67 -2229
rect 81 -2231 83 -2229
rect 89 -2231 91 -2229
rect 99 -2231 101 -2229
rect 175 -2231 177 -2229
rect 185 -2231 187 -2229
rect 201 -2231 203 -2229
rect 211 -2231 213 -2229
rect 227 -2231 229 -2229
rect 237 -2231 239 -2229
rect 245 -2231 247 -2229
rect 255 -2231 257 -2229
rect 271 -2231 273 -2229
rect 279 -2231 281 -2229
rect 289 -2231 291 -2229
rect 305 -2231 307 -2229
rect 315 -2231 317 -2229
rect 323 -2231 325 -2229
rect 333 -2231 335 -2229
rect 349 -2231 351 -2229
rect 357 -2231 359 -2229
rect 373 -2231 375 -2229
rect 389 -2231 391 -2229
rect 397 -2231 399 -2229
rect 407 -2231 409 -2229
rect 483 -2231 485 -2229
rect 493 -2231 495 -2229
rect 509 -2231 511 -2229
rect 519 -2231 521 -2229
rect 535 -2231 537 -2229
rect 545 -2231 547 -2229
rect 553 -2231 555 -2229
rect 563 -2231 565 -2229
rect 579 -2231 581 -2229
rect 587 -2231 589 -2229
rect 597 -2231 599 -2229
rect 613 -2231 615 -2229
rect 623 -2231 625 -2229
rect 631 -2231 633 -2229
rect 641 -2231 643 -2229
rect 657 -2231 659 -2229
rect 665 -2231 667 -2229
rect 681 -2231 683 -2229
rect 697 -2231 699 -2229
rect 705 -2231 707 -2229
rect 715 -2231 717 -2229
rect 791 -2231 793 -2229
rect 801 -2231 803 -2229
rect 817 -2231 819 -2229
rect 827 -2231 829 -2229
rect 843 -2231 845 -2229
rect 853 -2231 855 -2229
rect 861 -2231 863 -2229
rect 871 -2231 873 -2229
rect 887 -2231 889 -2229
rect 895 -2231 897 -2229
rect 905 -2231 907 -2229
rect 921 -2231 923 -2229
rect 931 -2231 933 -2229
rect 939 -2231 941 -2229
rect 949 -2231 951 -2229
rect 965 -2231 967 -2229
rect 973 -2231 975 -2229
rect 989 -2231 991 -2229
rect 1005 -2231 1007 -2229
rect 1013 -2231 1015 -2229
rect 1023 -2231 1025 -2229
rect -1229 -2307 -1227 -2239
rect -1219 -2307 -1217 -2239
rect -1203 -2307 -1201 -2239
rect -1193 -2307 -1191 -2239
rect -1185 -2307 -1183 -2239
rect -1175 -2307 -1173 -2239
rect -1159 -2307 -1157 -2239
rect -1151 -2307 -1149 -2239
rect -1141 -2307 -1139 -2239
rect -1057 -2307 -1055 -2239
rect -1047 -2307 -1045 -2239
rect -1031 -2307 -1029 -2239
rect -1021 -2307 -1019 -2239
rect -1005 -2307 -1003 -2239
rect -995 -2307 -993 -2239
rect -987 -2307 -985 -2239
rect -977 -2307 -975 -2239
rect -961 -2307 -959 -2239
rect -953 -2307 -951 -2239
rect -943 -2307 -941 -2239
rect -927 -2307 -925 -2239
rect -917 -2307 -915 -2239
rect -909 -2307 -907 -2239
rect -899 -2307 -897 -2239
rect -883 -2307 -881 -2239
rect -875 -2307 -873 -2239
rect -859 -2307 -857 -2239
rect -843 -2307 -841 -2239
rect -835 -2307 -833 -2239
rect -825 -2307 -823 -2239
rect -749 -2307 -747 -2239
rect -739 -2307 -737 -2239
rect -723 -2307 -721 -2239
rect -713 -2307 -711 -2239
rect -697 -2307 -695 -2239
rect -687 -2307 -685 -2239
rect -679 -2307 -677 -2239
rect -669 -2307 -667 -2239
rect -653 -2307 -651 -2239
rect -645 -2307 -643 -2239
rect -635 -2307 -633 -2239
rect -619 -2307 -617 -2239
rect -609 -2307 -607 -2239
rect -601 -2307 -599 -2239
rect -591 -2307 -589 -2239
rect -575 -2307 -573 -2239
rect -567 -2307 -565 -2239
rect -551 -2307 -549 -2239
rect -535 -2307 -533 -2239
rect -527 -2307 -525 -2239
rect -517 -2307 -515 -2239
rect -441 -2307 -439 -2239
rect -431 -2307 -429 -2239
rect -415 -2307 -413 -2239
rect -405 -2307 -403 -2239
rect -389 -2307 -387 -2239
rect -379 -2307 -377 -2239
rect -371 -2307 -369 -2239
rect -361 -2307 -359 -2239
rect -345 -2307 -343 -2239
rect -337 -2307 -335 -2239
rect -327 -2307 -325 -2239
rect -311 -2307 -309 -2239
rect -301 -2307 -299 -2239
rect -293 -2307 -291 -2239
rect -283 -2307 -281 -2239
rect -267 -2307 -265 -2239
rect -259 -2307 -257 -2239
rect -243 -2307 -241 -2239
rect -227 -2307 -225 -2239
rect -219 -2307 -217 -2239
rect -209 -2307 -207 -2239
rect -133 -2307 -131 -2239
rect -123 -2307 -121 -2239
rect -107 -2307 -105 -2239
rect -97 -2307 -95 -2239
rect -81 -2307 -79 -2239
rect -71 -2307 -69 -2239
rect -63 -2307 -61 -2239
rect -53 -2307 -51 -2239
rect -37 -2307 -35 -2239
rect -29 -2307 -27 -2239
rect -19 -2307 -17 -2239
rect -3 -2307 -1 -2239
rect 7 -2307 9 -2239
rect 15 -2307 17 -2239
rect 25 -2307 27 -2239
rect 41 -2307 43 -2239
rect 49 -2307 51 -2239
rect 65 -2307 67 -2239
rect 81 -2307 83 -2239
rect 89 -2307 91 -2239
rect 99 -2307 101 -2239
rect 175 -2307 177 -2239
rect 185 -2307 187 -2239
rect 201 -2307 203 -2239
rect 211 -2307 213 -2239
rect 227 -2307 229 -2239
rect 237 -2307 239 -2239
rect 245 -2307 247 -2239
rect 255 -2307 257 -2239
rect 271 -2307 273 -2239
rect 279 -2307 281 -2239
rect 289 -2307 291 -2239
rect 305 -2307 307 -2239
rect 315 -2307 317 -2239
rect 323 -2307 325 -2239
rect 333 -2307 335 -2239
rect 349 -2307 351 -2239
rect 357 -2307 359 -2239
rect 373 -2307 375 -2239
rect 389 -2307 391 -2239
rect 397 -2307 399 -2239
rect 407 -2307 409 -2239
rect 483 -2307 485 -2239
rect 493 -2307 495 -2239
rect 509 -2307 511 -2239
rect 519 -2307 521 -2239
rect 535 -2307 537 -2239
rect 545 -2307 547 -2239
rect 553 -2307 555 -2239
rect 563 -2307 565 -2239
rect 579 -2307 581 -2239
rect 587 -2307 589 -2239
rect 597 -2307 599 -2239
rect 613 -2307 615 -2239
rect 623 -2307 625 -2239
rect 631 -2307 633 -2239
rect 641 -2307 643 -2239
rect 657 -2307 659 -2239
rect 665 -2307 667 -2239
rect 681 -2307 683 -2239
rect 697 -2307 699 -2239
rect 705 -2307 707 -2239
rect 715 -2307 717 -2239
rect 791 -2307 793 -2239
rect 801 -2307 803 -2239
rect 817 -2307 819 -2239
rect 827 -2307 829 -2239
rect 843 -2307 845 -2239
rect 853 -2307 855 -2239
rect 861 -2307 863 -2239
rect 871 -2307 873 -2239
rect 887 -2307 889 -2239
rect 895 -2307 897 -2239
rect 905 -2307 907 -2239
rect 921 -2307 923 -2239
rect 931 -2307 933 -2239
rect 939 -2307 941 -2239
rect 949 -2307 951 -2239
rect 965 -2307 967 -2239
rect 973 -2307 975 -2239
rect 989 -2307 991 -2239
rect 1005 -2307 1007 -2239
rect 1013 -2307 1015 -2239
rect 1023 -2307 1025 -2239
rect -1229 -2313 -1227 -2311
rect -1219 -2313 -1217 -2311
rect -1203 -2313 -1201 -2311
rect -1193 -2313 -1191 -2311
rect -1185 -2313 -1183 -2311
rect -1175 -2313 -1173 -2311
rect -1159 -2313 -1157 -2311
rect -1151 -2313 -1149 -2311
rect -1141 -2313 -1139 -2311
rect -1057 -2313 -1055 -2311
rect -1047 -2313 -1045 -2311
rect -1031 -2313 -1029 -2311
rect -1021 -2313 -1019 -2311
rect -1005 -2313 -1003 -2311
rect -995 -2313 -993 -2311
rect -987 -2313 -985 -2311
rect -977 -2313 -975 -2311
rect -961 -2313 -959 -2311
rect -953 -2313 -951 -2311
rect -943 -2313 -941 -2311
rect -927 -2313 -925 -2311
rect -917 -2313 -915 -2311
rect -909 -2313 -907 -2311
rect -899 -2313 -897 -2311
rect -883 -2313 -881 -2311
rect -875 -2313 -873 -2311
rect -859 -2313 -857 -2311
rect -843 -2313 -841 -2311
rect -835 -2313 -833 -2311
rect -825 -2313 -823 -2311
rect -749 -2313 -747 -2311
rect -739 -2313 -737 -2311
rect -723 -2313 -721 -2311
rect -713 -2313 -711 -2311
rect -697 -2313 -695 -2311
rect -687 -2313 -685 -2311
rect -679 -2313 -677 -2311
rect -669 -2313 -667 -2311
rect -653 -2313 -651 -2311
rect -645 -2313 -643 -2311
rect -635 -2313 -633 -2311
rect -619 -2313 -617 -2311
rect -609 -2313 -607 -2311
rect -601 -2313 -599 -2311
rect -591 -2313 -589 -2311
rect -575 -2313 -573 -2311
rect -567 -2313 -565 -2311
rect -551 -2313 -549 -2311
rect -535 -2313 -533 -2311
rect -527 -2313 -525 -2311
rect -517 -2313 -515 -2311
rect -441 -2313 -439 -2311
rect -431 -2313 -429 -2311
rect -415 -2313 -413 -2311
rect -405 -2313 -403 -2311
rect -389 -2313 -387 -2311
rect -379 -2313 -377 -2311
rect -371 -2313 -369 -2311
rect -361 -2313 -359 -2311
rect -345 -2313 -343 -2311
rect -337 -2313 -335 -2311
rect -327 -2313 -325 -2311
rect -311 -2313 -309 -2311
rect -301 -2313 -299 -2311
rect -293 -2313 -291 -2311
rect -283 -2313 -281 -2311
rect -267 -2313 -265 -2311
rect -259 -2313 -257 -2311
rect -243 -2313 -241 -2311
rect -227 -2313 -225 -2311
rect -219 -2313 -217 -2311
rect -209 -2313 -207 -2311
rect -133 -2313 -131 -2311
rect -123 -2313 -121 -2311
rect -107 -2313 -105 -2311
rect -97 -2313 -95 -2311
rect -81 -2313 -79 -2311
rect -71 -2313 -69 -2311
rect -63 -2313 -61 -2311
rect -53 -2313 -51 -2311
rect -37 -2313 -35 -2311
rect -29 -2313 -27 -2311
rect -19 -2313 -17 -2311
rect -3 -2313 -1 -2311
rect 7 -2313 9 -2311
rect 15 -2313 17 -2311
rect 25 -2313 27 -2311
rect 41 -2313 43 -2311
rect 49 -2313 51 -2311
rect 65 -2313 67 -2311
rect 81 -2313 83 -2311
rect 89 -2313 91 -2311
rect 99 -2313 101 -2311
rect 175 -2313 177 -2311
rect 185 -2313 187 -2311
rect 201 -2313 203 -2311
rect 211 -2313 213 -2311
rect 227 -2313 229 -2311
rect 237 -2313 239 -2311
rect 245 -2313 247 -2311
rect 255 -2313 257 -2311
rect 271 -2313 273 -2311
rect 279 -2313 281 -2311
rect 289 -2313 291 -2311
rect 305 -2313 307 -2311
rect 315 -2313 317 -2311
rect 323 -2313 325 -2311
rect 333 -2313 335 -2311
rect 349 -2313 351 -2311
rect 357 -2313 359 -2311
rect 373 -2313 375 -2311
rect 389 -2313 391 -2311
rect 397 -2313 399 -2311
rect 407 -2313 409 -2311
rect 483 -2313 485 -2311
rect 493 -2313 495 -2311
rect 509 -2313 511 -2311
rect 519 -2313 521 -2311
rect 535 -2313 537 -2311
rect 545 -2313 547 -2311
rect 553 -2313 555 -2311
rect 563 -2313 565 -2311
rect 579 -2313 581 -2311
rect 587 -2313 589 -2311
rect 597 -2313 599 -2311
rect 613 -2313 615 -2311
rect 623 -2313 625 -2311
rect 631 -2313 633 -2311
rect 641 -2313 643 -2311
rect 657 -2313 659 -2311
rect 665 -2313 667 -2311
rect 681 -2313 683 -2311
rect 697 -2313 699 -2311
rect 705 -2313 707 -2311
rect 715 -2313 717 -2311
rect 791 -2313 793 -2311
rect 801 -2313 803 -2311
rect 817 -2313 819 -2311
rect 827 -2313 829 -2311
rect 843 -2313 845 -2311
rect 853 -2313 855 -2311
rect 861 -2313 863 -2311
rect 871 -2313 873 -2311
rect 887 -2313 889 -2311
rect 895 -2313 897 -2311
rect 905 -2313 907 -2311
rect 921 -2313 923 -2311
rect 931 -2313 933 -2311
rect 939 -2313 941 -2311
rect 949 -2313 951 -2311
rect 965 -2313 967 -2311
rect 973 -2313 975 -2311
rect 989 -2313 991 -2311
rect 1005 -2313 1007 -2311
rect 1013 -2313 1015 -2311
rect 1023 -2313 1025 -2311
rect -1304 -2363 -1302 -2361
rect -1296 -2363 -1294 -2361
rect -1286 -2363 -1284 -2361
rect -1057 -2363 -1055 -2361
rect -1049 -2363 -1047 -2361
rect -1039 -2363 -1037 -2361
rect -749 -2363 -747 -2361
rect -741 -2363 -739 -2361
rect -731 -2363 -729 -2361
rect -441 -2363 -439 -2361
rect -433 -2363 -431 -2361
rect -423 -2363 -421 -2361
rect -133 -2363 -131 -2361
rect -125 -2363 -123 -2361
rect -115 -2363 -113 -2361
rect 175 -2363 177 -2361
rect 183 -2363 185 -2361
rect 193 -2363 195 -2361
rect 483 -2363 485 -2361
rect 491 -2363 493 -2361
rect 501 -2363 503 -2361
rect 791 -2363 793 -2361
rect 799 -2363 801 -2361
rect 809 -2363 811 -2361
rect -1304 -2439 -1302 -2371
rect -1296 -2395 -1294 -2371
rect -1296 -2439 -1294 -2399
rect -1286 -2439 -1284 -2371
rect -1057 -2439 -1055 -2371
rect -1049 -2395 -1047 -2371
rect -1049 -2439 -1047 -2399
rect -1039 -2439 -1037 -2371
rect -749 -2439 -747 -2371
rect -741 -2395 -739 -2371
rect -741 -2439 -739 -2399
rect -731 -2439 -729 -2371
rect -441 -2439 -439 -2371
rect -433 -2395 -431 -2371
rect -433 -2439 -431 -2399
rect -423 -2439 -421 -2371
rect -133 -2439 -131 -2371
rect -125 -2395 -123 -2371
rect -125 -2439 -123 -2399
rect -115 -2439 -113 -2371
rect 175 -2439 177 -2371
rect 183 -2395 185 -2371
rect 183 -2439 185 -2399
rect 193 -2439 195 -2371
rect 483 -2439 485 -2371
rect 491 -2395 493 -2371
rect 491 -2439 493 -2399
rect 501 -2439 503 -2371
rect 791 -2439 793 -2371
rect 799 -2395 801 -2371
rect 799 -2439 801 -2399
rect 809 -2439 811 -2371
rect -1304 -2445 -1302 -2443
rect -1296 -2445 -1294 -2443
rect -1286 -2445 -1284 -2443
rect -1057 -2445 -1055 -2443
rect -1049 -2445 -1047 -2443
rect -1039 -2445 -1037 -2443
rect -749 -2445 -747 -2443
rect -741 -2445 -739 -2443
rect -731 -2445 -729 -2443
rect -441 -2445 -439 -2443
rect -433 -2445 -431 -2443
rect -423 -2445 -421 -2443
rect -133 -2445 -131 -2443
rect -125 -2445 -123 -2443
rect -115 -2445 -113 -2443
rect 175 -2445 177 -2443
rect 183 -2445 185 -2443
rect 193 -2445 195 -2443
rect 483 -2445 485 -2443
rect 491 -2445 493 -2443
rect 501 -2445 503 -2443
rect 791 -2445 793 -2443
rect 799 -2445 801 -2443
rect 809 -2445 811 -2443
rect -1229 -2522 -1227 -2520
rect -1219 -2522 -1217 -2520
rect -1203 -2522 -1201 -2520
rect -1193 -2522 -1191 -2520
rect -1185 -2522 -1183 -2520
rect -1175 -2522 -1173 -2520
rect -1159 -2522 -1157 -2520
rect -1151 -2522 -1149 -2520
rect -1141 -2522 -1139 -2520
rect -1057 -2522 -1055 -2520
rect -1047 -2522 -1045 -2520
rect -1031 -2522 -1029 -2520
rect -1021 -2522 -1019 -2520
rect -1005 -2522 -1003 -2520
rect -995 -2522 -993 -2520
rect -987 -2522 -985 -2520
rect -977 -2522 -975 -2520
rect -961 -2522 -959 -2520
rect -953 -2522 -951 -2520
rect -943 -2522 -941 -2520
rect -927 -2522 -925 -2520
rect -917 -2522 -915 -2520
rect -909 -2522 -907 -2520
rect -899 -2522 -897 -2520
rect -883 -2522 -881 -2520
rect -875 -2522 -873 -2520
rect -859 -2522 -857 -2520
rect -843 -2522 -841 -2520
rect -835 -2522 -833 -2520
rect -825 -2522 -823 -2520
rect -749 -2522 -747 -2520
rect -739 -2522 -737 -2520
rect -723 -2522 -721 -2520
rect -713 -2522 -711 -2520
rect -697 -2522 -695 -2520
rect -687 -2522 -685 -2520
rect -679 -2522 -677 -2520
rect -669 -2522 -667 -2520
rect -653 -2522 -651 -2520
rect -645 -2522 -643 -2520
rect -635 -2522 -633 -2520
rect -619 -2522 -617 -2520
rect -609 -2522 -607 -2520
rect -601 -2522 -599 -2520
rect -591 -2522 -589 -2520
rect -575 -2522 -573 -2520
rect -567 -2522 -565 -2520
rect -551 -2522 -549 -2520
rect -535 -2522 -533 -2520
rect -527 -2522 -525 -2520
rect -517 -2522 -515 -2520
rect -441 -2522 -439 -2520
rect -431 -2522 -429 -2520
rect -415 -2522 -413 -2520
rect -405 -2522 -403 -2520
rect -389 -2522 -387 -2520
rect -379 -2522 -377 -2520
rect -371 -2522 -369 -2520
rect -361 -2522 -359 -2520
rect -345 -2522 -343 -2520
rect -337 -2522 -335 -2520
rect -327 -2522 -325 -2520
rect -311 -2522 -309 -2520
rect -301 -2522 -299 -2520
rect -293 -2522 -291 -2520
rect -283 -2522 -281 -2520
rect -267 -2522 -265 -2520
rect -259 -2522 -257 -2520
rect -243 -2522 -241 -2520
rect -227 -2522 -225 -2520
rect -219 -2522 -217 -2520
rect -209 -2522 -207 -2520
rect -133 -2522 -131 -2520
rect -123 -2522 -121 -2520
rect -107 -2522 -105 -2520
rect -97 -2522 -95 -2520
rect -81 -2522 -79 -2520
rect -71 -2522 -69 -2520
rect -63 -2522 -61 -2520
rect -53 -2522 -51 -2520
rect -37 -2522 -35 -2520
rect -29 -2522 -27 -2520
rect -19 -2522 -17 -2520
rect -3 -2522 -1 -2520
rect 7 -2522 9 -2520
rect 15 -2522 17 -2520
rect 25 -2522 27 -2520
rect 41 -2522 43 -2520
rect 49 -2522 51 -2520
rect 65 -2522 67 -2520
rect 81 -2522 83 -2520
rect 89 -2522 91 -2520
rect 99 -2522 101 -2520
rect 175 -2522 177 -2520
rect 185 -2522 187 -2520
rect 201 -2522 203 -2520
rect 211 -2522 213 -2520
rect 227 -2522 229 -2520
rect 237 -2522 239 -2520
rect 245 -2522 247 -2520
rect 255 -2522 257 -2520
rect 271 -2522 273 -2520
rect 279 -2522 281 -2520
rect 289 -2522 291 -2520
rect 305 -2522 307 -2520
rect 315 -2522 317 -2520
rect 323 -2522 325 -2520
rect 333 -2522 335 -2520
rect 349 -2522 351 -2520
rect 357 -2522 359 -2520
rect 373 -2522 375 -2520
rect 389 -2522 391 -2520
rect 397 -2522 399 -2520
rect 407 -2522 409 -2520
rect 483 -2522 485 -2520
rect 493 -2522 495 -2520
rect 509 -2522 511 -2520
rect 519 -2522 521 -2520
rect 535 -2522 537 -2520
rect 545 -2522 547 -2520
rect 553 -2522 555 -2520
rect 563 -2522 565 -2520
rect 579 -2522 581 -2520
rect 587 -2522 589 -2520
rect 597 -2522 599 -2520
rect 613 -2522 615 -2520
rect 623 -2522 625 -2520
rect 631 -2522 633 -2520
rect 641 -2522 643 -2520
rect 657 -2522 659 -2520
rect 665 -2522 667 -2520
rect 681 -2522 683 -2520
rect 697 -2522 699 -2520
rect 705 -2522 707 -2520
rect 715 -2522 717 -2520
rect 791 -2522 793 -2520
rect 801 -2522 803 -2520
rect 817 -2522 819 -2520
rect 827 -2522 829 -2520
rect 843 -2522 845 -2520
rect 853 -2522 855 -2520
rect 861 -2522 863 -2520
rect 871 -2522 873 -2520
rect 887 -2522 889 -2520
rect 895 -2522 897 -2520
rect 905 -2522 907 -2520
rect 921 -2522 923 -2520
rect 931 -2522 933 -2520
rect 939 -2522 941 -2520
rect 949 -2522 951 -2520
rect 965 -2522 967 -2520
rect 973 -2522 975 -2520
rect 989 -2522 991 -2520
rect 1005 -2522 1007 -2520
rect 1013 -2522 1015 -2520
rect 1023 -2522 1025 -2520
rect -1229 -2598 -1227 -2530
rect -1219 -2598 -1217 -2530
rect -1203 -2598 -1201 -2530
rect -1193 -2598 -1191 -2530
rect -1185 -2598 -1183 -2530
rect -1175 -2598 -1173 -2530
rect -1159 -2598 -1157 -2530
rect -1151 -2598 -1149 -2530
rect -1141 -2598 -1139 -2530
rect -1057 -2598 -1055 -2530
rect -1047 -2598 -1045 -2530
rect -1031 -2598 -1029 -2530
rect -1021 -2598 -1019 -2530
rect -1005 -2598 -1003 -2530
rect -995 -2598 -993 -2530
rect -987 -2598 -985 -2530
rect -977 -2598 -975 -2530
rect -961 -2598 -959 -2530
rect -953 -2598 -951 -2530
rect -943 -2598 -941 -2530
rect -927 -2598 -925 -2530
rect -917 -2598 -915 -2530
rect -909 -2598 -907 -2530
rect -899 -2598 -897 -2530
rect -883 -2598 -881 -2530
rect -875 -2598 -873 -2530
rect -859 -2598 -857 -2530
rect -843 -2598 -841 -2530
rect -835 -2598 -833 -2530
rect -825 -2598 -823 -2530
rect -749 -2598 -747 -2530
rect -739 -2598 -737 -2530
rect -723 -2598 -721 -2530
rect -713 -2598 -711 -2530
rect -697 -2598 -695 -2530
rect -687 -2598 -685 -2530
rect -679 -2598 -677 -2530
rect -669 -2598 -667 -2530
rect -653 -2598 -651 -2530
rect -645 -2598 -643 -2530
rect -635 -2598 -633 -2530
rect -619 -2598 -617 -2530
rect -609 -2598 -607 -2530
rect -601 -2598 -599 -2530
rect -591 -2598 -589 -2530
rect -575 -2598 -573 -2530
rect -567 -2598 -565 -2530
rect -551 -2598 -549 -2530
rect -535 -2598 -533 -2530
rect -527 -2598 -525 -2530
rect -517 -2598 -515 -2530
rect -441 -2598 -439 -2530
rect -431 -2598 -429 -2530
rect -415 -2598 -413 -2530
rect -405 -2598 -403 -2530
rect -389 -2598 -387 -2530
rect -379 -2598 -377 -2530
rect -371 -2598 -369 -2530
rect -361 -2598 -359 -2530
rect -345 -2598 -343 -2530
rect -337 -2598 -335 -2530
rect -327 -2598 -325 -2530
rect -311 -2598 -309 -2530
rect -301 -2598 -299 -2530
rect -293 -2598 -291 -2530
rect -283 -2598 -281 -2530
rect -267 -2598 -265 -2530
rect -259 -2598 -257 -2530
rect -243 -2598 -241 -2530
rect -227 -2598 -225 -2530
rect -219 -2598 -217 -2530
rect -209 -2598 -207 -2530
rect -133 -2598 -131 -2530
rect -123 -2598 -121 -2530
rect -107 -2598 -105 -2530
rect -97 -2598 -95 -2530
rect -81 -2598 -79 -2530
rect -71 -2598 -69 -2530
rect -63 -2598 -61 -2530
rect -53 -2598 -51 -2530
rect -37 -2598 -35 -2530
rect -29 -2598 -27 -2530
rect -19 -2598 -17 -2530
rect -3 -2598 -1 -2530
rect 7 -2598 9 -2530
rect 15 -2598 17 -2530
rect 25 -2598 27 -2530
rect 41 -2598 43 -2530
rect 49 -2598 51 -2530
rect 65 -2598 67 -2530
rect 81 -2598 83 -2530
rect 89 -2598 91 -2530
rect 99 -2598 101 -2530
rect 175 -2598 177 -2530
rect 185 -2598 187 -2530
rect 201 -2598 203 -2530
rect 211 -2598 213 -2530
rect 227 -2598 229 -2530
rect 237 -2598 239 -2530
rect 245 -2598 247 -2530
rect 255 -2598 257 -2530
rect 271 -2598 273 -2530
rect 279 -2598 281 -2530
rect 289 -2598 291 -2530
rect 305 -2598 307 -2530
rect 315 -2598 317 -2530
rect 323 -2598 325 -2530
rect 333 -2598 335 -2530
rect 349 -2598 351 -2530
rect 357 -2598 359 -2530
rect 373 -2598 375 -2530
rect 389 -2598 391 -2530
rect 397 -2598 399 -2530
rect 407 -2598 409 -2530
rect 483 -2598 485 -2530
rect 493 -2598 495 -2530
rect 509 -2598 511 -2530
rect 519 -2598 521 -2530
rect 535 -2598 537 -2530
rect 545 -2598 547 -2530
rect 553 -2598 555 -2530
rect 563 -2598 565 -2530
rect 579 -2598 581 -2530
rect 587 -2598 589 -2530
rect 597 -2598 599 -2530
rect 613 -2598 615 -2530
rect 623 -2598 625 -2530
rect 631 -2598 633 -2530
rect 641 -2598 643 -2530
rect 657 -2598 659 -2530
rect 665 -2598 667 -2530
rect 681 -2598 683 -2530
rect 697 -2598 699 -2530
rect 705 -2598 707 -2530
rect 715 -2598 717 -2530
rect 791 -2598 793 -2530
rect 801 -2598 803 -2530
rect 817 -2598 819 -2530
rect 827 -2598 829 -2530
rect 843 -2598 845 -2530
rect 853 -2598 855 -2530
rect 861 -2598 863 -2530
rect 871 -2598 873 -2530
rect 887 -2598 889 -2530
rect 895 -2598 897 -2530
rect 905 -2598 907 -2530
rect 921 -2598 923 -2530
rect 931 -2598 933 -2530
rect 939 -2598 941 -2530
rect 949 -2598 951 -2530
rect 965 -2598 967 -2530
rect 973 -2598 975 -2530
rect 989 -2598 991 -2530
rect 1005 -2598 1007 -2530
rect 1013 -2598 1015 -2530
rect 1023 -2598 1025 -2530
rect -1229 -2604 -1227 -2602
rect -1219 -2604 -1217 -2602
rect -1203 -2604 -1201 -2602
rect -1193 -2604 -1191 -2602
rect -1185 -2604 -1183 -2602
rect -1175 -2604 -1173 -2602
rect -1159 -2604 -1157 -2602
rect -1151 -2604 -1149 -2602
rect -1141 -2604 -1139 -2602
rect -1057 -2604 -1055 -2602
rect -1047 -2604 -1045 -2602
rect -1031 -2604 -1029 -2602
rect -1021 -2604 -1019 -2602
rect -1005 -2604 -1003 -2602
rect -995 -2604 -993 -2602
rect -987 -2604 -985 -2602
rect -977 -2604 -975 -2602
rect -961 -2604 -959 -2602
rect -953 -2604 -951 -2602
rect -943 -2604 -941 -2602
rect -927 -2604 -925 -2602
rect -917 -2604 -915 -2602
rect -909 -2604 -907 -2602
rect -899 -2604 -897 -2602
rect -883 -2604 -881 -2602
rect -875 -2604 -873 -2602
rect -859 -2604 -857 -2602
rect -843 -2604 -841 -2602
rect -835 -2604 -833 -2602
rect -825 -2604 -823 -2602
rect -749 -2604 -747 -2602
rect -739 -2604 -737 -2602
rect -723 -2604 -721 -2602
rect -713 -2604 -711 -2602
rect -697 -2604 -695 -2602
rect -687 -2604 -685 -2602
rect -679 -2604 -677 -2602
rect -669 -2604 -667 -2602
rect -653 -2604 -651 -2602
rect -645 -2604 -643 -2602
rect -635 -2604 -633 -2602
rect -619 -2604 -617 -2602
rect -609 -2604 -607 -2602
rect -601 -2604 -599 -2602
rect -591 -2604 -589 -2602
rect -575 -2604 -573 -2602
rect -567 -2604 -565 -2602
rect -551 -2604 -549 -2602
rect -535 -2604 -533 -2602
rect -527 -2604 -525 -2602
rect -517 -2604 -515 -2602
rect -441 -2604 -439 -2602
rect -431 -2604 -429 -2602
rect -415 -2604 -413 -2602
rect -405 -2604 -403 -2602
rect -389 -2604 -387 -2602
rect -379 -2604 -377 -2602
rect -371 -2604 -369 -2602
rect -361 -2604 -359 -2602
rect -345 -2604 -343 -2602
rect -337 -2604 -335 -2602
rect -327 -2604 -325 -2602
rect -311 -2604 -309 -2602
rect -301 -2604 -299 -2602
rect -293 -2604 -291 -2602
rect -283 -2604 -281 -2602
rect -267 -2604 -265 -2602
rect -259 -2604 -257 -2602
rect -243 -2604 -241 -2602
rect -227 -2604 -225 -2602
rect -219 -2604 -217 -2602
rect -209 -2604 -207 -2602
rect -133 -2604 -131 -2602
rect -123 -2604 -121 -2602
rect -107 -2604 -105 -2602
rect -97 -2604 -95 -2602
rect -81 -2604 -79 -2602
rect -71 -2604 -69 -2602
rect -63 -2604 -61 -2602
rect -53 -2604 -51 -2602
rect -37 -2604 -35 -2602
rect -29 -2604 -27 -2602
rect -19 -2604 -17 -2602
rect -3 -2604 -1 -2602
rect 7 -2604 9 -2602
rect 15 -2604 17 -2602
rect 25 -2604 27 -2602
rect 41 -2604 43 -2602
rect 49 -2604 51 -2602
rect 65 -2604 67 -2602
rect 81 -2604 83 -2602
rect 89 -2604 91 -2602
rect 99 -2604 101 -2602
rect 175 -2604 177 -2602
rect 185 -2604 187 -2602
rect 201 -2604 203 -2602
rect 211 -2604 213 -2602
rect 227 -2604 229 -2602
rect 237 -2604 239 -2602
rect 245 -2604 247 -2602
rect 255 -2604 257 -2602
rect 271 -2604 273 -2602
rect 279 -2604 281 -2602
rect 289 -2604 291 -2602
rect 305 -2604 307 -2602
rect 315 -2604 317 -2602
rect 323 -2604 325 -2602
rect 333 -2604 335 -2602
rect 349 -2604 351 -2602
rect 357 -2604 359 -2602
rect 373 -2604 375 -2602
rect 389 -2604 391 -2602
rect 397 -2604 399 -2602
rect 407 -2604 409 -2602
rect 483 -2604 485 -2602
rect 493 -2604 495 -2602
rect 509 -2604 511 -2602
rect 519 -2604 521 -2602
rect 535 -2604 537 -2602
rect 545 -2604 547 -2602
rect 553 -2604 555 -2602
rect 563 -2604 565 -2602
rect 579 -2604 581 -2602
rect 587 -2604 589 -2602
rect 597 -2604 599 -2602
rect 613 -2604 615 -2602
rect 623 -2604 625 -2602
rect 631 -2604 633 -2602
rect 641 -2604 643 -2602
rect 657 -2604 659 -2602
rect 665 -2604 667 -2602
rect 681 -2604 683 -2602
rect 697 -2604 699 -2602
rect 705 -2604 707 -2602
rect 715 -2604 717 -2602
rect 791 -2604 793 -2602
rect 801 -2604 803 -2602
rect 817 -2604 819 -2602
rect 827 -2604 829 -2602
rect 843 -2604 845 -2602
rect 853 -2604 855 -2602
rect 861 -2604 863 -2602
rect 871 -2604 873 -2602
rect 887 -2604 889 -2602
rect 895 -2604 897 -2602
rect 905 -2604 907 -2602
rect 921 -2604 923 -2602
rect 931 -2604 933 -2602
rect 939 -2604 941 -2602
rect 949 -2604 951 -2602
rect 965 -2604 967 -2602
rect 973 -2604 975 -2602
rect 989 -2604 991 -2602
rect 1005 -2604 1007 -2602
rect 1013 -2604 1015 -2602
rect 1023 -2604 1025 -2602
rect -1304 -2654 -1302 -2652
rect -1296 -2654 -1294 -2652
rect -1286 -2654 -1284 -2652
rect -1057 -2654 -1055 -2652
rect -1049 -2654 -1047 -2652
rect -1039 -2654 -1037 -2652
rect -749 -2654 -747 -2652
rect -741 -2654 -739 -2652
rect -731 -2654 -729 -2652
rect -441 -2654 -439 -2652
rect -433 -2654 -431 -2652
rect -423 -2654 -421 -2652
rect -133 -2654 -131 -2652
rect -125 -2654 -123 -2652
rect -115 -2654 -113 -2652
rect 175 -2654 177 -2652
rect 183 -2654 185 -2652
rect 193 -2654 195 -2652
rect 483 -2654 485 -2652
rect 491 -2654 493 -2652
rect 501 -2654 503 -2652
rect 791 -2654 793 -2652
rect 799 -2654 801 -2652
rect 809 -2654 811 -2652
rect -1304 -2730 -1302 -2662
rect -1296 -2686 -1294 -2662
rect -1296 -2730 -1294 -2690
rect -1286 -2730 -1284 -2662
rect -1057 -2730 -1055 -2662
rect -1049 -2686 -1047 -2662
rect -1049 -2730 -1047 -2690
rect -1039 -2730 -1037 -2662
rect -749 -2730 -747 -2662
rect -741 -2686 -739 -2662
rect -741 -2730 -739 -2690
rect -731 -2730 -729 -2662
rect -441 -2730 -439 -2662
rect -433 -2686 -431 -2662
rect -433 -2730 -431 -2690
rect -423 -2730 -421 -2662
rect -133 -2730 -131 -2662
rect -125 -2686 -123 -2662
rect -125 -2730 -123 -2690
rect -115 -2730 -113 -2662
rect 175 -2730 177 -2662
rect 183 -2686 185 -2662
rect 183 -2730 185 -2690
rect 193 -2730 195 -2662
rect 483 -2730 485 -2662
rect 491 -2686 493 -2662
rect 491 -2730 493 -2690
rect 501 -2730 503 -2662
rect 791 -2730 793 -2662
rect 799 -2686 801 -2662
rect 799 -2730 801 -2690
rect 809 -2730 811 -2662
rect -1304 -2736 -1302 -2734
rect -1296 -2736 -1294 -2734
rect -1286 -2736 -1284 -2734
rect -1057 -2736 -1055 -2734
rect -1049 -2736 -1047 -2734
rect -1039 -2736 -1037 -2734
rect -749 -2736 -747 -2734
rect -741 -2736 -739 -2734
rect -731 -2736 -729 -2734
rect -441 -2736 -439 -2734
rect -433 -2736 -431 -2734
rect -423 -2736 -421 -2734
rect -133 -2736 -131 -2734
rect -125 -2736 -123 -2734
rect -115 -2736 -113 -2734
rect 175 -2736 177 -2734
rect 183 -2736 185 -2734
rect 193 -2736 195 -2734
rect 483 -2736 485 -2734
rect 491 -2736 493 -2734
rect 501 -2736 503 -2734
rect 791 -2736 793 -2734
rect 799 -2736 801 -2734
rect 809 -2736 811 -2734
rect -1229 -2813 -1227 -2811
rect -1219 -2813 -1217 -2811
rect -1203 -2813 -1201 -2811
rect -1193 -2813 -1191 -2811
rect -1185 -2813 -1183 -2811
rect -1175 -2813 -1173 -2811
rect -1159 -2813 -1157 -2811
rect -1151 -2813 -1149 -2811
rect -1141 -2813 -1139 -2811
rect -1057 -2813 -1055 -2811
rect -1047 -2813 -1045 -2811
rect -1031 -2813 -1029 -2811
rect -1021 -2813 -1019 -2811
rect -1005 -2813 -1003 -2811
rect -995 -2813 -993 -2811
rect -987 -2813 -985 -2811
rect -977 -2813 -975 -2811
rect -961 -2813 -959 -2811
rect -953 -2813 -951 -2811
rect -943 -2813 -941 -2811
rect -927 -2813 -925 -2811
rect -917 -2813 -915 -2811
rect -909 -2813 -907 -2811
rect -899 -2813 -897 -2811
rect -883 -2813 -881 -2811
rect -875 -2813 -873 -2811
rect -859 -2813 -857 -2811
rect -843 -2813 -841 -2811
rect -835 -2813 -833 -2811
rect -825 -2813 -823 -2811
rect -749 -2813 -747 -2811
rect -739 -2813 -737 -2811
rect -723 -2813 -721 -2811
rect -713 -2813 -711 -2811
rect -697 -2813 -695 -2811
rect -687 -2813 -685 -2811
rect -679 -2813 -677 -2811
rect -669 -2813 -667 -2811
rect -653 -2813 -651 -2811
rect -645 -2813 -643 -2811
rect -635 -2813 -633 -2811
rect -619 -2813 -617 -2811
rect -609 -2813 -607 -2811
rect -601 -2813 -599 -2811
rect -591 -2813 -589 -2811
rect -575 -2813 -573 -2811
rect -567 -2813 -565 -2811
rect -551 -2813 -549 -2811
rect -535 -2813 -533 -2811
rect -527 -2813 -525 -2811
rect -517 -2813 -515 -2811
rect -441 -2813 -439 -2811
rect -431 -2813 -429 -2811
rect -415 -2813 -413 -2811
rect -405 -2813 -403 -2811
rect -389 -2813 -387 -2811
rect -379 -2813 -377 -2811
rect -371 -2813 -369 -2811
rect -361 -2813 -359 -2811
rect -345 -2813 -343 -2811
rect -337 -2813 -335 -2811
rect -327 -2813 -325 -2811
rect -311 -2813 -309 -2811
rect -301 -2813 -299 -2811
rect -293 -2813 -291 -2811
rect -283 -2813 -281 -2811
rect -267 -2813 -265 -2811
rect -259 -2813 -257 -2811
rect -243 -2813 -241 -2811
rect -227 -2813 -225 -2811
rect -219 -2813 -217 -2811
rect -209 -2813 -207 -2811
rect -133 -2813 -131 -2811
rect -123 -2813 -121 -2811
rect -107 -2813 -105 -2811
rect -97 -2813 -95 -2811
rect -81 -2813 -79 -2811
rect -71 -2813 -69 -2811
rect -63 -2813 -61 -2811
rect -53 -2813 -51 -2811
rect -37 -2813 -35 -2811
rect -29 -2813 -27 -2811
rect -19 -2813 -17 -2811
rect -3 -2813 -1 -2811
rect 7 -2813 9 -2811
rect 15 -2813 17 -2811
rect 25 -2813 27 -2811
rect 41 -2813 43 -2811
rect 49 -2813 51 -2811
rect 65 -2813 67 -2811
rect 81 -2813 83 -2811
rect 89 -2813 91 -2811
rect 99 -2813 101 -2811
rect 175 -2813 177 -2811
rect 185 -2813 187 -2811
rect 201 -2813 203 -2811
rect 211 -2813 213 -2811
rect 227 -2813 229 -2811
rect 237 -2813 239 -2811
rect 245 -2813 247 -2811
rect 255 -2813 257 -2811
rect 271 -2813 273 -2811
rect 279 -2813 281 -2811
rect 289 -2813 291 -2811
rect 305 -2813 307 -2811
rect 315 -2813 317 -2811
rect 323 -2813 325 -2811
rect 333 -2813 335 -2811
rect 349 -2813 351 -2811
rect 357 -2813 359 -2811
rect 373 -2813 375 -2811
rect 389 -2813 391 -2811
rect 397 -2813 399 -2811
rect 407 -2813 409 -2811
rect 483 -2813 485 -2811
rect 493 -2813 495 -2811
rect 509 -2813 511 -2811
rect 519 -2813 521 -2811
rect 535 -2813 537 -2811
rect 545 -2813 547 -2811
rect 553 -2813 555 -2811
rect 563 -2813 565 -2811
rect 579 -2813 581 -2811
rect 587 -2813 589 -2811
rect 597 -2813 599 -2811
rect 613 -2813 615 -2811
rect 623 -2813 625 -2811
rect 631 -2813 633 -2811
rect 641 -2813 643 -2811
rect 657 -2813 659 -2811
rect 665 -2813 667 -2811
rect 681 -2813 683 -2811
rect 697 -2813 699 -2811
rect 705 -2813 707 -2811
rect 715 -2813 717 -2811
rect 791 -2813 793 -2811
rect 801 -2813 803 -2811
rect 817 -2813 819 -2811
rect 827 -2813 829 -2811
rect 843 -2813 845 -2811
rect 853 -2813 855 -2811
rect 861 -2813 863 -2811
rect 871 -2813 873 -2811
rect 887 -2813 889 -2811
rect 895 -2813 897 -2811
rect 905 -2813 907 -2811
rect 921 -2813 923 -2811
rect 931 -2813 933 -2811
rect 939 -2813 941 -2811
rect 949 -2813 951 -2811
rect 965 -2813 967 -2811
rect 973 -2813 975 -2811
rect 989 -2813 991 -2811
rect 1005 -2813 1007 -2811
rect 1013 -2813 1015 -2811
rect 1023 -2813 1025 -2811
rect -1229 -2889 -1227 -2821
rect -1219 -2889 -1217 -2821
rect -1203 -2889 -1201 -2821
rect -1193 -2889 -1191 -2821
rect -1185 -2889 -1183 -2821
rect -1175 -2889 -1173 -2821
rect -1159 -2889 -1157 -2821
rect -1151 -2889 -1149 -2821
rect -1141 -2889 -1139 -2821
rect -1057 -2889 -1055 -2821
rect -1047 -2889 -1045 -2821
rect -1031 -2889 -1029 -2821
rect -1021 -2889 -1019 -2821
rect -1005 -2889 -1003 -2821
rect -995 -2889 -993 -2821
rect -987 -2889 -985 -2821
rect -977 -2889 -975 -2821
rect -961 -2889 -959 -2821
rect -953 -2889 -951 -2821
rect -943 -2889 -941 -2821
rect -927 -2889 -925 -2821
rect -917 -2889 -915 -2821
rect -909 -2889 -907 -2821
rect -899 -2889 -897 -2821
rect -883 -2889 -881 -2821
rect -875 -2889 -873 -2821
rect -859 -2889 -857 -2821
rect -843 -2889 -841 -2821
rect -835 -2889 -833 -2821
rect -825 -2889 -823 -2821
rect -749 -2889 -747 -2821
rect -739 -2889 -737 -2821
rect -723 -2889 -721 -2821
rect -713 -2889 -711 -2821
rect -697 -2889 -695 -2821
rect -687 -2889 -685 -2821
rect -679 -2889 -677 -2821
rect -669 -2889 -667 -2821
rect -653 -2889 -651 -2821
rect -645 -2889 -643 -2821
rect -635 -2889 -633 -2821
rect -619 -2889 -617 -2821
rect -609 -2889 -607 -2821
rect -601 -2889 -599 -2821
rect -591 -2889 -589 -2821
rect -575 -2889 -573 -2821
rect -567 -2889 -565 -2821
rect -551 -2889 -549 -2821
rect -535 -2889 -533 -2821
rect -527 -2889 -525 -2821
rect -517 -2889 -515 -2821
rect -441 -2889 -439 -2821
rect -431 -2889 -429 -2821
rect -415 -2889 -413 -2821
rect -405 -2889 -403 -2821
rect -389 -2889 -387 -2821
rect -379 -2889 -377 -2821
rect -371 -2889 -369 -2821
rect -361 -2889 -359 -2821
rect -345 -2889 -343 -2821
rect -337 -2889 -335 -2821
rect -327 -2889 -325 -2821
rect -311 -2889 -309 -2821
rect -301 -2889 -299 -2821
rect -293 -2889 -291 -2821
rect -283 -2889 -281 -2821
rect -267 -2889 -265 -2821
rect -259 -2889 -257 -2821
rect -243 -2889 -241 -2821
rect -227 -2889 -225 -2821
rect -219 -2889 -217 -2821
rect -209 -2889 -207 -2821
rect -133 -2889 -131 -2821
rect -123 -2889 -121 -2821
rect -107 -2889 -105 -2821
rect -97 -2889 -95 -2821
rect -81 -2889 -79 -2821
rect -71 -2889 -69 -2821
rect -63 -2889 -61 -2821
rect -53 -2889 -51 -2821
rect -37 -2889 -35 -2821
rect -29 -2889 -27 -2821
rect -19 -2889 -17 -2821
rect -3 -2889 -1 -2821
rect 7 -2889 9 -2821
rect 15 -2889 17 -2821
rect 25 -2889 27 -2821
rect 41 -2889 43 -2821
rect 49 -2889 51 -2821
rect 65 -2889 67 -2821
rect 81 -2889 83 -2821
rect 89 -2889 91 -2821
rect 99 -2889 101 -2821
rect 175 -2889 177 -2821
rect 185 -2889 187 -2821
rect 201 -2889 203 -2821
rect 211 -2889 213 -2821
rect 227 -2889 229 -2821
rect 237 -2889 239 -2821
rect 245 -2889 247 -2821
rect 255 -2889 257 -2821
rect 271 -2889 273 -2821
rect 279 -2889 281 -2821
rect 289 -2889 291 -2821
rect 305 -2889 307 -2821
rect 315 -2889 317 -2821
rect 323 -2889 325 -2821
rect 333 -2889 335 -2821
rect 349 -2889 351 -2821
rect 357 -2889 359 -2821
rect 373 -2889 375 -2821
rect 389 -2889 391 -2821
rect 397 -2889 399 -2821
rect 407 -2889 409 -2821
rect 483 -2889 485 -2821
rect 493 -2889 495 -2821
rect 509 -2889 511 -2821
rect 519 -2889 521 -2821
rect 535 -2889 537 -2821
rect 545 -2889 547 -2821
rect 553 -2889 555 -2821
rect 563 -2889 565 -2821
rect 579 -2889 581 -2821
rect 587 -2889 589 -2821
rect 597 -2889 599 -2821
rect 613 -2889 615 -2821
rect 623 -2889 625 -2821
rect 631 -2889 633 -2821
rect 641 -2889 643 -2821
rect 657 -2889 659 -2821
rect 665 -2889 667 -2821
rect 681 -2889 683 -2821
rect 697 -2889 699 -2821
rect 705 -2889 707 -2821
rect 715 -2889 717 -2821
rect 791 -2889 793 -2821
rect 801 -2889 803 -2821
rect 817 -2889 819 -2821
rect 827 -2889 829 -2821
rect 843 -2889 845 -2821
rect 853 -2889 855 -2821
rect 861 -2889 863 -2821
rect 871 -2889 873 -2821
rect 887 -2889 889 -2821
rect 895 -2889 897 -2821
rect 905 -2889 907 -2821
rect 921 -2889 923 -2821
rect 931 -2889 933 -2821
rect 939 -2889 941 -2821
rect 949 -2889 951 -2821
rect 965 -2889 967 -2821
rect 973 -2889 975 -2821
rect 989 -2889 991 -2821
rect 1005 -2889 1007 -2821
rect 1013 -2889 1015 -2821
rect 1023 -2889 1025 -2821
rect -1229 -2895 -1227 -2893
rect -1219 -2895 -1217 -2893
rect -1203 -2895 -1201 -2893
rect -1193 -2895 -1191 -2893
rect -1185 -2895 -1183 -2893
rect -1175 -2895 -1173 -2893
rect -1159 -2895 -1157 -2893
rect -1151 -2895 -1149 -2893
rect -1141 -2895 -1139 -2893
rect -1057 -2895 -1055 -2893
rect -1047 -2895 -1045 -2893
rect -1031 -2895 -1029 -2893
rect -1021 -2895 -1019 -2893
rect -1005 -2895 -1003 -2893
rect -995 -2895 -993 -2893
rect -987 -2895 -985 -2893
rect -977 -2895 -975 -2893
rect -961 -2895 -959 -2893
rect -953 -2895 -951 -2893
rect -943 -2895 -941 -2893
rect -927 -2895 -925 -2893
rect -917 -2895 -915 -2893
rect -909 -2895 -907 -2893
rect -899 -2895 -897 -2893
rect -883 -2895 -881 -2893
rect -875 -2895 -873 -2893
rect -859 -2895 -857 -2893
rect -843 -2895 -841 -2893
rect -835 -2895 -833 -2893
rect -825 -2895 -823 -2893
rect -749 -2895 -747 -2893
rect -739 -2895 -737 -2893
rect -723 -2895 -721 -2893
rect -713 -2895 -711 -2893
rect -697 -2895 -695 -2893
rect -687 -2895 -685 -2893
rect -679 -2895 -677 -2893
rect -669 -2895 -667 -2893
rect -653 -2895 -651 -2893
rect -645 -2895 -643 -2893
rect -635 -2895 -633 -2893
rect -619 -2895 -617 -2893
rect -609 -2895 -607 -2893
rect -601 -2895 -599 -2893
rect -591 -2895 -589 -2893
rect -575 -2895 -573 -2893
rect -567 -2895 -565 -2893
rect -551 -2895 -549 -2893
rect -535 -2895 -533 -2893
rect -527 -2895 -525 -2893
rect -517 -2895 -515 -2893
rect -441 -2895 -439 -2893
rect -431 -2895 -429 -2893
rect -415 -2895 -413 -2893
rect -405 -2895 -403 -2893
rect -389 -2895 -387 -2893
rect -379 -2895 -377 -2893
rect -371 -2895 -369 -2893
rect -361 -2895 -359 -2893
rect -345 -2895 -343 -2893
rect -337 -2895 -335 -2893
rect -327 -2895 -325 -2893
rect -311 -2895 -309 -2893
rect -301 -2895 -299 -2893
rect -293 -2895 -291 -2893
rect -283 -2895 -281 -2893
rect -267 -2895 -265 -2893
rect -259 -2895 -257 -2893
rect -243 -2895 -241 -2893
rect -227 -2895 -225 -2893
rect -219 -2895 -217 -2893
rect -209 -2895 -207 -2893
rect -133 -2895 -131 -2893
rect -123 -2895 -121 -2893
rect -107 -2895 -105 -2893
rect -97 -2895 -95 -2893
rect -81 -2895 -79 -2893
rect -71 -2895 -69 -2893
rect -63 -2895 -61 -2893
rect -53 -2895 -51 -2893
rect -37 -2895 -35 -2893
rect -29 -2895 -27 -2893
rect -19 -2895 -17 -2893
rect -3 -2895 -1 -2893
rect 7 -2895 9 -2893
rect 15 -2895 17 -2893
rect 25 -2895 27 -2893
rect 41 -2895 43 -2893
rect 49 -2895 51 -2893
rect 65 -2895 67 -2893
rect 81 -2895 83 -2893
rect 89 -2895 91 -2893
rect 99 -2895 101 -2893
rect 175 -2895 177 -2893
rect 185 -2895 187 -2893
rect 201 -2895 203 -2893
rect 211 -2895 213 -2893
rect 227 -2895 229 -2893
rect 237 -2895 239 -2893
rect 245 -2895 247 -2893
rect 255 -2895 257 -2893
rect 271 -2895 273 -2893
rect 279 -2895 281 -2893
rect 289 -2895 291 -2893
rect 305 -2895 307 -2893
rect 315 -2895 317 -2893
rect 323 -2895 325 -2893
rect 333 -2895 335 -2893
rect 349 -2895 351 -2893
rect 357 -2895 359 -2893
rect 373 -2895 375 -2893
rect 389 -2895 391 -2893
rect 397 -2895 399 -2893
rect 407 -2895 409 -2893
rect 483 -2895 485 -2893
rect 493 -2895 495 -2893
rect 509 -2895 511 -2893
rect 519 -2895 521 -2893
rect 535 -2895 537 -2893
rect 545 -2895 547 -2893
rect 553 -2895 555 -2893
rect 563 -2895 565 -2893
rect 579 -2895 581 -2893
rect 587 -2895 589 -2893
rect 597 -2895 599 -2893
rect 613 -2895 615 -2893
rect 623 -2895 625 -2893
rect 631 -2895 633 -2893
rect 641 -2895 643 -2893
rect 657 -2895 659 -2893
rect 665 -2895 667 -2893
rect 681 -2895 683 -2893
rect 697 -2895 699 -2893
rect 705 -2895 707 -2893
rect 715 -2895 717 -2893
rect 791 -2895 793 -2893
rect 801 -2895 803 -2893
rect 817 -2895 819 -2893
rect 827 -2895 829 -2893
rect 843 -2895 845 -2893
rect 853 -2895 855 -2893
rect 861 -2895 863 -2893
rect 871 -2895 873 -2893
rect 887 -2895 889 -2893
rect 895 -2895 897 -2893
rect 905 -2895 907 -2893
rect 921 -2895 923 -2893
rect 931 -2895 933 -2893
rect 939 -2895 941 -2893
rect 949 -2895 951 -2893
rect 965 -2895 967 -2893
rect 973 -2895 975 -2893
rect 989 -2895 991 -2893
rect 1005 -2895 1007 -2893
rect 1013 -2895 1015 -2893
rect 1023 -2895 1025 -2893
rect -1304 -2945 -1302 -2943
rect -1296 -2945 -1294 -2943
rect -1286 -2945 -1284 -2943
rect -1057 -2945 -1055 -2943
rect -1049 -2945 -1047 -2943
rect -1039 -2945 -1037 -2943
rect -749 -2945 -747 -2943
rect -741 -2945 -739 -2943
rect -731 -2945 -729 -2943
rect -441 -2945 -439 -2943
rect -433 -2945 -431 -2943
rect -423 -2945 -421 -2943
rect -133 -2945 -131 -2943
rect -125 -2945 -123 -2943
rect -115 -2945 -113 -2943
rect 175 -2945 177 -2943
rect 183 -2945 185 -2943
rect 193 -2945 195 -2943
rect 483 -2945 485 -2943
rect 491 -2945 493 -2943
rect 501 -2945 503 -2943
rect 791 -2945 793 -2943
rect 799 -2945 801 -2943
rect 809 -2945 811 -2943
rect -1304 -3021 -1302 -2953
rect -1296 -2977 -1294 -2953
rect -1296 -3021 -1294 -2981
rect -1286 -3021 -1284 -2953
rect -1057 -3021 -1055 -2953
rect -1049 -2977 -1047 -2953
rect -1049 -3021 -1047 -2981
rect -1039 -3021 -1037 -2953
rect -749 -3021 -747 -2953
rect -741 -2977 -739 -2953
rect -741 -3021 -739 -2981
rect -731 -3021 -729 -2953
rect -441 -3021 -439 -2953
rect -433 -2977 -431 -2953
rect -433 -3021 -431 -2981
rect -423 -3021 -421 -2953
rect -133 -3021 -131 -2953
rect -125 -2977 -123 -2953
rect -125 -3021 -123 -2981
rect -115 -3021 -113 -2953
rect 175 -3021 177 -2953
rect 183 -2977 185 -2953
rect 183 -3021 185 -2981
rect 193 -3021 195 -2953
rect 483 -3021 485 -2953
rect 491 -2977 493 -2953
rect 491 -3021 493 -2981
rect 501 -3021 503 -2953
rect 791 -3021 793 -2953
rect 799 -2977 801 -2953
rect 799 -3021 801 -2981
rect 809 -3021 811 -2953
rect -1304 -3027 -1302 -3025
rect -1296 -3027 -1294 -3025
rect -1286 -3027 -1284 -3025
rect -1057 -3027 -1055 -3025
rect -1049 -3027 -1047 -3025
rect -1039 -3027 -1037 -3025
rect -749 -3027 -747 -3025
rect -741 -3027 -739 -3025
rect -731 -3027 -729 -3025
rect -441 -3027 -439 -3025
rect -433 -3027 -431 -3025
rect -423 -3027 -421 -3025
rect -133 -3027 -131 -3025
rect -125 -3027 -123 -3025
rect -115 -3027 -113 -3025
rect 175 -3027 177 -3025
rect 183 -3027 185 -3025
rect 193 -3027 195 -3025
rect 483 -3027 485 -3025
rect 491 -3027 493 -3025
rect 501 -3027 503 -3025
rect 791 -3027 793 -3025
rect 799 -3027 801 -3025
rect 809 -3027 811 -3025
rect -1229 -3104 -1227 -3102
rect -1219 -3104 -1217 -3102
rect -1203 -3104 -1201 -3102
rect -1193 -3104 -1191 -3102
rect -1185 -3104 -1183 -3102
rect -1175 -3104 -1173 -3102
rect -1159 -3104 -1157 -3102
rect -1151 -3104 -1149 -3102
rect -1141 -3104 -1139 -3102
rect -1057 -3104 -1055 -3102
rect -1047 -3104 -1045 -3102
rect -1031 -3104 -1029 -3102
rect -1021 -3104 -1019 -3102
rect -1005 -3104 -1003 -3102
rect -995 -3104 -993 -3102
rect -987 -3104 -985 -3102
rect -977 -3104 -975 -3102
rect -961 -3104 -959 -3102
rect -953 -3104 -951 -3102
rect -943 -3104 -941 -3102
rect -927 -3104 -925 -3102
rect -917 -3104 -915 -3102
rect -909 -3104 -907 -3102
rect -899 -3104 -897 -3102
rect -883 -3104 -881 -3102
rect -875 -3104 -873 -3102
rect -859 -3104 -857 -3102
rect -843 -3104 -841 -3102
rect -835 -3104 -833 -3102
rect -825 -3104 -823 -3102
rect -749 -3104 -747 -3102
rect -739 -3104 -737 -3102
rect -723 -3104 -721 -3102
rect -713 -3104 -711 -3102
rect -697 -3104 -695 -3102
rect -687 -3104 -685 -3102
rect -679 -3104 -677 -3102
rect -669 -3104 -667 -3102
rect -653 -3104 -651 -3102
rect -645 -3104 -643 -3102
rect -635 -3104 -633 -3102
rect -619 -3104 -617 -3102
rect -609 -3104 -607 -3102
rect -601 -3104 -599 -3102
rect -591 -3104 -589 -3102
rect -575 -3104 -573 -3102
rect -567 -3104 -565 -3102
rect -551 -3104 -549 -3102
rect -535 -3104 -533 -3102
rect -527 -3104 -525 -3102
rect -517 -3104 -515 -3102
rect -441 -3104 -439 -3102
rect -431 -3104 -429 -3102
rect -415 -3104 -413 -3102
rect -405 -3104 -403 -3102
rect -389 -3104 -387 -3102
rect -379 -3104 -377 -3102
rect -371 -3104 -369 -3102
rect -361 -3104 -359 -3102
rect -345 -3104 -343 -3102
rect -337 -3104 -335 -3102
rect -327 -3104 -325 -3102
rect -311 -3104 -309 -3102
rect -301 -3104 -299 -3102
rect -293 -3104 -291 -3102
rect -283 -3104 -281 -3102
rect -267 -3104 -265 -3102
rect -259 -3104 -257 -3102
rect -243 -3104 -241 -3102
rect -227 -3104 -225 -3102
rect -219 -3104 -217 -3102
rect -209 -3104 -207 -3102
rect -133 -3104 -131 -3102
rect -123 -3104 -121 -3102
rect -107 -3104 -105 -3102
rect -97 -3104 -95 -3102
rect -81 -3104 -79 -3102
rect -71 -3104 -69 -3102
rect -63 -3104 -61 -3102
rect -53 -3104 -51 -3102
rect -37 -3104 -35 -3102
rect -29 -3104 -27 -3102
rect -19 -3104 -17 -3102
rect -3 -3104 -1 -3102
rect 7 -3104 9 -3102
rect 15 -3104 17 -3102
rect 25 -3104 27 -3102
rect 41 -3104 43 -3102
rect 49 -3104 51 -3102
rect 65 -3104 67 -3102
rect 81 -3104 83 -3102
rect 89 -3104 91 -3102
rect 99 -3104 101 -3102
rect 175 -3104 177 -3102
rect 185 -3104 187 -3102
rect 201 -3104 203 -3102
rect 211 -3104 213 -3102
rect 227 -3104 229 -3102
rect 237 -3104 239 -3102
rect 245 -3104 247 -3102
rect 255 -3104 257 -3102
rect 271 -3104 273 -3102
rect 279 -3104 281 -3102
rect 289 -3104 291 -3102
rect 305 -3104 307 -3102
rect 315 -3104 317 -3102
rect 323 -3104 325 -3102
rect 333 -3104 335 -3102
rect 349 -3104 351 -3102
rect 357 -3104 359 -3102
rect 373 -3104 375 -3102
rect 389 -3104 391 -3102
rect 397 -3104 399 -3102
rect 407 -3104 409 -3102
rect 483 -3104 485 -3102
rect 493 -3104 495 -3102
rect 509 -3104 511 -3102
rect 519 -3104 521 -3102
rect 535 -3104 537 -3102
rect 545 -3104 547 -3102
rect 553 -3104 555 -3102
rect 563 -3104 565 -3102
rect 579 -3104 581 -3102
rect 587 -3104 589 -3102
rect 597 -3104 599 -3102
rect 613 -3104 615 -3102
rect 623 -3104 625 -3102
rect 631 -3104 633 -3102
rect 641 -3104 643 -3102
rect 657 -3104 659 -3102
rect 665 -3104 667 -3102
rect 681 -3104 683 -3102
rect 697 -3104 699 -3102
rect 705 -3104 707 -3102
rect 715 -3104 717 -3102
rect 791 -3104 793 -3102
rect 801 -3104 803 -3102
rect 817 -3104 819 -3102
rect 827 -3104 829 -3102
rect 843 -3104 845 -3102
rect 853 -3104 855 -3102
rect 861 -3104 863 -3102
rect 871 -3104 873 -3102
rect 887 -3104 889 -3102
rect 895 -3104 897 -3102
rect 905 -3104 907 -3102
rect 921 -3104 923 -3102
rect 931 -3104 933 -3102
rect 939 -3104 941 -3102
rect 949 -3104 951 -3102
rect 965 -3104 967 -3102
rect 973 -3104 975 -3102
rect 989 -3104 991 -3102
rect 1005 -3104 1007 -3102
rect 1013 -3104 1015 -3102
rect 1023 -3104 1025 -3102
rect -1229 -3180 -1227 -3112
rect -1219 -3180 -1217 -3112
rect -1203 -3180 -1201 -3112
rect -1193 -3180 -1191 -3112
rect -1185 -3180 -1183 -3112
rect -1175 -3180 -1173 -3112
rect -1159 -3180 -1157 -3112
rect -1151 -3180 -1149 -3112
rect -1141 -3180 -1139 -3112
rect -1057 -3180 -1055 -3112
rect -1047 -3180 -1045 -3112
rect -1031 -3180 -1029 -3112
rect -1021 -3180 -1019 -3112
rect -1005 -3180 -1003 -3112
rect -995 -3180 -993 -3112
rect -987 -3180 -985 -3112
rect -977 -3180 -975 -3112
rect -961 -3180 -959 -3112
rect -953 -3180 -951 -3112
rect -943 -3180 -941 -3112
rect -927 -3180 -925 -3112
rect -917 -3180 -915 -3112
rect -909 -3180 -907 -3112
rect -899 -3180 -897 -3112
rect -883 -3180 -881 -3112
rect -875 -3180 -873 -3112
rect -859 -3180 -857 -3112
rect -843 -3180 -841 -3112
rect -835 -3180 -833 -3112
rect -825 -3180 -823 -3112
rect -749 -3180 -747 -3112
rect -739 -3180 -737 -3112
rect -723 -3180 -721 -3112
rect -713 -3180 -711 -3112
rect -697 -3180 -695 -3112
rect -687 -3180 -685 -3112
rect -679 -3180 -677 -3112
rect -669 -3180 -667 -3112
rect -653 -3180 -651 -3112
rect -645 -3180 -643 -3112
rect -635 -3180 -633 -3112
rect -619 -3180 -617 -3112
rect -609 -3180 -607 -3112
rect -601 -3180 -599 -3112
rect -591 -3180 -589 -3112
rect -575 -3180 -573 -3112
rect -567 -3180 -565 -3112
rect -551 -3180 -549 -3112
rect -535 -3180 -533 -3112
rect -527 -3180 -525 -3112
rect -517 -3180 -515 -3112
rect -441 -3180 -439 -3112
rect -431 -3180 -429 -3112
rect -415 -3180 -413 -3112
rect -405 -3180 -403 -3112
rect -389 -3180 -387 -3112
rect -379 -3180 -377 -3112
rect -371 -3180 -369 -3112
rect -361 -3180 -359 -3112
rect -345 -3180 -343 -3112
rect -337 -3180 -335 -3112
rect -327 -3180 -325 -3112
rect -311 -3180 -309 -3112
rect -301 -3180 -299 -3112
rect -293 -3180 -291 -3112
rect -283 -3180 -281 -3112
rect -267 -3180 -265 -3112
rect -259 -3180 -257 -3112
rect -243 -3180 -241 -3112
rect -227 -3180 -225 -3112
rect -219 -3180 -217 -3112
rect -209 -3180 -207 -3112
rect -133 -3180 -131 -3112
rect -123 -3180 -121 -3112
rect -107 -3180 -105 -3112
rect -97 -3180 -95 -3112
rect -81 -3180 -79 -3112
rect -71 -3180 -69 -3112
rect -63 -3180 -61 -3112
rect -53 -3180 -51 -3112
rect -37 -3180 -35 -3112
rect -29 -3180 -27 -3112
rect -19 -3180 -17 -3112
rect -3 -3180 -1 -3112
rect 7 -3180 9 -3112
rect 15 -3180 17 -3112
rect 25 -3180 27 -3112
rect 41 -3180 43 -3112
rect 49 -3180 51 -3112
rect 65 -3180 67 -3112
rect 81 -3180 83 -3112
rect 89 -3180 91 -3112
rect 99 -3180 101 -3112
rect 175 -3180 177 -3112
rect 185 -3180 187 -3112
rect 201 -3180 203 -3112
rect 211 -3180 213 -3112
rect 227 -3180 229 -3112
rect 237 -3180 239 -3112
rect 245 -3180 247 -3112
rect 255 -3180 257 -3112
rect 271 -3180 273 -3112
rect 279 -3180 281 -3112
rect 289 -3180 291 -3112
rect 305 -3180 307 -3112
rect 315 -3180 317 -3112
rect 323 -3180 325 -3112
rect 333 -3180 335 -3112
rect 349 -3180 351 -3112
rect 357 -3180 359 -3112
rect 373 -3180 375 -3112
rect 389 -3180 391 -3112
rect 397 -3180 399 -3112
rect 407 -3180 409 -3112
rect 483 -3180 485 -3112
rect 493 -3180 495 -3112
rect 509 -3180 511 -3112
rect 519 -3180 521 -3112
rect 535 -3180 537 -3112
rect 545 -3180 547 -3112
rect 553 -3180 555 -3112
rect 563 -3180 565 -3112
rect 579 -3180 581 -3112
rect 587 -3180 589 -3112
rect 597 -3180 599 -3112
rect 613 -3180 615 -3112
rect 623 -3180 625 -3112
rect 631 -3180 633 -3112
rect 641 -3180 643 -3112
rect 657 -3180 659 -3112
rect 665 -3180 667 -3112
rect 681 -3180 683 -3112
rect 697 -3180 699 -3112
rect 705 -3180 707 -3112
rect 715 -3180 717 -3112
rect 791 -3180 793 -3112
rect 801 -3180 803 -3112
rect 817 -3180 819 -3112
rect 827 -3180 829 -3112
rect 843 -3180 845 -3112
rect 853 -3180 855 -3112
rect 861 -3180 863 -3112
rect 871 -3180 873 -3112
rect 887 -3180 889 -3112
rect 895 -3180 897 -3112
rect 905 -3180 907 -3112
rect 921 -3180 923 -3112
rect 931 -3180 933 -3112
rect 939 -3180 941 -3112
rect 949 -3180 951 -3112
rect 965 -3180 967 -3112
rect 973 -3180 975 -3112
rect 989 -3180 991 -3112
rect 1005 -3180 1007 -3112
rect 1013 -3180 1015 -3112
rect 1023 -3180 1025 -3112
rect -1229 -3186 -1227 -3184
rect -1219 -3186 -1217 -3184
rect -1203 -3186 -1201 -3184
rect -1193 -3186 -1191 -3184
rect -1185 -3186 -1183 -3184
rect -1175 -3186 -1173 -3184
rect -1159 -3186 -1157 -3184
rect -1151 -3186 -1149 -3184
rect -1141 -3186 -1139 -3184
rect -1057 -3186 -1055 -3184
rect -1047 -3186 -1045 -3184
rect -1031 -3186 -1029 -3184
rect -1021 -3186 -1019 -3184
rect -1005 -3186 -1003 -3184
rect -995 -3186 -993 -3184
rect -987 -3186 -985 -3184
rect -977 -3186 -975 -3184
rect -961 -3186 -959 -3184
rect -953 -3186 -951 -3184
rect -943 -3186 -941 -3184
rect -927 -3186 -925 -3184
rect -917 -3186 -915 -3184
rect -909 -3186 -907 -3184
rect -899 -3186 -897 -3184
rect -883 -3186 -881 -3184
rect -875 -3186 -873 -3184
rect -859 -3186 -857 -3184
rect -843 -3186 -841 -3184
rect -835 -3186 -833 -3184
rect -825 -3186 -823 -3184
rect -749 -3186 -747 -3184
rect -739 -3186 -737 -3184
rect -723 -3186 -721 -3184
rect -713 -3186 -711 -3184
rect -697 -3186 -695 -3184
rect -687 -3186 -685 -3184
rect -679 -3186 -677 -3184
rect -669 -3186 -667 -3184
rect -653 -3186 -651 -3184
rect -645 -3186 -643 -3184
rect -635 -3186 -633 -3184
rect -619 -3186 -617 -3184
rect -609 -3186 -607 -3184
rect -601 -3186 -599 -3184
rect -591 -3186 -589 -3184
rect -575 -3186 -573 -3184
rect -567 -3186 -565 -3184
rect -551 -3186 -549 -3184
rect -535 -3186 -533 -3184
rect -527 -3186 -525 -3184
rect -517 -3186 -515 -3184
rect -441 -3186 -439 -3184
rect -431 -3186 -429 -3184
rect -415 -3186 -413 -3184
rect -405 -3186 -403 -3184
rect -389 -3186 -387 -3184
rect -379 -3186 -377 -3184
rect -371 -3186 -369 -3184
rect -361 -3186 -359 -3184
rect -345 -3186 -343 -3184
rect -337 -3186 -335 -3184
rect -327 -3186 -325 -3184
rect -311 -3186 -309 -3184
rect -301 -3186 -299 -3184
rect -293 -3186 -291 -3184
rect -283 -3186 -281 -3184
rect -267 -3186 -265 -3184
rect -259 -3186 -257 -3184
rect -243 -3186 -241 -3184
rect -227 -3186 -225 -3184
rect -219 -3186 -217 -3184
rect -209 -3186 -207 -3184
rect -133 -3186 -131 -3184
rect -123 -3186 -121 -3184
rect -107 -3186 -105 -3184
rect -97 -3186 -95 -3184
rect -81 -3186 -79 -3184
rect -71 -3186 -69 -3184
rect -63 -3186 -61 -3184
rect -53 -3186 -51 -3184
rect -37 -3186 -35 -3184
rect -29 -3186 -27 -3184
rect -19 -3186 -17 -3184
rect -3 -3186 -1 -3184
rect 7 -3186 9 -3184
rect 15 -3186 17 -3184
rect 25 -3186 27 -3184
rect 41 -3186 43 -3184
rect 49 -3186 51 -3184
rect 65 -3186 67 -3184
rect 81 -3186 83 -3184
rect 89 -3186 91 -3184
rect 99 -3186 101 -3184
rect 175 -3186 177 -3184
rect 185 -3186 187 -3184
rect 201 -3186 203 -3184
rect 211 -3186 213 -3184
rect 227 -3186 229 -3184
rect 237 -3186 239 -3184
rect 245 -3186 247 -3184
rect 255 -3186 257 -3184
rect 271 -3186 273 -3184
rect 279 -3186 281 -3184
rect 289 -3186 291 -3184
rect 305 -3186 307 -3184
rect 315 -3186 317 -3184
rect 323 -3186 325 -3184
rect 333 -3186 335 -3184
rect 349 -3186 351 -3184
rect 357 -3186 359 -3184
rect 373 -3186 375 -3184
rect 389 -3186 391 -3184
rect 397 -3186 399 -3184
rect 407 -3186 409 -3184
rect 483 -3186 485 -3184
rect 493 -3186 495 -3184
rect 509 -3186 511 -3184
rect 519 -3186 521 -3184
rect 535 -3186 537 -3184
rect 545 -3186 547 -3184
rect 553 -3186 555 -3184
rect 563 -3186 565 -3184
rect 579 -3186 581 -3184
rect 587 -3186 589 -3184
rect 597 -3186 599 -3184
rect 613 -3186 615 -3184
rect 623 -3186 625 -3184
rect 631 -3186 633 -3184
rect 641 -3186 643 -3184
rect 657 -3186 659 -3184
rect 665 -3186 667 -3184
rect 681 -3186 683 -3184
rect 697 -3186 699 -3184
rect 705 -3186 707 -3184
rect 715 -3186 717 -3184
rect 791 -3186 793 -3184
rect 801 -3186 803 -3184
rect 817 -3186 819 -3184
rect 827 -3186 829 -3184
rect 843 -3186 845 -3184
rect 853 -3186 855 -3184
rect 861 -3186 863 -3184
rect 871 -3186 873 -3184
rect 887 -3186 889 -3184
rect 895 -3186 897 -3184
rect 905 -3186 907 -3184
rect 921 -3186 923 -3184
rect 931 -3186 933 -3184
rect 939 -3186 941 -3184
rect 949 -3186 951 -3184
rect 965 -3186 967 -3184
rect 973 -3186 975 -3184
rect 989 -3186 991 -3184
rect 1005 -3186 1007 -3184
rect 1013 -3186 1015 -3184
rect 1023 -3186 1025 -3184
<< ndiffusion >>
rect -1303 -1068 -1302 -1064
rect -1300 -1068 -1294 -1064
rect -1292 -1068 -1290 -1064
rect -1286 -1068 -1284 -1064
rect -1282 -1068 -1281 -1064
rect -1059 -1068 -1058 -1064
rect -1056 -1068 -1050 -1064
rect -1048 -1068 -1046 -1064
rect -1042 -1068 -1040 -1064
rect -1038 -1068 -1037 -1064
rect -750 -1068 -749 -1064
rect -747 -1068 -741 -1064
rect -739 -1068 -737 -1064
rect -733 -1068 -731 -1064
rect -729 -1068 -728 -1064
rect -442 -1068 -441 -1064
rect -439 -1068 -433 -1064
rect -431 -1068 -429 -1064
rect -425 -1068 -423 -1064
rect -421 -1068 -420 -1064
rect -135 -1068 -134 -1064
rect -132 -1068 -126 -1064
rect -124 -1068 -122 -1064
rect -118 -1068 -116 -1064
rect -114 -1068 -113 -1064
rect 174 -1068 175 -1064
rect 177 -1068 183 -1064
rect 185 -1068 187 -1064
rect 191 -1068 193 -1064
rect 195 -1068 196 -1064
rect 482 -1068 483 -1064
rect 485 -1068 491 -1064
rect 493 -1068 495 -1064
rect 499 -1068 501 -1064
rect 503 -1068 504 -1064
rect 790 -1068 791 -1064
rect 793 -1068 799 -1064
rect 801 -1068 803 -1064
rect 807 -1068 809 -1064
rect 811 -1068 812 -1064
rect -1305 -1218 -1304 -1214
rect -1302 -1218 -1296 -1214
rect -1294 -1218 -1292 -1214
rect -1288 -1218 -1286 -1214
rect -1284 -1218 -1283 -1214
rect -1058 -1218 -1057 -1214
rect -1055 -1218 -1049 -1214
rect -1047 -1218 -1045 -1214
rect -1041 -1218 -1039 -1214
rect -1037 -1218 -1036 -1214
rect -750 -1218 -749 -1214
rect -747 -1218 -741 -1214
rect -739 -1218 -737 -1214
rect -733 -1218 -731 -1214
rect -729 -1218 -728 -1214
rect -442 -1218 -441 -1214
rect -439 -1218 -433 -1214
rect -431 -1218 -429 -1214
rect -425 -1218 -423 -1214
rect -421 -1218 -420 -1214
rect -134 -1218 -133 -1214
rect -131 -1218 -125 -1214
rect -123 -1218 -121 -1214
rect -117 -1218 -115 -1214
rect -113 -1218 -112 -1214
rect 174 -1218 175 -1214
rect 177 -1218 183 -1214
rect 185 -1218 187 -1214
rect 191 -1218 193 -1214
rect 195 -1218 196 -1214
rect 482 -1218 483 -1214
rect 485 -1218 491 -1214
rect 493 -1218 495 -1214
rect 499 -1218 501 -1214
rect 503 -1218 504 -1214
rect 790 -1218 791 -1214
rect 793 -1218 799 -1214
rect 801 -1218 803 -1214
rect 807 -1218 809 -1214
rect 811 -1218 812 -1214
rect -1226 -1382 -1225 -1378
rect -1223 -1382 -1221 -1378
rect -1217 -1382 -1215 -1378
rect -1213 -1382 -1212 -1378
rect -1200 -1382 -1199 -1378
rect -1197 -1382 -1195 -1378
rect -1191 -1382 -1189 -1378
rect -1187 -1382 -1181 -1378
rect -1179 -1382 -1177 -1378
rect -1173 -1382 -1171 -1378
rect -1169 -1382 -1168 -1378
rect -1156 -1382 -1155 -1378
rect -1153 -1382 -1147 -1378
rect -1145 -1382 -1143 -1378
rect -1139 -1382 -1137 -1378
rect -1135 -1382 -1134 -1378
rect -1058 -1382 -1057 -1378
rect -1055 -1382 -1053 -1378
rect -1049 -1382 -1047 -1378
rect -1045 -1382 -1044 -1378
rect -1032 -1382 -1031 -1378
rect -1029 -1382 -1027 -1378
rect -1023 -1382 -1021 -1378
rect -1019 -1382 -1018 -1378
rect -1006 -1382 -1005 -1378
rect -1003 -1382 -1002 -1378
rect -998 -1382 -995 -1378
rect -993 -1382 -987 -1378
rect -985 -1382 -984 -1378
rect -980 -1382 -977 -1378
rect -975 -1382 -974 -1378
rect -962 -1382 -961 -1378
rect -959 -1382 -953 -1378
rect -951 -1382 -949 -1378
rect -945 -1382 -943 -1378
rect -941 -1382 -940 -1378
rect -928 -1382 -927 -1378
rect -925 -1382 -923 -1378
rect -919 -1382 -917 -1378
rect -915 -1382 -909 -1378
rect -907 -1382 -905 -1378
rect -901 -1382 -899 -1378
rect -897 -1382 -896 -1378
rect -884 -1382 -883 -1378
rect -881 -1382 -875 -1378
rect -873 -1382 -872 -1378
rect -860 -1382 -859 -1378
rect -857 -1382 -852 -1378
rect -848 -1382 -843 -1378
rect -841 -1382 -840 -1378
rect -836 -1382 -835 -1378
rect -833 -1382 -831 -1378
rect -827 -1382 -825 -1378
rect -823 -1382 -822 -1378
rect -750 -1382 -749 -1378
rect -747 -1382 -745 -1378
rect -741 -1382 -739 -1378
rect -737 -1382 -736 -1378
rect -724 -1382 -723 -1378
rect -721 -1382 -719 -1378
rect -715 -1382 -713 -1378
rect -711 -1382 -710 -1378
rect -698 -1382 -697 -1378
rect -695 -1382 -694 -1378
rect -690 -1382 -687 -1378
rect -685 -1382 -679 -1378
rect -677 -1382 -676 -1378
rect -672 -1382 -669 -1378
rect -667 -1382 -666 -1378
rect -654 -1382 -653 -1378
rect -651 -1382 -645 -1378
rect -643 -1382 -641 -1378
rect -637 -1382 -635 -1378
rect -633 -1382 -632 -1378
rect -620 -1382 -619 -1378
rect -617 -1382 -615 -1378
rect -611 -1382 -609 -1378
rect -607 -1382 -601 -1378
rect -599 -1382 -597 -1378
rect -593 -1382 -591 -1378
rect -589 -1382 -588 -1378
rect -576 -1382 -575 -1378
rect -573 -1382 -567 -1378
rect -565 -1382 -564 -1378
rect -552 -1382 -551 -1378
rect -549 -1382 -544 -1378
rect -540 -1382 -535 -1378
rect -533 -1382 -532 -1378
rect -528 -1382 -527 -1378
rect -525 -1382 -523 -1378
rect -519 -1382 -517 -1378
rect -515 -1382 -514 -1378
rect -442 -1382 -441 -1378
rect -439 -1382 -437 -1378
rect -433 -1382 -431 -1378
rect -429 -1382 -428 -1378
rect -416 -1382 -415 -1378
rect -413 -1382 -411 -1378
rect -407 -1382 -405 -1378
rect -403 -1382 -402 -1378
rect -390 -1382 -389 -1378
rect -387 -1382 -386 -1378
rect -382 -1382 -379 -1378
rect -377 -1382 -371 -1378
rect -369 -1382 -368 -1378
rect -364 -1382 -361 -1378
rect -359 -1382 -358 -1378
rect -346 -1382 -345 -1378
rect -343 -1382 -337 -1378
rect -335 -1382 -333 -1378
rect -329 -1382 -327 -1378
rect -325 -1382 -324 -1378
rect -312 -1382 -311 -1378
rect -309 -1382 -307 -1378
rect -303 -1382 -301 -1378
rect -299 -1382 -293 -1378
rect -291 -1382 -289 -1378
rect -285 -1382 -283 -1378
rect -281 -1382 -280 -1378
rect -268 -1382 -267 -1378
rect -265 -1382 -259 -1378
rect -257 -1382 -256 -1378
rect -244 -1382 -243 -1378
rect -241 -1382 -236 -1378
rect -232 -1382 -227 -1378
rect -225 -1382 -224 -1378
rect -220 -1382 -219 -1378
rect -217 -1382 -215 -1378
rect -211 -1382 -209 -1378
rect -207 -1382 -206 -1378
rect -134 -1382 -133 -1378
rect -131 -1382 -129 -1378
rect -125 -1382 -123 -1378
rect -121 -1382 -120 -1378
rect -108 -1382 -107 -1378
rect -105 -1382 -103 -1378
rect -99 -1382 -97 -1378
rect -95 -1382 -94 -1378
rect -82 -1382 -81 -1378
rect -79 -1382 -78 -1378
rect -74 -1382 -71 -1378
rect -69 -1382 -63 -1378
rect -61 -1382 -60 -1378
rect -56 -1382 -53 -1378
rect -51 -1382 -50 -1378
rect -38 -1382 -37 -1378
rect -35 -1382 -29 -1378
rect -27 -1382 -25 -1378
rect -21 -1382 -19 -1378
rect -17 -1382 -16 -1378
rect -4 -1382 -3 -1378
rect -1 -1382 1 -1378
rect 5 -1382 7 -1378
rect 9 -1382 15 -1378
rect 17 -1382 19 -1378
rect 23 -1382 25 -1378
rect 27 -1382 28 -1378
rect 40 -1382 41 -1378
rect 43 -1382 49 -1378
rect 51 -1382 52 -1378
rect 64 -1382 65 -1378
rect 67 -1382 72 -1378
rect 76 -1382 81 -1378
rect 83 -1382 84 -1378
rect 88 -1382 89 -1378
rect 91 -1382 93 -1378
rect 97 -1382 99 -1378
rect 101 -1382 102 -1378
rect 174 -1382 175 -1378
rect 177 -1382 179 -1378
rect 183 -1382 185 -1378
rect 187 -1382 188 -1378
rect 200 -1382 201 -1378
rect 203 -1382 205 -1378
rect 209 -1382 211 -1378
rect 213 -1382 214 -1378
rect 226 -1382 227 -1378
rect 229 -1382 230 -1378
rect 234 -1382 237 -1378
rect 239 -1382 245 -1378
rect 247 -1382 248 -1378
rect 252 -1382 255 -1378
rect 257 -1382 258 -1378
rect 270 -1382 271 -1378
rect 273 -1382 279 -1378
rect 281 -1382 283 -1378
rect 287 -1382 289 -1378
rect 291 -1382 292 -1378
rect 304 -1382 305 -1378
rect 307 -1382 309 -1378
rect 313 -1382 315 -1378
rect 317 -1382 323 -1378
rect 325 -1382 327 -1378
rect 331 -1382 333 -1378
rect 335 -1382 336 -1378
rect 348 -1382 349 -1378
rect 351 -1382 357 -1378
rect 359 -1382 360 -1378
rect 372 -1382 373 -1378
rect 375 -1382 380 -1378
rect 384 -1382 389 -1378
rect 391 -1382 392 -1378
rect 396 -1382 397 -1378
rect 399 -1382 401 -1378
rect 405 -1382 407 -1378
rect 409 -1382 410 -1378
rect 482 -1382 483 -1378
rect 485 -1382 487 -1378
rect 491 -1382 493 -1378
rect 495 -1382 496 -1378
rect 508 -1382 509 -1378
rect 511 -1382 513 -1378
rect 517 -1382 519 -1378
rect 521 -1382 522 -1378
rect 534 -1382 535 -1378
rect 537 -1382 538 -1378
rect 542 -1382 545 -1378
rect 547 -1382 553 -1378
rect 555 -1382 556 -1378
rect 560 -1382 563 -1378
rect 565 -1382 566 -1378
rect 578 -1382 579 -1378
rect 581 -1382 587 -1378
rect 589 -1382 591 -1378
rect 595 -1382 597 -1378
rect 599 -1382 600 -1378
rect 612 -1382 613 -1378
rect 615 -1382 617 -1378
rect 621 -1382 623 -1378
rect 625 -1382 631 -1378
rect 633 -1382 635 -1378
rect 639 -1382 641 -1378
rect 643 -1382 644 -1378
rect 656 -1382 657 -1378
rect 659 -1382 665 -1378
rect 667 -1382 668 -1378
rect 680 -1382 681 -1378
rect 683 -1382 688 -1378
rect 692 -1382 697 -1378
rect 699 -1382 700 -1378
rect 704 -1382 705 -1378
rect 707 -1382 709 -1378
rect 713 -1382 715 -1378
rect 717 -1382 718 -1378
rect 788 -1382 789 -1378
rect 791 -1382 793 -1378
rect 797 -1382 799 -1378
rect 801 -1382 802 -1378
rect 814 -1382 815 -1378
rect 817 -1382 819 -1378
rect 823 -1382 825 -1378
rect 827 -1382 833 -1378
rect 835 -1382 837 -1378
rect 841 -1382 843 -1378
rect 845 -1382 846 -1378
rect 858 -1382 859 -1378
rect 861 -1382 867 -1378
rect 869 -1382 871 -1378
rect 875 -1382 877 -1378
rect 879 -1382 880 -1378
rect -1305 -1539 -1304 -1535
rect -1302 -1539 -1296 -1535
rect -1294 -1539 -1292 -1535
rect -1288 -1539 -1286 -1535
rect -1284 -1539 -1283 -1535
rect -1058 -1539 -1057 -1535
rect -1055 -1539 -1049 -1535
rect -1047 -1539 -1045 -1535
rect -1041 -1539 -1039 -1535
rect -1037 -1539 -1036 -1535
rect -750 -1539 -749 -1535
rect -747 -1539 -741 -1535
rect -739 -1539 -737 -1535
rect -733 -1539 -731 -1535
rect -729 -1539 -728 -1535
rect -442 -1539 -441 -1535
rect -439 -1539 -433 -1535
rect -431 -1539 -429 -1535
rect -425 -1539 -423 -1535
rect -421 -1539 -420 -1535
rect -134 -1539 -133 -1535
rect -131 -1539 -125 -1535
rect -123 -1539 -121 -1535
rect -117 -1539 -115 -1535
rect -113 -1539 -112 -1535
rect 174 -1539 175 -1535
rect 177 -1539 183 -1535
rect 185 -1539 187 -1535
rect 191 -1539 193 -1535
rect 195 -1539 196 -1535
rect 482 -1539 483 -1535
rect 485 -1539 491 -1535
rect 493 -1539 495 -1535
rect 499 -1539 501 -1535
rect 503 -1539 504 -1535
rect 790 -1539 791 -1535
rect 793 -1539 799 -1535
rect 801 -1539 803 -1535
rect 807 -1539 809 -1535
rect 811 -1539 812 -1535
rect -1230 -1698 -1229 -1694
rect -1227 -1698 -1225 -1694
rect -1221 -1698 -1219 -1694
rect -1217 -1698 -1216 -1694
rect -1204 -1698 -1203 -1694
rect -1201 -1698 -1199 -1694
rect -1195 -1698 -1193 -1694
rect -1191 -1698 -1185 -1694
rect -1183 -1698 -1181 -1694
rect -1177 -1698 -1175 -1694
rect -1173 -1698 -1172 -1694
rect -1160 -1698 -1159 -1694
rect -1157 -1698 -1151 -1694
rect -1149 -1698 -1147 -1694
rect -1143 -1698 -1141 -1694
rect -1139 -1698 -1138 -1694
rect -1058 -1698 -1057 -1694
rect -1055 -1698 -1053 -1694
rect -1049 -1698 -1047 -1694
rect -1045 -1698 -1044 -1694
rect -1032 -1698 -1031 -1694
rect -1029 -1698 -1027 -1694
rect -1023 -1698 -1021 -1694
rect -1019 -1698 -1018 -1694
rect -1006 -1698 -1005 -1694
rect -1003 -1698 -1002 -1694
rect -998 -1698 -995 -1694
rect -993 -1698 -987 -1694
rect -985 -1698 -984 -1694
rect -980 -1698 -977 -1694
rect -975 -1698 -974 -1694
rect -962 -1698 -961 -1694
rect -959 -1698 -953 -1694
rect -951 -1698 -949 -1694
rect -945 -1698 -943 -1694
rect -941 -1698 -940 -1694
rect -928 -1698 -927 -1694
rect -925 -1698 -923 -1694
rect -919 -1698 -917 -1694
rect -915 -1698 -909 -1694
rect -907 -1698 -905 -1694
rect -901 -1698 -899 -1694
rect -897 -1698 -896 -1694
rect -884 -1698 -883 -1694
rect -881 -1698 -875 -1694
rect -873 -1698 -872 -1694
rect -860 -1698 -859 -1694
rect -857 -1698 -852 -1694
rect -848 -1698 -843 -1694
rect -841 -1698 -840 -1694
rect -836 -1698 -835 -1694
rect -833 -1698 -831 -1694
rect -827 -1698 -825 -1694
rect -823 -1698 -822 -1694
rect -750 -1698 -749 -1694
rect -747 -1698 -745 -1694
rect -741 -1698 -739 -1694
rect -737 -1698 -736 -1694
rect -724 -1698 -723 -1694
rect -721 -1698 -719 -1694
rect -715 -1698 -713 -1694
rect -711 -1698 -710 -1694
rect -698 -1698 -697 -1694
rect -695 -1698 -694 -1694
rect -690 -1698 -687 -1694
rect -685 -1698 -679 -1694
rect -677 -1698 -676 -1694
rect -672 -1698 -669 -1694
rect -667 -1698 -666 -1694
rect -654 -1698 -653 -1694
rect -651 -1698 -645 -1694
rect -643 -1698 -641 -1694
rect -637 -1698 -635 -1694
rect -633 -1698 -632 -1694
rect -620 -1698 -619 -1694
rect -617 -1698 -615 -1694
rect -611 -1698 -609 -1694
rect -607 -1698 -601 -1694
rect -599 -1698 -597 -1694
rect -593 -1698 -591 -1694
rect -589 -1698 -588 -1694
rect -576 -1698 -575 -1694
rect -573 -1698 -567 -1694
rect -565 -1698 -564 -1694
rect -552 -1698 -551 -1694
rect -549 -1698 -544 -1694
rect -540 -1698 -535 -1694
rect -533 -1698 -532 -1694
rect -528 -1698 -527 -1694
rect -525 -1698 -523 -1694
rect -519 -1698 -517 -1694
rect -515 -1698 -514 -1694
rect -442 -1698 -441 -1694
rect -439 -1698 -437 -1694
rect -433 -1698 -431 -1694
rect -429 -1698 -428 -1694
rect -416 -1698 -415 -1694
rect -413 -1698 -411 -1694
rect -407 -1698 -405 -1694
rect -403 -1698 -402 -1694
rect -390 -1698 -389 -1694
rect -387 -1698 -386 -1694
rect -382 -1698 -379 -1694
rect -377 -1698 -371 -1694
rect -369 -1698 -368 -1694
rect -364 -1698 -361 -1694
rect -359 -1698 -358 -1694
rect -346 -1698 -345 -1694
rect -343 -1698 -337 -1694
rect -335 -1698 -333 -1694
rect -329 -1698 -327 -1694
rect -325 -1698 -324 -1694
rect -312 -1698 -311 -1694
rect -309 -1698 -307 -1694
rect -303 -1698 -301 -1694
rect -299 -1698 -293 -1694
rect -291 -1698 -289 -1694
rect -285 -1698 -283 -1694
rect -281 -1698 -280 -1694
rect -268 -1698 -267 -1694
rect -265 -1698 -259 -1694
rect -257 -1698 -256 -1694
rect -244 -1698 -243 -1694
rect -241 -1698 -236 -1694
rect -232 -1698 -227 -1694
rect -225 -1698 -224 -1694
rect -220 -1698 -219 -1694
rect -217 -1698 -215 -1694
rect -211 -1698 -209 -1694
rect -207 -1698 -206 -1694
rect -134 -1698 -133 -1694
rect -131 -1698 -129 -1694
rect -125 -1698 -123 -1694
rect -121 -1698 -120 -1694
rect -108 -1698 -107 -1694
rect -105 -1698 -103 -1694
rect -99 -1698 -97 -1694
rect -95 -1698 -94 -1694
rect -82 -1698 -81 -1694
rect -79 -1698 -78 -1694
rect -74 -1698 -71 -1694
rect -69 -1698 -63 -1694
rect -61 -1698 -60 -1694
rect -56 -1698 -53 -1694
rect -51 -1698 -50 -1694
rect -38 -1698 -37 -1694
rect -35 -1698 -29 -1694
rect -27 -1698 -25 -1694
rect -21 -1698 -19 -1694
rect -17 -1698 -16 -1694
rect -4 -1698 -3 -1694
rect -1 -1698 1 -1694
rect 5 -1698 7 -1694
rect 9 -1698 15 -1694
rect 17 -1698 19 -1694
rect 23 -1698 25 -1694
rect 27 -1698 28 -1694
rect 40 -1698 41 -1694
rect 43 -1698 49 -1694
rect 51 -1698 52 -1694
rect 64 -1698 65 -1694
rect 67 -1698 72 -1694
rect 76 -1698 81 -1694
rect 83 -1698 84 -1694
rect 88 -1698 89 -1694
rect 91 -1698 93 -1694
rect 97 -1698 99 -1694
rect 101 -1698 102 -1694
rect 174 -1698 175 -1694
rect 177 -1698 179 -1694
rect 183 -1698 185 -1694
rect 187 -1698 188 -1694
rect 200 -1698 201 -1694
rect 203 -1698 205 -1694
rect 209 -1698 211 -1694
rect 213 -1698 214 -1694
rect 226 -1698 227 -1694
rect 229 -1698 230 -1694
rect 234 -1698 237 -1694
rect 239 -1698 245 -1694
rect 247 -1698 248 -1694
rect 252 -1698 255 -1694
rect 257 -1698 258 -1694
rect 270 -1698 271 -1694
rect 273 -1698 279 -1694
rect 281 -1698 283 -1694
rect 287 -1698 289 -1694
rect 291 -1698 292 -1694
rect 304 -1698 305 -1694
rect 307 -1698 309 -1694
rect 313 -1698 315 -1694
rect 317 -1698 323 -1694
rect 325 -1698 327 -1694
rect 331 -1698 333 -1694
rect 335 -1698 336 -1694
rect 348 -1698 349 -1694
rect 351 -1698 357 -1694
rect 359 -1698 360 -1694
rect 372 -1698 373 -1694
rect 375 -1698 380 -1694
rect 384 -1698 389 -1694
rect 391 -1698 392 -1694
rect 396 -1698 397 -1694
rect 399 -1698 401 -1694
rect 405 -1698 407 -1694
rect 409 -1698 410 -1694
rect 482 -1698 483 -1694
rect 485 -1698 487 -1694
rect 491 -1698 493 -1694
rect 495 -1698 496 -1694
rect 508 -1698 509 -1694
rect 511 -1698 513 -1694
rect 517 -1698 519 -1694
rect 521 -1698 522 -1694
rect 534 -1698 535 -1694
rect 537 -1698 538 -1694
rect 542 -1698 545 -1694
rect 547 -1698 553 -1694
rect 555 -1698 556 -1694
rect 560 -1698 563 -1694
rect 565 -1698 566 -1694
rect 578 -1698 579 -1694
rect 581 -1698 587 -1694
rect 589 -1698 591 -1694
rect 595 -1698 597 -1694
rect 599 -1698 600 -1694
rect 612 -1698 613 -1694
rect 615 -1698 617 -1694
rect 621 -1698 623 -1694
rect 625 -1698 631 -1694
rect 633 -1698 635 -1694
rect 639 -1698 641 -1694
rect 643 -1698 644 -1694
rect 656 -1698 657 -1694
rect 659 -1698 665 -1694
rect 667 -1698 668 -1694
rect 680 -1698 681 -1694
rect 683 -1698 688 -1694
rect 692 -1698 697 -1694
rect 699 -1698 700 -1694
rect 704 -1698 705 -1694
rect 707 -1698 709 -1694
rect 713 -1698 715 -1694
rect 717 -1698 718 -1694
rect 790 -1698 791 -1694
rect 793 -1698 795 -1694
rect 799 -1698 801 -1694
rect 803 -1698 804 -1694
rect 816 -1698 817 -1694
rect 819 -1698 821 -1694
rect 825 -1698 827 -1694
rect 829 -1698 830 -1694
rect 842 -1698 843 -1694
rect 845 -1698 846 -1694
rect 850 -1698 853 -1694
rect 855 -1698 861 -1694
rect 863 -1698 864 -1694
rect 868 -1698 871 -1694
rect 873 -1698 874 -1694
rect 886 -1698 887 -1694
rect 889 -1698 895 -1694
rect 897 -1698 899 -1694
rect 903 -1698 905 -1694
rect 907 -1698 908 -1694
rect 920 -1698 921 -1694
rect 923 -1698 925 -1694
rect 929 -1698 931 -1694
rect 933 -1698 939 -1694
rect 941 -1698 943 -1694
rect 947 -1698 949 -1694
rect 951 -1698 952 -1694
rect 964 -1698 965 -1694
rect 967 -1698 973 -1694
rect 975 -1698 976 -1694
rect 988 -1698 989 -1694
rect 991 -1698 996 -1694
rect 1000 -1698 1005 -1694
rect 1007 -1698 1008 -1694
rect 1012 -1698 1013 -1694
rect 1015 -1698 1017 -1694
rect 1021 -1698 1023 -1694
rect 1025 -1698 1026 -1694
rect -1305 -1830 -1304 -1826
rect -1302 -1830 -1296 -1826
rect -1294 -1830 -1292 -1826
rect -1288 -1830 -1286 -1826
rect -1284 -1830 -1283 -1826
rect -1058 -1830 -1057 -1826
rect -1055 -1830 -1049 -1826
rect -1047 -1830 -1045 -1826
rect -1041 -1830 -1039 -1826
rect -1037 -1830 -1036 -1826
rect -750 -1830 -749 -1826
rect -747 -1830 -741 -1826
rect -739 -1830 -737 -1826
rect -733 -1830 -731 -1826
rect -729 -1830 -728 -1826
rect -442 -1830 -441 -1826
rect -439 -1830 -433 -1826
rect -431 -1830 -429 -1826
rect -425 -1830 -423 -1826
rect -421 -1830 -420 -1826
rect -134 -1830 -133 -1826
rect -131 -1830 -125 -1826
rect -123 -1830 -121 -1826
rect -117 -1830 -115 -1826
rect -113 -1830 -112 -1826
rect 174 -1830 175 -1826
rect 177 -1830 183 -1826
rect 185 -1830 187 -1826
rect 191 -1830 193 -1826
rect 195 -1830 196 -1826
rect 482 -1830 483 -1826
rect 485 -1830 491 -1826
rect 493 -1830 495 -1826
rect 499 -1830 501 -1826
rect 503 -1830 504 -1826
rect 790 -1830 791 -1826
rect 793 -1830 799 -1826
rect 801 -1830 803 -1826
rect 807 -1830 809 -1826
rect 811 -1830 812 -1826
rect -1230 -1989 -1229 -1985
rect -1227 -1989 -1225 -1985
rect -1221 -1989 -1219 -1985
rect -1217 -1989 -1216 -1985
rect -1204 -1989 -1203 -1985
rect -1201 -1989 -1199 -1985
rect -1195 -1989 -1193 -1985
rect -1191 -1989 -1185 -1985
rect -1183 -1989 -1181 -1985
rect -1177 -1989 -1175 -1985
rect -1173 -1989 -1172 -1985
rect -1160 -1989 -1159 -1985
rect -1157 -1989 -1151 -1985
rect -1149 -1989 -1147 -1985
rect -1143 -1989 -1141 -1985
rect -1139 -1989 -1138 -1985
rect -1058 -1989 -1057 -1985
rect -1055 -1989 -1053 -1985
rect -1049 -1989 -1047 -1985
rect -1045 -1989 -1044 -1985
rect -1032 -1989 -1031 -1985
rect -1029 -1989 -1027 -1985
rect -1023 -1989 -1021 -1985
rect -1019 -1989 -1018 -1985
rect -1006 -1989 -1005 -1985
rect -1003 -1989 -1002 -1985
rect -998 -1989 -995 -1985
rect -993 -1989 -987 -1985
rect -985 -1989 -984 -1985
rect -980 -1989 -977 -1985
rect -975 -1989 -974 -1985
rect -962 -1989 -961 -1985
rect -959 -1989 -953 -1985
rect -951 -1989 -949 -1985
rect -945 -1989 -943 -1985
rect -941 -1989 -940 -1985
rect -928 -1989 -927 -1985
rect -925 -1989 -923 -1985
rect -919 -1989 -917 -1985
rect -915 -1989 -909 -1985
rect -907 -1989 -905 -1985
rect -901 -1989 -899 -1985
rect -897 -1989 -896 -1985
rect -884 -1989 -883 -1985
rect -881 -1989 -875 -1985
rect -873 -1989 -872 -1985
rect -860 -1989 -859 -1985
rect -857 -1989 -852 -1985
rect -848 -1989 -843 -1985
rect -841 -1989 -840 -1985
rect -836 -1989 -835 -1985
rect -833 -1989 -831 -1985
rect -827 -1989 -825 -1985
rect -823 -1989 -822 -1985
rect -750 -1989 -749 -1985
rect -747 -1989 -745 -1985
rect -741 -1989 -739 -1985
rect -737 -1989 -736 -1985
rect -724 -1989 -723 -1985
rect -721 -1989 -719 -1985
rect -715 -1989 -713 -1985
rect -711 -1989 -710 -1985
rect -698 -1989 -697 -1985
rect -695 -1989 -694 -1985
rect -690 -1989 -687 -1985
rect -685 -1989 -679 -1985
rect -677 -1989 -676 -1985
rect -672 -1989 -669 -1985
rect -667 -1989 -666 -1985
rect -654 -1989 -653 -1985
rect -651 -1989 -645 -1985
rect -643 -1989 -641 -1985
rect -637 -1989 -635 -1985
rect -633 -1989 -632 -1985
rect -620 -1989 -619 -1985
rect -617 -1989 -615 -1985
rect -611 -1989 -609 -1985
rect -607 -1989 -601 -1985
rect -599 -1989 -597 -1985
rect -593 -1989 -591 -1985
rect -589 -1989 -588 -1985
rect -576 -1989 -575 -1985
rect -573 -1989 -567 -1985
rect -565 -1989 -564 -1985
rect -552 -1989 -551 -1985
rect -549 -1989 -544 -1985
rect -540 -1989 -535 -1985
rect -533 -1989 -532 -1985
rect -528 -1989 -527 -1985
rect -525 -1989 -523 -1985
rect -519 -1989 -517 -1985
rect -515 -1989 -514 -1985
rect -442 -1989 -441 -1985
rect -439 -1989 -437 -1985
rect -433 -1989 -431 -1985
rect -429 -1989 -428 -1985
rect -416 -1989 -415 -1985
rect -413 -1989 -411 -1985
rect -407 -1989 -405 -1985
rect -403 -1989 -402 -1985
rect -390 -1989 -389 -1985
rect -387 -1989 -386 -1985
rect -382 -1989 -379 -1985
rect -377 -1989 -371 -1985
rect -369 -1989 -368 -1985
rect -364 -1989 -361 -1985
rect -359 -1989 -358 -1985
rect -346 -1989 -345 -1985
rect -343 -1989 -337 -1985
rect -335 -1989 -333 -1985
rect -329 -1989 -327 -1985
rect -325 -1989 -324 -1985
rect -312 -1989 -311 -1985
rect -309 -1989 -307 -1985
rect -303 -1989 -301 -1985
rect -299 -1989 -293 -1985
rect -291 -1989 -289 -1985
rect -285 -1989 -283 -1985
rect -281 -1989 -280 -1985
rect -268 -1989 -267 -1985
rect -265 -1989 -259 -1985
rect -257 -1989 -256 -1985
rect -244 -1989 -243 -1985
rect -241 -1989 -236 -1985
rect -232 -1989 -227 -1985
rect -225 -1989 -224 -1985
rect -220 -1989 -219 -1985
rect -217 -1989 -215 -1985
rect -211 -1989 -209 -1985
rect -207 -1989 -206 -1985
rect -134 -1989 -133 -1985
rect -131 -1989 -129 -1985
rect -125 -1989 -123 -1985
rect -121 -1989 -120 -1985
rect -108 -1989 -107 -1985
rect -105 -1989 -103 -1985
rect -99 -1989 -97 -1985
rect -95 -1989 -94 -1985
rect -82 -1989 -81 -1985
rect -79 -1989 -78 -1985
rect -74 -1989 -71 -1985
rect -69 -1989 -63 -1985
rect -61 -1989 -60 -1985
rect -56 -1989 -53 -1985
rect -51 -1989 -50 -1985
rect -38 -1989 -37 -1985
rect -35 -1989 -29 -1985
rect -27 -1989 -25 -1985
rect -21 -1989 -19 -1985
rect -17 -1989 -16 -1985
rect -4 -1989 -3 -1985
rect -1 -1989 1 -1985
rect 5 -1989 7 -1985
rect 9 -1989 15 -1985
rect 17 -1989 19 -1985
rect 23 -1989 25 -1985
rect 27 -1989 28 -1985
rect 40 -1989 41 -1985
rect 43 -1989 49 -1985
rect 51 -1989 52 -1985
rect 64 -1989 65 -1985
rect 67 -1989 72 -1985
rect 76 -1989 81 -1985
rect 83 -1989 84 -1985
rect 88 -1989 89 -1985
rect 91 -1989 93 -1985
rect 97 -1989 99 -1985
rect 101 -1989 102 -1985
rect 174 -1989 175 -1985
rect 177 -1989 179 -1985
rect 183 -1989 185 -1985
rect 187 -1989 188 -1985
rect 200 -1989 201 -1985
rect 203 -1989 205 -1985
rect 209 -1989 211 -1985
rect 213 -1989 214 -1985
rect 226 -1989 227 -1985
rect 229 -1989 230 -1985
rect 234 -1989 237 -1985
rect 239 -1989 245 -1985
rect 247 -1989 248 -1985
rect 252 -1989 255 -1985
rect 257 -1989 258 -1985
rect 270 -1989 271 -1985
rect 273 -1989 279 -1985
rect 281 -1989 283 -1985
rect 287 -1989 289 -1985
rect 291 -1989 292 -1985
rect 304 -1989 305 -1985
rect 307 -1989 309 -1985
rect 313 -1989 315 -1985
rect 317 -1989 323 -1985
rect 325 -1989 327 -1985
rect 331 -1989 333 -1985
rect 335 -1989 336 -1985
rect 348 -1989 349 -1985
rect 351 -1989 357 -1985
rect 359 -1989 360 -1985
rect 372 -1989 373 -1985
rect 375 -1989 380 -1985
rect 384 -1989 389 -1985
rect 391 -1989 392 -1985
rect 396 -1989 397 -1985
rect 399 -1989 401 -1985
rect 405 -1989 407 -1985
rect 409 -1989 410 -1985
rect 482 -1989 483 -1985
rect 485 -1989 487 -1985
rect 491 -1989 493 -1985
rect 495 -1989 496 -1985
rect 508 -1989 509 -1985
rect 511 -1989 513 -1985
rect 517 -1989 519 -1985
rect 521 -1989 522 -1985
rect 534 -1989 535 -1985
rect 537 -1989 538 -1985
rect 542 -1989 545 -1985
rect 547 -1989 553 -1985
rect 555 -1989 556 -1985
rect 560 -1989 563 -1985
rect 565 -1989 566 -1985
rect 578 -1989 579 -1985
rect 581 -1989 587 -1985
rect 589 -1989 591 -1985
rect 595 -1989 597 -1985
rect 599 -1989 600 -1985
rect 612 -1989 613 -1985
rect 615 -1989 617 -1985
rect 621 -1989 623 -1985
rect 625 -1989 631 -1985
rect 633 -1989 635 -1985
rect 639 -1989 641 -1985
rect 643 -1989 644 -1985
rect 656 -1989 657 -1985
rect 659 -1989 665 -1985
rect 667 -1989 668 -1985
rect 680 -1989 681 -1985
rect 683 -1989 688 -1985
rect 692 -1989 697 -1985
rect 699 -1989 700 -1985
rect 704 -1989 705 -1985
rect 707 -1989 709 -1985
rect 713 -1989 715 -1985
rect 717 -1989 718 -1985
rect 790 -1989 791 -1985
rect 793 -1989 795 -1985
rect 799 -1989 801 -1985
rect 803 -1989 804 -1985
rect 816 -1989 817 -1985
rect 819 -1989 821 -1985
rect 825 -1989 827 -1985
rect 829 -1989 830 -1985
rect 842 -1989 843 -1985
rect 845 -1989 846 -1985
rect 850 -1989 853 -1985
rect 855 -1989 861 -1985
rect 863 -1989 864 -1985
rect 868 -1989 871 -1985
rect 873 -1989 874 -1985
rect 886 -1989 887 -1985
rect 889 -1989 895 -1985
rect 897 -1989 899 -1985
rect 903 -1989 905 -1985
rect 907 -1989 908 -1985
rect 920 -1989 921 -1985
rect 923 -1989 925 -1985
rect 929 -1989 931 -1985
rect 933 -1989 939 -1985
rect 941 -1989 943 -1985
rect 947 -1989 949 -1985
rect 951 -1989 952 -1985
rect 964 -1989 965 -1985
rect 967 -1989 973 -1985
rect 975 -1989 976 -1985
rect 988 -1989 989 -1985
rect 991 -1989 996 -1985
rect 1000 -1989 1005 -1985
rect 1007 -1989 1008 -1985
rect 1012 -1989 1013 -1985
rect 1015 -1989 1017 -1985
rect 1021 -1989 1023 -1985
rect 1025 -1989 1026 -1985
rect -1305 -2152 -1304 -2148
rect -1302 -2152 -1296 -2148
rect -1294 -2152 -1292 -2148
rect -1288 -2152 -1286 -2148
rect -1284 -2152 -1283 -2148
rect -1058 -2152 -1057 -2148
rect -1055 -2152 -1049 -2148
rect -1047 -2152 -1045 -2148
rect -1041 -2152 -1039 -2148
rect -1037 -2152 -1036 -2148
rect -750 -2152 -749 -2148
rect -747 -2152 -741 -2148
rect -739 -2152 -737 -2148
rect -733 -2152 -731 -2148
rect -729 -2152 -728 -2148
rect -442 -2152 -441 -2148
rect -439 -2152 -433 -2148
rect -431 -2152 -429 -2148
rect -425 -2152 -423 -2148
rect -421 -2152 -420 -2148
rect -134 -2152 -133 -2148
rect -131 -2152 -125 -2148
rect -123 -2152 -121 -2148
rect -117 -2152 -115 -2148
rect -113 -2152 -112 -2148
rect 174 -2152 175 -2148
rect 177 -2152 183 -2148
rect 185 -2152 187 -2148
rect 191 -2152 193 -2148
rect 195 -2152 196 -2148
rect 482 -2152 483 -2148
rect 485 -2152 491 -2148
rect 493 -2152 495 -2148
rect 499 -2152 501 -2148
rect 503 -2152 504 -2148
rect 790 -2152 791 -2148
rect 793 -2152 799 -2148
rect 801 -2152 803 -2148
rect 807 -2152 809 -2148
rect 811 -2152 812 -2148
rect -1230 -2311 -1229 -2307
rect -1227 -2311 -1225 -2307
rect -1221 -2311 -1219 -2307
rect -1217 -2311 -1216 -2307
rect -1204 -2311 -1203 -2307
rect -1201 -2311 -1199 -2307
rect -1195 -2311 -1193 -2307
rect -1191 -2311 -1185 -2307
rect -1183 -2311 -1181 -2307
rect -1177 -2311 -1175 -2307
rect -1173 -2311 -1172 -2307
rect -1160 -2311 -1159 -2307
rect -1157 -2311 -1151 -2307
rect -1149 -2311 -1147 -2307
rect -1143 -2311 -1141 -2307
rect -1139 -2311 -1138 -2307
rect -1058 -2311 -1057 -2307
rect -1055 -2311 -1053 -2307
rect -1049 -2311 -1047 -2307
rect -1045 -2311 -1044 -2307
rect -1032 -2311 -1031 -2307
rect -1029 -2311 -1027 -2307
rect -1023 -2311 -1021 -2307
rect -1019 -2311 -1018 -2307
rect -1006 -2311 -1005 -2307
rect -1003 -2311 -1002 -2307
rect -998 -2311 -995 -2307
rect -993 -2311 -987 -2307
rect -985 -2311 -984 -2307
rect -980 -2311 -977 -2307
rect -975 -2311 -974 -2307
rect -962 -2311 -961 -2307
rect -959 -2311 -953 -2307
rect -951 -2311 -949 -2307
rect -945 -2311 -943 -2307
rect -941 -2311 -940 -2307
rect -928 -2311 -927 -2307
rect -925 -2311 -923 -2307
rect -919 -2311 -917 -2307
rect -915 -2311 -909 -2307
rect -907 -2311 -905 -2307
rect -901 -2311 -899 -2307
rect -897 -2311 -896 -2307
rect -884 -2311 -883 -2307
rect -881 -2311 -875 -2307
rect -873 -2311 -872 -2307
rect -860 -2311 -859 -2307
rect -857 -2311 -852 -2307
rect -848 -2311 -843 -2307
rect -841 -2311 -840 -2307
rect -836 -2311 -835 -2307
rect -833 -2311 -831 -2307
rect -827 -2311 -825 -2307
rect -823 -2311 -822 -2307
rect -750 -2311 -749 -2307
rect -747 -2311 -745 -2307
rect -741 -2311 -739 -2307
rect -737 -2311 -736 -2307
rect -724 -2311 -723 -2307
rect -721 -2311 -719 -2307
rect -715 -2311 -713 -2307
rect -711 -2311 -710 -2307
rect -698 -2311 -697 -2307
rect -695 -2311 -694 -2307
rect -690 -2311 -687 -2307
rect -685 -2311 -679 -2307
rect -677 -2311 -676 -2307
rect -672 -2311 -669 -2307
rect -667 -2311 -666 -2307
rect -654 -2311 -653 -2307
rect -651 -2311 -645 -2307
rect -643 -2311 -641 -2307
rect -637 -2311 -635 -2307
rect -633 -2311 -632 -2307
rect -620 -2311 -619 -2307
rect -617 -2311 -615 -2307
rect -611 -2311 -609 -2307
rect -607 -2311 -601 -2307
rect -599 -2311 -597 -2307
rect -593 -2311 -591 -2307
rect -589 -2311 -588 -2307
rect -576 -2311 -575 -2307
rect -573 -2311 -567 -2307
rect -565 -2311 -564 -2307
rect -552 -2311 -551 -2307
rect -549 -2311 -544 -2307
rect -540 -2311 -535 -2307
rect -533 -2311 -532 -2307
rect -528 -2311 -527 -2307
rect -525 -2311 -523 -2307
rect -519 -2311 -517 -2307
rect -515 -2311 -514 -2307
rect -442 -2311 -441 -2307
rect -439 -2311 -437 -2307
rect -433 -2311 -431 -2307
rect -429 -2311 -428 -2307
rect -416 -2311 -415 -2307
rect -413 -2311 -411 -2307
rect -407 -2311 -405 -2307
rect -403 -2311 -402 -2307
rect -390 -2311 -389 -2307
rect -387 -2311 -386 -2307
rect -382 -2311 -379 -2307
rect -377 -2311 -371 -2307
rect -369 -2311 -368 -2307
rect -364 -2311 -361 -2307
rect -359 -2311 -358 -2307
rect -346 -2311 -345 -2307
rect -343 -2311 -337 -2307
rect -335 -2311 -333 -2307
rect -329 -2311 -327 -2307
rect -325 -2311 -324 -2307
rect -312 -2311 -311 -2307
rect -309 -2311 -307 -2307
rect -303 -2311 -301 -2307
rect -299 -2311 -293 -2307
rect -291 -2311 -289 -2307
rect -285 -2311 -283 -2307
rect -281 -2311 -280 -2307
rect -268 -2311 -267 -2307
rect -265 -2311 -259 -2307
rect -257 -2311 -256 -2307
rect -244 -2311 -243 -2307
rect -241 -2311 -236 -2307
rect -232 -2311 -227 -2307
rect -225 -2311 -224 -2307
rect -220 -2311 -219 -2307
rect -217 -2311 -215 -2307
rect -211 -2311 -209 -2307
rect -207 -2311 -206 -2307
rect -134 -2311 -133 -2307
rect -131 -2311 -129 -2307
rect -125 -2311 -123 -2307
rect -121 -2311 -120 -2307
rect -108 -2311 -107 -2307
rect -105 -2311 -103 -2307
rect -99 -2311 -97 -2307
rect -95 -2311 -94 -2307
rect -82 -2311 -81 -2307
rect -79 -2311 -78 -2307
rect -74 -2311 -71 -2307
rect -69 -2311 -63 -2307
rect -61 -2311 -60 -2307
rect -56 -2311 -53 -2307
rect -51 -2311 -50 -2307
rect -38 -2311 -37 -2307
rect -35 -2311 -29 -2307
rect -27 -2311 -25 -2307
rect -21 -2311 -19 -2307
rect -17 -2311 -16 -2307
rect -4 -2311 -3 -2307
rect -1 -2311 1 -2307
rect 5 -2311 7 -2307
rect 9 -2311 15 -2307
rect 17 -2311 19 -2307
rect 23 -2311 25 -2307
rect 27 -2311 28 -2307
rect 40 -2311 41 -2307
rect 43 -2311 49 -2307
rect 51 -2311 52 -2307
rect 64 -2311 65 -2307
rect 67 -2311 72 -2307
rect 76 -2311 81 -2307
rect 83 -2311 84 -2307
rect 88 -2311 89 -2307
rect 91 -2311 93 -2307
rect 97 -2311 99 -2307
rect 101 -2311 102 -2307
rect 174 -2311 175 -2307
rect 177 -2311 179 -2307
rect 183 -2311 185 -2307
rect 187 -2311 188 -2307
rect 200 -2311 201 -2307
rect 203 -2311 205 -2307
rect 209 -2311 211 -2307
rect 213 -2311 214 -2307
rect 226 -2311 227 -2307
rect 229 -2311 230 -2307
rect 234 -2311 237 -2307
rect 239 -2311 245 -2307
rect 247 -2311 248 -2307
rect 252 -2311 255 -2307
rect 257 -2311 258 -2307
rect 270 -2311 271 -2307
rect 273 -2311 279 -2307
rect 281 -2311 283 -2307
rect 287 -2311 289 -2307
rect 291 -2311 292 -2307
rect 304 -2311 305 -2307
rect 307 -2311 309 -2307
rect 313 -2311 315 -2307
rect 317 -2311 323 -2307
rect 325 -2311 327 -2307
rect 331 -2311 333 -2307
rect 335 -2311 336 -2307
rect 348 -2311 349 -2307
rect 351 -2311 357 -2307
rect 359 -2311 360 -2307
rect 372 -2311 373 -2307
rect 375 -2311 380 -2307
rect 384 -2311 389 -2307
rect 391 -2311 392 -2307
rect 396 -2311 397 -2307
rect 399 -2311 401 -2307
rect 405 -2311 407 -2307
rect 409 -2311 410 -2307
rect 482 -2311 483 -2307
rect 485 -2311 487 -2307
rect 491 -2311 493 -2307
rect 495 -2311 496 -2307
rect 508 -2311 509 -2307
rect 511 -2311 513 -2307
rect 517 -2311 519 -2307
rect 521 -2311 522 -2307
rect 534 -2311 535 -2307
rect 537 -2311 538 -2307
rect 542 -2311 545 -2307
rect 547 -2311 553 -2307
rect 555 -2311 556 -2307
rect 560 -2311 563 -2307
rect 565 -2311 566 -2307
rect 578 -2311 579 -2307
rect 581 -2311 587 -2307
rect 589 -2311 591 -2307
rect 595 -2311 597 -2307
rect 599 -2311 600 -2307
rect 612 -2311 613 -2307
rect 615 -2311 617 -2307
rect 621 -2311 623 -2307
rect 625 -2311 631 -2307
rect 633 -2311 635 -2307
rect 639 -2311 641 -2307
rect 643 -2311 644 -2307
rect 656 -2311 657 -2307
rect 659 -2311 665 -2307
rect 667 -2311 668 -2307
rect 680 -2311 681 -2307
rect 683 -2311 688 -2307
rect 692 -2311 697 -2307
rect 699 -2311 700 -2307
rect 704 -2311 705 -2307
rect 707 -2311 709 -2307
rect 713 -2311 715 -2307
rect 717 -2311 718 -2307
rect 790 -2311 791 -2307
rect 793 -2311 795 -2307
rect 799 -2311 801 -2307
rect 803 -2311 804 -2307
rect 816 -2311 817 -2307
rect 819 -2311 821 -2307
rect 825 -2311 827 -2307
rect 829 -2311 830 -2307
rect 842 -2311 843 -2307
rect 845 -2311 846 -2307
rect 850 -2311 853 -2307
rect 855 -2311 861 -2307
rect 863 -2311 864 -2307
rect 868 -2311 871 -2307
rect 873 -2311 874 -2307
rect 886 -2311 887 -2307
rect 889 -2311 895 -2307
rect 897 -2311 899 -2307
rect 903 -2311 905 -2307
rect 907 -2311 908 -2307
rect 920 -2311 921 -2307
rect 923 -2311 925 -2307
rect 929 -2311 931 -2307
rect 933 -2311 939 -2307
rect 941 -2311 943 -2307
rect 947 -2311 949 -2307
rect 951 -2311 952 -2307
rect 964 -2311 965 -2307
rect 967 -2311 973 -2307
rect 975 -2311 976 -2307
rect 988 -2311 989 -2307
rect 991 -2311 996 -2307
rect 1000 -2311 1005 -2307
rect 1007 -2311 1008 -2307
rect 1012 -2311 1013 -2307
rect 1015 -2311 1017 -2307
rect 1021 -2311 1023 -2307
rect 1025 -2311 1026 -2307
rect -1305 -2443 -1304 -2439
rect -1302 -2443 -1296 -2439
rect -1294 -2443 -1292 -2439
rect -1288 -2443 -1286 -2439
rect -1284 -2443 -1283 -2439
rect -1058 -2443 -1057 -2439
rect -1055 -2443 -1049 -2439
rect -1047 -2443 -1045 -2439
rect -1041 -2443 -1039 -2439
rect -1037 -2443 -1036 -2439
rect -750 -2443 -749 -2439
rect -747 -2443 -741 -2439
rect -739 -2443 -737 -2439
rect -733 -2443 -731 -2439
rect -729 -2443 -728 -2439
rect -442 -2443 -441 -2439
rect -439 -2443 -433 -2439
rect -431 -2443 -429 -2439
rect -425 -2443 -423 -2439
rect -421 -2443 -420 -2439
rect -134 -2443 -133 -2439
rect -131 -2443 -125 -2439
rect -123 -2443 -121 -2439
rect -117 -2443 -115 -2439
rect -113 -2443 -112 -2439
rect 174 -2443 175 -2439
rect 177 -2443 183 -2439
rect 185 -2443 187 -2439
rect 191 -2443 193 -2439
rect 195 -2443 196 -2439
rect 482 -2443 483 -2439
rect 485 -2443 491 -2439
rect 493 -2443 495 -2439
rect 499 -2443 501 -2439
rect 503 -2443 504 -2439
rect 790 -2443 791 -2439
rect 793 -2443 799 -2439
rect 801 -2443 803 -2439
rect 807 -2443 809 -2439
rect 811 -2443 812 -2439
rect -1230 -2602 -1229 -2598
rect -1227 -2602 -1225 -2598
rect -1221 -2602 -1219 -2598
rect -1217 -2602 -1216 -2598
rect -1204 -2602 -1203 -2598
rect -1201 -2602 -1199 -2598
rect -1195 -2602 -1193 -2598
rect -1191 -2602 -1185 -2598
rect -1183 -2602 -1181 -2598
rect -1177 -2602 -1175 -2598
rect -1173 -2602 -1172 -2598
rect -1160 -2602 -1159 -2598
rect -1157 -2602 -1151 -2598
rect -1149 -2602 -1147 -2598
rect -1143 -2602 -1141 -2598
rect -1139 -2602 -1138 -2598
rect -1058 -2602 -1057 -2598
rect -1055 -2602 -1053 -2598
rect -1049 -2602 -1047 -2598
rect -1045 -2602 -1044 -2598
rect -1032 -2602 -1031 -2598
rect -1029 -2602 -1027 -2598
rect -1023 -2602 -1021 -2598
rect -1019 -2602 -1018 -2598
rect -1006 -2602 -1005 -2598
rect -1003 -2602 -1002 -2598
rect -998 -2602 -995 -2598
rect -993 -2602 -987 -2598
rect -985 -2602 -984 -2598
rect -980 -2602 -977 -2598
rect -975 -2602 -974 -2598
rect -962 -2602 -961 -2598
rect -959 -2602 -953 -2598
rect -951 -2602 -949 -2598
rect -945 -2602 -943 -2598
rect -941 -2602 -940 -2598
rect -928 -2602 -927 -2598
rect -925 -2602 -923 -2598
rect -919 -2602 -917 -2598
rect -915 -2602 -909 -2598
rect -907 -2602 -905 -2598
rect -901 -2602 -899 -2598
rect -897 -2602 -896 -2598
rect -884 -2602 -883 -2598
rect -881 -2602 -875 -2598
rect -873 -2602 -872 -2598
rect -860 -2602 -859 -2598
rect -857 -2602 -852 -2598
rect -848 -2602 -843 -2598
rect -841 -2602 -840 -2598
rect -836 -2602 -835 -2598
rect -833 -2602 -831 -2598
rect -827 -2602 -825 -2598
rect -823 -2602 -822 -2598
rect -750 -2602 -749 -2598
rect -747 -2602 -745 -2598
rect -741 -2602 -739 -2598
rect -737 -2602 -736 -2598
rect -724 -2602 -723 -2598
rect -721 -2602 -719 -2598
rect -715 -2602 -713 -2598
rect -711 -2602 -710 -2598
rect -698 -2602 -697 -2598
rect -695 -2602 -694 -2598
rect -690 -2602 -687 -2598
rect -685 -2602 -679 -2598
rect -677 -2602 -676 -2598
rect -672 -2602 -669 -2598
rect -667 -2602 -666 -2598
rect -654 -2602 -653 -2598
rect -651 -2602 -645 -2598
rect -643 -2602 -641 -2598
rect -637 -2602 -635 -2598
rect -633 -2602 -632 -2598
rect -620 -2602 -619 -2598
rect -617 -2602 -615 -2598
rect -611 -2602 -609 -2598
rect -607 -2602 -601 -2598
rect -599 -2602 -597 -2598
rect -593 -2602 -591 -2598
rect -589 -2602 -588 -2598
rect -576 -2602 -575 -2598
rect -573 -2602 -567 -2598
rect -565 -2602 -564 -2598
rect -552 -2602 -551 -2598
rect -549 -2602 -544 -2598
rect -540 -2602 -535 -2598
rect -533 -2602 -532 -2598
rect -528 -2602 -527 -2598
rect -525 -2602 -523 -2598
rect -519 -2602 -517 -2598
rect -515 -2602 -514 -2598
rect -442 -2602 -441 -2598
rect -439 -2602 -437 -2598
rect -433 -2602 -431 -2598
rect -429 -2602 -428 -2598
rect -416 -2602 -415 -2598
rect -413 -2602 -411 -2598
rect -407 -2602 -405 -2598
rect -403 -2602 -402 -2598
rect -390 -2602 -389 -2598
rect -387 -2602 -386 -2598
rect -382 -2602 -379 -2598
rect -377 -2602 -371 -2598
rect -369 -2602 -368 -2598
rect -364 -2602 -361 -2598
rect -359 -2602 -358 -2598
rect -346 -2602 -345 -2598
rect -343 -2602 -337 -2598
rect -335 -2602 -333 -2598
rect -329 -2602 -327 -2598
rect -325 -2602 -324 -2598
rect -312 -2602 -311 -2598
rect -309 -2602 -307 -2598
rect -303 -2602 -301 -2598
rect -299 -2602 -293 -2598
rect -291 -2602 -289 -2598
rect -285 -2602 -283 -2598
rect -281 -2602 -280 -2598
rect -268 -2602 -267 -2598
rect -265 -2602 -259 -2598
rect -257 -2602 -256 -2598
rect -244 -2602 -243 -2598
rect -241 -2602 -236 -2598
rect -232 -2602 -227 -2598
rect -225 -2602 -224 -2598
rect -220 -2602 -219 -2598
rect -217 -2602 -215 -2598
rect -211 -2602 -209 -2598
rect -207 -2602 -206 -2598
rect -134 -2602 -133 -2598
rect -131 -2602 -129 -2598
rect -125 -2602 -123 -2598
rect -121 -2602 -120 -2598
rect -108 -2602 -107 -2598
rect -105 -2602 -103 -2598
rect -99 -2602 -97 -2598
rect -95 -2602 -94 -2598
rect -82 -2602 -81 -2598
rect -79 -2602 -78 -2598
rect -74 -2602 -71 -2598
rect -69 -2602 -63 -2598
rect -61 -2602 -60 -2598
rect -56 -2602 -53 -2598
rect -51 -2602 -50 -2598
rect -38 -2602 -37 -2598
rect -35 -2602 -29 -2598
rect -27 -2602 -25 -2598
rect -21 -2602 -19 -2598
rect -17 -2602 -16 -2598
rect -4 -2602 -3 -2598
rect -1 -2602 1 -2598
rect 5 -2602 7 -2598
rect 9 -2602 15 -2598
rect 17 -2602 19 -2598
rect 23 -2602 25 -2598
rect 27 -2602 28 -2598
rect 40 -2602 41 -2598
rect 43 -2602 49 -2598
rect 51 -2602 52 -2598
rect 64 -2602 65 -2598
rect 67 -2602 72 -2598
rect 76 -2602 81 -2598
rect 83 -2602 84 -2598
rect 88 -2602 89 -2598
rect 91 -2602 93 -2598
rect 97 -2602 99 -2598
rect 101 -2602 102 -2598
rect 174 -2602 175 -2598
rect 177 -2602 179 -2598
rect 183 -2602 185 -2598
rect 187 -2602 188 -2598
rect 200 -2602 201 -2598
rect 203 -2602 205 -2598
rect 209 -2602 211 -2598
rect 213 -2602 214 -2598
rect 226 -2602 227 -2598
rect 229 -2602 230 -2598
rect 234 -2602 237 -2598
rect 239 -2602 245 -2598
rect 247 -2602 248 -2598
rect 252 -2602 255 -2598
rect 257 -2602 258 -2598
rect 270 -2602 271 -2598
rect 273 -2602 279 -2598
rect 281 -2602 283 -2598
rect 287 -2602 289 -2598
rect 291 -2602 292 -2598
rect 304 -2602 305 -2598
rect 307 -2602 309 -2598
rect 313 -2602 315 -2598
rect 317 -2602 323 -2598
rect 325 -2602 327 -2598
rect 331 -2602 333 -2598
rect 335 -2602 336 -2598
rect 348 -2602 349 -2598
rect 351 -2602 357 -2598
rect 359 -2602 360 -2598
rect 372 -2602 373 -2598
rect 375 -2602 380 -2598
rect 384 -2602 389 -2598
rect 391 -2602 392 -2598
rect 396 -2602 397 -2598
rect 399 -2602 401 -2598
rect 405 -2602 407 -2598
rect 409 -2602 410 -2598
rect 482 -2602 483 -2598
rect 485 -2602 487 -2598
rect 491 -2602 493 -2598
rect 495 -2602 496 -2598
rect 508 -2602 509 -2598
rect 511 -2602 513 -2598
rect 517 -2602 519 -2598
rect 521 -2602 522 -2598
rect 534 -2602 535 -2598
rect 537 -2602 538 -2598
rect 542 -2602 545 -2598
rect 547 -2602 553 -2598
rect 555 -2602 556 -2598
rect 560 -2602 563 -2598
rect 565 -2602 566 -2598
rect 578 -2602 579 -2598
rect 581 -2602 587 -2598
rect 589 -2602 591 -2598
rect 595 -2602 597 -2598
rect 599 -2602 600 -2598
rect 612 -2602 613 -2598
rect 615 -2602 617 -2598
rect 621 -2602 623 -2598
rect 625 -2602 631 -2598
rect 633 -2602 635 -2598
rect 639 -2602 641 -2598
rect 643 -2602 644 -2598
rect 656 -2602 657 -2598
rect 659 -2602 665 -2598
rect 667 -2602 668 -2598
rect 680 -2602 681 -2598
rect 683 -2602 688 -2598
rect 692 -2602 697 -2598
rect 699 -2602 700 -2598
rect 704 -2602 705 -2598
rect 707 -2602 709 -2598
rect 713 -2602 715 -2598
rect 717 -2602 718 -2598
rect 790 -2602 791 -2598
rect 793 -2602 795 -2598
rect 799 -2602 801 -2598
rect 803 -2602 804 -2598
rect 816 -2602 817 -2598
rect 819 -2602 821 -2598
rect 825 -2602 827 -2598
rect 829 -2602 830 -2598
rect 842 -2602 843 -2598
rect 845 -2602 846 -2598
rect 850 -2602 853 -2598
rect 855 -2602 861 -2598
rect 863 -2602 864 -2598
rect 868 -2602 871 -2598
rect 873 -2602 874 -2598
rect 886 -2602 887 -2598
rect 889 -2602 895 -2598
rect 897 -2602 899 -2598
rect 903 -2602 905 -2598
rect 907 -2602 908 -2598
rect 920 -2602 921 -2598
rect 923 -2602 925 -2598
rect 929 -2602 931 -2598
rect 933 -2602 939 -2598
rect 941 -2602 943 -2598
rect 947 -2602 949 -2598
rect 951 -2602 952 -2598
rect 964 -2602 965 -2598
rect 967 -2602 973 -2598
rect 975 -2602 976 -2598
rect 988 -2602 989 -2598
rect 991 -2602 996 -2598
rect 1000 -2602 1005 -2598
rect 1007 -2602 1008 -2598
rect 1012 -2602 1013 -2598
rect 1015 -2602 1017 -2598
rect 1021 -2602 1023 -2598
rect 1025 -2602 1026 -2598
rect -1305 -2734 -1304 -2730
rect -1302 -2734 -1296 -2730
rect -1294 -2734 -1292 -2730
rect -1288 -2734 -1286 -2730
rect -1284 -2734 -1283 -2730
rect -1058 -2734 -1057 -2730
rect -1055 -2734 -1049 -2730
rect -1047 -2734 -1045 -2730
rect -1041 -2734 -1039 -2730
rect -1037 -2734 -1036 -2730
rect -750 -2734 -749 -2730
rect -747 -2734 -741 -2730
rect -739 -2734 -737 -2730
rect -733 -2734 -731 -2730
rect -729 -2734 -728 -2730
rect -442 -2734 -441 -2730
rect -439 -2734 -433 -2730
rect -431 -2734 -429 -2730
rect -425 -2734 -423 -2730
rect -421 -2734 -420 -2730
rect -134 -2734 -133 -2730
rect -131 -2734 -125 -2730
rect -123 -2734 -121 -2730
rect -117 -2734 -115 -2730
rect -113 -2734 -112 -2730
rect 174 -2734 175 -2730
rect 177 -2734 183 -2730
rect 185 -2734 187 -2730
rect 191 -2734 193 -2730
rect 195 -2734 196 -2730
rect 482 -2734 483 -2730
rect 485 -2734 491 -2730
rect 493 -2734 495 -2730
rect 499 -2734 501 -2730
rect 503 -2734 504 -2730
rect 790 -2734 791 -2730
rect 793 -2734 799 -2730
rect 801 -2734 803 -2730
rect 807 -2734 809 -2730
rect 811 -2734 812 -2730
rect -1230 -2893 -1229 -2889
rect -1227 -2893 -1225 -2889
rect -1221 -2893 -1219 -2889
rect -1217 -2893 -1216 -2889
rect -1204 -2893 -1203 -2889
rect -1201 -2893 -1199 -2889
rect -1195 -2893 -1193 -2889
rect -1191 -2893 -1185 -2889
rect -1183 -2893 -1181 -2889
rect -1177 -2893 -1175 -2889
rect -1173 -2893 -1172 -2889
rect -1160 -2893 -1159 -2889
rect -1157 -2893 -1151 -2889
rect -1149 -2893 -1147 -2889
rect -1143 -2893 -1141 -2889
rect -1139 -2893 -1138 -2889
rect -1058 -2893 -1057 -2889
rect -1055 -2893 -1053 -2889
rect -1049 -2893 -1047 -2889
rect -1045 -2893 -1044 -2889
rect -1032 -2893 -1031 -2889
rect -1029 -2893 -1027 -2889
rect -1023 -2893 -1021 -2889
rect -1019 -2893 -1018 -2889
rect -1006 -2893 -1005 -2889
rect -1003 -2893 -1002 -2889
rect -998 -2893 -995 -2889
rect -993 -2893 -987 -2889
rect -985 -2893 -984 -2889
rect -980 -2893 -977 -2889
rect -975 -2893 -974 -2889
rect -962 -2893 -961 -2889
rect -959 -2893 -953 -2889
rect -951 -2893 -949 -2889
rect -945 -2893 -943 -2889
rect -941 -2893 -940 -2889
rect -928 -2893 -927 -2889
rect -925 -2893 -923 -2889
rect -919 -2893 -917 -2889
rect -915 -2893 -909 -2889
rect -907 -2893 -905 -2889
rect -901 -2893 -899 -2889
rect -897 -2893 -896 -2889
rect -884 -2893 -883 -2889
rect -881 -2893 -875 -2889
rect -873 -2893 -872 -2889
rect -860 -2893 -859 -2889
rect -857 -2893 -852 -2889
rect -848 -2893 -843 -2889
rect -841 -2893 -840 -2889
rect -836 -2893 -835 -2889
rect -833 -2893 -831 -2889
rect -827 -2893 -825 -2889
rect -823 -2893 -822 -2889
rect -750 -2893 -749 -2889
rect -747 -2893 -745 -2889
rect -741 -2893 -739 -2889
rect -737 -2893 -736 -2889
rect -724 -2893 -723 -2889
rect -721 -2893 -719 -2889
rect -715 -2893 -713 -2889
rect -711 -2893 -710 -2889
rect -698 -2893 -697 -2889
rect -695 -2893 -694 -2889
rect -690 -2893 -687 -2889
rect -685 -2893 -679 -2889
rect -677 -2893 -676 -2889
rect -672 -2893 -669 -2889
rect -667 -2893 -666 -2889
rect -654 -2893 -653 -2889
rect -651 -2893 -645 -2889
rect -643 -2893 -641 -2889
rect -637 -2893 -635 -2889
rect -633 -2893 -632 -2889
rect -620 -2893 -619 -2889
rect -617 -2893 -615 -2889
rect -611 -2893 -609 -2889
rect -607 -2893 -601 -2889
rect -599 -2893 -597 -2889
rect -593 -2893 -591 -2889
rect -589 -2893 -588 -2889
rect -576 -2893 -575 -2889
rect -573 -2893 -567 -2889
rect -565 -2893 -564 -2889
rect -552 -2893 -551 -2889
rect -549 -2893 -544 -2889
rect -540 -2893 -535 -2889
rect -533 -2893 -532 -2889
rect -528 -2893 -527 -2889
rect -525 -2893 -523 -2889
rect -519 -2893 -517 -2889
rect -515 -2893 -514 -2889
rect -442 -2893 -441 -2889
rect -439 -2893 -437 -2889
rect -433 -2893 -431 -2889
rect -429 -2893 -428 -2889
rect -416 -2893 -415 -2889
rect -413 -2893 -411 -2889
rect -407 -2893 -405 -2889
rect -403 -2893 -402 -2889
rect -390 -2893 -389 -2889
rect -387 -2893 -386 -2889
rect -382 -2893 -379 -2889
rect -377 -2893 -371 -2889
rect -369 -2893 -368 -2889
rect -364 -2893 -361 -2889
rect -359 -2893 -358 -2889
rect -346 -2893 -345 -2889
rect -343 -2893 -337 -2889
rect -335 -2893 -333 -2889
rect -329 -2893 -327 -2889
rect -325 -2893 -324 -2889
rect -312 -2893 -311 -2889
rect -309 -2893 -307 -2889
rect -303 -2893 -301 -2889
rect -299 -2893 -293 -2889
rect -291 -2893 -289 -2889
rect -285 -2893 -283 -2889
rect -281 -2893 -280 -2889
rect -268 -2893 -267 -2889
rect -265 -2893 -259 -2889
rect -257 -2893 -256 -2889
rect -244 -2893 -243 -2889
rect -241 -2893 -236 -2889
rect -232 -2893 -227 -2889
rect -225 -2893 -224 -2889
rect -220 -2893 -219 -2889
rect -217 -2893 -215 -2889
rect -211 -2893 -209 -2889
rect -207 -2893 -206 -2889
rect -134 -2893 -133 -2889
rect -131 -2893 -129 -2889
rect -125 -2893 -123 -2889
rect -121 -2893 -120 -2889
rect -108 -2893 -107 -2889
rect -105 -2893 -103 -2889
rect -99 -2893 -97 -2889
rect -95 -2893 -94 -2889
rect -82 -2893 -81 -2889
rect -79 -2893 -78 -2889
rect -74 -2893 -71 -2889
rect -69 -2893 -63 -2889
rect -61 -2893 -60 -2889
rect -56 -2893 -53 -2889
rect -51 -2893 -50 -2889
rect -38 -2893 -37 -2889
rect -35 -2893 -29 -2889
rect -27 -2893 -25 -2889
rect -21 -2893 -19 -2889
rect -17 -2893 -16 -2889
rect -4 -2893 -3 -2889
rect -1 -2893 1 -2889
rect 5 -2893 7 -2889
rect 9 -2893 15 -2889
rect 17 -2893 19 -2889
rect 23 -2893 25 -2889
rect 27 -2893 28 -2889
rect 40 -2893 41 -2889
rect 43 -2893 49 -2889
rect 51 -2893 52 -2889
rect 64 -2893 65 -2889
rect 67 -2893 72 -2889
rect 76 -2893 81 -2889
rect 83 -2893 84 -2889
rect 88 -2893 89 -2889
rect 91 -2893 93 -2889
rect 97 -2893 99 -2889
rect 101 -2893 102 -2889
rect 174 -2893 175 -2889
rect 177 -2893 179 -2889
rect 183 -2893 185 -2889
rect 187 -2893 188 -2889
rect 200 -2893 201 -2889
rect 203 -2893 205 -2889
rect 209 -2893 211 -2889
rect 213 -2893 214 -2889
rect 226 -2893 227 -2889
rect 229 -2893 230 -2889
rect 234 -2893 237 -2889
rect 239 -2893 245 -2889
rect 247 -2893 248 -2889
rect 252 -2893 255 -2889
rect 257 -2893 258 -2889
rect 270 -2893 271 -2889
rect 273 -2893 279 -2889
rect 281 -2893 283 -2889
rect 287 -2893 289 -2889
rect 291 -2893 292 -2889
rect 304 -2893 305 -2889
rect 307 -2893 309 -2889
rect 313 -2893 315 -2889
rect 317 -2893 323 -2889
rect 325 -2893 327 -2889
rect 331 -2893 333 -2889
rect 335 -2893 336 -2889
rect 348 -2893 349 -2889
rect 351 -2893 357 -2889
rect 359 -2893 360 -2889
rect 372 -2893 373 -2889
rect 375 -2893 380 -2889
rect 384 -2893 389 -2889
rect 391 -2893 392 -2889
rect 396 -2893 397 -2889
rect 399 -2893 401 -2889
rect 405 -2893 407 -2889
rect 409 -2893 410 -2889
rect 482 -2893 483 -2889
rect 485 -2893 487 -2889
rect 491 -2893 493 -2889
rect 495 -2893 496 -2889
rect 508 -2893 509 -2889
rect 511 -2893 513 -2889
rect 517 -2893 519 -2889
rect 521 -2893 522 -2889
rect 534 -2893 535 -2889
rect 537 -2893 538 -2889
rect 542 -2893 545 -2889
rect 547 -2893 553 -2889
rect 555 -2893 556 -2889
rect 560 -2893 563 -2889
rect 565 -2893 566 -2889
rect 578 -2893 579 -2889
rect 581 -2893 587 -2889
rect 589 -2893 591 -2889
rect 595 -2893 597 -2889
rect 599 -2893 600 -2889
rect 612 -2893 613 -2889
rect 615 -2893 617 -2889
rect 621 -2893 623 -2889
rect 625 -2893 631 -2889
rect 633 -2893 635 -2889
rect 639 -2893 641 -2889
rect 643 -2893 644 -2889
rect 656 -2893 657 -2889
rect 659 -2893 665 -2889
rect 667 -2893 668 -2889
rect 680 -2893 681 -2889
rect 683 -2893 688 -2889
rect 692 -2893 697 -2889
rect 699 -2893 700 -2889
rect 704 -2893 705 -2889
rect 707 -2893 709 -2889
rect 713 -2893 715 -2889
rect 717 -2893 718 -2889
rect 790 -2893 791 -2889
rect 793 -2893 795 -2889
rect 799 -2893 801 -2889
rect 803 -2893 804 -2889
rect 816 -2893 817 -2889
rect 819 -2893 821 -2889
rect 825 -2893 827 -2889
rect 829 -2893 830 -2889
rect 842 -2893 843 -2889
rect 845 -2893 846 -2889
rect 850 -2893 853 -2889
rect 855 -2893 861 -2889
rect 863 -2893 864 -2889
rect 868 -2893 871 -2889
rect 873 -2893 874 -2889
rect 886 -2893 887 -2889
rect 889 -2893 895 -2889
rect 897 -2893 899 -2889
rect 903 -2893 905 -2889
rect 907 -2893 908 -2889
rect 920 -2893 921 -2889
rect 923 -2893 925 -2889
rect 929 -2893 931 -2889
rect 933 -2893 939 -2889
rect 941 -2893 943 -2889
rect 947 -2893 949 -2889
rect 951 -2893 952 -2889
rect 964 -2893 965 -2889
rect 967 -2893 973 -2889
rect 975 -2893 976 -2889
rect 988 -2893 989 -2889
rect 991 -2893 996 -2889
rect 1000 -2893 1005 -2889
rect 1007 -2893 1008 -2889
rect 1012 -2893 1013 -2889
rect 1015 -2893 1017 -2889
rect 1021 -2893 1023 -2889
rect 1025 -2893 1026 -2889
rect -1305 -3025 -1304 -3021
rect -1302 -3025 -1296 -3021
rect -1294 -3025 -1292 -3021
rect -1288 -3025 -1286 -3021
rect -1284 -3025 -1283 -3021
rect -1058 -3025 -1057 -3021
rect -1055 -3025 -1049 -3021
rect -1047 -3025 -1045 -3021
rect -1041 -3025 -1039 -3021
rect -1037 -3025 -1036 -3021
rect -750 -3025 -749 -3021
rect -747 -3025 -741 -3021
rect -739 -3025 -737 -3021
rect -733 -3025 -731 -3021
rect -729 -3025 -728 -3021
rect -442 -3025 -441 -3021
rect -439 -3025 -433 -3021
rect -431 -3025 -429 -3021
rect -425 -3025 -423 -3021
rect -421 -3025 -420 -3021
rect -134 -3025 -133 -3021
rect -131 -3025 -125 -3021
rect -123 -3025 -121 -3021
rect -117 -3025 -115 -3021
rect -113 -3025 -112 -3021
rect 174 -3025 175 -3021
rect 177 -3025 183 -3021
rect 185 -3025 187 -3021
rect 191 -3025 193 -3021
rect 195 -3025 196 -3021
rect 482 -3025 483 -3021
rect 485 -3025 491 -3021
rect 493 -3025 495 -3021
rect 499 -3025 501 -3021
rect 503 -3025 504 -3021
rect 790 -3025 791 -3021
rect 793 -3025 799 -3021
rect 801 -3025 803 -3021
rect 807 -3025 809 -3021
rect 811 -3025 812 -3021
rect -1230 -3184 -1229 -3180
rect -1227 -3184 -1225 -3180
rect -1221 -3184 -1219 -3180
rect -1217 -3184 -1216 -3180
rect -1204 -3184 -1203 -3180
rect -1201 -3184 -1199 -3180
rect -1195 -3184 -1193 -3180
rect -1191 -3184 -1185 -3180
rect -1183 -3184 -1181 -3180
rect -1177 -3184 -1175 -3180
rect -1173 -3184 -1172 -3180
rect -1160 -3184 -1159 -3180
rect -1157 -3184 -1151 -3180
rect -1149 -3184 -1147 -3180
rect -1143 -3184 -1141 -3180
rect -1139 -3184 -1138 -3180
rect -1058 -3184 -1057 -3180
rect -1055 -3184 -1053 -3180
rect -1049 -3184 -1047 -3180
rect -1045 -3184 -1044 -3180
rect -1032 -3184 -1031 -3180
rect -1029 -3184 -1027 -3180
rect -1023 -3184 -1021 -3180
rect -1019 -3184 -1018 -3180
rect -1006 -3184 -1005 -3180
rect -1003 -3184 -1002 -3180
rect -998 -3184 -995 -3180
rect -993 -3184 -987 -3180
rect -985 -3184 -984 -3180
rect -980 -3184 -977 -3180
rect -975 -3184 -974 -3180
rect -962 -3184 -961 -3180
rect -959 -3184 -953 -3180
rect -951 -3184 -949 -3180
rect -945 -3184 -943 -3180
rect -941 -3184 -940 -3180
rect -928 -3184 -927 -3180
rect -925 -3184 -923 -3180
rect -919 -3184 -917 -3180
rect -915 -3184 -909 -3180
rect -907 -3184 -905 -3180
rect -901 -3184 -899 -3180
rect -897 -3184 -896 -3180
rect -884 -3184 -883 -3180
rect -881 -3184 -875 -3180
rect -873 -3184 -872 -3180
rect -860 -3184 -859 -3180
rect -857 -3184 -852 -3180
rect -848 -3184 -843 -3180
rect -841 -3184 -840 -3180
rect -836 -3184 -835 -3180
rect -833 -3184 -831 -3180
rect -827 -3184 -825 -3180
rect -823 -3184 -822 -3180
rect -750 -3184 -749 -3180
rect -747 -3184 -745 -3180
rect -741 -3184 -739 -3180
rect -737 -3184 -736 -3180
rect -724 -3184 -723 -3180
rect -721 -3184 -719 -3180
rect -715 -3184 -713 -3180
rect -711 -3184 -710 -3180
rect -698 -3184 -697 -3180
rect -695 -3184 -694 -3180
rect -690 -3184 -687 -3180
rect -685 -3184 -679 -3180
rect -677 -3184 -676 -3180
rect -672 -3184 -669 -3180
rect -667 -3184 -666 -3180
rect -654 -3184 -653 -3180
rect -651 -3184 -645 -3180
rect -643 -3184 -641 -3180
rect -637 -3184 -635 -3180
rect -633 -3184 -632 -3180
rect -620 -3184 -619 -3180
rect -617 -3184 -615 -3180
rect -611 -3184 -609 -3180
rect -607 -3184 -601 -3180
rect -599 -3184 -597 -3180
rect -593 -3184 -591 -3180
rect -589 -3184 -588 -3180
rect -576 -3184 -575 -3180
rect -573 -3184 -567 -3180
rect -565 -3184 -564 -3180
rect -552 -3184 -551 -3180
rect -549 -3184 -544 -3180
rect -540 -3184 -535 -3180
rect -533 -3184 -532 -3180
rect -528 -3184 -527 -3180
rect -525 -3184 -523 -3180
rect -519 -3184 -517 -3180
rect -515 -3184 -514 -3180
rect -442 -3184 -441 -3180
rect -439 -3184 -437 -3180
rect -433 -3184 -431 -3180
rect -429 -3184 -428 -3180
rect -416 -3184 -415 -3180
rect -413 -3184 -411 -3180
rect -407 -3184 -405 -3180
rect -403 -3184 -402 -3180
rect -390 -3184 -389 -3180
rect -387 -3184 -386 -3180
rect -382 -3184 -379 -3180
rect -377 -3184 -371 -3180
rect -369 -3184 -368 -3180
rect -364 -3184 -361 -3180
rect -359 -3184 -358 -3180
rect -346 -3184 -345 -3180
rect -343 -3184 -337 -3180
rect -335 -3184 -333 -3180
rect -329 -3184 -327 -3180
rect -325 -3184 -324 -3180
rect -312 -3184 -311 -3180
rect -309 -3184 -307 -3180
rect -303 -3184 -301 -3180
rect -299 -3184 -293 -3180
rect -291 -3184 -289 -3180
rect -285 -3184 -283 -3180
rect -281 -3184 -280 -3180
rect -268 -3184 -267 -3180
rect -265 -3184 -259 -3180
rect -257 -3184 -256 -3180
rect -244 -3184 -243 -3180
rect -241 -3184 -236 -3180
rect -232 -3184 -227 -3180
rect -225 -3184 -224 -3180
rect -220 -3184 -219 -3180
rect -217 -3184 -215 -3180
rect -211 -3184 -209 -3180
rect -207 -3184 -206 -3180
rect -134 -3184 -133 -3180
rect -131 -3184 -129 -3180
rect -125 -3184 -123 -3180
rect -121 -3184 -120 -3180
rect -108 -3184 -107 -3180
rect -105 -3184 -103 -3180
rect -99 -3184 -97 -3180
rect -95 -3184 -94 -3180
rect -82 -3184 -81 -3180
rect -79 -3184 -78 -3180
rect -74 -3184 -71 -3180
rect -69 -3184 -63 -3180
rect -61 -3184 -60 -3180
rect -56 -3184 -53 -3180
rect -51 -3184 -50 -3180
rect -38 -3184 -37 -3180
rect -35 -3184 -29 -3180
rect -27 -3184 -25 -3180
rect -21 -3184 -19 -3180
rect -17 -3184 -16 -3180
rect -4 -3184 -3 -3180
rect -1 -3184 1 -3180
rect 5 -3184 7 -3180
rect 9 -3184 15 -3180
rect 17 -3184 19 -3180
rect 23 -3184 25 -3180
rect 27 -3184 28 -3180
rect 40 -3184 41 -3180
rect 43 -3184 49 -3180
rect 51 -3184 52 -3180
rect 64 -3184 65 -3180
rect 67 -3184 72 -3180
rect 76 -3184 81 -3180
rect 83 -3184 84 -3180
rect 88 -3184 89 -3180
rect 91 -3184 93 -3180
rect 97 -3184 99 -3180
rect 101 -3184 102 -3180
rect 174 -3184 175 -3180
rect 177 -3184 179 -3180
rect 183 -3184 185 -3180
rect 187 -3184 188 -3180
rect 200 -3184 201 -3180
rect 203 -3184 205 -3180
rect 209 -3184 211 -3180
rect 213 -3184 214 -3180
rect 226 -3184 227 -3180
rect 229 -3184 230 -3180
rect 234 -3184 237 -3180
rect 239 -3184 245 -3180
rect 247 -3184 248 -3180
rect 252 -3184 255 -3180
rect 257 -3184 258 -3180
rect 270 -3184 271 -3180
rect 273 -3184 279 -3180
rect 281 -3184 283 -3180
rect 287 -3184 289 -3180
rect 291 -3184 292 -3180
rect 304 -3184 305 -3180
rect 307 -3184 309 -3180
rect 313 -3184 315 -3180
rect 317 -3184 323 -3180
rect 325 -3184 327 -3180
rect 331 -3184 333 -3180
rect 335 -3184 336 -3180
rect 348 -3184 349 -3180
rect 351 -3184 357 -3180
rect 359 -3184 360 -3180
rect 372 -3184 373 -3180
rect 375 -3184 380 -3180
rect 384 -3184 389 -3180
rect 391 -3184 392 -3180
rect 396 -3184 397 -3180
rect 399 -3184 401 -3180
rect 405 -3184 407 -3180
rect 409 -3184 410 -3180
rect 482 -3184 483 -3180
rect 485 -3184 487 -3180
rect 491 -3184 493 -3180
rect 495 -3184 496 -3180
rect 508 -3184 509 -3180
rect 511 -3184 513 -3180
rect 517 -3184 519 -3180
rect 521 -3184 522 -3180
rect 534 -3184 535 -3180
rect 537 -3184 538 -3180
rect 542 -3184 545 -3180
rect 547 -3184 553 -3180
rect 555 -3184 556 -3180
rect 560 -3184 563 -3180
rect 565 -3184 566 -3180
rect 578 -3184 579 -3180
rect 581 -3184 587 -3180
rect 589 -3184 591 -3180
rect 595 -3184 597 -3180
rect 599 -3184 600 -3180
rect 612 -3184 613 -3180
rect 615 -3184 617 -3180
rect 621 -3184 623 -3180
rect 625 -3184 631 -3180
rect 633 -3184 635 -3180
rect 639 -3184 641 -3180
rect 643 -3184 644 -3180
rect 656 -3184 657 -3180
rect 659 -3184 665 -3180
rect 667 -3184 668 -3180
rect 680 -3184 681 -3180
rect 683 -3184 688 -3180
rect 692 -3184 697 -3180
rect 699 -3184 700 -3180
rect 704 -3184 705 -3180
rect 707 -3184 709 -3180
rect 713 -3184 715 -3180
rect 717 -3184 718 -3180
rect 790 -3184 791 -3180
rect 793 -3184 795 -3180
rect 799 -3184 801 -3180
rect 803 -3184 804 -3180
rect 816 -3184 817 -3180
rect 819 -3184 821 -3180
rect 825 -3184 827 -3180
rect 829 -3184 830 -3180
rect 842 -3184 843 -3180
rect 845 -3184 846 -3180
rect 850 -3184 853 -3180
rect 855 -3184 861 -3180
rect 863 -3184 864 -3180
rect 868 -3184 871 -3180
rect 873 -3184 874 -3180
rect 886 -3184 887 -3180
rect 889 -3184 895 -3180
rect 897 -3184 899 -3180
rect 903 -3184 905 -3180
rect 907 -3184 908 -3180
rect 920 -3184 921 -3180
rect 923 -3184 925 -3180
rect 929 -3184 931 -3180
rect 933 -3184 939 -3180
rect 941 -3184 943 -3180
rect 947 -3184 949 -3180
rect 951 -3184 952 -3180
rect 964 -3184 965 -3180
rect 967 -3184 973 -3180
rect 975 -3184 976 -3180
rect 988 -3184 989 -3180
rect 991 -3184 996 -3180
rect 1000 -3184 1005 -3180
rect 1007 -3184 1008 -3180
rect 1012 -3184 1013 -3180
rect 1015 -3184 1017 -3180
rect 1021 -3184 1023 -3180
rect 1025 -3184 1026 -3180
<< pdiffusion >>
rect -1303 -996 -1302 -988
rect -1300 -996 -1299 -988
rect -1295 -996 -1294 -988
rect -1292 -996 -1290 -988
rect -1286 -996 -1284 -988
rect -1282 -996 -1281 -988
rect -1059 -996 -1058 -988
rect -1056 -996 -1055 -988
rect -1051 -996 -1050 -988
rect -1048 -996 -1046 -988
rect -1042 -996 -1040 -988
rect -1038 -996 -1037 -988
rect -750 -996 -749 -988
rect -747 -996 -746 -988
rect -742 -996 -741 -988
rect -739 -996 -737 -988
rect -733 -996 -731 -988
rect -729 -996 -728 -988
rect -442 -996 -441 -988
rect -439 -996 -438 -988
rect -434 -996 -433 -988
rect -431 -996 -429 -988
rect -425 -996 -423 -988
rect -421 -996 -420 -988
rect -135 -996 -134 -988
rect -132 -996 -131 -988
rect -127 -996 -126 -988
rect -124 -996 -122 -988
rect -118 -996 -116 -988
rect -114 -996 -113 -988
rect 174 -996 175 -988
rect 177 -996 178 -988
rect 182 -996 183 -988
rect 185 -996 187 -988
rect 191 -996 193 -988
rect 195 -996 196 -988
rect 482 -996 483 -988
rect 485 -996 486 -988
rect 490 -996 491 -988
rect 493 -996 495 -988
rect 499 -996 501 -988
rect 503 -996 504 -988
rect 790 -996 791 -988
rect 793 -996 794 -988
rect 798 -996 799 -988
rect 801 -996 803 -988
rect 807 -996 809 -988
rect 811 -996 812 -988
rect -1305 -1146 -1304 -1138
rect -1302 -1146 -1301 -1138
rect -1297 -1146 -1296 -1138
rect -1294 -1146 -1292 -1138
rect -1288 -1146 -1286 -1138
rect -1284 -1146 -1283 -1138
rect -1058 -1146 -1057 -1138
rect -1055 -1146 -1054 -1138
rect -1050 -1146 -1049 -1138
rect -1047 -1146 -1045 -1138
rect -1041 -1146 -1039 -1138
rect -1037 -1146 -1036 -1138
rect -750 -1146 -749 -1138
rect -747 -1146 -746 -1138
rect -742 -1146 -741 -1138
rect -739 -1146 -737 -1138
rect -733 -1146 -731 -1138
rect -729 -1146 -728 -1138
rect -442 -1146 -441 -1138
rect -439 -1146 -438 -1138
rect -434 -1146 -433 -1138
rect -431 -1146 -429 -1138
rect -425 -1146 -423 -1138
rect -421 -1146 -420 -1138
rect -134 -1146 -133 -1138
rect -131 -1146 -130 -1138
rect -126 -1146 -125 -1138
rect -123 -1146 -121 -1138
rect -117 -1146 -115 -1138
rect -113 -1146 -112 -1138
rect 174 -1146 175 -1138
rect 177 -1146 178 -1138
rect 182 -1146 183 -1138
rect 185 -1146 187 -1138
rect 191 -1146 193 -1138
rect 195 -1146 196 -1138
rect 482 -1146 483 -1138
rect 485 -1146 486 -1138
rect 490 -1146 491 -1138
rect 493 -1146 495 -1138
rect 499 -1146 501 -1138
rect 503 -1146 504 -1138
rect 790 -1146 791 -1138
rect 793 -1146 794 -1138
rect 798 -1146 799 -1138
rect 801 -1146 803 -1138
rect 807 -1146 809 -1138
rect 811 -1146 812 -1138
rect -1226 -1310 -1225 -1302
rect -1223 -1310 -1221 -1302
rect -1217 -1310 -1215 -1302
rect -1213 -1310 -1212 -1302
rect -1200 -1310 -1199 -1302
rect -1197 -1310 -1189 -1302
rect -1187 -1310 -1186 -1302
rect -1182 -1310 -1181 -1302
rect -1179 -1310 -1171 -1302
rect -1169 -1310 -1164 -1302
rect -1160 -1310 -1155 -1302
rect -1153 -1310 -1152 -1302
rect -1148 -1310 -1147 -1302
rect -1145 -1310 -1143 -1302
rect -1139 -1310 -1137 -1302
rect -1135 -1310 -1134 -1302
rect -1058 -1310 -1057 -1302
rect -1055 -1310 -1053 -1302
rect -1049 -1310 -1047 -1302
rect -1045 -1310 -1044 -1302
rect -1032 -1310 -1031 -1302
rect -1029 -1310 -1027 -1302
rect -1023 -1310 -1021 -1302
rect -1019 -1310 -1018 -1302
rect -1006 -1310 -1005 -1302
rect -1003 -1310 -995 -1302
rect -993 -1310 -992 -1302
rect -988 -1310 -987 -1302
rect -985 -1310 -977 -1302
rect -975 -1310 -970 -1302
rect -966 -1310 -961 -1302
rect -959 -1310 -958 -1302
rect -954 -1310 -953 -1302
rect -951 -1310 -949 -1302
rect -945 -1310 -943 -1302
rect -941 -1310 -940 -1302
rect -928 -1310 -927 -1302
rect -925 -1310 -917 -1302
rect -915 -1310 -914 -1302
rect -910 -1310 -909 -1302
rect -907 -1310 -899 -1302
rect -897 -1310 -892 -1302
rect -888 -1310 -883 -1302
rect -881 -1310 -880 -1302
rect -876 -1310 -875 -1302
rect -873 -1310 -868 -1302
rect -864 -1310 -859 -1302
rect -857 -1310 -856 -1302
rect -844 -1310 -843 -1302
rect -841 -1310 -835 -1302
rect -833 -1310 -831 -1302
rect -827 -1310 -825 -1302
rect -823 -1310 -822 -1302
rect -750 -1310 -749 -1302
rect -747 -1310 -745 -1302
rect -741 -1310 -739 -1302
rect -737 -1310 -736 -1302
rect -724 -1310 -723 -1302
rect -721 -1310 -719 -1302
rect -715 -1310 -713 -1302
rect -711 -1310 -710 -1302
rect -698 -1310 -697 -1302
rect -695 -1310 -687 -1302
rect -685 -1310 -684 -1302
rect -680 -1310 -679 -1302
rect -677 -1310 -669 -1302
rect -667 -1310 -662 -1302
rect -658 -1310 -653 -1302
rect -651 -1310 -650 -1302
rect -646 -1310 -645 -1302
rect -643 -1310 -641 -1302
rect -637 -1310 -635 -1302
rect -633 -1310 -632 -1302
rect -620 -1310 -619 -1302
rect -617 -1310 -609 -1302
rect -607 -1310 -606 -1302
rect -602 -1310 -601 -1302
rect -599 -1310 -591 -1302
rect -589 -1310 -584 -1302
rect -580 -1310 -575 -1302
rect -573 -1310 -572 -1302
rect -568 -1310 -567 -1302
rect -565 -1310 -560 -1302
rect -556 -1310 -551 -1302
rect -549 -1310 -548 -1302
rect -536 -1310 -535 -1302
rect -533 -1310 -527 -1302
rect -525 -1310 -523 -1302
rect -519 -1310 -517 -1302
rect -515 -1310 -514 -1302
rect -442 -1310 -441 -1302
rect -439 -1310 -437 -1302
rect -433 -1310 -431 -1302
rect -429 -1310 -428 -1302
rect -416 -1310 -415 -1302
rect -413 -1310 -411 -1302
rect -407 -1310 -405 -1302
rect -403 -1310 -402 -1302
rect -390 -1310 -389 -1302
rect -387 -1310 -379 -1302
rect -377 -1310 -376 -1302
rect -372 -1310 -371 -1302
rect -369 -1310 -361 -1302
rect -359 -1310 -354 -1302
rect -350 -1310 -345 -1302
rect -343 -1310 -342 -1302
rect -338 -1310 -337 -1302
rect -335 -1310 -333 -1302
rect -329 -1310 -327 -1302
rect -325 -1310 -324 -1302
rect -312 -1310 -311 -1302
rect -309 -1310 -301 -1302
rect -299 -1310 -298 -1302
rect -294 -1310 -293 -1302
rect -291 -1310 -283 -1302
rect -281 -1310 -276 -1302
rect -272 -1310 -267 -1302
rect -265 -1310 -264 -1302
rect -260 -1310 -259 -1302
rect -257 -1310 -252 -1302
rect -248 -1310 -243 -1302
rect -241 -1310 -240 -1302
rect -228 -1310 -227 -1302
rect -225 -1310 -219 -1302
rect -217 -1310 -215 -1302
rect -211 -1310 -209 -1302
rect -207 -1310 -206 -1302
rect -134 -1310 -133 -1302
rect -131 -1310 -129 -1302
rect -125 -1310 -123 -1302
rect -121 -1310 -120 -1302
rect -108 -1310 -107 -1302
rect -105 -1310 -103 -1302
rect -99 -1310 -97 -1302
rect -95 -1310 -94 -1302
rect -82 -1310 -81 -1302
rect -79 -1310 -71 -1302
rect -69 -1310 -68 -1302
rect -64 -1310 -63 -1302
rect -61 -1310 -53 -1302
rect -51 -1310 -46 -1302
rect -42 -1310 -37 -1302
rect -35 -1310 -34 -1302
rect -30 -1310 -29 -1302
rect -27 -1310 -25 -1302
rect -21 -1310 -19 -1302
rect -17 -1310 -16 -1302
rect -4 -1310 -3 -1302
rect -1 -1310 7 -1302
rect 9 -1310 10 -1302
rect 14 -1310 15 -1302
rect 17 -1310 25 -1302
rect 27 -1310 32 -1302
rect 36 -1310 41 -1302
rect 43 -1310 44 -1302
rect 48 -1310 49 -1302
rect 51 -1310 56 -1302
rect 60 -1310 65 -1302
rect 67 -1310 68 -1302
rect 80 -1310 81 -1302
rect 83 -1310 89 -1302
rect 91 -1310 93 -1302
rect 97 -1310 99 -1302
rect 101 -1310 102 -1302
rect 174 -1310 175 -1302
rect 177 -1310 179 -1302
rect 183 -1310 185 -1302
rect 187 -1310 188 -1302
rect 200 -1310 201 -1302
rect 203 -1310 205 -1302
rect 209 -1310 211 -1302
rect 213 -1310 214 -1302
rect 226 -1310 227 -1302
rect 229 -1310 237 -1302
rect 239 -1310 240 -1302
rect 244 -1310 245 -1302
rect 247 -1310 255 -1302
rect 257 -1310 262 -1302
rect 266 -1310 271 -1302
rect 273 -1310 274 -1302
rect 278 -1310 279 -1302
rect 281 -1310 283 -1302
rect 287 -1310 289 -1302
rect 291 -1310 292 -1302
rect 304 -1310 305 -1302
rect 307 -1310 315 -1302
rect 317 -1310 318 -1302
rect 322 -1310 323 -1302
rect 325 -1310 333 -1302
rect 335 -1310 340 -1302
rect 344 -1310 349 -1302
rect 351 -1310 352 -1302
rect 356 -1310 357 -1302
rect 359 -1310 364 -1302
rect 368 -1310 373 -1302
rect 375 -1310 376 -1302
rect 388 -1310 389 -1302
rect 391 -1310 397 -1302
rect 399 -1310 401 -1302
rect 405 -1310 407 -1302
rect 409 -1310 410 -1302
rect 482 -1310 483 -1302
rect 485 -1310 487 -1302
rect 491 -1310 493 -1302
rect 495 -1310 496 -1302
rect 508 -1310 509 -1302
rect 511 -1310 513 -1302
rect 517 -1310 519 -1302
rect 521 -1310 522 -1302
rect 534 -1310 535 -1302
rect 537 -1310 545 -1302
rect 547 -1310 548 -1302
rect 552 -1310 553 -1302
rect 555 -1310 563 -1302
rect 565 -1310 570 -1302
rect 574 -1310 579 -1302
rect 581 -1310 582 -1302
rect 586 -1310 587 -1302
rect 589 -1310 591 -1302
rect 595 -1310 597 -1302
rect 599 -1310 600 -1302
rect 612 -1310 613 -1302
rect 615 -1310 623 -1302
rect 625 -1310 626 -1302
rect 630 -1310 631 -1302
rect 633 -1310 641 -1302
rect 643 -1310 648 -1302
rect 652 -1310 657 -1302
rect 659 -1310 660 -1302
rect 664 -1310 665 -1302
rect 667 -1310 672 -1302
rect 676 -1310 681 -1302
rect 683 -1310 684 -1302
rect 696 -1310 697 -1302
rect 699 -1310 705 -1302
rect 707 -1310 709 -1302
rect 713 -1310 715 -1302
rect 717 -1310 718 -1302
rect 788 -1310 789 -1302
rect 791 -1310 793 -1302
rect 797 -1310 799 -1302
rect 801 -1310 802 -1302
rect 814 -1310 815 -1302
rect 817 -1310 825 -1302
rect 827 -1310 828 -1302
rect 832 -1310 833 -1302
rect 835 -1310 843 -1302
rect 845 -1310 850 -1302
rect 854 -1310 859 -1302
rect 861 -1310 862 -1302
rect 866 -1310 867 -1302
rect 869 -1310 871 -1302
rect 875 -1310 877 -1302
rect 879 -1310 880 -1302
rect -1305 -1467 -1304 -1459
rect -1302 -1467 -1301 -1459
rect -1297 -1467 -1296 -1459
rect -1294 -1467 -1292 -1459
rect -1288 -1467 -1286 -1459
rect -1284 -1467 -1283 -1459
rect -1058 -1467 -1057 -1459
rect -1055 -1467 -1054 -1459
rect -1050 -1467 -1049 -1459
rect -1047 -1467 -1045 -1459
rect -1041 -1467 -1039 -1459
rect -1037 -1467 -1036 -1459
rect -750 -1467 -749 -1459
rect -747 -1467 -746 -1459
rect -742 -1467 -741 -1459
rect -739 -1467 -737 -1459
rect -733 -1467 -731 -1459
rect -729 -1467 -728 -1459
rect -442 -1467 -441 -1459
rect -439 -1467 -438 -1459
rect -434 -1467 -433 -1459
rect -431 -1467 -429 -1459
rect -425 -1467 -423 -1459
rect -421 -1467 -420 -1459
rect -134 -1467 -133 -1459
rect -131 -1467 -130 -1459
rect -126 -1467 -125 -1459
rect -123 -1467 -121 -1459
rect -117 -1467 -115 -1459
rect -113 -1467 -112 -1459
rect 174 -1467 175 -1459
rect 177 -1467 178 -1459
rect 182 -1467 183 -1459
rect 185 -1467 187 -1459
rect 191 -1467 193 -1459
rect 195 -1467 196 -1459
rect 482 -1467 483 -1459
rect 485 -1467 486 -1459
rect 490 -1467 491 -1459
rect 493 -1467 495 -1459
rect 499 -1467 501 -1459
rect 503 -1467 504 -1459
rect 790 -1467 791 -1459
rect 793 -1467 794 -1459
rect 798 -1467 799 -1459
rect 801 -1467 803 -1459
rect 807 -1467 809 -1459
rect 811 -1467 812 -1459
rect -1230 -1626 -1229 -1618
rect -1227 -1626 -1225 -1618
rect -1221 -1626 -1219 -1618
rect -1217 -1626 -1216 -1618
rect -1204 -1626 -1203 -1618
rect -1201 -1626 -1193 -1618
rect -1191 -1626 -1190 -1618
rect -1186 -1626 -1185 -1618
rect -1183 -1626 -1175 -1618
rect -1173 -1626 -1168 -1618
rect -1164 -1626 -1159 -1618
rect -1157 -1626 -1156 -1618
rect -1152 -1626 -1151 -1618
rect -1149 -1626 -1147 -1618
rect -1143 -1626 -1141 -1618
rect -1139 -1626 -1138 -1618
rect -1058 -1626 -1057 -1618
rect -1055 -1626 -1053 -1618
rect -1049 -1626 -1047 -1618
rect -1045 -1626 -1044 -1618
rect -1032 -1626 -1031 -1618
rect -1029 -1626 -1027 -1618
rect -1023 -1626 -1021 -1618
rect -1019 -1626 -1018 -1618
rect -1006 -1626 -1005 -1618
rect -1003 -1626 -995 -1618
rect -993 -1626 -992 -1618
rect -988 -1626 -987 -1618
rect -985 -1626 -977 -1618
rect -975 -1626 -970 -1618
rect -966 -1626 -961 -1618
rect -959 -1626 -958 -1618
rect -954 -1626 -953 -1618
rect -951 -1626 -949 -1618
rect -945 -1626 -943 -1618
rect -941 -1626 -940 -1618
rect -928 -1626 -927 -1618
rect -925 -1626 -917 -1618
rect -915 -1626 -914 -1618
rect -910 -1626 -909 -1618
rect -907 -1626 -899 -1618
rect -897 -1626 -892 -1618
rect -888 -1626 -883 -1618
rect -881 -1626 -880 -1618
rect -876 -1626 -875 -1618
rect -873 -1626 -868 -1618
rect -864 -1626 -859 -1618
rect -857 -1626 -856 -1618
rect -844 -1626 -843 -1618
rect -841 -1626 -835 -1618
rect -833 -1626 -831 -1618
rect -827 -1626 -825 -1618
rect -823 -1626 -822 -1618
rect -750 -1626 -749 -1618
rect -747 -1626 -745 -1618
rect -741 -1626 -739 -1618
rect -737 -1626 -736 -1618
rect -724 -1626 -723 -1618
rect -721 -1626 -719 -1618
rect -715 -1626 -713 -1618
rect -711 -1626 -710 -1618
rect -698 -1626 -697 -1618
rect -695 -1626 -687 -1618
rect -685 -1626 -684 -1618
rect -680 -1626 -679 -1618
rect -677 -1626 -669 -1618
rect -667 -1626 -662 -1618
rect -658 -1626 -653 -1618
rect -651 -1626 -650 -1618
rect -646 -1626 -645 -1618
rect -643 -1626 -641 -1618
rect -637 -1626 -635 -1618
rect -633 -1626 -632 -1618
rect -620 -1626 -619 -1618
rect -617 -1626 -609 -1618
rect -607 -1626 -606 -1618
rect -602 -1626 -601 -1618
rect -599 -1626 -591 -1618
rect -589 -1626 -584 -1618
rect -580 -1626 -575 -1618
rect -573 -1626 -572 -1618
rect -568 -1626 -567 -1618
rect -565 -1626 -560 -1618
rect -556 -1626 -551 -1618
rect -549 -1626 -548 -1618
rect -536 -1626 -535 -1618
rect -533 -1626 -527 -1618
rect -525 -1626 -523 -1618
rect -519 -1626 -517 -1618
rect -515 -1626 -514 -1618
rect -442 -1626 -441 -1618
rect -439 -1626 -437 -1618
rect -433 -1626 -431 -1618
rect -429 -1626 -428 -1618
rect -416 -1626 -415 -1618
rect -413 -1626 -411 -1618
rect -407 -1626 -405 -1618
rect -403 -1626 -402 -1618
rect -390 -1626 -389 -1618
rect -387 -1626 -379 -1618
rect -377 -1626 -376 -1618
rect -372 -1626 -371 -1618
rect -369 -1626 -361 -1618
rect -359 -1626 -354 -1618
rect -350 -1626 -345 -1618
rect -343 -1626 -342 -1618
rect -338 -1626 -337 -1618
rect -335 -1626 -333 -1618
rect -329 -1626 -327 -1618
rect -325 -1626 -324 -1618
rect -312 -1626 -311 -1618
rect -309 -1626 -301 -1618
rect -299 -1626 -298 -1618
rect -294 -1626 -293 -1618
rect -291 -1626 -283 -1618
rect -281 -1626 -276 -1618
rect -272 -1626 -267 -1618
rect -265 -1626 -264 -1618
rect -260 -1626 -259 -1618
rect -257 -1626 -252 -1618
rect -248 -1626 -243 -1618
rect -241 -1626 -240 -1618
rect -228 -1626 -227 -1618
rect -225 -1626 -219 -1618
rect -217 -1626 -215 -1618
rect -211 -1626 -209 -1618
rect -207 -1626 -206 -1618
rect -134 -1626 -133 -1618
rect -131 -1626 -129 -1618
rect -125 -1626 -123 -1618
rect -121 -1626 -120 -1618
rect -108 -1626 -107 -1618
rect -105 -1626 -103 -1618
rect -99 -1626 -97 -1618
rect -95 -1626 -94 -1618
rect -82 -1626 -81 -1618
rect -79 -1626 -71 -1618
rect -69 -1626 -68 -1618
rect -64 -1626 -63 -1618
rect -61 -1626 -53 -1618
rect -51 -1626 -46 -1618
rect -42 -1626 -37 -1618
rect -35 -1626 -34 -1618
rect -30 -1626 -29 -1618
rect -27 -1626 -25 -1618
rect -21 -1626 -19 -1618
rect -17 -1626 -16 -1618
rect -4 -1626 -3 -1618
rect -1 -1626 7 -1618
rect 9 -1626 10 -1618
rect 14 -1626 15 -1618
rect 17 -1626 25 -1618
rect 27 -1626 32 -1618
rect 36 -1626 41 -1618
rect 43 -1626 44 -1618
rect 48 -1626 49 -1618
rect 51 -1626 56 -1618
rect 60 -1626 65 -1618
rect 67 -1626 68 -1618
rect 80 -1626 81 -1618
rect 83 -1626 89 -1618
rect 91 -1626 93 -1618
rect 97 -1626 99 -1618
rect 101 -1626 102 -1618
rect 174 -1626 175 -1618
rect 177 -1626 179 -1618
rect 183 -1626 185 -1618
rect 187 -1626 188 -1618
rect 200 -1626 201 -1618
rect 203 -1626 205 -1618
rect 209 -1626 211 -1618
rect 213 -1626 214 -1618
rect 226 -1626 227 -1618
rect 229 -1626 237 -1618
rect 239 -1626 240 -1618
rect 244 -1626 245 -1618
rect 247 -1626 255 -1618
rect 257 -1626 262 -1618
rect 266 -1626 271 -1618
rect 273 -1626 274 -1618
rect 278 -1626 279 -1618
rect 281 -1626 283 -1618
rect 287 -1626 289 -1618
rect 291 -1626 292 -1618
rect 304 -1626 305 -1618
rect 307 -1626 315 -1618
rect 317 -1626 318 -1618
rect 322 -1626 323 -1618
rect 325 -1626 333 -1618
rect 335 -1626 340 -1618
rect 344 -1626 349 -1618
rect 351 -1626 352 -1618
rect 356 -1626 357 -1618
rect 359 -1626 364 -1618
rect 368 -1626 373 -1618
rect 375 -1626 376 -1618
rect 388 -1626 389 -1618
rect 391 -1626 397 -1618
rect 399 -1626 401 -1618
rect 405 -1626 407 -1618
rect 409 -1626 410 -1618
rect 482 -1626 483 -1618
rect 485 -1626 487 -1618
rect 491 -1626 493 -1618
rect 495 -1626 496 -1618
rect 508 -1626 509 -1618
rect 511 -1626 513 -1618
rect 517 -1626 519 -1618
rect 521 -1626 522 -1618
rect 534 -1626 535 -1618
rect 537 -1626 545 -1618
rect 547 -1626 548 -1618
rect 552 -1626 553 -1618
rect 555 -1626 563 -1618
rect 565 -1626 570 -1618
rect 574 -1626 579 -1618
rect 581 -1626 582 -1618
rect 586 -1626 587 -1618
rect 589 -1626 591 -1618
rect 595 -1626 597 -1618
rect 599 -1626 600 -1618
rect 612 -1626 613 -1618
rect 615 -1626 623 -1618
rect 625 -1626 626 -1618
rect 630 -1626 631 -1618
rect 633 -1626 641 -1618
rect 643 -1626 648 -1618
rect 652 -1626 657 -1618
rect 659 -1626 660 -1618
rect 664 -1626 665 -1618
rect 667 -1626 672 -1618
rect 676 -1626 681 -1618
rect 683 -1626 684 -1618
rect 696 -1626 697 -1618
rect 699 -1626 705 -1618
rect 707 -1626 709 -1618
rect 713 -1626 715 -1618
rect 717 -1626 718 -1618
rect 790 -1626 791 -1618
rect 793 -1626 795 -1618
rect 799 -1626 801 -1618
rect 803 -1626 804 -1618
rect 816 -1626 817 -1618
rect 819 -1626 821 -1618
rect 825 -1626 827 -1618
rect 829 -1626 830 -1618
rect 842 -1626 843 -1618
rect 845 -1626 853 -1618
rect 855 -1626 856 -1618
rect 860 -1626 861 -1618
rect 863 -1626 871 -1618
rect 873 -1626 878 -1618
rect 882 -1626 887 -1618
rect 889 -1626 890 -1618
rect 894 -1626 895 -1618
rect 897 -1626 899 -1618
rect 903 -1626 905 -1618
rect 907 -1626 908 -1618
rect 920 -1626 921 -1618
rect 923 -1626 931 -1618
rect 933 -1626 934 -1618
rect 938 -1626 939 -1618
rect 941 -1626 949 -1618
rect 951 -1626 956 -1618
rect 960 -1626 965 -1618
rect 967 -1626 968 -1618
rect 972 -1626 973 -1618
rect 975 -1626 980 -1618
rect 984 -1626 989 -1618
rect 991 -1626 992 -1618
rect 1004 -1626 1005 -1618
rect 1007 -1626 1013 -1618
rect 1015 -1626 1017 -1618
rect 1021 -1626 1023 -1618
rect 1025 -1626 1026 -1618
rect -1305 -1758 -1304 -1750
rect -1302 -1758 -1301 -1750
rect -1297 -1758 -1296 -1750
rect -1294 -1758 -1292 -1750
rect -1288 -1758 -1286 -1750
rect -1284 -1758 -1283 -1750
rect -1058 -1758 -1057 -1750
rect -1055 -1758 -1054 -1750
rect -1050 -1758 -1049 -1750
rect -1047 -1758 -1045 -1750
rect -1041 -1758 -1039 -1750
rect -1037 -1758 -1036 -1750
rect -750 -1758 -749 -1750
rect -747 -1758 -746 -1750
rect -742 -1758 -741 -1750
rect -739 -1758 -737 -1750
rect -733 -1758 -731 -1750
rect -729 -1758 -728 -1750
rect -442 -1758 -441 -1750
rect -439 -1758 -438 -1750
rect -434 -1758 -433 -1750
rect -431 -1758 -429 -1750
rect -425 -1758 -423 -1750
rect -421 -1758 -420 -1750
rect -134 -1758 -133 -1750
rect -131 -1758 -130 -1750
rect -126 -1758 -125 -1750
rect -123 -1758 -121 -1750
rect -117 -1758 -115 -1750
rect -113 -1758 -112 -1750
rect 174 -1758 175 -1750
rect 177 -1758 178 -1750
rect 182 -1758 183 -1750
rect 185 -1758 187 -1750
rect 191 -1758 193 -1750
rect 195 -1758 196 -1750
rect 482 -1758 483 -1750
rect 485 -1758 486 -1750
rect 490 -1758 491 -1750
rect 493 -1758 495 -1750
rect 499 -1758 501 -1750
rect 503 -1758 504 -1750
rect 790 -1758 791 -1750
rect 793 -1758 794 -1750
rect 798 -1758 799 -1750
rect 801 -1758 803 -1750
rect 807 -1758 809 -1750
rect 811 -1758 812 -1750
rect -1230 -1917 -1229 -1909
rect -1227 -1917 -1225 -1909
rect -1221 -1917 -1219 -1909
rect -1217 -1917 -1216 -1909
rect -1204 -1917 -1203 -1909
rect -1201 -1917 -1193 -1909
rect -1191 -1917 -1190 -1909
rect -1186 -1917 -1185 -1909
rect -1183 -1917 -1175 -1909
rect -1173 -1917 -1168 -1909
rect -1164 -1917 -1159 -1909
rect -1157 -1917 -1156 -1909
rect -1152 -1917 -1151 -1909
rect -1149 -1917 -1147 -1909
rect -1143 -1917 -1141 -1909
rect -1139 -1917 -1138 -1909
rect -1058 -1917 -1057 -1909
rect -1055 -1917 -1053 -1909
rect -1049 -1917 -1047 -1909
rect -1045 -1917 -1044 -1909
rect -1032 -1917 -1031 -1909
rect -1029 -1917 -1027 -1909
rect -1023 -1917 -1021 -1909
rect -1019 -1917 -1018 -1909
rect -1006 -1917 -1005 -1909
rect -1003 -1917 -995 -1909
rect -993 -1917 -992 -1909
rect -988 -1917 -987 -1909
rect -985 -1917 -977 -1909
rect -975 -1917 -970 -1909
rect -966 -1917 -961 -1909
rect -959 -1917 -958 -1909
rect -954 -1917 -953 -1909
rect -951 -1917 -949 -1909
rect -945 -1917 -943 -1909
rect -941 -1917 -940 -1909
rect -928 -1917 -927 -1909
rect -925 -1917 -917 -1909
rect -915 -1917 -914 -1909
rect -910 -1917 -909 -1909
rect -907 -1917 -899 -1909
rect -897 -1917 -892 -1909
rect -888 -1917 -883 -1909
rect -881 -1917 -880 -1909
rect -876 -1917 -875 -1909
rect -873 -1917 -868 -1909
rect -864 -1917 -859 -1909
rect -857 -1917 -856 -1909
rect -844 -1917 -843 -1909
rect -841 -1917 -835 -1909
rect -833 -1917 -831 -1909
rect -827 -1917 -825 -1909
rect -823 -1917 -822 -1909
rect -750 -1917 -749 -1909
rect -747 -1917 -745 -1909
rect -741 -1917 -739 -1909
rect -737 -1917 -736 -1909
rect -724 -1917 -723 -1909
rect -721 -1917 -719 -1909
rect -715 -1917 -713 -1909
rect -711 -1917 -710 -1909
rect -698 -1917 -697 -1909
rect -695 -1917 -687 -1909
rect -685 -1917 -684 -1909
rect -680 -1917 -679 -1909
rect -677 -1917 -669 -1909
rect -667 -1917 -662 -1909
rect -658 -1917 -653 -1909
rect -651 -1917 -650 -1909
rect -646 -1917 -645 -1909
rect -643 -1917 -641 -1909
rect -637 -1917 -635 -1909
rect -633 -1917 -632 -1909
rect -620 -1917 -619 -1909
rect -617 -1917 -609 -1909
rect -607 -1917 -606 -1909
rect -602 -1917 -601 -1909
rect -599 -1917 -591 -1909
rect -589 -1917 -584 -1909
rect -580 -1917 -575 -1909
rect -573 -1917 -572 -1909
rect -568 -1917 -567 -1909
rect -565 -1917 -560 -1909
rect -556 -1917 -551 -1909
rect -549 -1917 -548 -1909
rect -536 -1917 -535 -1909
rect -533 -1917 -527 -1909
rect -525 -1917 -523 -1909
rect -519 -1917 -517 -1909
rect -515 -1917 -514 -1909
rect -442 -1917 -441 -1909
rect -439 -1917 -437 -1909
rect -433 -1917 -431 -1909
rect -429 -1917 -428 -1909
rect -416 -1917 -415 -1909
rect -413 -1917 -411 -1909
rect -407 -1917 -405 -1909
rect -403 -1917 -402 -1909
rect -390 -1917 -389 -1909
rect -387 -1917 -379 -1909
rect -377 -1917 -376 -1909
rect -372 -1917 -371 -1909
rect -369 -1917 -361 -1909
rect -359 -1917 -354 -1909
rect -350 -1917 -345 -1909
rect -343 -1917 -342 -1909
rect -338 -1917 -337 -1909
rect -335 -1917 -333 -1909
rect -329 -1917 -327 -1909
rect -325 -1917 -324 -1909
rect -312 -1917 -311 -1909
rect -309 -1917 -301 -1909
rect -299 -1917 -298 -1909
rect -294 -1917 -293 -1909
rect -291 -1917 -283 -1909
rect -281 -1917 -276 -1909
rect -272 -1917 -267 -1909
rect -265 -1917 -264 -1909
rect -260 -1917 -259 -1909
rect -257 -1917 -252 -1909
rect -248 -1917 -243 -1909
rect -241 -1917 -240 -1909
rect -228 -1917 -227 -1909
rect -225 -1917 -219 -1909
rect -217 -1917 -215 -1909
rect -211 -1917 -209 -1909
rect -207 -1917 -206 -1909
rect -134 -1917 -133 -1909
rect -131 -1917 -129 -1909
rect -125 -1917 -123 -1909
rect -121 -1917 -120 -1909
rect -108 -1917 -107 -1909
rect -105 -1917 -103 -1909
rect -99 -1917 -97 -1909
rect -95 -1917 -94 -1909
rect -82 -1917 -81 -1909
rect -79 -1917 -71 -1909
rect -69 -1917 -68 -1909
rect -64 -1917 -63 -1909
rect -61 -1917 -53 -1909
rect -51 -1917 -46 -1909
rect -42 -1917 -37 -1909
rect -35 -1917 -34 -1909
rect -30 -1917 -29 -1909
rect -27 -1917 -25 -1909
rect -21 -1917 -19 -1909
rect -17 -1917 -16 -1909
rect -4 -1917 -3 -1909
rect -1 -1917 7 -1909
rect 9 -1917 10 -1909
rect 14 -1917 15 -1909
rect 17 -1917 25 -1909
rect 27 -1917 32 -1909
rect 36 -1917 41 -1909
rect 43 -1917 44 -1909
rect 48 -1917 49 -1909
rect 51 -1917 56 -1909
rect 60 -1917 65 -1909
rect 67 -1917 68 -1909
rect 80 -1917 81 -1909
rect 83 -1917 89 -1909
rect 91 -1917 93 -1909
rect 97 -1917 99 -1909
rect 101 -1917 102 -1909
rect 174 -1917 175 -1909
rect 177 -1917 179 -1909
rect 183 -1917 185 -1909
rect 187 -1917 188 -1909
rect 200 -1917 201 -1909
rect 203 -1917 205 -1909
rect 209 -1917 211 -1909
rect 213 -1917 214 -1909
rect 226 -1917 227 -1909
rect 229 -1917 237 -1909
rect 239 -1917 240 -1909
rect 244 -1917 245 -1909
rect 247 -1917 255 -1909
rect 257 -1917 262 -1909
rect 266 -1917 271 -1909
rect 273 -1917 274 -1909
rect 278 -1917 279 -1909
rect 281 -1917 283 -1909
rect 287 -1917 289 -1909
rect 291 -1917 292 -1909
rect 304 -1917 305 -1909
rect 307 -1917 315 -1909
rect 317 -1917 318 -1909
rect 322 -1917 323 -1909
rect 325 -1917 333 -1909
rect 335 -1917 340 -1909
rect 344 -1917 349 -1909
rect 351 -1917 352 -1909
rect 356 -1917 357 -1909
rect 359 -1917 364 -1909
rect 368 -1917 373 -1909
rect 375 -1917 376 -1909
rect 388 -1917 389 -1909
rect 391 -1917 397 -1909
rect 399 -1917 401 -1909
rect 405 -1917 407 -1909
rect 409 -1917 410 -1909
rect 482 -1917 483 -1909
rect 485 -1917 487 -1909
rect 491 -1917 493 -1909
rect 495 -1917 496 -1909
rect 508 -1917 509 -1909
rect 511 -1917 513 -1909
rect 517 -1917 519 -1909
rect 521 -1917 522 -1909
rect 534 -1917 535 -1909
rect 537 -1917 545 -1909
rect 547 -1917 548 -1909
rect 552 -1917 553 -1909
rect 555 -1917 563 -1909
rect 565 -1917 570 -1909
rect 574 -1917 579 -1909
rect 581 -1917 582 -1909
rect 586 -1917 587 -1909
rect 589 -1917 591 -1909
rect 595 -1917 597 -1909
rect 599 -1917 600 -1909
rect 612 -1917 613 -1909
rect 615 -1917 623 -1909
rect 625 -1917 626 -1909
rect 630 -1917 631 -1909
rect 633 -1917 641 -1909
rect 643 -1917 648 -1909
rect 652 -1917 657 -1909
rect 659 -1917 660 -1909
rect 664 -1917 665 -1909
rect 667 -1917 672 -1909
rect 676 -1917 681 -1909
rect 683 -1917 684 -1909
rect 696 -1917 697 -1909
rect 699 -1917 705 -1909
rect 707 -1917 709 -1909
rect 713 -1917 715 -1909
rect 717 -1917 718 -1909
rect 790 -1917 791 -1909
rect 793 -1917 795 -1909
rect 799 -1917 801 -1909
rect 803 -1917 804 -1909
rect 816 -1917 817 -1909
rect 819 -1917 821 -1909
rect 825 -1917 827 -1909
rect 829 -1917 830 -1909
rect 842 -1917 843 -1909
rect 845 -1917 853 -1909
rect 855 -1917 856 -1909
rect 860 -1917 861 -1909
rect 863 -1917 871 -1909
rect 873 -1917 878 -1909
rect 882 -1917 887 -1909
rect 889 -1917 890 -1909
rect 894 -1917 895 -1909
rect 897 -1917 899 -1909
rect 903 -1917 905 -1909
rect 907 -1917 908 -1909
rect 920 -1917 921 -1909
rect 923 -1917 931 -1909
rect 933 -1917 934 -1909
rect 938 -1917 939 -1909
rect 941 -1917 949 -1909
rect 951 -1917 956 -1909
rect 960 -1917 965 -1909
rect 967 -1917 968 -1909
rect 972 -1917 973 -1909
rect 975 -1917 980 -1909
rect 984 -1917 989 -1909
rect 991 -1917 992 -1909
rect 1004 -1917 1005 -1909
rect 1007 -1917 1013 -1909
rect 1015 -1917 1017 -1909
rect 1021 -1917 1023 -1909
rect 1025 -1917 1026 -1909
rect -1305 -2080 -1304 -2072
rect -1302 -2080 -1301 -2072
rect -1297 -2080 -1296 -2072
rect -1294 -2080 -1292 -2072
rect -1288 -2080 -1286 -2072
rect -1284 -2080 -1283 -2072
rect -1058 -2080 -1057 -2072
rect -1055 -2080 -1054 -2072
rect -1050 -2080 -1049 -2072
rect -1047 -2080 -1045 -2072
rect -1041 -2080 -1039 -2072
rect -1037 -2080 -1036 -2072
rect -750 -2080 -749 -2072
rect -747 -2080 -746 -2072
rect -742 -2080 -741 -2072
rect -739 -2080 -737 -2072
rect -733 -2080 -731 -2072
rect -729 -2080 -728 -2072
rect -442 -2080 -441 -2072
rect -439 -2080 -438 -2072
rect -434 -2080 -433 -2072
rect -431 -2080 -429 -2072
rect -425 -2080 -423 -2072
rect -421 -2080 -420 -2072
rect -134 -2080 -133 -2072
rect -131 -2080 -130 -2072
rect -126 -2080 -125 -2072
rect -123 -2080 -121 -2072
rect -117 -2080 -115 -2072
rect -113 -2080 -112 -2072
rect 174 -2080 175 -2072
rect 177 -2080 178 -2072
rect 182 -2080 183 -2072
rect 185 -2080 187 -2072
rect 191 -2080 193 -2072
rect 195 -2080 196 -2072
rect 482 -2080 483 -2072
rect 485 -2080 486 -2072
rect 490 -2080 491 -2072
rect 493 -2080 495 -2072
rect 499 -2080 501 -2072
rect 503 -2080 504 -2072
rect 790 -2080 791 -2072
rect 793 -2080 794 -2072
rect 798 -2080 799 -2072
rect 801 -2080 803 -2072
rect 807 -2080 809 -2072
rect 811 -2080 812 -2072
rect -1230 -2239 -1229 -2231
rect -1227 -2239 -1225 -2231
rect -1221 -2239 -1219 -2231
rect -1217 -2239 -1216 -2231
rect -1204 -2239 -1203 -2231
rect -1201 -2239 -1193 -2231
rect -1191 -2239 -1190 -2231
rect -1186 -2239 -1185 -2231
rect -1183 -2239 -1175 -2231
rect -1173 -2239 -1168 -2231
rect -1164 -2239 -1159 -2231
rect -1157 -2239 -1156 -2231
rect -1152 -2239 -1151 -2231
rect -1149 -2239 -1147 -2231
rect -1143 -2239 -1141 -2231
rect -1139 -2239 -1138 -2231
rect -1058 -2239 -1057 -2231
rect -1055 -2239 -1053 -2231
rect -1049 -2239 -1047 -2231
rect -1045 -2239 -1044 -2231
rect -1032 -2239 -1031 -2231
rect -1029 -2239 -1027 -2231
rect -1023 -2239 -1021 -2231
rect -1019 -2239 -1018 -2231
rect -1006 -2239 -1005 -2231
rect -1003 -2239 -995 -2231
rect -993 -2239 -992 -2231
rect -988 -2239 -987 -2231
rect -985 -2239 -977 -2231
rect -975 -2239 -970 -2231
rect -966 -2239 -961 -2231
rect -959 -2239 -958 -2231
rect -954 -2239 -953 -2231
rect -951 -2239 -949 -2231
rect -945 -2239 -943 -2231
rect -941 -2239 -940 -2231
rect -928 -2239 -927 -2231
rect -925 -2239 -917 -2231
rect -915 -2239 -914 -2231
rect -910 -2239 -909 -2231
rect -907 -2239 -899 -2231
rect -897 -2239 -892 -2231
rect -888 -2239 -883 -2231
rect -881 -2239 -880 -2231
rect -876 -2239 -875 -2231
rect -873 -2239 -868 -2231
rect -864 -2239 -859 -2231
rect -857 -2239 -856 -2231
rect -844 -2239 -843 -2231
rect -841 -2239 -835 -2231
rect -833 -2239 -831 -2231
rect -827 -2239 -825 -2231
rect -823 -2239 -822 -2231
rect -750 -2239 -749 -2231
rect -747 -2239 -745 -2231
rect -741 -2239 -739 -2231
rect -737 -2239 -736 -2231
rect -724 -2239 -723 -2231
rect -721 -2239 -719 -2231
rect -715 -2239 -713 -2231
rect -711 -2239 -710 -2231
rect -698 -2239 -697 -2231
rect -695 -2239 -687 -2231
rect -685 -2239 -684 -2231
rect -680 -2239 -679 -2231
rect -677 -2239 -669 -2231
rect -667 -2239 -662 -2231
rect -658 -2239 -653 -2231
rect -651 -2239 -650 -2231
rect -646 -2239 -645 -2231
rect -643 -2239 -641 -2231
rect -637 -2239 -635 -2231
rect -633 -2239 -632 -2231
rect -620 -2239 -619 -2231
rect -617 -2239 -609 -2231
rect -607 -2239 -606 -2231
rect -602 -2239 -601 -2231
rect -599 -2239 -591 -2231
rect -589 -2239 -584 -2231
rect -580 -2239 -575 -2231
rect -573 -2239 -572 -2231
rect -568 -2239 -567 -2231
rect -565 -2239 -560 -2231
rect -556 -2239 -551 -2231
rect -549 -2239 -548 -2231
rect -536 -2239 -535 -2231
rect -533 -2239 -527 -2231
rect -525 -2239 -523 -2231
rect -519 -2239 -517 -2231
rect -515 -2239 -514 -2231
rect -442 -2239 -441 -2231
rect -439 -2239 -437 -2231
rect -433 -2239 -431 -2231
rect -429 -2239 -428 -2231
rect -416 -2239 -415 -2231
rect -413 -2239 -411 -2231
rect -407 -2239 -405 -2231
rect -403 -2239 -402 -2231
rect -390 -2239 -389 -2231
rect -387 -2239 -379 -2231
rect -377 -2239 -376 -2231
rect -372 -2239 -371 -2231
rect -369 -2239 -361 -2231
rect -359 -2239 -354 -2231
rect -350 -2239 -345 -2231
rect -343 -2239 -342 -2231
rect -338 -2239 -337 -2231
rect -335 -2239 -333 -2231
rect -329 -2239 -327 -2231
rect -325 -2239 -324 -2231
rect -312 -2239 -311 -2231
rect -309 -2239 -301 -2231
rect -299 -2239 -298 -2231
rect -294 -2239 -293 -2231
rect -291 -2239 -283 -2231
rect -281 -2239 -276 -2231
rect -272 -2239 -267 -2231
rect -265 -2239 -264 -2231
rect -260 -2239 -259 -2231
rect -257 -2239 -252 -2231
rect -248 -2239 -243 -2231
rect -241 -2239 -240 -2231
rect -228 -2239 -227 -2231
rect -225 -2239 -219 -2231
rect -217 -2239 -215 -2231
rect -211 -2239 -209 -2231
rect -207 -2239 -206 -2231
rect -134 -2239 -133 -2231
rect -131 -2239 -129 -2231
rect -125 -2239 -123 -2231
rect -121 -2239 -120 -2231
rect -108 -2239 -107 -2231
rect -105 -2239 -103 -2231
rect -99 -2239 -97 -2231
rect -95 -2239 -94 -2231
rect -82 -2239 -81 -2231
rect -79 -2239 -71 -2231
rect -69 -2239 -68 -2231
rect -64 -2239 -63 -2231
rect -61 -2239 -53 -2231
rect -51 -2239 -46 -2231
rect -42 -2239 -37 -2231
rect -35 -2239 -34 -2231
rect -30 -2239 -29 -2231
rect -27 -2239 -25 -2231
rect -21 -2239 -19 -2231
rect -17 -2239 -16 -2231
rect -4 -2239 -3 -2231
rect -1 -2239 7 -2231
rect 9 -2239 10 -2231
rect 14 -2239 15 -2231
rect 17 -2239 25 -2231
rect 27 -2239 32 -2231
rect 36 -2239 41 -2231
rect 43 -2239 44 -2231
rect 48 -2239 49 -2231
rect 51 -2239 56 -2231
rect 60 -2239 65 -2231
rect 67 -2239 68 -2231
rect 80 -2239 81 -2231
rect 83 -2239 89 -2231
rect 91 -2239 93 -2231
rect 97 -2239 99 -2231
rect 101 -2239 102 -2231
rect 174 -2239 175 -2231
rect 177 -2239 179 -2231
rect 183 -2239 185 -2231
rect 187 -2239 188 -2231
rect 200 -2239 201 -2231
rect 203 -2239 205 -2231
rect 209 -2239 211 -2231
rect 213 -2239 214 -2231
rect 226 -2239 227 -2231
rect 229 -2239 237 -2231
rect 239 -2239 240 -2231
rect 244 -2239 245 -2231
rect 247 -2239 255 -2231
rect 257 -2239 262 -2231
rect 266 -2239 271 -2231
rect 273 -2239 274 -2231
rect 278 -2239 279 -2231
rect 281 -2239 283 -2231
rect 287 -2239 289 -2231
rect 291 -2239 292 -2231
rect 304 -2239 305 -2231
rect 307 -2239 315 -2231
rect 317 -2239 318 -2231
rect 322 -2239 323 -2231
rect 325 -2239 333 -2231
rect 335 -2239 340 -2231
rect 344 -2239 349 -2231
rect 351 -2239 352 -2231
rect 356 -2239 357 -2231
rect 359 -2239 364 -2231
rect 368 -2239 373 -2231
rect 375 -2239 376 -2231
rect 388 -2239 389 -2231
rect 391 -2239 397 -2231
rect 399 -2239 401 -2231
rect 405 -2239 407 -2231
rect 409 -2239 410 -2231
rect 482 -2239 483 -2231
rect 485 -2239 487 -2231
rect 491 -2239 493 -2231
rect 495 -2239 496 -2231
rect 508 -2239 509 -2231
rect 511 -2239 513 -2231
rect 517 -2239 519 -2231
rect 521 -2239 522 -2231
rect 534 -2239 535 -2231
rect 537 -2239 545 -2231
rect 547 -2239 548 -2231
rect 552 -2239 553 -2231
rect 555 -2239 563 -2231
rect 565 -2239 570 -2231
rect 574 -2239 579 -2231
rect 581 -2239 582 -2231
rect 586 -2239 587 -2231
rect 589 -2239 591 -2231
rect 595 -2239 597 -2231
rect 599 -2239 600 -2231
rect 612 -2239 613 -2231
rect 615 -2239 623 -2231
rect 625 -2239 626 -2231
rect 630 -2239 631 -2231
rect 633 -2239 641 -2231
rect 643 -2239 648 -2231
rect 652 -2239 657 -2231
rect 659 -2239 660 -2231
rect 664 -2239 665 -2231
rect 667 -2239 672 -2231
rect 676 -2239 681 -2231
rect 683 -2239 684 -2231
rect 696 -2239 697 -2231
rect 699 -2239 705 -2231
rect 707 -2239 709 -2231
rect 713 -2239 715 -2231
rect 717 -2239 718 -2231
rect 790 -2239 791 -2231
rect 793 -2239 795 -2231
rect 799 -2239 801 -2231
rect 803 -2239 804 -2231
rect 816 -2239 817 -2231
rect 819 -2239 821 -2231
rect 825 -2239 827 -2231
rect 829 -2239 830 -2231
rect 842 -2239 843 -2231
rect 845 -2239 853 -2231
rect 855 -2239 856 -2231
rect 860 -2239 861 -2231
rect 863 -2239 871 -2231
rect 873 -2239 878 -2231
rect 882 -2239 887 -2231
rect 889 -2239 890 -2231
rect 894 -2239 895 -2231
rect 897 -2239 899 -2231
rect 903 -2239 905 -2231
rect 907 -2239 908 -2231
rect 920 -2239 921 -2231
rect 923 -2239 931 -2231
rect 933 -2239 934 -2231
rect 938 -2239 939 -2231
rect 941 -2239 949 -2231
rect 951 -2239 956 -2231
rect 960 -2239 965 -2231
rect 967 -2239 968 -2231
rect 972 -2239 973 -2231
rect 975 -2239 980 -2231
rect 984 -2239 989 -2231
rect 991 -2239 992 -2231
rect 1004 -2239 1005 -2231
rect 1007 -2239 1013 -2231
rect 1015 -2239 1017 -2231
rect 1021 -2239 1023 -2231
rect 1025 -2239 1026 -2231
rect -1305 -2371 -1304 -2363
rect -1302 -2371 -1301 -2363
rect -1297 -2371 -1296 -2363
rect -1294 -2371 -1292 -2363
rect -1288 -2371 -1286 -2363
rect -1284 -2371 -1283 -2363
rect -1058 -2371 -1057 -2363
rect -1055 -2371 -1054 -2363
rect -1050 -2371 -1049 -2363
rect -1047 -2371 -1045 -2363
rect -1041 -2371 -1039 -2363
rect -1037 -2371 -1036 -2363
rect -750 -2371 -749 -2363
rect -747 -2371 -746 -2363
rect -742 -2371 -741 -2363
rect -739 -2371 -737 -2363
rect -733 -2371 -731 -2363
rect -729 -2371 -728 -2363
rect -442 -2371 -441 -2363
rect -439 -2371 -438 -2363
rect -434 -2371 -433 -2363
rect -431 -2371 -429 -2363
rect -425 -2371 -423 -2363
rect -421 -2371 -420 -2363
rect -134 -2371 -133 -2363
rect -131 -2371 -130 -2363
rect -126 -2371 -125 -2363
rect -123 -2371 -121 -2363
rect -117 -2371 -115 -2363
rect -113 -2371 -112 -2363
rect 174 -2371 175 -2363
rect 177 -2371 178 -2363
rect 182 -2371 183 -2363
rect 185 -2371 187 -2363
rect 191 -2371 193 -2363
rect 195 -2371 196 -2363
rect 482 -2371 483 -2363
rect 485 -2371 486 -2363
rect 490 -2371 491 -2363
rect 493 -2371 495 -2363
rect 499 -2371 501 -2363
rect 503 -2371 504 -2363
rect 790 -2371 791 -2363
rect 793 -2371 794 -2363
rect 798 -2371 799 -2363
rect 801 -2371 803 -2363
rect 807 -2371 809 -2363
rect 811 -2371 812 -2363
rect -1230 -2530 -1229 -2522
rect -1227 -2530 -1225 -2522
rect -1221 -2530 -1219 -2522
rect -1217 -2530 -1216 -2522
rect -1204 -2530 -1203 -2522
rect -1201 -2530 -1193 -2522
rect -1191 -2530 -1190 -2522
rect -1186 -2530 -1185 -2522
rect -1183 -2530 -1175 -2522
rect -1173 -2530 -1168 -2522
rect -1164 -2530 -1159 -2522
rect -1157 -2530 -1156 -2522
rect -1152 -2530 -1151 -2522
rect -1149 -2530 -1147 -2522
rect -1143 -2530 -1141 -2522
rect -1139 -2530 -1138 -2522
rect -1058 -2530 -1057 -2522
rect -1055 -2530 -1053 -2522
rect -1049 -2530 -1047 -2522
rect -1045 -2530 -1044 -2522
rect -1032 -2530 -1031 -2522
rect -1029 -2530 -1027 -2522
rect -1023 -2530 -1021 -2522
rect -1019 -2530 -1018 -2522
rect -1006 -2530 -1005 -2522
rect -1003 -2530 -995 -2522
rect -993 -2530 -992 -2522
rect -988 -2530 -987 -2522
rect -985 -2530 -977 -2522
rect -975 -2530 -970 -2522
rect -966 -2530 -961 -2522
rect -959 -2530 -958 -2522
rect -954 -2530 -953 -2522
rect -951 -2530 -949 -2522
rect -945 -2530 -943 -2522
rect -941 -2530 -940 -2522
rect -928 -2530 -927 -2522
rect -925 -2530 -917 -2522
rect -915 -2530 -914 -2522
rect -910 -2530 -909 -2522
rect -907 -2530 -899 -2522
rect -897 -2530 -892 -2522
rect -888 -2530 -883 -2522
rect -881 -2530 -880 -2522
rect -876 -2530 -875 -2522
rect -873 -2530 -868 -2522
rect -864 -2530 -859 -2522
rect -857 -2530 -856 -2522
rect -844 -2530 -843 -2522
rect -841 -2530 -835 -2522
rect -833 -2530 -831 -2522
rect -827 -2530 -825 -2522
rect -823 -2530 -822 -2522
rect -750 -2530 -749 -2522
rect -747 -2530 -745 -2522
rect -741 -2530 -739 -2522
rect -737 -2530 -736 -2522
rect -724 -2530 -723 -2522
rect -721 -2530 -719 -2522
rect -715 -2530 -713 -2522
rect -711 -2530 -710 -2522
rect -698 -2530 -697 -2522
rect -695 -2530 -687 -2522
rect -685 -2530 -684 -2522
rect -680 -2530 -679 -2522
rect -677 -2530 -669 -2522
rect -667 -2530 -662 -2522
rect -658 -2530 -653 -2522
rect -651 -2530 -650 -2522
rect -646 -2530 -645 -2522
rect -643 -2530 -641 -2522
rect -637 -2530 -635 -2522
rect -633 -2530 -632 -2522
rect -620 -2530 -619 -2522
rect -617 -2530 -609 -2522
rect -607 -2530 -606 -2522
rect -602 -2530 -601 -2522
rect -599 -2530 -591 -2522
rect -589 -2530 -584 -2522
rect -580 -2530 -575 -2522
rect -573 -2530 -572 -2522
rect -568 -2530 -567 -2522
rect -565 -2530 -560 -2522
rect -556 -2530 -551 -2522
rect -549 -2530 -548 -2522
rect -536 -2530 -535 -2522
rect -533 -2530 -527 -2522
rect -525 -2530 -523 -2522
rect -519 -2530 -517 -2522
rect -515 -2530 -514 -2522
rect -442 -2530 -441 -2522
rect -439 -2530 -437 -2522
rect -433 -2530 -431 -2522
rect -429 -2530 -428 -2522
rect -416 -2530 -415 -2522
rect -413 -2530 -411 -2522
rect -407 -2530 -405 -2522
rect -403 -2530 -402 -2522
rect -390 -2530 -389 -2522
rect -387 -2530 -379 -2522
rect -377 -2530 -376 -2522
rect -372 -2530 -371 -2522
rect -369 -2530 -361 -2522
rect -359 -2530 -354 -2522
rect -350 -2530 -345 -2522
rect -343 -2530 -342 -2522
rect -338 -2530 -337 -2522
rect -335 -2530 -333 -2522
rect -329 -2530 -327 -2522
rect -325 -2530 -324 -2522
rect -312 -2530 -311 -2522
rect -309 -2530 -301 -2522
rect -299 -2530 -298 -2522
rect -294 -2530 -293 -2522
rect -291 -2530 -283 -2522
rect -281 -2530 -276 -2522
rect -272 -2530 -267 -2522
rect -265 -2530 -264 -2522
rect -260 -2530 -259 -2522
rect -257 -2530 -252 -2522
rect -248 -2530 -243 -2522
rect -241 -2530 -240 -2522
rect -228 -2530 -227 -2522
rect -225 -2530 -219 -2522
rect -217 -2530 -215 -2522
rect -211 -2530 -209 -2522
rect -207 -2530 -206 -2522
rect -134 -2530 -133 -2522
rect -131 -2530 -129 -2522
rect -125 -2530 -123 -2522
rect -121 -2530 -120 -2522
rect -108 -2530 -107 -2522
rect -105 -2530 -103 -2522
rect -99 -2530 -97 -2522
rect -95 -2530 -94 -2522
rect -82 -2530 -81 -2522
rect -79 -2530 -71 -2522
rect -69 -2530 -68 -2522
rect -64 -2530 -63 -2522
rect -61 -2530 -53 -2522
rect -51 -2530 -46 -2522
rect -42 -2530 -37 -2522
rect -35 -2530 -34 -2522
rect -30 -2530 -29 -2522
rect -27 -2530 -25 -2522
rect -21 -2530 -19 -2522
rect -17 -2530 -16 -2522
rect -4 -2530 -3 -2522
rect -1 -2530 7 -2522
rect 9 -2530 10 -2522
rect 14 -2530 15 -2522
rect 17 -2530 25 -2522
rect 27 -2530 32 -2522
rect 36 -2530 41 -2522
rect 43 -2530 44 -2522
rect 48 -2530 49 -2522
rect 51 -2530 56 -2522
rect 60 -2530 65 -2522
rect 67 -2530 68 -2522
rect 80 -2530 81 -2522
rect 83 -2530 89 -2522
rect 91 -2530 93 -2522
rect 97 -2530 99 -2522
rect 101 -2530 102 -2522
rect 174 -2530 175 -2522
rect 177 -2530 179 -2522
rect 183 -2530 185 -2522
rect 187 -2530 188 -2522
rect 200 -2530 201 -2522
rect 203 -2530 205 -2522
rect 209 -2530 211 -2522
rect 213 -2530 214 -2522
rect 226 -2530 227 -2522
rect 229 -2530 237 -2522
rect 239 -2530 240 -2522
rect 244 -2530 245 -2522
rect 247 -2530 255 -2522
rect 257 -2530 262 -2522
rect 266 -2530 271 -2522
rect 273 -2530 274 -2522
rect 278 -2530 279 -2522
rect 281 -2530 283 -2522
rect 287 -2530 289 -2522
rect 291 -2530 292 -2522
rect 304 -2530 305 -2522
rect 307 -2530 315 -2522
rect 317 -2530 318 -2522
rect 322 -2530 323 -2522
rect 325 -2530 333 -2522
rect 335 -2530 340 -2522
rect 344 -2530 349 -2522
rect 351 -2530 352 -2522
rect 356 -2530 357 -2522
rect 359 -2530 364 -2522
rect 368 -2530 373 -2522
rect 375 -2530 376 -2522
rect 388 -2530 389 -2522
rect 391 -2530 397 -2522
rect 399 -2530 401 -2522
rect 405 -2530 407 -2522
rect 409 -2530 410 -2522
rect 482 -2530 483 -2522
rect 485 -2530 487 -2522
rect 491 -2530 493 -2522
rect 495 -2530 496 -2522
rect 508 -2530 509 -2522
rect 511 -2530 513 -2522
rect 517 -2530 519 -2522
rect 521 -2530 522 -2522
rect 534 -2530 535 -2522
rect 537 -2530 545 -2522
rect 547 -2530 548 -2522
rect 552 -2530 553 -2522
rect 555 -2530 563 -2522
rect 565 -2530 570 -2522
rect 574 -2530 579 -2522
rect 581 -2530 582 -2522
rect 586 -2530 587 -2522
rect 589 -2530 591 -2522
rect 595 -2530 597 -2522
rect 599 -2530 600 -2522
rect 612 -2530 613 -2522
rect 615 -2530 623 -2522
rect 625 -2530 626 -2522
rect 630 -2530 631 -2522
rect 633 -2530 641 -2522
rect 643 -2530 648 -2522
rect 652 -2530 657 -2522
rect 659 -2530 660 -2522
rect 664 -2530 665 -2522
rect 667 -2530 672 -2522
rect 676 -2530 681 -2522
rect 683 -2530 684 -2522
rect 696 -2530 697 -2522
rect 699 -2530 705 -2522
rect 707 -2530 709 -2522
rect 713 -2530 715 -2522
rect 717 -2530 718 -2522
rect 790 -2530 791 -2522
rect 793 -2530 795 -2522
rect 799 -2530 801 -2522
rect 803 -2530 804 -2522
rect 816 -2530 817 -2522
rect 819 -2530 821 -2522
rect 825 -2530 827 -2522
rect 829 -2530 830 -2522
rect 842 -2530 843 -2522
rect 845 -2530 853 -2522
rect 855 -2530 856 -2522
rect 860 -2530 861 -2522
rect 863 -2530 871 -2522
rect 873 -2530 878 -2522
rect 882 -2530 887 -2522
rect 889 -2530 890 -2522
rect 894 -2530 895 -2522
rect 897 -2530 899 -2522
rect 903 -2530 905 -2522
rect 907 -2530 908 -2522
rect 920 -2530 921 -2522
rect 923 -2530 931 -2522
rect 933 -2530 934 -2522
rect 938 -2530 939 -2522
rect 941 -2530 949 -2522
rect 951 -2530 956 -2522
rect 960 -2530 965 -2522
rect 967 -2530 968 -2522
rect 972 -2530 973 -2522
rect 975 -2530 980 -2522
rect 984 -2530 989 -2522
rect 991 -2530 992 -2522
rect 1004 -2530 1005 -2522
rect 1007 -2530 1013 -2522
rect 1015 -2530 1017 -2522
rect 1021 -2530 1023 -2522
rect 1025 -2530 1026 -2522
rect -1305 -2662 -1304 -2654
rect -1302 -2662 -1301 -2654
rect -1297 -2662 -1296 -2654
rect -1294 -2662 -1292 -2654
rect -1288 -2662 -1286 -2654
rect -1284 -2662 -1283 -2654
rect -1058 -2662 -1057 -2654
rect -1055 -2662 -1054 -2654
rect -1050 -2662 -1049 -2654
rect -1047 -2662 -1045 -2654
rect -1041 -2662 -1039 -2654
rect -1037 -2662 -1036 -2654
rect -750 -2662 -749 -2654
rect -747 -2662 -746 -2654
rect -742 -2662 -741 -2654
rect -739 -2662 -737 -2654
rect -733 -2662 -731 -2654
rect -729 -2662 -728 -2654
rect -442 -2662 -441 -2654
rect -439 -2662 -438 -2654
rect -434 -2662 -433 -2654
rect -431 -2662 -429 -2654
rect -425 -2662 -423 -2654
rect -421 -2662 -420 -2654
rect -134 -2662 -133 -2654
rect -131 -2662 -130 -2654
rect -126 -2662 -125 -2654
rect -123 -2662 -121 -2654
rect -117 -2662 -115 -2654
rect -113 -2662 -112 -2654
rect 174 -2662 175 -2654
rect 177 -2662 178 -2654
rect 182 -2662 183 -2654
rect 185 -2662 187 -2654
rect 191 -2662 193 -2654
rect 195 -2662 196 -2654
rect 482 -2662 483 -2654
rect 485 -2662 486 -2654
rect 490 -2662 491 -2654
rect 493 -2662 495 -2654
rect 499 -2662 501 -2654
rect 503 -2662 504 -2654
rect 790 -2662 791 -2654
rect 793 -2662 794 -2654
rect 798 -2662 799 -2654
rect 801 -2662 803 -2654
rect 807 -2662 809 -2654
rect 811 -2662 812 -2654
rect -1230 -2821 -1229 -2813
rect -1227 -2821 -1225 -2813
rect -1221 -2821 -1219 -2813
rect -1217 -2821 -1216 -2813
rect -1204 -2821 -1203 -2813
rect -1201 -2821 -1193 -2813
rect -1191 -2821 -1190 -2813
rect -1186 -2821 -1185 -2813
rect -1183 -2821 -1175 -2813
rect -1173 -2821 -1168 -2813
rect -1164 -2821 -1159 -2813
rect -1157 -2821 -1156 -2813
rect -1152 -2821 -1151 -2813
rect -1149 -2821 -1147 -2813
rect -1143 -2821 -1141 -2813
rect -1139 -2821 -1138 -2813
rect -1058 -2821 -1057 -2813
rect -1055 -2821 -1053 -2813
rect -1049 -2821 -1047 -2813
rect -1045 -2821 -1044 -2813
rect -1032 -2821 -1031 -2813
rect -1029 -2821 -1027 -2813
rect -1023 -2821 -1021 -2813
rect -1019 -2821 -1018 -2813
rect -1006 -2821 -1005 -2813
rect -1003 -2821 -995 -2813
rect -993 -2821 -992 -2813
rect -988 -2821 -987 -2813
rect -985 -2821 -977 -2813
rect -975 -2821 -970 -2813
rect -966 -2821 -961 -2813
rect -959 -2821 -958 -2813
rect -954 -2821 -953 -2813
rect -951 -2821 -949 -2813
rect -945 -2821 -943 -2813
rect -941 -2821 -940 -2813
rect -928 -2821 -927 -2813
rect -925 -2821 -917 -2813
rect -915 -2821 -914 -2813
rect -910 -2821 -909 -2813
rect -907 -2821 -899 -2813
rect -897 -2821 -892 -2813
rect -888 -2821 -883 -2813
rect -881 -2821 -880 -2813
rect -876 -2821 -875 -2813
rect -873 -2821 -868 -2813
rect -864 -2821 -859 -2813
rect -857 -2821 -856 -2813
rect -844 -2821 -843 -2813
rect -841 -2821 -835 -2813
rect -833 -2821 -831 -2813
rect -827 -2821 -825 -2813
rect -823 -2821 -822 -2813
rect -750 -2821 -749 -2813
rect -747 -2821 -745 -2813
rect -741 -2821 -739 -2813
rect -737 -2821 -736 -2813
rect -724 -2821 -723 -2813
rect -721 -2821 -719 -2813
rect -715 -2821 -713 -2813
rect -711 -2821 -710 -2813
rect -698 -2821 -697 -2813
rect -695 -2821 -687 -2813
rect -685 -2821 -684 -2813
rect -680 -2821 -679 -2813
rect -677 -2821 -669 -2813
rect -667 -2821 -662 -2813
rect -658 -2821 -653 -2813
rect -651 -2821 -650 -2813
rect -646 -2821 -645 -2813
rect -643 -2821 -641 -2813
rect -637 -2821 -635 -2813
rect -633 -2821 -632 -2813
rect -620 -2821 -619 -2813
rect -617 -2821 -609 -2813
rect -607 -2821 -606 -2813
rect -602 -2821 -601 -2813
rect -599 -2821 -591 -2813
rect -589 -2821 -584 -2813
rect -580 -2821 -575 -2813
rect -573 -2821 -572 -2813
rect -568 -2821 -567 -2813
rect -565 -2821 -560 -2813
rect -556 -2821 -551 -2813
rect -549 -2821 -548 -2813
rect -536 -2821 -535 -2813
rect -533 -2821 -527 -2813
rect -525 -2821 -523 -2813
rect -519 -2821 -517 -2813
rect -515 -2821 -514 -2813
rect -442 -2821 -441 -2813
rect -439 -2821 -437 -2813
rect -433 -2821 -431 -2813
rect -429 -2821 -428 -2813
rect -416 -2821 -415 -2813
rect -413 -2821 -411 -2813
rect -407 -2821 -405 -2813
rect -403 -2821 -402 -2813
rect -390 -2821 -389 -2813
rect -387 -2821 -379 -2813
rect -377 -2821 -376 -2813
rect -372 -2821 -371 -2813
rect -369 -2821 -361 -2813
rect -359 -2821 -354 -2813
rect -350 -2821 -345 -2813
rect -343 -2821 -342 -2813
rect -338 -2821 -337 -2813
rect -335 -2821 -333 -2813
rect -329 -2821 -327 -2813
rect -325 -2821 -324 -2813
rect -312 -2821 -311 -2813
rect -309 -2821 -301 -2813
rect -299 -2821 -298 -2813
rect -294 -2821 -293 -2813
rect -291 -2821 -283 -2813
rect -281 -2821 -276 -2813
rect -272 -2821 -267 -2813
rect -265 -2821 -264 -2813
rect -260 -2821 -259 -2813
rect -257 -2821 -252 -2813
rect -248 -2821 -243 -2813
rect -241 -2821 -240 -2813
rect -228 -2821 -227 -2813
rect -225 -2821 -219 -2813
rect -217 -2821 -215 -2813
rect -211 -2821 -209 -2813
rect -207 -2821 -206 -2813
rect -134 -2821 -133 -2813
rect -131 -2821 -129 -2813
rect -125 -2821 -123 -2813
rect -121 -2821 -120 -2813
rect -108 -2821 -107 -2813
rect -105 -2821 -103 -2813
rect -99 -2821 -97 -2813
rect -95 -2821 -94 -2813
rect -82 -2821 -81 -2813
rect -79 -2821 -71 -2813
rect -69 -2821 -68 -2813
rect -64 -2821 -63 -2813
rect -61 -2821 -53 -2813
rect -51 -2821 -46 -2813
rect -42 -2821 -37 -2813
rect -35 -2821 -34 -2813
rect -30 -2821 -29 -2813
rect -27 -2821 -25 -2813
rect -21 -2821 -19 -2813
rect -17 -2821 -16 -2813
rect -4 -2821 -3 -2813
rect -1 -2821 7 -2813
rect 9 -2821 10 -2813
rect 14 -2821 15 -2813
rect 17 -2821 25 -2813
rect 27 -2821 32 -2813
rect 36 -2821 41 -2813
rect 43 -2821 44 -2813
rect 48 -2821 49 -2813
rect 51 -2821 56 -2813
rect 60 -2821 65 -2813
rect 67 -2821 68 -2813
rect 80 -2821 81 -2813
rect 83 -2821 89 -2813
rect 91 -2821 93 -2813
rect 97 -2821 99 -2813
rect 101 -2821 102 -2813
rect 174 -2821 175 -2813
rect 177 -2821 179 -2813
rect 183 -2821 185 -2813
rect 187 -2821 188 -2813
rect 200 -2821 201 -2813
rect 203 -2821 205 -2813
rect 209 -2821 211 -2813
rect 213 -2821 214 -2813
rect 226 -2821 227 -2813
rect 229 -2821 237 -2813
rect 239 -2821 240 -2813
rect 244 -2821 245 -2813
rect 247 -2821 255 -2813
rect 257 -2821 262 -2813
rect 266 -2821 271 -2813
rect 273 -2821 274 -2813
rect 278 -2821 279 -2813
rect 281 -2821 283 -2813
rect 287 -2821 289 -2813
rect 291 -2821 292 -2813
rect 304 -2821 305 -2813
rect 307 -2821 315 -2813
rect 317 -2821 318 -2813
rect 322 -2821 323 -2813
rect 325 -2821 333 -2813
rect 335 -2821 340 -2813
rect 344 -2821 349 -2813
rect 351 -2821 352 -2813
rect 356 -2821 357 -2813
rect 359 -2821 364 -2813
rect 368 -2821 373 -2813
rect 375 -2821 376 -2813
rect 388 -2821 389 -2813
rect 391 -2821 397 -2813
rect 399 -2821 401 -2813
rect 405 -2821 407 -2813
rect 409 -2821 410 -2813
rect 482 -2821 483 -2813
rect 485 -2821 487 -2813
rect 491 -2821 493 -2813
rect 495 -2821 496 -2813
rect 508 -2821 509 -2813
rect 511 -2821 513 -2813
rect 517 -2821 519 -2813
rect 521 -2821 522 -2813
rect 534 -2821 535 -2813
rect 537 -2821 545 -2813
rect 547 -2821 548 -2813
rect 552 -2821 553 -2813
rect 555 -2821 563 -2813
rect 565 -2821 570 -2813
rect 574 -2821 579 -2813
rect 581 -2821 582 -2813
rect 586 -2821 587 -2813
rect 589 -2821 591 -2813
rect 595 -2821 597 -2813
rect 599 -2821 600 -2813
rect 612 -2821 613 -2813
rect 615 -2821 623 -2813
rect 625 -2821 626 -2813
rect 630 -2821 631 -2813
rect 633 -2821 641 -2813
rect 643 -2821 648 -2813
rect 652 -2821 657 -2813
rect 659 -2821 660 -2813
rect 664 -2821 665 -2813
rect 667 -2821 672 -2813
rect 676 -2821 681 -2813
rect 683 -2821 684 -2813
rect 696 -2821 697 -2813
rect 699 -2821 705 -2813
rect 707 -2821 709 -2813
rect 713 -2821 715 -2813
rect 717 -2821 718 -2813
rect 790 -2821 791 -2813
rect 793 -2821 795 -2813
rect 799 -2821 801 -2813
rect 803 -2821 804 -2813
rect 816 -2821 817 -2813
rect 819 -2821 821 -2813
rect 825 -2821 827 -2813
rect 829 -2821 830 -2813
rect 842 -2821 843 -2813
rect 845 -2821 853 -2813
rect 855 -2821 856 -2813
rect 860 -2821 861 -2813
rect 863 -2821 871 -2813
rect 873 -2821 878 -2813
rect 882 -2821 887 -2813
rect 889 -2821 890 -2813
rect 894 -2821 895 -2813
rect 897 -2821 899 -2813
rect 903 -2821 905 -2813
rect 907 -2821 908 -2813
rect 920 -2821 921 -2813
rect 923 -2821 931 -2813
rect 933 -2821 934 -2813
rect 938 -2821 939 -2813
rect 941 -2821 949 -2813
rect 951 -2821 956 -2813
rect 960 -2821 965 -2813
rect 967 -2821 968 -2813
rect 972 -2821 973 -2813
rect 975 -2821 980 -2813
rect 984 -2821 989 -2813
rect 991 -2821 992 -2813
rect 1004 -2821 1005 -2813
rect 1007 -2821 1013 -2813
rect 1015 -2821 1017 -2813
rect 1021 -2821 1023 -2813
rect 1025 -2821 1026 -2813
rect -1305 -2953 -1304 -2945
rect -1302 -2953 -1301 -2945
rect -1297 -2953 -1296 -2945
rect -1294 -2953 -1292 -2945
rect -1288 -2953 -1286 -2945
rect -1284 -2953 -1283 -2945
rect -1058 -2953 -1057 -2945
rect -1055 -2953 -1054 -2945
rect -1050 -2953 -1049 -2945
rect -1047 -2953 -1045 -2945
rect -1041 -2953 -1039 -2945
rect -1037 -2953 -1036 -2945
rect -750 -2953 -749 -2945
rect -747 -2953 -746 -2945
rect -742 -2953 -741 -2945
rect -739 -2953 -737 -2945
rect -733 -2953 -731 -2945
rect -729 -2953 -728 -2945
rect -442 -2953 -441 -2945
rect -439 -2953 -438 -2945
rect -434 -2953 -433 -2945
rect -431 -2953 -429 -2945
rect -425 -2953 -423 -2945
rect -421 -2953 -420 -2945
rect -134 -2953 -133 -2945
rect -131 -2953 -130 -2945
rect -126 -2953 -125 -2945
rect -123 -2953 -121 -2945
rect -117 -2953 -115 -2945
rect -113 -2953 -112 -2945
rect 174 -2953 175 -2945
rect 177 -2953 178 -2945
rect 182 -2953 183 -2945
rect 185 -2953 187 -2945
rect 191 -2953 193 -2945
rect 195 -2953 196 -2945
rect 482 -2953 483 -2945
rect 485 -2953 486 -2945
rect 490 -2953 491 -2945
rect 493 -2953 495 -2945
rect 499 -2953 501 -2945
rect 503 -2953 504 -2945
rect 790 -2953 791 -2945
rect 793 -2953 794 -2945
rect 798 -2953 799 -2945
rect 801 -2953 803 -2945
rect 807 -2953 809 -2945
rect 811 -2953 812 -2945
rect -1230 -3112 -1229 -3104
rect -1227 -3112 -1225 -3104
rect -1221 -3112 -1219 -3104
rect -1217 -3112 -1216 -3104
rect -1204 -3112 -1203 -3104
rect -1201 -3112 -1193 -3104
rect -1191 -3112 -1190 -3104
rect -1186 -3112 -1185 -3104
rect -1183 -3112 -1175 -3104
rect -1173 -3112 -1168 -3104
rect -1164 -3112 -1159 -3104
rect -1157 -3112 -1156 -3104
rect -1152 -3112 -1151 -3104
rect -1149 -3112 -1147 -3104
rect -1143 -3112 -1141 -3104
rect -1139 -3112 -1138 -3104
rect -1058 -3112 -1057 -3104
rect -1055 -3112 -1053 -3104
rect -1049 -3112 -1047 -3104
rect -1045 -3112 -1044 -3104
rect -1032 -3112 -1031 -3104
rect -1029 -3112 -1027 -3104
rect -1023 -3112 -1021 -3104
rect -1019 -3112 -1018 -3104
rect -1006 -3112 -1005 -3104
rect -1003 -3112 -995 -3104
rect -993 -3112 -992 -3104
rect -988 -3112 -987 -3104
rect -985 -3112 -977 -3104
rect -975 -3112 -970 -3104
rect -966 -3112 -961 -3104
rect -959 -3112 -958 -3104
rect -954 -3112 -953 -3104
rect -951 -3112 -949 -3104
rect -945 -3112 -943 -3104
rect -941 -3112 -940 -3104
rect -928 -3112 -927 -3104
rect -925 -3112 -917 -3104
rect -915 -3112 -914 -3104
rect -910 -3112 -909 -3104
rect -907 -3112 -899 -3104
rect -897 -3112 -892 -3104
rect -888 -3112 -883 -3104
rect -881 -3112 -880 -3104
rect -876 -3112 -875 -3104
rect -873 -3112 -868 -3104
rect -864 -3112 -859 -3104
rect -857 -3112 -856 -3104
rect -844 -3112 -843 -3104
rect -841 -3112 -835 -3104
rect -833 -3112 -831 -3104
rect -827 -3112 -825 -3104
rect -823 -3112 -822 -3104
rect -750 -3112 -749 -3104
rect -747 -3112 -745 -3104
rect -741 -3112 -739 -3104
rect -737 -3112 -736 -3104
rect -724 -3112 -723 -3104
rect -721 -3112 -719 -3104
rect -715 -3112 -713 -3104
rect -711 -3112 -710 -3104
rect -698 -3112 -697 -3104
rect -695 -3112 -687 -3104
rect -685 -3112 -684 -3104
rect -680 -3112 -679 -3104
rect -677 -3112 -669 -3104
rect -667 -3112 -662 -3104
rect -658 -3112 -653 -3104
rect -651 -3112 -650 -3104
rect -646 -3112 -645 -3104
rect -643 -3112 -641 -3104
rect -637 -3112 -635 -3104
rect -633 -3112 -632 -3104
rect -620 -3112 -619 -3104
rect -617 -3112 -609 -3104
rect -607 -3112 -606 -3104
rect -602 -3112 -601 -3104
rect -599 -3112 -591 -3104
rect -589 -3112 -584 -3104
rect -580 -3112 -575 -3104
rect -573 -3112 -572 -3104
rect -568 -3112 -567 -3104
rect -565 -3112 -560 -3104
rect -556 -3112 -551 -3104
rect -549 -3112 -548 -3104
rect -536 -3112 -535 -3104
rect -533 -3112 -527 -3104
rect -525 -3112 -523 -3104
rect -519 -3112 -517 -3104
rect -515 -3112 -514 -3104
rect -442 -3112 -441 -3104
rect -439 -3112 -437 -3104
rect -433 -3112 -431 -3104
rect -429 -3112 -428 -3104
rect -416 -3112 -415 -3104
rect -413 -3112 -411 -3104
rect -407 -3112 -405 -3104
rect -403 -3112 -402 -3104
rect -390 -3112 -389 -3104
rect -387 -3112 -379 -3104
rect -377 -3112 -376 -3104
rect -372 -3112 -371 -3104
rect -369 -3112 -361 -3104
rect -359 -3112 -354 -3104
rect -350 -3112 -345 -3104
rect -343 -3112 -342 -3104
rect -338 -3112 -337 -3104
rect -335 -3112 -333 -3104
rect -329 -3112 -327 -3104
rect -325 -3112 -324 -3104
rect -312 -3112 -311 -3104
rect -309 -3112 -301 -3104
rect -299 -3112 -298 -3104
rect -294 -3112 -293 -3104
rect -291 -3112 -283 -3104
rect -281 -3112 -276 -3104
rect -272 -3112 -267 -3104
rect -265 -3112 -264 -3104
rect -260 -3112 -259 -3104
rect -257 -3112 -252 -3104
rect -248 -3112 -243 -3104
rect -241 -3112 -240 -3104
rect -228 -3112 -227 -3104
rect -225 -3112 -219 -3104
rect -217 -3112 -215 -3104
rect -211 -3112 -209 -3104
rect -207 -3112 -206 -3104
rect -134 -3112 -133 -3104
rect -131 -3112 -129 -3104
rect -125 -3112 -123 -3104
rect -121 -3112 -120 -3104
rect -108 -3112 -107 -3104
rect -105 -3112 -103 -3104
rect -99 -3112 -97 -3104
rect -95 -3112 -94 -3104
rect -82 -3112 -81 -3104
rect -79 -3112 -71 -3104
rect -69 -3112 -68 -3104
rect -64 -3112 -63 -3104
rect -61 -3112 -53 -3104
rect -51 -3112 -46 -3104
rect -42 -3112 -37 -3104
rect -35 -3112 -34 -3104
rect -30 -3112 -29 -3104
rect -27 -3112 -25 -3104
rect -21 -3112 -19 -3104
rect -17 -3112 -16 -3104
rect -4 -3112 -3 -3104
rect -1 -3112 7 -3104
rect 9 -3112 10 -3104
rect 14 -3112 15 -3104
rect 17 -3112 25 -3104
rect 27 -3112 32 -3104
rect 36 -3112 41 -3104
rect 43 -3112 44 -3104
rect 48 -3112 49 -3104
rect 51 -3112 56 -3104
rect 60 -3112 65 -3104
rect 67 -3112 68 -3104
rect 80 -3112 81 -3104
rect 83 -3112 89 -3104
rect 91 -3112 93 -3104
rect 97 -3112 99 -3104
rect 101 -3112 102 -3104
rect 174 -3112 175 -3104
rect 177 -3112 179 -3104
rect 183 -3112 185 -3104
rect 187 -3112 188 -3104
rect 200 -3112 201 -3104
rect 203 -3112 205 -3104
rect 209 -3112 211 -3104
rect 213 -3112 214 -3104
rect 226 -3112 227 -3104
rect 229 -3112 237 -3104
rect 239 -3112 240 -3104
rect 244 -3112 245 -3104
rect 247 -3112 255 -3104
rect 257 -3112 262 -3104
rect 266 -3112 271 -3104
rect 273 -3112 274 -3104
rect 278 -3112 279 -3104
rect 281 -3112 283 -3104
rect 287 -3112 289 -3104
rect 291 -3112 292 -3104
rect 304 -3112 305 -3104
rect 307 -3112 315 -3104
rect 317 -3112 318 -3104
rect 322 -3112 323 -3104
rect 325 -3112 333 -3104
rect 335 -3112 340 -3104
rect 344 -3112 349 -3104
rect 351 -3112 352 -3104
rect 356 -3112 357 -3104
rect 359 -3112 364 -3104
rect 368 -3112 373 -3104
rect 375 -3112 376 -3104
rect 388 -3112 389 -3104
rect 391 -3112 397 -3104
rect 399 -3112 401 -3104
rect 405 -3112 407 -3104
rect 409 -3112 410 -3104
rect 482 -3112 483 -3104
rect 485 -3112 487 -3104
rect 491 -3112 493 -3104
rect 495 -3112 496 -3104
rect 508 -3112 509 -3104
rect 511 -3112 513 -3104
rect 517 -3112 519 -3104
rect 521 -3112 522 -3104
rect 534 -3112 535 -3104
rect 537 -3112 545 -3104
rect 547 -3112 548 -3104
rect 552 -3112 553 -3104
rect 555 -3112 563 -3104
rect 565 -3112 570 -3104
rect 574 -3112 579 -3104
rect 581 -3112 582 -3104
rect 586 -3112 587 -3104
rect 589 -3112 591 -3104
rect 595 -3112 597 -3104
rect 599 -3112 600 -3104
rect 612 -3112 613 -3104
rect 615 -3112 623 -3104
rect 625 -3112 626 -3104
rect 630 -3112 631 -3104
rect 633 -3112 641 -3104
rect 643 -3112 648 -3104
rect 652 -3112 657 -3104
rect 659 -3112 660 -3104
rect 664 -3112 665 -3104
rect 667 -3112 672 -3104
rect 676 -3112 681 -3104
rect 683 -3112 684 -3104
rect 696 -3112 697 -3104
rect 699 -3112 705 -3104
rect 707 -3112 709 -3104
rect 713 -3112 715 -3104
rect 717 -3112 718 -3104
rect 790 -3112 791 -3104
rect 793 -3112 795 -3104
rect 799 -3112 801 -3104
rect 803 -3112 804 -3104
rect 816 -3112 817 -3104
rect 819 -3112 821 -3104
rect 825 -3112 827 -3104
rect 829 -3112 830 -3104
rect 842 -3112 843 -3104
rect 845 -3112 853 -3104
rect 855 -3112 856 -3104
rect 860 -3112 861 -3104
rect 863 -3112 871 -3104
rect 873 -3112 878 -3104
rect 882 -3112 887 -3104
rect 889 -3112 890 -3104
rect 894 -3112 895 -3104
rect 897 -3112 899 -3104
rect 903 -3112 905 -3104
rect 907 -3112 908 -3104
rect 920 -3112 921 -3104
rect 923 -3112 931 -3104
rect 933 -3112 934 -3104
rect 938 -3112 939 -3104
rect 941 -3112 949 -3104
rect 951 -3112 956 -3104
rect 960 -3112 965 -3104
rect 967 -3112 968 -3104
rect 972 -3112 973 -3104
rect 975 -3112 980 -3104
rect 984 -3112 989 -3104
rect 991 -3112 992 -3104
rect 1004 -3112 1005 -3104
rect 1007 -3112 1013 -3104
rect 1015 -3112 1017 -3104
rect 1021 -3112 1023 -3104
rect 1025 -3112 1026 -3104
<< metal1 >>
rect -1319 -1012 -1315 -948
rect -1307 -988 -1303 -984
rect -1290 -988 -1286 -984
rect -1299 -999 -1295 -996
rect -1299 -1003 -1284 -999
rect -1319 -1016 -1306 -1012
rect -1319 -1162 -1315 -1016
rect -1288 -1042 -1284 -1003
rect -1288 -1057 -1284 -1046
rect -1307 -1061 -1284 -1057
rect -1307 -1064 -1303 -1061
rect -1281 -1064 -1277 -996
rect -1076 -1012 -1072 -948
rect -1063 -988 -1059 -984
rect -1046 -988 -1042 -984
rect -1055 -999 -1051 -996
rect -1055 -1003 -1040 -999
rect -1076 -1016 -1062 -1012
rect -1290 -1072 -1286 -1068
rect -1309 -1138 -1305 -1134
rect -1292 -1138 -1288 -1134
rect -1301 -1149 -1297 -1146
rect -1301 -1153 -1286 -1149
rect -1319 -1166 -1308 -1162
rect -1319 -1483 -1315 -1166
rect -1290 -1192 -1286 -1153
rect -1290 -1207 -1286 -1196
rect -1309 -1211 -1286 -1207
rect -1309 -1214 -1305 -1211
rect -1283 -1214 -1279 -1146
rect -1292 -1222 -1288 -1218
rect -1283 -1357 -1279 -1218
rect -1251 -1350 -1247 -1040
rect -1221 -1302 -1217 -1298
rect -1204 -1302 -1200 -1298
rect -1164 -1302 -1160 -1298
rect -1143 -1302 -1139 -1298
rect -1230 -1343 -1226 -1310
rect -1230 -1378 -1226 -1347
rect -1212 -1337 -1208 -1310
rect -1212 -1341 -1203 -1337
rect -1212 -1378 -1208 -1341
rect -1186 -1364 -1182 -1310
rect -1186 -1371 -1182 -1368
rect -1152 -1371 -1148 -1310
rect -1134 -1342 -1130 -1310
rect -1204 -1378 -1200 -1375
rect -1195 -1375 -1182 -1371
rect -1195 -1378 -1191 -1375
rect -1168 -1378 -1164 -1375
rect -1160 -1375 -1141 -1371
rect -1160 -1378 -1156 -1375
rect -1134 -1378 -1130 -1346
rect -1103 -1349 -1099 -1187
rect -1091 -1334 -1087 -1032
rect -1076 -1162 -1072 -1016
rect -1044 -1044 -1040 -1003
rect -1044 -1057 -1040 -1048
rect -1063 -1061 -1040 -1057
rect -1037 -1036 -1033 -996
rect -768 -1012 -764 -949
rect -754 -988 -750 -984
rect -737 -988 -733 -984
rect -746 -999 -742 -996
rect -746 -1003 -731 -999
rect -768 -1016 -753 -1012
rect -1063 -1064 -1059 -1061
rect -1037 -1064 -1033 -1040
rect -1046 -1072 -1042 -1068
rect -1062 -1138 -1058 -1134
rect -1045 -1138 -1041 -1134
rect -1054 -1149 -1050 -1146
rect -1054 -1153 -1039 -1149
rect -1076 -1166 -1061 -1162
rect -1221 -1386 -1217 -1382
rect -1177 -1386 -1173 -1382
rect -1143 -1386 -1139 -1382
rect -1309 -1459 -1305 -1455
rect -1292 -1459 -1288 -1455
rect -1301 -1470 -1297 -1467
rect -1301 -1474 -1286 -1470
rect -1319 -1487 -1308 -1483
rect -1319 -1774 -1315 -1487
rect -1290 -1513 -1286 -1474
rect -1290 -1528 -1286 -1517
rect -1309 -1532 -1286 -1528
rect -1309 -1535 -1305 -1532
rect -1283 -1535 -1279 -1467
rect -1292 -1543 -1288 -1539
rect -1283 -1673 -1279 -1539
rect -1257 -1666 -1253 -1397
rect -1225 -1618 -1221 -1614
rect -1208 -1618 -1204 -1614
rect -1168 -1618 -1164 -1614
rect -1147 -1618 -1143 -1614
rect -1234 -1659 -1230 -1626
rect -1234 -1694 -1230 -1663
rect -1216 -1653 -1212 -1626
rect -1216 -1657 -1207 -1653
rect -1216 -1694 -1212 -1657
rect -1190 -1680 -1186 -1626
rect -1190 -1687 -1186 -1684
rect -1156 -1687 -1152 -1626
rect -1138 -1658 -1134 -1626
rect -1113 -1650 -1109 -1404
rect -1076 -1483 -1072 -1166
rect -1043 -1192 -1039 -1153
rect -1043 -1207 -1039 -1196
rect -1062 -1211 -1039 -1207
rect -1036 -1183 -1032 -1146
rect -1062 -1214 -1058 -1211
rect -1036 -1214 -1032 -1187
rect -1045 -1222 -1041 -1218
rect -1053 -1302 -1049 -1298
rect -1027 -1302 -1023 -1298
rect -1010 -1302 -1006 -1298
rect -970 -1302 -966 -1298
rect -949 -1302 -945 -1298
rect -932 -1302 -928 -1298
rect -892 -1302 -888 -1298
rect -868 -1302 -864 -1298
rect -831 -1302 -827 -1298
rect -1062 -1327 -1058 -1310
rect -1062 -1378 -1058 -1331
rect -1044 -1320 -1040 -1310
rect -1044 -1378 -1040 -1324
rect -1036 -1349 -1032 -1310
rect -1018 -1342 -1014 -1310
rect -1036 -1378 -1032 -1353
rect -1018 -1378 -1014 -1346
rect -992 -1334 -988 -1310
rect -992 -1371 -988 -1338
rect -958 -1371 -954 -1310
rect -940 -1327 -936 -1310
rect -1010 -1378 -1006 -1375
rect -1002 -1375 -988 -1371
rect -1002 -1378 -998 -1375
rect -974 -1378 -970 -1375
rect -966 -1375 -947 -1371
rect -966 -1378 -962 -1375
rect -940 -1378 -936 -1331
rect -914 -1342 -910 -1310
rect -914 -1371 -910 -1346
rect -880 -1364 -876 -1310
rect -880 -1368 -863 -1364
rect -932 -1378 -928 -1375
rect -923 -1375 -910 -1371
rect -923 -1378 -919 -1375
rect -896 -1378 -892 -1375
rect -872 -1378 -868 -1368
rect -856 -1371 -852 -1310
rect -848 -1364 -844 -1310
rect -822 -1334 -818 -1310
rect -848 -1368 -829 -1364
rect -864 -1375 -847 -1371
rect -864 -1378 -860 -1375
rect -840 -1378 -836 -1368
rect -822 -1378 -818 -1338
rect -1053 -1386 -1049 -1382
rect -1027 -1386 -1023 -1382
rect -984 -1386 -980 -1382
rect -949 -1386 -945 -1382
rect -905 -1386 -901 -1382
rect -888 -1386 -884 -1382
rect -852 -1386 -848 -1382
rect -831 -1386 -827 -1382
rect -815 -1393 -811 -1346
rect -795 -1349 -791 -1187
rect -782 -1334 -778 -1040
rect -768 -1162 -764 -1016
rect -735 -1044 -731 -1003
rect -735 -1057 -731 -1048
rect -754 -1061 -731 -1057
rect -728 -1028 -724 -996
rect -460 -1012 -456 -948
rect -446 -988 -442 -984
rect -429 -988 -425 -984
rect -438 -999 -434 -996
rect -438 -1003 -423 -999
rect -460 -1016 -445 -1012
rect -754 -1064 -750 -1061
rect -728 -1064 -724 -1032
rect -737 -1072 -733 -1068
rect -754 -1138 -750 -1134
rect -737 -1138 -733 -1134
rect -746 -1149 -742 -1146
rect -746 -1153 -731 -1149
rect -768 -1166 -753 -1162
rect -1062 -1459 -1058 -1455
rect -1045 -1459 -1041 -1455
rect -1054 -1470 -1050 -1467
rect -1054 -1474 -1039 -1470
rect -1076 -1487 -1061 -1483
rect -1208 -1694 -1204 -1691
rect -1199 -1691 -1186 -1687
rect -1199 -1694 -1195 -1691
rect -1172 -1694 -1168 -1691
rect -1164 -1691 -1145 -1687
rect -1164 -1694 -1160 -1691
rect -1138 -1694 -1134 -1662
rect -1095 -1665 -1091 -1508
rect -1225 -1702 -1221 -1698
rect -1181 -1702 -1177 -1698
rect -1147 -1702 -1143 -1698
rect -1309 -1750 -1305 -1746
rect -1292 -1750 -1288 -1746
rect -1301 -1761 -1297 -1758
rect -1301 -1765 -1286 -1761
rect -1319 -1778 -1308 -1774
rect -1319 -2096 -1315 -1778
rect -1290 -1804 -1286 -1765
rect -1290 -1819 -1286 -1808
rect -1309 -1823 -1286 -1819
rect -1309 -1826 -1305 -1823
rect -1283 -1826 -1279 -1758
rect -1292 -1834 -1288 -1830
rect -1283 -1964 -1279 -1830
rect -1257 -1957 -1253 -1713
rect -1225 -1909 -1221 -1905
rect -1208 -1909 -1204 -1905
rect -1168 -1909 -1164 -1905
rect -1147 -1909 -1143 -1905
rect -1234 -1950 -1230 -1917
rect -1234 -1985 -1230 -1954
rect -1216 -1944 -1212 -1917
rect -1216 -1948 -1207 -1944
rect -1216 -1985 -1212 -1948
rect -1190 -1971 -1186 -1917
rect -1190 -1978 -1186 -1975
rect -1156 -1978 -1152 -1917
rect -1138 -1949 -1134 -1917
rect -1106 -1941 -1102 -1799
rect -1208 -1985 -1204 -1982
rect -1199 -1982 -1186 -1978
rect -1199 -1985 -1195 -1982
rect -1172 -1985 -1168 -1982
rect -1164 -1982 -1145 -1978
rect -1164 -1985 -1160 -1982
rect -1138 -1985 -1134 -1953
rect -1090 -1956 -1086 -1720
rect -1076 -1774 -1072 -1487
rect -1043 -1513 -1039 -1474
rect -1043 -1528 -1039 -1517
rect -1062 -1532 -1039 -1528
rect -1036 -1504 -1032 -1467
rect -1062 -1535 -1058 -1532
rect -1036 -1535 -1032 -1508
rect -1045 -1543 -1041 -1539
rect -1053 -1618 -1049 -1614
rect -1027 -1618 -1023 -1614
rect -1010 -1618 -1006 -1614
rect -970 -1618 -966 -1614
rect -949 -1618 -945 -1614
rect -932 -1618 -928 -1614
rect -892 -1618 -888 -1614
rect -868 -1618 -864 -1614
rect -831 -1618 -827 -1614
rect -1062 -1643 -1058 -1626
rect -1062 -1694 -1058 -1647
rect -1044 -1636 -1040 -1626
rect -1044 -1694 -1040 -1640
rect -1036 -1665 -1032 -1626
rect -1018 -1658 -1014 -1626
rect -1036 -1694 -1032 -1669
rect -1018 -1694 -1014 -1662
rect -992 -1650 -988 -1626
rect -992 -1687 -988 -1654
rect -958 -1687 -954 -1626
rect -940 -1643 -936 -1626
rect -1010 -1694 -1006 -1691
rect -1002 -1691 -988 -1687
rect -1002 -1694 -998 -1691
rect -974 -1694 -970 -1691
rect -966 -1691 -947 -1687
rect -966 -1694 -962 -1691
rect -940 -1694 -936 -1647
rect -914 -1658 -910 -1626
rect -914 -1687 -910 -1662
rect -880 -1680 -876 -1626
rect -880 -1684 -863 -1680
rect -932 -1694 -928 -1691
rect -923 -1691 -910 -1687
rect -923 -1694 -919 -1691
rect -896 -1694 -892 -1691
rect -872 -1694 -868 -1684
rect -856 -1687 -852 -1626
rect -848 -1680 -844 -1626
rect -822 -1650 -818 -1626
rect -848 -1684 -829 -1680
rect -864 -1691 -847 -1687
rect -864 -1694 -860 -1691
rect -840 -1694 -836 -1684
rect -822 -1694 -818 -1654
rect -1053 -1702 -1049 -1698
rect -1027 -1702 -1023 -1698
rect -984 -1702 -980 -1698
rect -949 -1702 -945 -1698
rect -905 -1702 -901 -1698
rect -888 -1702 -884 -1698
rect -852 -1702 -848 -1698
rect -831 -1702 -827 -1698
rect -814 -1709 -810 -1662
rect -795 -1665 -791 -1508
rect -782 -1650 -778 -1411
rect -768 -1483 -764 -1166
rect -735 -1192 -731 -1153
rect -735 -1207 -731 -1196
rect -754 -1211 -731 -1207
rect -728 -1183 -724 -1146
rect -754 -1214 -750 -1211
rect -728 -1214 -724 -1187
rect -737 -1222 -733 -1218
rect -745 -1302 -741 -1298
rect -719 -1302 -715 -1298
rect -702 -1302 -698 -1298
rect -662 -1302 -658 -1298
rect -641 -1302 -637 -1298
rect -624 -1302 -620 -1298
rect -584 -1302 -580 -1298
rect -560 -1302 -556 -1298
rect -523 -1302 -519 -1298
rect -754 -1327 -750 -1310
rect -754 -1378 -750 -1331
rect -736 -1320 -732 -1310
rect -736 -1378 -732 -1324
rect -728 -1349 -724 -1310
rect -710 -1342 -706 -1310
rect -728 -1378 -724 -1353
rect -710 -1378 -706 -1346
rect -684 -1334 -680 -1310
rect -684 -1371 -680 -1338
rect -650 -1371 -646 -1310
rect -632 -1327 -628 -1310
rect -702 -1378 -698 -1375
rect -694 -1375 -680 -1371
rect -694 -1378 -690 -1375
rect -666 -1378 -662 -1375
rect -658 -1375 -639 -1371
rect -658 -1378 -654 -1375
rect -632 -1378 -628 -1331
rect -606 -1342 -602 -1310
rect -606 -1371 -602 -1346
rect -572 -1364 -568 -1310
rect -572 -1368 -555 -1364
rect -624 -1378 -620 -1375
rect -615 -1375 -602 -1371
rect -615 -1378 -611 -1375
rect -588 -1378 -584 -1375
rect -564 -1378 -560 -1368
rect -548 -1371 -544 -1310
rect -540 -1364 -536 -1310
rect -514 -1334 -510 -1310
rect -540 -1368 -521 -1364
rect -556 -1375 -539 -1371
rect -556 -1378 -552 -1375
rect -532 -1378 -528 -1368
rect -514 -1378 -510 -1338
rect -745 -1386 -741 -1382
rect -719 -1386 -715 -1382
rect -676 -1386 -672 -1382
rect -641 -1386 -637 -1382
rect -597 -1386 -593 -1382
rect -580 -1386 -576 -1382
rect -544 -1386 -540 -1382
rect -523 -1386 -519 -1382
rect -505 -1400 -501 -1346
rect -494 -1349 -490 -1187
rect -471 -1334 -467 -1032
rect -460 -1162 -456 -1016
rect -427 -1044 -423 -1003
rect -427 -1057 -423 -1048
rect -446 -1061 -423 -1057
rect -420 -1036 -416 -996
rect -152 -1012 -148 -948
rect -139 -988 -135 -984
rect -122 -988 -118 -984
rect -131 -999 -127 -996
rect -131 -1003 -116 -999
rect -152 -1016 -138 -1012
rect -446 -1064 -442 -1061
rect -420 -1064 -416 -1040
rect -429 -1072 -425 -1068
rect -446 -1138 -442 -1134
rect -429 -1138 -425 -1134
rect -438 -1149 -434 -1146
rect -438 -1153 -423 -1149
rect -460 -1166 -445 -1162
rect -754 -1459 -750 -1455
rect -737 -1459 -733 -1455
rect -746 -1470 -742 -1467
rect -746 -1474 -731 -1470
rect -768 -1487 -753 -1483
rect -1062 -1750 -1058 -1746
rect -1045 -1750 -1041 -1746
rect -1054 -1761 -1050 -1758
rect -1054 -1765 -1039 -1761
rect -1076 -1778 -1061 -1774
rect -1225 -1993 -1221 -1989
rect -1181 -1993 -1177 -1989
rect -1147 -1993 -1143 -1989
rect -1309 -2072 -1305 -2068
rect -1292 -2072 -1288 -2068
rect -1301 -2083 -1297 -2080
rect -1301 -2087 -1286 -2083
rect -1319 -2100 -1308 -2096
rect -1319 -2387 -1315 -2100
rect -1290 -2126 -1286 -2087
rect -1290 -2141 -1286 -2130
rect -1309 -2145 -1286 -2141
rect -1309 -2148 -1305 -2145
rect -1283 -2148 -1279 -2080
rect -1292 -2156 -1288 -2152
rect -1283 -2286 -1279 -2152
rect -1257 -2279 -1253 -2004
rect -1225 -2231 -1221 -2227
rect -1208 -2231 -1204 -2227
rect -1168 -2231 -1164 -2227
rect -1147 -2231 -1143 -2227
rect -1234 -2272 -1230 -2239
rect -1234 -2307 -1230 -2276
rect -1216 -2266 -1212 -2239
rect -1216 -2270 -1207 -2266
rect -1216 -2307 -1212 -2270
rect -1190 -2293 -1186 -2239
rect -1190 -2300 -1186 -2297
rect -1156 -2300 -1152 -2239
rect -1138 -2271 -1134 -2239
rect -1106 -2263 -1102 -2121
rect -1208 -2307 -1204 -2304
rect -1199 -2304 -1186 -2300
rect -1199 -2307 -1195 -2304
rect -1172 -2307 -1168 -2304
rect -1164 -2304 -1145 -2300
rect -1164 -2307 -1160 -2304
rect -1138 -2307 -1134 -2275
rect -1090 -2278 -1086 -2011
rect -1076 -2096 -1072 -1778
rect -1043 -1804 -1039 -1765
rect -1043 -1819 -1039 -1808
rect -1062 -1823 -1039 -1819
rect -1036 -1795 -1032 -1758
rect -1062 -1826 -1058 -1823
rect -1036 -1826 -1032 -1799
rect -1045 -1834 -1041 -1830
rect -1053 -1909 -1049 -1905
rect -1027 -1909 -1023 -1905
rect -1010 -1909 -1006 -1905
rect -970 -1909 -966 -1905
rect -949 -1909 -945 -1905
rect -932 -1909 -928 -1905
rect -892 -1909 -888 -1905
rect -868 -1909 -864 -1905
rect -831 -1909 -827 -1905
rect -1062 -1934 -1058 -1917
rect -1062 -1985 -1058 -1938
rect -1044 -1927 -1040 -1917
rect -1044 -1985 -1040 -1931
rect -1036 -1956 -1032 -1917
rect -1018 -1949 -1014 -1917
rect -1036 -1985 -1032 -1960
rect -1018 -1985 -1014 -1953
rect -992 -1941 -988 -1917
rect -992 -1978 -988 -1945
rect -958 -1978 -954 -1917
rect -940 -1934 -936 -1917
rect -1010 -1985 -1006 -1982
rect -1002 -1982 -988 -1978
rect -1002 -1985 -998 -1982
rect -974 -1985 -970 -1982
rect -966 -1982 -947 -1978
rect -966 -1985 -962 -1982
rect -940 -1985 -936 -1938
rect -914 -1949 -910 -1917
rect -914 -1978 -910 -1953
rect -880 -1971 -876 -1917
rect -880 -1975 -863 -1971
rect -932 -1985 -928 -1982
rect -923 -1982 -910 -1978
rect -923 -1985 -919 -1982
rect -896 -1985 -892 -1982
rect -872 -1985 -868 -1975
rect -856 -1978 -852 -1917
rect -848 -1971 -844 -1917
rect -822 -1941 -818 -1917
rect -848 -1975 -829 -1971
rect -864 -1982 -847 -1978
rect -864 -1985 -860 -1982
rect -840 -1985 -836 -1975
rect -822 -1985 -818 -1945
rect -1053 -1993 -1049 -1989
rect -1027 -1993 -1023 -1989
rect -984 -1993 -980 -1989
rect -949 -1993 -945 -1989
rect -905 -1993 -901 -1989
rect -888 -1993 -884 -1989
rect -852 -1993 -848 -1989
rect -831 -1993 -827 -1989
rect -815 -2000 -811 -1953
rect -793 -1956 -789 -1799
rect -780 -1941 -776 -1713
rect -768 -1774 -764 -1487
rect -735 -1513 -731 -1474
rect -735 -1528 -731 -1517
rect -754 -1532 -731 -1528
rect -728 -1504 -724 -1467
rect -754 -1535 -750 -1532
rect -728 -1535 -724 -1508
rect -737 -1543 -733 -1539
rect -745 -1618 -741 -1614
rect -719 -1618 -715 -1614
rect -702 -1618 -698 -1614
rect -662 -1618 -658 -1614
rect -641 -1618 -637 -1614
rect -624 -1618 -620 -1614
rect -584 -1618 -580 -1614
rect -560 -1618 -556 -1614
rect -523 -1618 -519 -1614
rect -754 -1643 -750 -1626
rect -754 -1694 -750 -1647
rect -736 -1636 -732 -1626
rect -736 -1694 -732 -1640
rect -728 -1665 -724 -1626
rect -710 -1658 -706 -1626
rect -728 -1694 -724 -1669
rect -710 -1694 -706 -1662
rect -684 -1650 -680 -1626
rect -684 -1687 -680 -1654
rect -650 -1687 -646 -1626
rect -632 -1643 -628 -1626
rect -702 -1694 -698 -1691
rect -694 -1691 -680 -1687
rect -694 -1694 -690 -1691
rect -666 -1694 -662 -1691
rect -658 -1691 -639 -1687
rect -658 -1694 -654 -1691
rect -632 -1694 -628 -1647
rect -606 -1658 -602 -1626
rect -606 -1687 -602 -1662
rect -572 -1680 -568 -1626
rect -572 -1684 -555 -1680
rect -624 -1694 -620 -1691
rect -615 -1691 -602 -1687
rect -615 -1694 -611 -1691
rect -588 -1694 -584 -1691
rect -564 -1694 -560 -1684
rect -548 -1687 -544 -1626
rect -540 -1680 -536 -1626
rect -514 -1647 -510 -1626
rect -540 -1684 -521 -1680
rect -556 -1691 -539 -1687
rect -556 -1694 -552 -1691
rect -532 -1694 -528 -1684
rect -514 -1694 -510 -1651
rect -745 -1702 -741 -1698
rect -719 -1702 -715 -1698
rect -676 -1702 -672 -1698
rect -641 -1702 -637 -1698
rect -597 -1702 -593 -1698
rect -580 -1702 -576 -1698
rect -544 -1702 -540 -1698
rect -523 -1702 -519 -1698
rect -505 -1716 -501 -1662
rect -489 -1665 -485 -1508
rect -471 -1650 -467 -1404
rect -460 -1483 -456 -1166
rect -427 -1192 -423 -1153
rect -427 -1207 -423 -1196
rect -446 -1211 -423 -1207
rect -420 -1183 -416 -1146
rect -446 -1214 -442 -1211
rect -420 -1214 -416 -1187
rect -429 -1222 -425 -1218
rect -437 -1302 -433 -1298
rect -411 -1302 -407 -1298
rect -394 -1302 -390 -1298
rect -354 -1302 -350 -1298
rect -333 -1302 -329 -1298
rect -316 -1302 -312 -1298
rect -276 -1302 -272 -1298
rect -252 -1302 -248 -1298
rect -215 -1302 -211 -1298
rect -446 -1327 -442 -1310
rect -446 -1378 -442 -1331
rect -428 -1320 -424 -1310
rect -428 -1378 -424 -1324
rect -420 -1349 -416 -1310
rect -402 -1342 -398 -1310
rect -420 -1378 -416 -1353
rect -402 -1378 -398 -1346
rect -376 -1334 -372 -1310
rect -376 -1371 -372 -1338
rect -342 -1371 -338 -1310
rect -324 -1327 -320 -1310
rect -394 -1378 -390 -1375
rect -386 -1375 -372 -1371
rect -386 -1378 -382 -1375
rect -358 -1378 -354 -1375
rect -350 -1375 -331 -1371
rect -350 -1378 -346 -1375
rect -324 -1378 -320 -1331
rect -298 -1342 -294 -1310
rect -298 -1371 -294 -1346
rect -264 -1364 -260 -1310
rect -264 -1368 -247 -1364
rect -316 -1378 -312 -1375
rect -307 -1375 -294 -1371
rect -307 -1378 -303 -1375
rect -280 -1378 -276 -1375
rect -256 -1378 -252 -1368
rect -240 -1371 -236 -1310
rect -232 -1364 -228 -1310
rect -206 -1334 -202 -1310
rect -232 -1368 -213 -1364
rect -248 -1375 -231 -1371
rect -248 -1378 -244 -1375
rect -224 -1378 -220 -1368
rect -206 -1378 -202 -1338
rect -437 -1386 -433 -1382
rect -411 -1386 -407 -1382
rect -368 -1386 -364 -1382
rect -333 -1386 -329 -1382
rect -289 -1386 -285 -1382
rect -272 -1386 -268 -1382
rect -236 -1386 -232 -1382
rect -215 -1386 -211 -1382
rect -198 -1407 -194 -1346
rect -186 -1349 -182 -1187
rect -170 -1334 -166 -1040
rect -152 -1162 -148 -1016
rect -120 -1057 -116 -1003
rect -139 -1061 -120 -1057
rect -113 -1028 -109 -996
rect 156 -1012 160 -948
rect 170 -988 174 -984
rect 187 -988 191 -984
rect 178 -999 182 -996
rect 178 -1003 193 -999
rect 156 -1016 171 -1012
rect -139 -1064 -135 -1061
rect -113 -1064 -109 -1032
rect -122 -1072 -118 -1068
rect -138 -1138 -134 -1134
rect -121 -1138 -117 -1134
rect -130 -1149 -126 -1146
rect -130 -1153 -115 -1149
rect -152 -1166 -137 -1162
rect -446 -1459 -442 -1455
rect -429 -1459 -425 -1455
rect -438 -1470 -434 -1467
rect -438 -1474 -423 -1470
rect -460 -1487 -445 -1483
rect -754 -1750 -750 -1746
rect -737 -1750 -733 -1746
rect -746 -1761 -742 -1758
rect -746 -1765 -731 -1761
rect -768 -1778 -753 -1774
rect -1062 -2072 -1058 -2068
rect -1045 -2072 -1041 -2068
rect -1054 -2083 -1050 -2080
rect -1054 -2087 -1039 -2083
rect -1076 -2100 -1061 -2096
rect -1225 -2315 -1221 -2311
rect -1181 -2315 -1177 -2311
rect -1147 -2315 -1143 -2311
rect -1309 -2363 -1305 -2359
rect -1292 -2363 -1288 -2359
rect -1301 -2374 -1297 -2371
rect -1301 -2378 -1286 -2374
rect -1319 -2391 -1308 -2387
rect -1319 -2678 -1315 -2391
rect -1290 -2417 -1286 -2378
rect -1290 -2432 -1286 -2421
rect -1309 -2436 -1286 -2432
rect -1309 -2439 -1305 -2436
rect -1283 -2439 -1279 -2371
rect -1292 -2447 -1288 -2443
rect -1283 -2577 -1279 -2443
rect -1257 -2570 -1253 -2326
rect -1225 -2522 -1221 -2518
rect -1208 -2522 -1204 -2518
rect -1168 -2522 -1164 -2518
rect -1147 -2522 -1143 -2518
rect -1234 -2563 -1230 -2530
rect -1234 -2598 -1230 -2567
rect -1216 -2557 -1212 -2530
rect -1216 -2561 -1207 -2557
rect -1216 -2598 -1212 -2561
rect -1190 -2584 -1186 -2530
rect -1190 -2591 -1186 -2588
rect -1156 -2591 -1152 -2530
rect -1138 -2562 -1134 -2530
rect -1106 -2554 -1102 -2412
rect -1208 -2598 -1204 -2595
rect -1199 -2595 -1186 -2591
rect -1199 -2598 -1195 -2595
rect -1172 -2598 -1168 -2595
rect -1164 -2595 -1145 -2591
rect -1164 -2598 -1160 -2595
rect -1138 -2598 -1134 -2566
rect -1090 -2569 -1086 -2333
rect -1076 -2387 -1072 -2100
rect -1043 -2126 -1039 -2087
rect -1043 -2141 -1039 -2130
rect -1062 -2145 -1039 -2141
rect -1036 -2117 -1032 -2080
rect -1062 -2148 -1058 -2145
rect -1036 -2148 -1032 -2121
rect -1045 -2156 -1041 -2152
rect -1053 -2231 -1049 -2227
rect -1027 -2231 -1023 -2227
rect -1010 -2231 -1006 -2227
rect -970 -2231 -966 -2227
rect -949 -2231 -945 -2227
rect -932 -2231 -928 -2227
rect -892 -2231 -888 -2227
rect -868 -2231 -864 -2227
rect -831 -2231 -827 -2227
rect -1062 -2256 -1058 -2239
rect -1062 -2307 -1058 -2260
rect -1044 -2249 -1040 -2239
rect -1044 -2307 -1040 -2253
rect -1036 -2278 -1032 -2239
rect -1018 -2271 -1014 -2239
rect -1036 -2307 -1032 -2282
rect -1018 -2307 -1014 -2275
rect -992 -2263 -988 -2239
rect -992 -2300 -988 -2267
rect -958 -2300 -954 -2239
rect -940 -2256 -936 -2239
rect -1010 -2307 -1006 -2304
rect -1002 -2304 -988 -2300
rect -1002 -2307 -998 -2304
rect -974 -2307 -970 -2304
rect -966 -2304 -947 -2300
rect -966 -2307 -962 -2304
rect -940 -2307 -936 -2260
rect -914 -2271 -910 -2239
rect -914 -2300 -910 -2275
rect -880 -2293 -876 -2239
rect -880 -2297 -863 -2293
rect -932 -2307 -928 -2304
rect -923 -2304 -910 -2300
rect -923 -2307 -919 -2304
rect -896 -2307 -892 -2304
rect -872 -2307 -868 -2297
rect -856 -2300 -852 -2239
rect -848 -2293 -844 -2239
rect -822 -2263 -818 -2239
rect -848 -2297 -829 -2293
rect -864 -2304 -847 -2300
rect -864 -2307 -860 -2304
rect -840 -2307 -836 -2297
rect -822 -2307 -818 -2267
rect -1053 -2315 -1049 -2311
rect -1027 -2315 -1023 -2311
rect -984 -2315 -980 -2311
rect -949 -2315 -945 -2311
rect -905 -2315 -901 -2311
rect -888 -2315 -884 -2311
rect -852 -2315 -848 -2311
rect -831 -2315 -827 -2311
rect -814 -2322 -810 -2275
rect -793 -2278 -789 -2121
rect -780 -2263 -776 -2004
rect -768 -2096 -764 -1778
rect -735 -1804 -731 -1765
rect -735 -1819 -731 -1808
rect -754 -1823 -731 -1819
rect -728 -1795 -724 -1758
rect -754 -1826 -750 -1823
rect -728 -1826 -724 -1799
rect -737 -1834 -733 -1830
rect -745 -1909 -741 -1905
rect -719 -1909 -715 -1905
rect -702 -1909 -698 -1905
rect -662 -1909 -658 -1905
rect -641 -1909 -637 -1905
rect -624 -1909 -620 -1905
rect -584 -1909 -580 -1905
rect -560 -1909 -556 -1905
rect -523 -1909 -519 -1905
rect -754 -1934 -750 -1917
rect -754 -1985 -750 -1938
rect -736 -1927 -732 -1917
rect -736 -1985 -732 -1931
rect -728 -1956 -724 -1917
rect -710 -1949 -706 -1917
rect -728 -1985 -724 -1960
rect -710 -1985 -706 -1953
rect -684 -1941 -680 -1917
rect -684 -1978 -680 -1945
rect -650 -1978 -646 -1917
rect -632 -1934 -628 -1917
rect -702 -1985 -698 -1982
rect -694 -1982 -680 -1978
rect -694 -1985 -690 -1982
rect -666 -1985 -662 -1982
rect -658 -1982 -639 -1978
rect -658 -1985 -654 -1982
rect -632 -1985 -628 -1938
rect -606 -1949 -602 -1917
rect -606 -1978 -602 -1953
rect -572 -1971 -568 -1917
rect -572 -1975 -555 -1971
rect -624 -1985 -620 -1982
rect -615 -1982 -602 -1978
rect -615 -1985 -611 -1982
rect -588 -1985 -584 -1982
rect -564 -1985 -560 -1975
rect -548 -1978 -544 -1917
rect -540 -1971 -536 -1917
rect -514 -1940 -510 -1917
rect -540 -1975 -521 -1971
rect -556 -1982 -539 -1978
rect -556 -1985 -552 -1982
rect -532 -1985 -528 -1975
rect -514 -1985 -510 -1944
rect -745 -1993 -741 -1989
rect -719 -1993 -715 -1989
rect -676 -1993 -672 -1989
rect -641 -1993 -637 -1989
rect -597 -1993 -593 -1989
rect -580 -1993 -576 -1989
rect -544 -1993 -540 -1989
rect -523 -1993 -519 -1989
rect -506 -2007 -502 -1953
rect -490 -1956 -486 -1799
rect -476 -1941 -472 -1720
rect -460 -1774 -456 -1487
rect -427 -1513 -423 -1474
rect -427 -1528 -423 -1517
rect -446 -1532 -423 -1528
rect -420 -1504 -416 -1467
rect -446 -1535 -442 -1532
rect -420 -1535 -416 -1508
rect -429 -1543 -425 -1539
rect -437 -1618 -433 -1614
rect -411 -1618 -407 -1614
rect -394 -1618 -390 -1614
rect -354 -1618 -350 -1614
rect -333 -1618 -329 -1614
rect -316 -1618 -312 -1614
rect -276 -1618 -272 -1614
rect -252 -1618 -248 -1614
rect -215 -1618 -211 -1614
rect -446 -1643 -442 -1626
rect -446 -1694 -442 -1647
rect -428 -1636 -424 -1626
rect -428 -1694 -424 -1640
rect -420 -1665 -416 -1626
rect -402 -1658 -398 -1626
rect -420 -1694 -416 -1669
rect -402 -1694 -398 -1662
rect -376 -1650 -372 -1626
rect -376 -1687 -372 -1654
rect -342 -1687 -338 -1626
rect -324 -1643 -320 -1626
rect -394 -1694 -390 -1691
rect -386 -1691 -372 -1687
rect -386 -1694 -382 -1691
rect -358 -1694 -354 -1691
rect -350 -1691 -331 -1687
rect -350 -1694 -346 -1691
rect -324 -1694 -320 -1647
rect -298 -1658 -294 -1626
rect -298 -1687 -294 -1662
rect -264 -1680 -260 -1626
rect -264 -1684 -247 -1680
rect -316 -1694 -312 -1691
rect -307 -1691 -294 -1687
rect -307 -1694 -303 -1691
rect -280 -1694 -276 -1691
rect -256 -1694 -252 -1684
rect -240 -1687 -236 -1626
rect -232 -1680 -228 -1626
rect -206 -1650 -202 -1626
rect -232 -1684 -213 -1680
rect -248 -1691 -231 -1687
rect -248 -1694 -244 -1691
rect -224 -1694 -220 -1684
rect -206 -1694 -202 -1654
rect -437 -1702 -433 -1698
rect -411 -1702 -407 -1698
rect -368 -1702 -364 -1698
rect -333 -1702 -329 -1698
rect -289 -1702 -285 -1698
rect -272 -1702 -268 -1698
rect -236 -1702 -232 -1698
rect -215 -1702 -211 -1698
rect -198 -1709 -194 -1662
rect -184 -1665 -180 -1508
rect -170 -1650 -166 -1411
rect -152 -1483 -148 -1166
rect -119 -1192 -115 -1153
rect -119 -1207 -115 -1196
rect -138 -1211 -115 -1207
rect -112 -1183 -108 -1146
rect -138 -1214 -134 -1211
rect -112 -1214 -108 -1187
rect -121 -1222 -117 -1218
rect -129 -1302 -125 -1298
rect -103 -1302 -99 -1298
rect -86 -1302 -82 -1298
rect -46 -1302 -42 -1298
rect -25 -1302 -21 -1298
rect -8 -1302 -4 -1298
rect 32 -1302 36 -1298
rect 56 -1302 60 -1298
rect 93 -1302 97 -1298
rect -138 -1327 -134 -1310
rect -138 -1378 -134 -1331
rect -120 -1320 -116 -1310
rect -120 -1378 -116 -1324
rect -112 -1349 -108 -1310
rect -94 -1342 -90 -1310
rect -112 -1378 -108 -1353
rect -94 -1378 -90 -1346
rect -68 -1334 -64 -1310
rect -68 -1371 -64 -1338
rect -34 -1371 -30 -1310
rect -16 -1327 -12 -1310
rect -86 -1378 -82 -1375
rect -78 -1375 -64 -1371
rect -78 -1378 -74 -1375
rect -50 -1378 -46 -1375
rect -42 -1375 -23 -1371
rect -42 -1378 -38 -1375
rect -16 -1378 -12 -1331
rect 10 -1342 14 -1310
rect 10 -1371 14 -1346
rect 44 -1364 48 -1310
rect 44 -1368 61 -1364
rect -8 -1378 -4 -1375
rect 1 -1375 14 -1371
rect 1 -1378 5 -1375
rect 28 -1378 32 -1375
rect 52 -1378 56 -1368
rect 68 -1371 72 -1310
rect 76 -1364 80 -1310
rect 102 -1334 106 -1310
rect 76 -1368 95 -1364
rect 60 -1375 77 -1371
rect 60 -1378 64 -1375
rect 84 -1378 88 -1368
rect 102 -1378 106 -1338
rect -129 -1386 -125 -1382
rect -103 -1386 -99 -1382
rect -60 -1386 -56 -1382
rect -25 -1386 -21 -1382
rect 19 -1386 23 -1382
rect 36 -1386 40 -1382
rect 72 -1386 76 -1382
rect 93 -1386 97 -1382
rect 109 -1400 113 -1346
rect 122 -1349 126 -1187
rect 145 -1334 149 -1032
rect 156 -1162 160 -1016
rect 189 -1057 193 -1003
rect 170 -1061 189 -1057
rect 196 -1036 200 -996
rect 464 -1012 468 -948
rect 478 -988 482 -984
rect 495 -988 499 -984
rect 486 -999 490 -996
rect 486 -1003 501 -999
rect 464 -1016 479 -1012
rect 170 -1064 174 -1061
rect 196 -1064 200 -1040
rect 187 -1072 191 -1068
rect 170 -1138 174 -1134
rect 187 -1138 191 -1134
rect 178 -1149 182 -1146
rect 178 -1153 193 -1149
rect 156 -1166 171 -1162
rect -138 -1459 -134 -1455
rect -121 -1459 -117 -1455
rect -130 -1470 -126 -1467
rect -130 -1474 -115 -1470
rect -152 -1487 -137 -1483
rect -446 -1750 -442 -1746
rect -429 -1750 -425 -1746
rect -438 -1761 -434 -1758
rect -438 -1765 -423 -1761
rect -460 -1778 -445 -1774
rect -754 -2072 -750 -2068
rect -737 -2072 -733 -2068
rect -746 -2083 -742 -2080
rect -746 -2087 -731 -2083
rect -768 -2100 -753 -2096
rect -1062 -2363 -1058 -2359
rect -1045 -2363 -1041 -2359
rect -1054 -2374 -1050 -2371
rect -1054 -2378 -1039 -2374
rect -1076 -2391 -1061 -2387
rect -1225 -2606 -1221 -2602
rect -1181 -2606 -1177 -2602
rect -1147 -2606 -1143 -2602
rect -1309 -2654 -1305 -2650
rect -1292 -2654 -1288 -2650
rect -1301 -2665 -1297 -2662
rect -1301 -2669 -1286 -2665
rect -1319 -2682 -1308 -2678
rect -1319 -2969 -1315 -2682
rect -1290 -2708 -1286 -2669
rect -1290 -2723 -1286 -2712
rect -1309 -2727 -1286 -2723
rect -1309 -2730 -1305 -2727
rect -1283 -2730 -1279 -2662
rect -1292 -2738 -1288 -2734
rect -1283 -2868 -1279 -2734
rect -1257 -2861 -1253 -2617
rect -1225 -2813 -1221 -2809
rect -1208 -2813 -1204 -2809
rect -1168 -2813 -1164 -2809
rect -1147 -2813 -1143 -2809
rect -1234 -2854 -1230 -2821
rect -1234 -2889 -1230 -2858
rect -1216 -2848 -1212 -2821
rect -1216 -2852 -1207 -2848
rect -1216 -2889 -1212 -2852
rect -1190 -2875 -1186 -2821
rect -1190 -2882 -1186 -2879
rect -1156 -2882 -1152 -2821
rect -1138 -2853 -1134 -2821
rect -1106 -2845 -1102 -2703
rect -1208 -2889 -1204 -2886
rect -1199 -2886 -1186 -2882
rect -1199 -2889 -1195 -2886
rect -1172 -2889 -1168 -2886
rect -1164 -2886 -1145 -2882
rect -1164 -2889 -1160 -2886
rect -1138 -2889 -1134 -2857
rect -1090 -2860 -1086 -2624
rect -1076 -2678 -1072 -2391
rect -1043 -2417 -1039 -2378
rect -1043 -2432 -1039 -2421
rect -1062 -2436 -1039 -2432
rect -1036 -2408 -1032 -2371
rect -1062 -2439 -1058 -2436
rect -1036 -2439 -1032 -2412
rect -1045 -2447 -1041 -2443
rect -1053 -2522 -1049 -2518
rect -1027 -2522 -1023 -2518
rect -1010 -2522 -1006 -2518
rect -970 -2522 -966 -2518
rect -949 -2522 -945 -2518
rect -932 -2522 -928 -2518
rect -892 -2522 -888 -2518
rect -868 -2522 -864 -2518
rect -831 -2522 -827 -2518
rect -1062 -2547 -1058 -2530
rect -1062 -2598 -1058 -2551
rect -1044 -2540 -1040 -2530
rect -1044 -2598 -1040 -2544
rect -1036 -2569 -1032 -2530
rect -1018 -2562 -1014 -2530
rect -1036 -2598 -1032 -2573
rect -1018 -2598 -1014 -2566
rect -992 -2554 -988 -2530
rect -992 -2591 -988 -2558
rect -958 -2591 -954 -2530
rect -940 -2547 -936 -2530
rect -1010 -2598 -1006 -2595
rect -1002 -2595 -988 -2591
rect -1002 -2598 -998 -2595
rect -974 -2598 -970 -2595
rect -966 -2595 -947 -2591
rect -966 -2598 -962 -2595
rect -940 -2598 -936 -2551
rect -914 -2562 -910 -2530
rect -914 -2591 -910 -2566
rect -880 -2584 -876 -2530
rect -880 -2588 -863 -2584
rect -932 -2598 -928 -2595
rect -923 -2595 -910 -2591
rect -923 -2598 -919 -2595
rect -896 -2598 -892 -2595
rect -872 -2598 -868 -2588
rect -856 -2591 -852 -2530
rect -848 -2584 -844 -2530
rect -822 -2554 -818 -2530
rect -848 -2588 -829 -2584
rect -864 -2595 -847 -2591
rect -864 -2598 -860 -2595
rect -840 -2598 -836 -2588
rect -822 -2598 -818 -2558
rect -1053 -2606 -1049 -2602
rect -1027 -2606 -1023 -2602
rect -984 -2606 -980 -2602
rect -949 -2606 -945 -2602
rect -905 -2606 -901 -2602
rect -888 -2606 -884 -2602
rect -852 -2606 -848 -2602
rect -831 -2606 -827 -2602
rect -814 -2613 -810 -2566
rect -793 -2569 -789 -2412
rect -780 -2554 -776 -2326
rect -768 -2387 -764 -2100
rect -735 -2126 -731 -2087
rect -735 -2141 -731 -2130
rect -754 -2145 -731 -2141
rect -728 -2117 -724 -2080
rect -754 -2148 -750 -2145
rect -728 -2148 -724 -2121
rect -737 -2156 -733 -2152
rect -745 -2231 -741 -2227
rect -719 -2231 -715 -2227
rect -702 -2231 -698 -2227
rect -662 -2231 -658 -2227
rect -641 -2231 -637 -2227
rect -624 -2231 -620 -2227
rect -584 -2231 -580 -2227
rect -560 -2231 -556 -2227
rect -523 -2231 -519 -2227
rect -754 -2256 -750 -2239
rect -754 -2307 -750 -2260
rect -736 -2249 -732 -2239
rect -736 -2307 -732 -2253
rect -728 -2278 -724 -2239
rect -710 -2271 -706 -2239
rect -728 -2307 -724 -2282
rect -710 -2307 -706 -2275
rect -684 -2263 -680 -2239
rect -684 -2300 -680 -2267
rect -650 -2300 -646 -2239
rect -632 -2256 -628 -2239
rect -702 -2307 -698 -2304
rect -694 -2304 -680 -2300
rect -694 -2307 -690 -2304
rect -666 -2307 -662 -2304
rect -658 -2304 -639 -2300
rect -658 -2307 -654 -2304
rect -632 -2307 -628 -2260
rect -606 -2271 -602 -2239
rect -606 -2300 -602 -2275
rect -572 -2293 -568 -2239
rect -572 -2297 -555 -2293
rect -624 -2307 -620 -2304
rect -615 -2304 -602 -2300
rect -615 -2307 -611 -2304
rect -588 -2307 -584 -2304
rect -564 -2307 -560 -2297
rect -548 -2300 -544 -2239
rect -540 -2293 -536 -2239
rect -514 -2262 -510 -2239
rect -540 -2297 -521 -2293
rect -556 -2304 -539 -2300
rect -556 -2307 -552 -2304
rect -532 -2307 -528 -2297
rect -514 -2307 -510 -2266
rect -745 -2315 -741 -2311
rect -719 -2315 -715 -2311
rect -676 -2315 -672 -2311
rect -641 -2315 -637 -2311
rect -597 -2315 -593 -2311
rect -580 -2315 -576 -2311
rect -544 -2315 -540 -2311
rect -523 -2315 -519 -2311
rect -505 -2329 -501 -2275
rect -490 -2278 -486 -2121
rect -476 -2263 -472 -2011
rect -460 -2096 -456 -1778
rect -427 -1804 -423 -1765
rect -427 -1819 -423 -1808
rect -446 -1823 -423 -1819
rect -420 -1795 -416 -1758
rect -446 -1826 -442 -1823
rect -420 -1826 -416 -1799
rect -429 -1834 -425 -1830
rect -437 -1909 -433 -1905
rect -411 -1909 -407 -1905
rect -394 -1909 -390 -1905
rect -354 -1909 -350 -1905
rect -333 -1909 -329 -1905
rect -316 -1909 -312 -1905
rect -276 -1909 -272 -1905
rect -252 -1909 -248 -1905
rect -215 -1909 -211 -1905
rect -446 -1934 -442 -1917
rect -446 -1985 -442 -1938
rect -428 -1927 -424 -1917
rect -428 -1985 -424 -1931
rect -420 -1956 -416 -1917
rect -402 -1949 -398 -1917
rect -420 -1985 -416 -1960
rect -402 -1985 -398 -1953
rect -376 -1941 -372 -1917
rect -376 -1978 -372 -1945
rect -342 -1978 -338 -1917
rect -324 -1934 -320 -1917
rect -394 -1985 -390 -1982
rect -386 -1982 -372 -1978
rect -386 -1985 -382 -1982
rect -358 -1985 -354 -1982
rect -350 -1982 -331 -1978
rect -350 -1985 -346 -1982
rect -324 -1985 -320 -1938
rect -298 -1949 -294 -1917
rect -298 -1978 -294 -1953
rect -264 -1971 -260 -1917
rect -264 -1975 -247 -1971
rect -316 -1985 -312 -1982
rect -307 -1982 -294 -1978
rect -307 -1985 -303 -1982
rect -280 -1985 -276 -1982
rect -256 -1985 -252 -1975
rect -240 -1978 -236 -1917
rect -232 -1971 -228 -1917
rect -206 -1941 -202 -1917
rect -232 -1975 -213 -1971
rect -248 -1982 -231 -1978
rect -248 -1985 -244 -1982
rect -224 -1985 -220 -1975
rect -206 -1985 -202 -1945
rect -437 -1993 -433 -1989
rect -411 -1993 -407 -1989
rect -368 -1993 -364 -1989
rect -333 -1993 -329 -1989
rect -289 -1993 -285 -1989
rect -272 -1993 -268 -1989
rect -236 -1993 -232 -1989
rect -215 -1993 -211 -1989
rect -199 -2000 -195 -1953
rect -180 -1956 -176 -1799
rect -166 -1941 -162 -1713
rect -152 -1774 -148 -1487
rect -119 -1513 -115 -1474
rect -119 -1528 -115 -1517
rect -138 -1532 -115 -1528
rect -112 -1504 -108 -1467
rect -138 -1535 -134 -1532
rect -112 -1535 -108 -1508
rect -121 -1543 -117 -1539
rect -129 -1618 -125 -1614
rect -103 -1618 -99 -1614
rect -86 -1618 -82 -1614
rect -46 -1618 -42 -1614
rect -25 -1618 -21 -1614
rect -8 -1618 -4 -1614
rect 32 -1618 36 -1614
rect 56 -1618 60 -1614
rect 93 -1618 97 -1614
rect -138 -1643 -134 -1626
rect -138 -1694 -134 -1647
rect -120 -1636 -116 -1626
rect -120 -1694 -116 -1640
rect -112 -1665 -108 -1626
rect -94 -1658 -90 -1626
rect -112 -1694 -108 -1669
rect -94 -1694 -90 -1662
rect -68 -1650 -64 -1626
rect -68 -1687 -64 -1654
rect -34 -1687 -30 -1626
rect -16 -1643 -12 -1626
rect -86 -1694 -82 -1691
rect -78 -1691 -64 -1687
rect -78 -1694 -74 -1691
rect -50 -1694 -46 -1691
rect -42 -1691 -23 -1687
rect -42 -1694 -38 -1691
rect -16 -1694 -12 -1647
rect 10 -1658 14 -1626
rect 10 -1687 14 -1662
rect 44 -1680 48 -1626
rect 44 -1684 61 -1680
rect -8 -1694 -4 -1691
rect 1 -1691 14 -1687
rect 1 -1694 5 -1691
rect 28 -1694 32 -1691
rect 52 -1694 56 -1684
rect 68 -1687 72 -1626
rect 76 -1680 80 -1626
rect 102 -1650 106 -1626
rect 76 -1684 95 -1680
rect 60 -1691 77 -1687
rect 60 -1694 64 -1691
rect 84 -1694 88 -1684
rect 102 -1694 106 -1654
rect -129 -1702 -125 -1698
rect -103 -1702 -99 -1698
rect -60 -1702 -56 -1698
rect -25 -1702 -21 -1698
rect 19 -1702 23 -1698
rect 36 -1702 40 -1698
rect 72 -1702 76 -1698
rect 93 -1702 97 -1698
rect 111 -1716 115 -1662
rect 126 -1665 130 -1508
rect 145 -1650 149 -1404
rect 156 -1483 160 -1166
rect 189 -1192 193 -1153
rect 189 -1207 193 -1196
rect 170 -1211 193 -1207
rect 196 -1183 200 -1146
rect 170 -1214 174 -1211
rect 196 -1214 200 -1187
rect 187 -1222 191 -1218
rect 179 -1302 183 -1298
rect 205 -1302 209 -1298
rect 222 -1302 226 -1298
rect 262 -1302 266 -1298
rect 283 -1302 287 -1298
rect 300 -1302 304 -1298
rect 340 -1302 344 -1298
rect 364 -1302 368 -1298
rect 401 -1302 405 -1298
rect 170 -1327 174 -1310
rect 170 -1378 174 -1331
rect 188 -1320 192 -1310
rect 188 -1378 192 -1324
rect 196 -1349 200 -1310
rect 214 -1342 218 -1310
rect 196 -1378 200 -1353
rect 214 -1378 218 -1346
rect 240 -1334 244 -1310
rect 240 -1371 244 -1338
rect 274 -1371 278 -1310
rect 292 -1327 296 -1310
rect 222 -1378 226 -1375
rect 230 -1375 244 -1371
rect 230 -1378 234 -1375
rect 258 -1378 262 -1375
rect 266 -1375 285 -1371
rect 266 -1378 270 -1375
rect 292 -1378 296 -1331
rect 318 -1342 322 -1310
rect 318 -1371 322 -1346
rect 352 -1364 356 -1310
rect 352 -1368 369 -1364
rect 300 -1378 304 -1375
rect 309 -1375 322 -1371
rect 309 -1378 313 -1375
rect 336 -1378 340 -1375
rect 360 -1378 364 -1368
rect 376 -1371 380 -1310
rect 384 -1364 388 -1310
rect 410 -1334 414 -1310
rect 384 -1368 403 -1364
rect 368 -1375 385 -1371
rect 368 -1378 372 -1375
rect 392 -1378 396 -1368
rect 410 -1378 414 -1338
rect 179 -1386 183 -1382
rect 205 -1386 209 -1382
rect 248 -1386 252 -1382
rect 283 -1386 287 -1382
rect 327 -1386 331 -1382
rect 344 -1386 348 -1382
rect 380 -1386 384 -1382
rect 401 -1386 405 -1382
rect 417 -1407 421 -1346
rect 430 -1349 434 -1187
rect 446 -1334 450 -1040
rect 464 -1162 468 -1016
rect 497 -1057 501 -1003
rect 478 -1061 497 -1057
rect 504 -1028 508 -996
rect 478 -1064 482 -1061
rect 504 -1064 508 -1032
rect 772 -1012 776 -948
rect 786 -988 790 -984
rect 803 -988 807 -984
rect 794 -999 798 -996
rect 794 -1003 809 -999
rect 772 -1016 787 -1012
rect 495 -1072 499 -1068
rect 478 -1138 482 -1134
rect 495 -1138 499 -1134
rect 486 -1149 490 -1146
rect 486 -1153 501 -1149
rect 464 -1166 479 -1162
rect 170 -1459 174 -1455
rect 187 -1459 191 -1455
rect 178 -1470 182 -1467
rect 178 -1474 193 -1470
rect 156 -1487 171 -1483
rect -138 -1750 -134 -1746
rect -121 -1750 -117 -1746
rect -130 -1761 -126 -1758
rect -130 -1765 -115 -1761
rect -152 -1778 -137 -1774
rect -446 -2072 -442 -2068
rect -429 -2072 -425 -2068
rect -438 -2083 -434 -2080
rect -438 -2087 -423 -2083
rect -460 -2100 -445 -2096
rect -754 -2363 -750 -2359
rect -737 -2363 -733 -2359
rect -746 -2374 -742 -2371
rect -746 -2378 -731 -2374
rect -768 -2391 -753 -2387
rect -1062 -2654 -1058 -2650
rect -1045 -2654 -1041 -2650
rect -1054 -2665 -1050 -2662
rect -1054 -2669 -1039 -2665
rect -1076 -2682 -1061 -2678
rect -1225 -2897 -1221 -2893
rect -1181 -2897 -1177 -2893
rect -1147 -2897 -1143 -2893
rect -1309 -2945 -1305 -2941
rect -1292 -2945 -1288 -2941
rect -1301 -2956 -1297 -2953
rect -1301 -2960 -1286 -2956
rect -1319 -2973 -1308 -2969
rect -1290 -2999 -1286 -2960
rect -1290 -3014 -1286 -3003
rect -1309 -3018 -1286 -3014
rect -1309 -3021 -1305 -3018
rect -1283 -3021 -1279 -2953
rect -1292 -3029 -1288 -3025
rect -1283 -3159 -1279 -3025
rect -1257 -3152 -1253 -2908
rect -1225 -3104 -1221 -3100
rect -1208 -3104 -1204 -3100
rect -1168 -3104 -1164 -3100
rect -1147 -3104 -1143 -3100
rect -1234 -3145 -1230 -3112
rect -1234 -3180 -1230 -3149
rect -1216 -3139 -1212 -3112
rect -1216 -3143 -1207 -3139
rect -1216 -3180 -1212 -3143
rect -1190 -3166 -1186 -3112
rect -1190 -3173 -1186 -3170
rect -1156 -3173 -1152 -3112
rect -1138 -3144 -1134 -3112
rect -1106 -3136 -1102 -2994
rect -1208 -3180 -1204 -3177
rect -1199 -3177 -1186 -3173
rect -1199 -3180 -1195 -3177
rect -1172 -3180 -1168 -3177
rect -1164 -3177 -1145 -3173
rect -1164 -3180 -1160 -3177
rect -1138 -3180 -1134 -3148
rect -1090 -3151 -1086 -2915
rect -1076 -2969 -1072 -2682
rect -1043 -2708 -1039 -2669
rect -1043 -2723 -1039 -2712
rect -1062 -2727 -1039 -2723
rect -1036 -2699 -1032 -2662
rect -1062 -2730 -1058 -2727
rect -1036 -2730 -1032 -2703
rect -1045 -2738 -1041 -2734
rect -1053 -2813 -1049 -2809
rect -1027 -2813 -1023 -2809
rect -1010 -2813 -1006 -2809
rect -970 -2813 -966 -2809
rect -949 -2813 -945 -2809
rect -932 -2813 -928 -2809
rect -892 -2813 -888 -2809
rect -868 -2813 -864 -2809
rect -831 -2813 -827 -2809
rect -1062 -2838 -1058 -2821
rect -1062 -2889 -1058 -2842
rect -1044 -2831 -1040 -2821
rect -1044 -2889 -1040 -2835
rect -1036 -2860 -1032 -2821
rect -1018 -2853 -1014 -2821
rect -1036 -2889 -1032 -2864
rect -1018 -2889 -1014 -2857
rect -992 -2845 -988 -2821
rect -992 -2882 -988 -2849
rect -958 -2882 -954 -2821
rect -940 -2838 -936 -2821
rect -1010 -2889 -1006 -2886
rect -1002 -2886 -988 -2882
rect -1002 -2889 -998 -2886
rect -974 -2889 -970 -2886
rect -966 -2886 -947 -2882
rect -966 -2889 -962 -2886
rect -940 -2889 -936 -2842
rect -914 -2853 -910 -2821
rect -914 -2882 -910 -2857
rect -880 -2875 -876 -2821
rect -880 -2879 -863 -2875
rect -932 -2889 -928 -2886
rect -923 -2886 -910 -2882
rect -923 -2889 -919 -2886
rect -896 -2889 -892 -2886
rect -872 -2889 -868 -2879
rect -856 -2882 -852 -2821
rect -848 -2875 -844 -2821
rect -822 -2845 -818 -2821
rect -848 -2879 -829 -2875
rect -864 -2886 -847 -2882
rect -864 -2889 -860 -2886
rect -840 -2889 -836 -2879
rect -822 -2889 -818 -2849
rect -1053 -2897 -1049 -2893
rect -1027 -2897 -1023 -2893
rect -984 -2897 -980 -2893
rect -949 -2897 -945 -2893
rect -905 -2897 -901 -2893
rect -888 -2897 -884 -2893
rect -852 -2897 -848 -2893
rect -831 -2897 -827 -2893
rect -814 -2904 -810 -2857
rect -793 -2860 -789 -2703
rect -780 -2845 -776 -2617
rect -768 -2678 -764 -2391
rect -735 -2417 -731 -2378
rect -735 -2432 -731 -2421
rect -754 -2436 -731 -2432
rect -728 -2408 -724 -2371
rect -754 -2439 -750 -2436
rect -728 -2439 -724 -2412
rect -737 -2447 -733 -2443
rect -745 -2522 -741 -2518
rect -719 -2522 -715 -2518
rect -702 -2522 -698 -2518
rect -662 -2522 -658 -2518
rect -641 -2522 -637 -2518
rect -624 -2522 -620 -2518
rect -584 -2522 -580 -2518
rect -560 -2522 -556 -2518
rect -523 -2522 -519 -2518
rect -754 -2547 -750 -2530
rect -754 -2598 -750 -2551
rect -736 -2540 -732 -2530
rect -736 -2598 -732 -2544
rect -728 -2569 -724 -2530
rect -710 -2562 -706 -2530
rect -728 -2598 -724 -2573
rect -710 -2598 -706 -2566
rect -684 -2554 -680 -2530
rect -684 -2591 -680 -2558
rect -650 -2591 -646 -2530
rect -632 -2547 -628 -2530
rect -702 -2598 -698 -2595
rect -694 -2595 -680 -2591
rect -694 -2598 -690 -2595
rect -666 -2598 -662 -2595
rect -658 -2595 -639 -2591
rect -658 -2598 -654 -2595
rect -632 -2598 -628 -2551
rect -606 -2562 -602 -2530
rect -606 -2591 -602 -2566
rect -572 -2584 -568 -2530
rect -572 -2588 -555 -2584
rect -624 -2598 -620 -2595
rect -615 -2595 -602 -2591
rect -615 -2598 -611 -2595
rect -588 -2598 -584 -2595
rect -564 -2598 -560 -2588
rect -548 -2591 -544 -2530
rect -540 -2584 -536 -2530
rect -514 -2553 -510 -2530
rect -540 -2588 -521 -2584
rect -556 -2595 -539 -2591
rect -556 -2598 -552 -2595
rect -532 -2598 -528 -2588
rect -514 -2598 -510 -2557
rect -745 -2606 -741 -2602
rect -719 -2606 -715 -2602
rect -676 -2606 -672 -2602
rect -641 -2606 -637 -2602
rect -597 -2606 -593 -2602
rect -580 -2606 -576 -2602
rect -544 -2606 -540 -2602
rect -523 -2606 -519 -2602
rect -505 -2620 -501 -2566
rect -490 -2569 -486 -2412
rect -476 -2554 -472 -2333
rect -460 -2387 -456 -2100
rect -427 -2126 -423 -2087
rect -427 -2141 -423 -2130
rect -446 -2145 -423 -2141
rect -420 -2117 -416 -2080
rect -446 -2148 -442 -2145
rect -420 -2148 -416 -2121
rect -429 -2156 -425 -2152
rect -437 -2231 -433 -2227
rect -411 -2231 -407 -2227
rect -394 -2231 -390 -2227
rect -354 -2231 -350 -2227
rect -333 -2231 -329 -2227
rect -316 -2231 -312 -2227
rect -276 -2231 -272 -2227
rect -252 -2231 -248 -2227
rect -215 -2231 -211 -2227
rect -446 -2256 -442 -2239
rect -446 -2307 -442 -2260
rect -428 -2249 -424 -2239
rect -428 -2307 -424 -2253
rect -420 -2278 -416 -2239
rect -402 -2271 -398 -2239
rect -420 -2307 -416 -2282
rect -402 -2307 -398 -2275
rect -376 -2263 -372 -2239
rect -376 -2300 -372 -2267
rect -342 -2300 -338 -2239
rect -324 -2256 -320 -2239
rect -394 -2307 -390 -2304
rect -386 -2304 -372 -2300
rect -386 -2307 -382 -2304
rect -358 -2307 -354 -2304
rect -350 -2304 -331 -2300
rect -350 -2307 -346 -2304
rect -324 -2307 -320 -2260
rect -298 -2271 -294 -2239
rect -298 -2300 -294 -2275
rect -264 -2293 -260 -2239
rect -264 -2297 -247 -2293
rect -316 -2307 -312 -2304
rect -307 -2304 -294 -2300
rect -307 -2307 -303 -2304
rect -280 -2307 -276 -2304
rect -256 -2307 -252 -2297
rect -240 -2300 -236 -2239
rect -232 -2293 -228 -2239
rect -206 -2263 -202 -2239
rect -232 -2297 -213 -2293
rect -248 -2304 -231 -2300
rect -248 -2307 -244 -2304
rect -224 -2307 -220 -2297
rect -206 -2307 -202 -2267
rect -437 -2315 -433 -2311
rect -411 -2315 -407 -2311
rect -368 -2315 -364 -2311
rect -333 -2315 -329 -2311
rect -289 -2315 -285 -2311
rect -272 -2315 -268 -2311
rect -236 -2315 -232 -2311
rect -215 -2315 -211 -2311
rect -198 -2322 -194 -2275
rect -180 -2278 -176 -2121
rect -166 -2263 -162 -2004
rect -152 -2096 -148 -1778
rect -119 -1804 -115 -1765
rect -119 -1819 -115 -1808
rect -138 -1823 -115 -1819
rect -112 -1795 -108 -1758
rect -138 -1826 -134 -1823
rect -112 -1826 -108 -1799
rect -121 -1834 -117 -1830
rect -129 -1909 -125 -1905
rect -103 -1909 -99 -1905
rect -86 -1909 -82 -1905
rect -46 -1909 -42 -1905
rect -25 -1909 -21 -1905
rect -8 -1909 -4 -1905
rect 32 -1909 36 -1905
rect 56 -1909 60 -1905
rect 93 -1909 97 -1905
rect -138 -1934 -134 -1917
rect -138 -1985 -134 -1938
rect -120 -1927 -116 -1917
rect -120 -1985 -116 -1931
rect -112 -1956 -108 -1917
rect -94 -1949 -90 -1917
rect -112 -1985 -108 -1960
rect -94 -1985 -90 -1953
rect -68 -1941 -64 -1917
rect -68 -1978 -64 -1945
rect -34 -1978 -30 -1917
rect -16 -1934 -12 -1917
rect -86 -1985 -82 -1982
rect -78 -1982 -64 -1978
rect -78 -1985 -74 -1982
rect -50 -1985 -46 -1982
rect -42 -1982 -23 -1978
rect -42 -1985 -38 -1982
rect -16 -1985 -12 -1938
rect 10 -1949 14 -1917
rect 10 -1978 14 -1953
rect 44 -1971 48 -1917
rect 44 -1975 61 -1971
rect -8 -1985 -4 -1982
rect 1 -1982 14 -1978
rect 1 -1985 5 -1982
rect 28 -1985 32 -1982
rect 52 -1985 56 -1975
rect 68 -1978 72 -1917
rect 76 -1971 80 -1917
rect 102 -1941 106 -1917
rect 76 -1975 95 -1971
rect 60 -1982 77 -1978
rect 60 -1985 64 -1982
rect 84 -1985 88 -1975
rect 102 -1985 106 -1945
rect -129 -1993 -125 -1989
rect -103 -1993 -99 -1989
rect -60 -1993 -56 -1989
rect -25 -1993 -21 -1989
rect 19 -1993 23 -1989
rect 36 -1993 40 -1989
rect 72 -1993 76 -1989
rect 93 -1993 97 -1989
rect 112 -2007 116 -1953
rect 126 -1956 130 -1799
rect 140 -1941 144 -1720
rect 156 -1774 160 -1487
rect 189 -1513 193 -1474
rect 189 -1528 193 -1517
rect 170 -1532 193 -1528
rect 196 -1504 200 -1467
rect 170 -1535 174 -1532
rect 196 -1535 200 -1508
rect 187 -1543 191 -1539
rect 179 -1618 183 -1614
rect 205 -1618 209 -1614
rect 222 -1618 226 -1614
rect 262 -1618 266 -1614
rect 283 -1618 287 -1614
rect 300 -1618 304 -1614
rect 340 -1618 344 -1614
rect 364 -1618 368 -1614
rect 401 -1618 405 -1614
rect 170 -1643 174 -1626
rect 170 -1694 174 -1647
rect 188 -1636 192 -1626
rect 188 -1694 192 -1640
rect 196 -1665 200 -1626
rect 214 -1658 218 -1626
rect 196 -1694 200 -1669
rect 214 -1694 218 -1662
rect 240 -1650 244 -1626
rect 240 -1687 244 -1654
rect 274 -1687 278 -1626
rect 292 -1643 296 -1626
rect 222 -1694 226 -1691
rect 230 -1691 244 -1687
rect 230 -1694 234 -1691
rect 258 -1694 262 -1691
rect 266 -1691 285 -1687
rect 266 -1694 270 -1691
rect 292 -1694 296 -1647
rect 318 -1658 322 -1626
rect 318 -1687 322 -1662
rect 352 -1680 356 -1626
rect 352 -1684 369 -1680
rect 300 -1694 304 -1691
rect 309 -1691 322 -1687
rect 309 -1694 313 -1691
rect 336 -1694 340 -1691
rect 360 -1694 364 -1684
rect 376 -1687 380 -1626
rect 384 -1680 388 -1626
rect 410 -1650 414 -1626
rect 384 -1684 403 -1680
rect 368 -1691 385 -1687
rect 368 -1694 372 -1691
rect 392 -1694 396 -1684
rect 410 -1694 414 -1654
rect 179 -1702 183 -1698
rect 205 -1702 209 -1698
rect 248 -1702 252 -1698
rect 283 -1702 287 -1698
rect 327 -1702 331 -1698
rect 344 -1702 348 -1698
rect 380 -1702 384 -1698
rect 401 -1702 405 -1698
rect 418 -1709 422 -1662
rect 434 -1665 438 -1508
rect 448 -1650 452 -1411
rect 464 -1483 468 -1166
rect 497 -1192 501 -1153
rect 497 -1207 501 -1196
rect 478 -1211 501 -1207
rect 504 -1183 508 -1146
rect 772 -1162 776 -1016
rect 805 -1057 809 -1003
rect 786 -1061 805 -1057
rect 812 -1036 816 -996
rect 786 -1064 790 -1061
rect 812 -1064 816 -1040
rect 803 -1072 807 -1068
rect 786 -1138 790 -1134
rect 803 -1138 807 -1134
rect 794 -1149 798 -1146
rect 794 -1153 809 -1149
rect 772 -1166 787 -1162
rect 478 -1214 482 -1211
rect 504 -1214 508 -1187
rect 495 -1222 499 -1218
rect 487 -1302 491 -1298
rect 513 -1302 517 -1298
rect 530 -1302 534 -1298
rect 570 -1302 574 -1298
rect 591 -1302 595 -1298
rect 608 -1302 612 -1298
rect 648 -1302 652 -1298
rect 672 -1302 676 -1298
rect 709 -1302 713 -1298
rect 478 -1327 482 -1310
rect 478 -1378 482 -1331
rect 496 -1320 500 -1310
rect 496 -1378 500 -1324
rect 504 -1349 508 -1310
rect 522 -1342 526 -1310
rect 504 -1378 508 -1353
rect 522 -1378 526 -1346
rect 548 -1334 552 -1310
rect 548 -1371 552 -1338
rect 582 -1371 586 -1310
rect 600 -1327 604 -1310
rect 530 -1378 534 -1375
rect 538 -1375 552 -1371
rect 538 -1378 542 -1375
rect 566 -1378 570 -1375
rect 574 -1375 593 -1371
rect 574 -1378 578 -1375
rect 600 -1378 604 -1331
rect 626 -1342 630 -1310
rect 626 -1371 630 -1346
rect 660 -1364 664 -1310
rect 660 -1368 677 -1364
rect 608 -1378 612 -1375
rect 617 -1375 630 -1371
rect 617 -1378 621 -1375
rect 644 -1378 648 -1375
rect 668 -1378 672 -1368
rect 684 -1371 688 -1310
rect 692 -1364 696 -1310
rect 718 -1350 722 -1310
rect 692 -1368 711 -1364
rect 676 -1375 693 -1371
rect 676 -1378 680 -1375
rect 700 -1378 704 -1368
rect 718 -1378 722 -1354
rect 487 -1386 491 -1382
rect 513 -1386 517 -1382
rect 556 -1386 560 -1382
rect 591 -1386 595 -1382
rect 635 -1386 639 -1382
rect 652 -1386 656 -1382
rect 688 -1386 692 -1382
rect 709 -1386 713 -1382
rect 725 -1400 729 -1346
rect 738 -1357 742 -1187
rect 478 -1459 482 -1455
rect 495 -1459 499 -1455
rect 486 -1470 490 -1467
rect 486 -1474 501 -1470
rect 464 -1487 479 -1483
rect 170 -1750 174 -1746
rect 187 -1750 191 -1746
rect 178 -1761 182 -1758
rect 178 -1765 193 -1761
rect 156 -1778 171 -1774
rect -138 -2072 -134 -2068
rect -121 -2072 -117 -2068
rect -130 -2083 -126 -2080
rect -130 -2087 -115 -2083
rect -152 -2100 -137 -2096
rect -446 -2363 -442 -2359
rect -429 -2363 -425 -2359
rect -438 -2374 -434 -2371
rect -438 -2378 -423 -2374
rect -460 -2391 -445 -2387
rect -754 -2654 -750 -2650
rect -737 -2654 -733 -2650
rect -746 -2665 -742 -2662
rect -746 -2669 -731 -2665
rect -768 -2682 -753 -2678
rect -1062 -2945 -1058 -2941
rect -1045 -2945 -1041 -2941
rect -1054 -2956 -1050 -2953
rect -1054 -2960 -1039 -2956
rect -1076 -2973 -1061 -2969
rect -1043 -2999 -1039 -2960
rect -1043 -3014 -1039 -3003
rect -1062 -3018 -1039 -3014
rect -1036 -2990 -1032 -2953
rect -1062 -3021 -1058 -3018
rect -1036 -3021 -1032 -2994
rect -1045 -3029 -1041 -3025
rect -1225 -3188 -1221 -3184
rect -1181 -3188 -1177 -3184
rect -1147 -3188 -1143 -3184
rect -1076 -3192 -1072 -3096
rect -1053 -3104 -1049 -3100
rect -1027 -3104 -1023 -3100
rect -1010 -3104 -1006 -3100
rect -970 -3104 -966 -3100
rect -949 -3104 -945 -3100
rect -932 -3104 -928 -3100
rect -892 -3104 -888 -3100
rect -868 -3104 -864 -3100
rect -831 -3104 -827 -3100
rect -1062 -3129 -1058 -3112
rect -1062 -3180 -1058 -3133
rect -1044 -3122 -1040 -3112
rect -1044 -3180 -1040 -3126
rect -1036 -3151 -1032 -3112
rect -1018 -3144 -1014 -3112
rect -1036 -3180 -1032 -3155
rect -1018 -3180 -1014 -3148
rect -992 -3136 -988 -3112
rect -992 -3173 -988 -3140
rect -958 -3173 -954 -3112
rect -940 -3129 -936 -3112
rect -1010 -3180 -1006 -3177
rect -1002 -3177 -988 -3173
rect -1002 -3180 -998 -3177
rect -974 -3180 -970 -3177
rect -966 -3177 -947 -3173
rect -966 -3180 -962 -3177
rect -940 -3180 -936 -3133
rect -914 -3144 -910 -3112
rect -914 -3173 -910 -3148
rect -880 -3166 -876 -3112
rect -880 -3170 -863 -3166
rect -932 -3180 -928 -3177
rect -923 -3177 -910 -3173
rect -923 -3180 -919 -3177
rect -896 -3180 -892 -3177
rect -872 -3180 -868 -3170
rect -856 -3173 -852 -3112
rect -848 -3166 -844 -3112
rect -822 -3136 -818 -3112
rect -848 -3170 -829 -3166
rect -864 -3177 -847 -3173
rect -864 -3180 -860 -3177
rect -840 -3180 -836 -3170
rect -822 -3180 -818 -3140
rect -793 -3151 -789 -2994
rect -780 -3136 -776 -2908
rect -768 -2969 -764 -2682
rect -735 -2708 -731 -2669
rect -735 -2723 -731 -2712
rect -754 -2727 -731 -2723
rect -728 -2699 -724 -2662
rect -754 -2730 -750 -2727
rect -728 -2730 -724 -2703
rect -737 -2738 -733 -2734
rect -745 -2813 -741 -2809
rect -719 -2813 -715 -2809
rect -702 -2813 -698 -2809
rect -662 -2813 -658 -2809
rect -641 -2813 -637 -2809
rect -624 -2813 -620 -2809
rect -584 -2813 -580 -2809
rect -560 -2813 -556 -2809
rect -523 -2813 -519 -2809
rect -754 -2838 -750 -2821
rect -754 -2889 -750 -2842
rect -736 -2831 -732 -2821
rect -736 -2889 -732 -2835
rect -728 -2860 -724 -2821
rect -710 -2853 -706 -2821
rect -728 -2889 -724 -2864
rect -710 -2889 -706 -2857
rect -684 -2845 -680 -2821
rect -684 -2882 -680 -2849
rect -650 -2882 -646 -2821
rect -632 -2838 -628 -2821
rect -702 -2889 -698 -2886
rect -694 -2886 -680 -2882
rect -694 -2889 -690 -2886
rect -666 -2889 -662 -2886
rect -658 -2886 -639 -2882
rect -658 -2889 -654 -2886
rect -632 -2889 -628 -2842
rect -606 -2853 -602 -2821
rect -606 -2882 -602 -2857
rect -572 -2875 -568 -2821
rect -572 -2879 -555 -2875
rect -624 -2889 -620 -2886
rect -615 -2886 -602 -2882
rect -615 -2889 -611 -2886
rect -588 -2889 -584 -2886
rect -564 -2889 -560 -2879
rect -548 -2882 -544 -2821
rect -540 -2875 -536 -2821
rect -514 -2844 -510 -2821
rect -540 -2879 -521 -2875
rect -556 -2886 -539 -2882
rect -556 -2889 -552 -2886
rect -532 -2889 -528 -2879
rect -514 -2889 -510 -2848
rect -745 -2897 -741 -2893
rect -719 -2897 -715 -2893
rect -676 -2897 -672 -2893
rect -641 -2897 -637 -2893
rect -597 -2897 -593 -2893
rect -580 -2897 -576 -2893
rect -544 -2897 -540 -2893
rect -523 -2897 -519 -2893
rect -505 -2911 -501 -2857
rect -490 -2860 -486 -2703
rect -476 -2845 -472 -2624
rect -460 -2678 -456 -2391
rect -427 -2417 -423 -2378
rect -427 -2432 -423 -2421
rect -446 -2436 -423 -2432
rect -420 -2408 -416 -2371
rect -446 -2439 -442 -2436
rect -420 -2439 -416 -2412
rect -429 -2447 -425 -2443
rect -437 -2522 -433 -2518
rect -411 -2522 -407 -2518
rect -394 -2522 -390 -2518
rect -354 -2522 -350 -2518
rect -333 -2522 -329 -2518
rect -316 -2522 -312 -2518
rect -276 -2522 -272 -2518
rect -252 -2522 -248 -2518
rect -215 -2522 -211 -2518
rect -446 -2547 -442 -2530
rect -446 -2598 -442 -2551
rect -428 -2540 -424 -2530
rect -428 -2598 -424 -2544
rect -420 -2569 -416 -2530
rect -402 -2562 -398 -2530
rect -420 -2598 -416 -2573
rect -402 -2598 -398 -2566
rect -376 -2554 -372 -2530
rect -376 -2591 -372 -2558
rect -342 -2591 -338 -2530
rect -324 -2547 -320 -2530
rect -394 -2598 -390 -2595
rect -386 -2595 -372 -2591
rect -386 -2598 -382 -2595
rect -358 -2598 -354 -2595
rect -350 -2595 -331 -2591
rect -350 -2598 -346 -2595
rect -324 -2598 -320 -2551
rect -298 -2562 -294 -2530
rect -298 -2591 -294 -2566
rect -264 -2584 -260 -2530
rect -264 -2588 -247 -2584
rect -316 -2598 -312 -2595
rect -307 -2595 -294 -2591
rect -307 -2598 -303 -2595
rect -280 -2598 -276 -2595
rect -256 -2598 -252 -2588
rect -240 -2591 -236 -2530
rect -232 -2584 -228 -2530
rect -206 -2554 -202 -2530
rect -232 -2588 -213 -2584
rect -248 -2595 -231 -2591
rect -248 -2598 -244 -2595
rect -224 -2598 -220 -2588
rect -206 -2598 -202 -2558
rect -437 -2606 -433 -2602
rect -411 -2606 -407 -2602
rect -368 -2606 -364 -2602
rect -333 -2606 -329 -2602
rect -289 -2606 -285 -2602
rect -272 -2606 -268 -2602
rect -236 -2606 -232 -2602
rect -215 -2606 -211 -2602
rect -198 -2613 -194 -2566
rect -180 -2569 -176 -2412
rect -166 -2554 -162 -2326
rect -152 -2387 -148 -2100
rect -119 -2126 -115 -2087
rect -119 -2141 -115 -2130
rect -138 -2145 -115 -2141
rect -112 -2117 -108 -2080
rect -138 -2148 -134 -2145
rect -112 -2148 -108 -2121
rect -121 -2156 -117 -2152
rect -129 -2231 -125 -2227
rect -103 -2231 -99 -2227
rect -86 -2231 -82 -2227
rect -46 -2231 -42 -2227
rect -25 -2231 -21 -2227
rect -8 -2231 -4 -2227
rect 32 -2231 36 -2227
rect 56 -2231 60 -2227
rect 93 -2231 97 -2227
rect -138 -2256 -134 -2239
rect -138 -2307 -134 -2260
rect -120 -2249 -116 -2239
rect -120 -2307 -116 -2253
rect -112 -2278 -108 -2239
rect -94 -2271 -90 -2239
rect -112 -2307 -108 -2282
rect -94 -2307 -90 -2275
rect -68 -2263 -64 -2239
rect -68 -2300 -64 -2267
rect -34 -2300 -30 -2239
rect -16 -2256 -12 -2239
rect -86 -2307 -82 -2304
rect -78 -2304 -64 -2300
rect -78 -2307 -74 -2304
rect -50 -2307 -46 -2304
rect -42 -2304 -23 -2300
rect -42 -2307 -38 -2304
rect -16 -2307 -12 -2260
rect 10 -2271 14 -2239
rect 10 -2300 14 -2275
rect 44 -2293 48 -2239
rect 44 -2297 61 -2293
rect -8 -2307 -4 -2304
rect 1 -2304 14 -2300
rect 1 -2307 5 -2304
rect 28 -2307 32 -2304
rect 52 -2307 56 -2297
rect 68 -2300 72 -2239
rect 76 -2293 80 -2239
rect 102 -2263 106 -2239
rect 76 -2297 95 -2293
rect 60 -2304 77 -2300
rect 60 -2307 64 -2304
rect 84 -2307 88 -2297
rect 102 -2307 106 -2267
rect -129 -2315 -125 -2311
rect -103 -2315 -99 -2311
rect -60 -2315 -56 -2311
rect -25 -2315 -21 -2311
rect 19 -2315 23 -2311
rect 36 -2315 40 -2311
rect 72 -2315 76 -2311
rect 93 -2315 97 -2311
rect 111 -2329 115 -2275
rect 126 -2278 130 -2121
rect 140 -2263 144 -2011
rect 156 -2096 160 -1778
rect 189 -1804 193 -1765
rect 189 -1819 193 -1808
rect 170 -1823 193 -1819
rect 196 -1795 200 -1758
rect 170 -1826 174 -1823
rect 196 -1826 200 -1799
rect 187 -1834 191 -1830
rect 179 -1909 183 -1905
rect 205 -1909 209 -1905
rect 222 -1909 226 -1905
rect 262 -1909 266 -1905
rect 283 -1909 287 -1905
rect 300 -1909 304 -1905
rect 340 -1909 344 -1905
rect 364 -1909 368 -1905
rect 401 -1909 405 -1905
rect 170 -1934 174 -1917
rect 170 -1985 174 -1938
rect 188 -1927 192 -1917
rect 188 -1985 192 -1931
rect 196 -1956 200 -1917
rect 214 -1949 218 -1917
rect 196 -1985 200 -1960
rect 214 -1985 218 -1953
rect 240 -1941 244 -1917
rect 240 -1978 244 -1945
rect 274 -1978 278 -1917
rect 292 -1934 296 -1917
rect 222 -1985 226 -1982
rect 230 -1982 244 -1978
rect 230 -1985 234 -1982
rect 258 -1985 262 -1982
rect 266 -1982 285 -1978
rect 266 -1985 270 -1982
rect 292 -1985 296 -1938
rect 318 -1949 322 -1917
rect 318 -1978 322 -1953
rect 352 -1971 356 -1917
rect 352 -1975 369 -1971
rect 300 -1985 304 -1982
rect 309 -1982 322 -1978
rect 309 -1985 313 -1982
rect 336 -1985 340 -1982
rect 360 -1985 364 -1975
rect 376 -1978 380 -1917
rect 384 -1971 388 -1917
rect 410 -1941 414 -1917
rect 384 -1975 403 -1971
rect 368 -1982 385 -1978
rect 368 -1985 372 -1982
rect 392 -1985 396 -1975
rect 410 -1985 414 -1945
rect 179 -1993 183 -1989
rect 205 -1993 209 -1989
rect 248 -1993 252 -1989
rect 283 -1993 287 -1989
rect 327 -1993 331 -1989
rect 344 -1993 348 -1989
rect 380 -1993 384 -1989
rect 401 -1993 405 -1989
rect 417 -2000 421 -1953
rect 435 -1956 439 -1799
rect 449 -1941 453 -1713
rect 464 -1774 468 -1487
rect 497 -1513 501 -1474
rect 497 -1528 501 -1517
rect 478 -1532 501 -1528
rect 504 -1504 508 -1467
rect 478 -1535 482 -1532
rect 504 -1535 508 -1508
rect 495 -1543 499 -1539
rect 487 -1618 491 -1614
rect 513 -1618 517 -1614
rect 530 -1618 534 -1614
rect 570 -1618 574 -1614
rect 591 -1618 595 -1614
rect 608 -1618 612 -1614
rect 648 -1618 652 -1614
rect 672 -1618 676 -1614
rect 709 -1618 713 -1614
rect 478 -1643 482 -1626
rect 478 -1694 482 -1647
rect 496 -1636 500 -1626
rect 496 -1694 500 -1640
rect 504 -1665 508 -1626
rect 522 -1658 526 -1626
rect 504 -1694 508 -1669
rect 522 -1694 526 -1662
rect 548 -1650 552 -1626
rect 548 -1687 552 -1654
rect 582 -1687 586 -1626
rect 600 -1643 604 -1626
rect 530 -1694 534 -1691
rect 538 -1691 552 -1687
rect 538 -1694 542 -1691
rect 566 -1694 570 -1691
rect 574 -1691 593 -1687
rect 574 -1694 578 -1691
rect 600 -1694 604 -1647
rect 626 -1658 630 -1626
rect 626 -1687 630 -1662
rect 660 -1680 664 -1626
rect 660 -1684 677 -1680
rect 608 -1694 612 -1691
rect 617 -1691 630 -1687
rect 617 -1694 621 -1691
rect 644 -1694 648 -1691
rect 668 -1694 672 -1684
rect 684 -1687 688 -1626
rect 692 -1680 696 -1626
rect 718 -1648 722 -1626
rect 718 -1666 722 -1652
rect 742 -1650 746 -1508
rect 692 -1684 711 -1680
rect 676 -1691 693 -1687
rect 676 -1694 680 -1691
rect 700 -1694 704 -1684
rect 718 -1694 722 -1670
rect 487 -1702 491 -1698
rect 513 -1702 517 -1698
rect 556 -1702 560 -1698
rect 591 -1702 595 -1698
rect 635 -1702 639 -1698
rect 652 -1702 656 -1698
rect 688 -1702 692 -1698
rect 709 -1702 713 -1698
rect 726 -1716 730 -1662
rect 759 -1665 763 -1404
rect 772 -1483 776 -1166
rect 805 -1192 809 -1153
rect 805 -1207 809 -1196
rect 786 -1211 809 -1207
rect 812 -1183 816 -1146
rect 786 -1214 790 -1211
rect 812 -1214 816 -1187
rect 803 -1222 807 -1218
rect 793 -1302 797 -1298
rect 810 -1302 814 -1298
rect 850 -1302 854 -1298
rect 871 -1302 875 -1298
rect 784 -1343 788 -1310
rect 784 -1378 788 -1347
rect 802 -1337 806 -1310
rect 802 -1341 811 -1337
rect 802 -1378 806 -1341
rect 828 -1364 832 -1310
rect 828 -1371 832 -1368
rect 862 -1371 866 -1310
rect 880 -1342 884 -1310
rect 884 -1346 908 -1342
rect 810 -1378 814 -1375
rect 819 -1375 832 -1371
rect 819 -1378 823 -1375
rect 846 -1378 850 -1375
rect 854 -1375 873 -1371
rect 854 -1378 858 -1375
rect 880 -1378 884 -1346
rect 793 -1386 797 -1382
rect 837 -1386 841 -1382
rect 871 -1386 875 -1382
rect 897 -1407 901 -1368
rect 904 -1400 908 -1346
rect 786 -1459 790 -1455
rect 803 -1459 807 -1455
rect 794 -1470 798 -1467
rect 794 -1474 809 -1470
rect 772 -1487 787 -1483
rect 478 -1750 482 -1746
rect 495 -1750 499 -1746
rect 486 -1761 490 -1758
rect 486 -1765 501 -1761
rect 464 -1778 479 -1774
rect 170 -2072 174 -2068
rect 187 -2072 191 -2068
rect 178 -2083 182 -2080
rect 178 -2087 193 -2083
rect 156 -2100 171 -2096
rect -138 -2363 -134 -2359
rect -121 -2363 -117 -2359
rect -130 -2374 -126 -2371
rect -130 -2378 -115 -2374
rect -152 -2391 -137 -2387
rect -446 -2654 -442 -2650
rect -429 -2654 -425 -2650
rect -438 -2665 -434 -2662
rect -438 -2669 -423 -2665
rect -460 -2682 -445 -2678
rect -754 -2945 -750 -2941
rect -737 -2945 -733 -2941
rect -746 -2956 -742 -2953
rect -746 -2960 -731 -2956
rect -768 -2973 -753 -2969
rect -735 -2999 -731 -2960
rect -735 -3014 -731 -3003
rect -754 -3018 -731 -3014
rect -728 -2990 -724 -2953
rect -754 -3021 -750 -3018
rect -728 -3021 -724 -2994
rect -737 -3029 -733 -3025
rect -745 -3104 -741 -3100
rect -719 -3104 -715 -3100
rect -702 -3104 -698 -3100
rect -662 -3104 -658 -3100
rect -641 -3104 -637 -3100
rect -624 -3104 -620 -3100
rect -584 -3104 -580 -3100
rect -560 -3104 -556 -3100
rect -523 -3104 -519 -3100
rect -754 -3129 -750 -3112
rect -754 -3180 -750 -3133
rect -736 -3122 -732 -3112
rect -736 -3180 -732 -3126
rect -728 -3151 -724 -3112
rect -710 -3144 -706 -3112
rect -728 -3180 -724 -3155
rect -710 -3180 -706 -3148
rect -684 -3136 -680 -3112
rect -684 -3173 -680 -3140
rect -650 -3173 -646 -3112
rect -632 -3129 -628 -3112
rect -702 -3180 -698 -3177
rect -694 -3177 -680 -3173
rect -694 -3180 -690 -3177
rect -666 -3180 -662 -3177
rect -658 -3177 -639 -3173
rect -658 -3180 -654 -3177
rect -632 -3180 -628 -3133
rect -606 -3144 -602 -3112
rect -606 -3173 -602 -3148
rect -572 -3166 -568 -3112
rect -572 -3170 -555 -3166
rect -624 -3180 -620 -3177
rect -615 -3177 -602 -3173
rect -615 -3180 -611 -3177
rect -588 -3180 -584 -3177
rect -564 -3180 -560 -3170
rect -548 -3173 -544 -3112
rect -540 -3166 -536 -3112
rect -514 -3135 -510 -3112
rect -540 -3170 -521 -3166
rect -556 -3177 -539 -3173
rect -556 -3180 -552 -3177
rect -532 -3180 -528 -3170
rect -514 -3180 -510 -3139
rect -490 -3151 -486 -2994
rect -476 -3136 -472 -2915
rect -460 -2969 -456 -2682
rect -427 -2708 -423 -2669
rect -427 -2723 -423 -2712
rect -446 -2727 -423 -2723
rect -420 -2699 -416 -2662
rect -446 -2730 -442 -2727
rect -420 -2730 -416 -2703
rect -429 -2738 -425 -2734
rect -437 -2813 -433 -2809
rect -411 -2813 -407 -2809
rect -394 -2813 -390 -2809
rect -354 -2813 -350 -2809
rect -333 -2813 -329 -2809
rect -316 -2813 -312 -2809
rect -276 -2813 -272 -2809
rect -252 -2813 -248 -2809
rect -215 -2813 -211 -2809
rect -446 -2838 -442 -2821
rect -446 -2889 -442 -2842
rect -428 -2831 -424 -2821
rect -428 -2889 -424 -2835
rect -420 -2860 -416 -2821
rect -402 -2853 -398 -2821
rect -420 -2889 -416 -2864
rect -402 -2889 -398 -2857
rect -376 -2845 -372 -2821
rect -376 -2882 -372 -2849
rect -342 -2882 -338 -2821
rect -324 -2838 -320 -2821
rect -394 -2889 -390 -2886
rect -386 -2886 -372 -2882
rect -386 -2889 -382 -2886
rect -358 -2889 -354 -2886
rect -350 -2886 -331 -2882
rect -350 -2889 -346 -2886
rect -324 -2889 -320 -2842
rect -298 -2853 -294 -2821
rect -298 -2882 -294 -2857
rect -264 -2875 -260 -2821
rect -264 -2879 -247 -2875
rect -316 -2889 -312 -2886
rect -307 -2886 -294 -2882
rect -307 -2889 -303 -2886
rect -280 -2889 -276 -2886
rect -256 -2889 -252 -2879
rect -240 -2882 -236 -2821
rect -232 -2875 -228 -2821
rect -206 -2845 -202 -2821
rect -232 -2879 -213 -2875
rect -248 -2886 -231 -2882
rect -248 -2889 -244 -2886
rect -224 -2889 -220 -2879
rect -206 -2889 -202 -2849
rect -437 -2897 -433 -2893
rect -411 -2897 -407 -2893
rect -368 -2897 -364 -2893
rect -333 -2897 -329 -2893
rect -289 -2897 -285 -2893
rect -272 -2897 -268 -2893
rect -236 -2897 -232 -2893
rect -215 -2897 -211 -2893
rect -198 -2904 -194 -2857
rect -180 -2860 -176 -2703
rect -166 -2845 -162 -2617
rect -152 -2678 -148 -2391
rect -119 -2417 -115 -2378
rect -119 -2432 -115 -2421
rect -138 -2436 -115 -2432
rect -112 -2408 -108 -2371
rect -138 -2439 -134 -2436
rect -112 -2439 -108 -2412
rect -121 -2447 -117 -2443
rect -129 -2522 -125 -2518
rect -103 -2522 -99 -2518
rect -86 -2522 -82 -2518
rect -46 -2522 -42 -2518
rect -25 -2522 -21 -2518
rect -8 -2522 -4 -2518
rect 32 -2522 36 -2518
rect 56 -2522 60 -2518
rect 93 -2522 97 -2518
rect -138 -2547 -134 -2530
rect -138 -2598 -134 -2551
rect -120 -2540 -116 -2530
rect -120 -2598 -116 -2544
rect -112 -2569 -108 -2530
rect -94 -2562 -90 -2530
rect -112 -2598 -108 -2573
rect -94 -2598 -90 -2566
rect -68 -2554 -64 -2530
rect -68 -2591 -64 -2558
rect -34 -2591 -30 -2530
rect -16 -2547 -12 -2530
rect -86 -2598 -82 -2595
rect -78 -2595 -64 -2591
rect -78 -2598 -74 -2595
rect -50 -2598 -46 -2595
rect -42 -2595 -23 -2591
rect -42 -2598 -38 -2595
rect -16 -2598 -12 -2551
rect 10 -2562 14 -2530
rect 10 -2591 14 -2566
rect 44 -2584 48 -2530
rect 44 -2588 61 -2584
rect -8 -2598 -4 -2595
rect 1 -2595 14 -2591
rect 1 -2598 5 -2595
rect 28 -2598 32 -2595
rect 52 -2598 56 -2588
rect 68 -2591 72 -2530
rect 76 -2584 80 -2530
rect 102 -2554 106 -2530
rect 76 -2588 95 -2584
rect 60 -2595 77 -2591
rect 60 -2598 64 -2595
rect 84 -2598 88 -2588
rect 102 -2598 106 -2558
rect -129 -2606 -125 -2602
rect -103 -2606 -99 -2602
rect -60 -2606 -56 -2602
rect -25 -2606 -21 -2602
rect 19 -2606 23 -2602
rect 36 -2606 40 -2602
rect 72 -2606 76 -2602
rect 93 -2606 97 -2602
rect 111 -2620 115 -2566
rect 126 -2569 130 -2412
rect 140 -2554 144 -2333
rect 156 -2387 160 -2100
rect 189 -2126 193 -2087
rect 189 -2141 193 -2130
rect 170 -2145 193 -2141
rect 196 -2117 200 -2080
rect 170 -2148 174 -2145
rect 196 -2148 200 -2121
rect 187 -2156 191 -2152
rect 434 -2223 438 -2121
rect 448 -2223 452 -2004
rect 464 -2096 468 -1778
rect 497 -1804 501 -1765
rect 497 -1819 501 -1808
rect 478 -1823 501 -1819
rect 504 -1795 508 -1758
rect 478 -1826 482 -1823
rect 504 -1826 508 -1799
rect 495 -1834 499 -1830
rect 487 -1909 491 -1905
rect 513 -1909 517 -1905
rect 530 -1909 534 -1905
rect 570 -1909 574 -1905
rect 591 -1909 595 -1905
rect 608 -1909 612 -1905
rect 648 -1909 652 -1905
rect 672 -1909 676 -1905
rect 709 -1909 713 -1905
rect 478 -1934 482 -1917
rect 478 -1985 482 -1938
rect 496 -1927 500 -1917
rect 496 -1985 500 -1931
rect 504 -1956 508 -1917
rect 522 -1949 526 -1917
rect 504 -1985 508 -1960
rect 522 -1985 526 -1953
rect 548 -1941 552 -1917
rect 548 -1978 552 -1945
rect 582 -1978 586 -1917
rect 600 -1934 604 -1917
rect 530 -1985 534 -1982
rect 538 -1982 552 -1978
rect 538 -1985 542 -1982
rect 566 -1985 570 -1982
rect 574 -1982 593 -1978
rect 574 -1985 578 -1982
rect 600 -1985 604 -1938
rect 626 -1949 630 -1917
rect 626 -1978 630 -1953
rect 660 -1971 664 -1917
rect 660 -1975 677 -1971
rect 608 -1985 612 -1982
rect 617 -1982 630 -1978
rect 617 -1985 621 -1982
rect 644 -1985 648 -1982
rect 668 -1985 672 -1975
rect 684 -1978 688 -1917
rect 692 -1971 696 -1917
rect 718 -1939 722 -1917
rect 718 -1957 722 -1943
rect 742 -1941 746 -1799
rect 692 -1975 711 -1971
rect 676 -1982 693 -1978
rect 676 -1985 680 -1982
rect 700 -1985 704 -1975
rect 718 -1985 722 -1961
rect 487 -1993 491 -1989
rect 513 -1993 517 -1989
rect 556 -1993 560 -1989
rect 591 -1993 595 -1989
rect 635 -1993 639 -1989
rect 652 -1993 656 -1989
rect 688 -1993 692 -1989
rect 709 -1993 713 -1989
rect 728 -2007 732 -1953
rect 759 -1956 763 -1720
rect 772 -1774 776 -1487
rect 805 -1513 809 -1474
rect 805 -1528 809 -1517
rect 786 -1532 809 -1528
rect 812 -1504 816 -1467
rect 786 -1535 790 -1532
rect 812 -1535 816 -1508
rect 803 -1543 807 -1539
rect 795 -1618 799 -1614
rect 821 -1618 825 -1614
rect 838 -1618 842 -1614
rect 878 -1618 882 -1614
rect 899 -1618 903 -1614
rect 916 -1618 920 -1614
rect 956 -1618 960 -1614
rect 980 -1618 984 -1614
rect 1017 -1618 1021 -1614
rect 786 -1643 790 -1626
rect 786 -1694 790 -1647
rect 804 -1636 808 -1626
rect 804 -1694 808 -1640
rect 812 -1665 816 -1626
rect 830 -1658 834 -1626
rect 812 -1694 816 -1669
rect 830 -1694 834 -1662
rect 856 -1650 860 -1626
rect 856 -1687 860 -1654
rect 890 -1687 894 -1626
rect 908 -1643 912 -1626
rect 838 -1694 842 -1691
rect 846 -1691 860 -1687
rect 846 -1694 850 -1691
rect 874 -1694 878 -1691
rect 882 -1691 901 -1687
rect 882 -1694 886 -1691
rect 908 -1694 912 -1647
rect 934 -1658 938 -1626
rect 934 -1687 938 -1662
rect 968 -1680 972 -1626
rect 968 -1684 985 -1680
rect 916 -1694 920 -1691
rect 925 -1691 938 -1687
rect 925 -1694 929 -1691
rect 952 -1694 956 -1691
rect 976 -1694 980 -1684
rect 992 -1687 996 -1626
rect 1000 -1680 1004 -1626
rect 1000 -1684 1019 -1680
rect 984 -1691 1001 -1687
rect 984 -1694 988 -1691
rect 1008 -1694 1012 -1684
rect 1026 -1694 1030 -1626
rect 795 -1702 799 -1698
rect 821 -1702 825 -1698
rect 864 -1702 868 -1698
rect 899 -1702 903 -1698
rect 943 -1702 947 -1698
rect 960 -1702 964 -1698
rect 996 -1702 1000 -1698
rect 1017 -1702 1021 -1698
rect 1026 -1716 1030 -1698
rect 1041 -1709 1045 -1662
rect 786 -1750 790 -1746
rect 803 -1750 807 -1746
rect 794 -1761 798 -1758
rect 794 -1765 809 -1761
rect 772 -1778 787 -1774
rect 478 -2072 482 -2068
rect 495 -2072 499 -2068
rect 486 -2083 490 -2080
rect 486 -2087 501 -2083
rect 464 -2100 479 -2096
rect 179 -2231 183 -2227
rect 205 -2231 209 -2227
rect 222 -2231 226 -2227
rect 262 -2231 266 -2227
rect 283 -2231 287 -2227
rect 300 -2231 304 -2227
rect 340 -2231 344 -2227
rect 364 -2231 368 -2227
rect 401 -2231 405 -2227
rect 170 -2256 174 -2239
rect 170 -2307 174 -2260
rect 188 -2249 192 -2239
rect 188 -2307 192 -2253
rect 196 -2278 200 -2239
rect 214 -2271 218 -2239
rect 196 -2307 200 -2282
rect 214 -2307 218 -2275
rect 240 -2263 244 -2239
rect 240 -2300 244 -2267
rect 274 -2300 278 -2239
rect 292 -2256 296 -2239
rect 222 -2307 226 -2304
rect 230 -2304 244 -2300
rect 230 -2307 234 -2304
rect 258 -2307 262 -2304
rect 266 -2304 285 -2300
rect 266 -2307 270 -2304
rect 292 -2307 296 -2260
rect 318 -2271 322 -2239
rect 318 -2300 322 -2275
rect 352 -2293 356 -2239
rect 352 -2297 369 -2293
rect 300 -2307 304 -2304
rect 309 -2304 322 -2300
rect 309 -2307 313 -2304
rect 336 -2307 340 -2304
rect 360 -2307 364 -2297
rect 376 -2300 380 -2239
rect 384 -2293 388 -2239
rect 410 -2263 414 -2239
rect 384 -2297 403 -2293
rect 368 -2304 385 -2300
rect 368 -2307 372 -2304
rect 392 -2307 396 -2297
rect 410 -2307 414 -2267
rect 179 -2315 183 -2311
rect 205 -2315 209 -2311
rect 248 -2315 252 -2311
rect 283 -2315 287 -2311
rect 327 -2315 331 -2311
rect 344 -2315 348 -2311
rect 380 -2315 384 -2311
rect 401 -2315 405 -2311
rect 418 -2322 422 -2275
rect 435 -2278 439 -2223
rect 449 -2263 453 -2223
rect 170 -2363 174 -2359
rect 187 -2363 191 -2359
rect 178 -2374 182 -2371
rect 178 -2378 193 -2374
rect 156 -2391 171 -2387
rect -138 -2654 -134 -2650
rect -121 -2654 -117 -2650
rect -130 -2665 -126 -2662
rect -130 -2669 -115 -2665
rect -152 -2682 -137 -2678
rect -446 -2945 -442 -2941
rect -429 -2945 -425 -2941
rect -438 -2956 -434 -2953
rect -438 -2960 -423 -2956
rect -460 -2973 -445 -2969
rect -427 -2999 -423 -2960
rect -427 -3014 -423 -3003
rect -446 -3018 -423 -3014
rect -420 -2990 -416 -2953
rect -446 -3021 -442 -3018
rect -420 -3021 -416 -2994
rect -429 -3029 -425 -3025
rect -1053 -3188 -1049 -3184
rect -1027 -3188 -1023 -3184
rect -984 -3188 -980 -3184
rect -949 -3188 -945 -3184
rect -905 -3188 -901 -3184
rect -888 -3188 -884 -3184
rect -852 -3188 -848 -3184
rect -831 -3188 -827 -3184
rect -745 -3188 -741 -3184
rect -719 -3188 -715 -3184
rect -676 -3188 -672 -3184
rect -641 -3188 -637 -3184
rect -597 -3188 -593 -3184
rect -580 -3188 -576 -3184
rect -544 -3188 -540 -3184
rect -523 -3188 -519 -3184
rect -460 -3192 -456 -3096
rect -437 -3104 -433 -3100
rect -411 -3104 -407 -3100
rect -394 -3104 -390 -3100
rect -354 -3104 -350 -3100
rect -333 -3104 -329 -3100
rect -316 -3104 -312 -3100
rect -276 -3104 -272 -3100
rect -252 -3104 -248 -3100
rect -215 -3104 -211 -3100
rect -446 -3129 -442 -3112
rect -446 -3180 -442 -3133
rect -428 -3122 -424 -3112
rect -428 -3180 -424 -3126
rect -420 -3151 -416 -3112
rect -402 -3144 -398 -3112
rect -420 -3180 -416 -3155
rect -402 -3180 -398 -3148
rect -376 -3136 -372 -3112
rect -376 -3173 -372 -3140
rect -342 -3173 -338 -3112
rect -324 -3129 -320 -3112
rect -394 -3180 -390 -3177
rect -386 -3177 -372 -3173
rect -386 -3180 -382 -3177
rect -358 -3180 -354 -3177
rect -350 -3177 -331 -3173
rect -350 -3180 -346 -3177
rect -324 -3180 -320 -3133
rect -298 -3144 -294 -3112
rect -298 -3173 -294 -3148
rect -264 -3166 -260 -3112
rect -264 -3170 -247 -3166
rect -316 -3180 -312 -3177
rect -307 -3177 -294 -3173
rect -307 -3180 -303 -3177
rect -280 -3180 -276 -3177
rect -256 -3180 -252 -3170
rect -240 -3173 -236 -3112
rect -232 -3166 -228 -3112
rect -206 -3136 -202 -3112
rect -232 -3170 -213 -3166
rect -248 -3177 -231 -3173
rect -248 -3180 -244 -3177
rect -224 -3180 -220 -3170
rect -206 -3180 -202 -3140
rect -180 -3151 -176 -2994
rect -169 -3136 -165 -2908
rect -152 -2969 -148 -2682
rect -119 -2708 -115 -2669
rect -119 -2723 -115 -2712
rect -138 -2727 -115 -2723
rect -112 -2699 -108 -2662
rect -138 -2730 -134 -2727
rect -112 -2730 -108 -2703
rect -121 -2738 -117 -2734
rect -129 -2813 -125 -2809
rect -103 -2813 -99 -2809
rect -86 -2813 -82 -2809
rect -46 -2813 -42 -2809
rect -25 -2813 -21 -2809
rect -8 -2813 -4 -2809
rect 32 -2813 36 -2809
rect 56 -2813 60 -2809
rect 93 -2813 97 -2809
rect -138 -2838 -134 -2821
rect -138 -2889 -134 -2842
rect -120 -2831 -116 -2821
rect -120 -2889 -116 -2835
rect -112 -2860 -108 -2821
rect -94 -2853 -90 -2821
rect -112 -2889 -108 -2864
rect -94 -2889 -90 -2857
rect -68 -2845 -64 -2821
rect -68 -2882 -64 -2849
rect -34 -2882 -30 -2821
rect -16 -2838 -12 -2821
rect -86 -2889 -82 -2886
rect -78 -2886 -64 -2882
rect -78 -2889 -74 -2886
rect -50 -2889 -46 -2886
rect -42 -2886 -23 -2882
rect -42 -2889 -38 -2886
rect -16 -2889 -12 -2842
rect 10 -2853 14 -2821
rect 10 -2882 14 -2857
rect 44 -2875 48 -2821
rect 44 -2879 61 -2875
rect -8 -2889 -4 -2886
rect 1 -2886 14 -2882
rect 1 -2889 5 -2886
rect 28 -2889 32 -2886
rect 52 -2889 56 -2879
rect 68 -2882 72 -2821
rect 76 -2875 80 -2821
rect 102 -2845 106 -2821
rect 76 -2879 95 -2875
rect 60 -2886 77 -2882
rect 60 -2889 64 -2886
rect 84 -2889 88 -2879
rect 102 -2889 106 -2849
rect -129 -2897 -125 -2893
rect -103 -2897 -99 -2893
rect -60 -2897 -56 -2893
rect -25 -2897 -21 -2893
rect 19 -2897 23 -2893
rect 36 -2897 40 -2893
rect 72 -2897 76 -2893
rect 93 -2897 97 -2893
rect 111 -2911 115 -2857
rect 126 -2860 130 -2703
rect 140 -2845 144 -2624
rect 156 -2678 160 -2391
rect 189 -2417 193 -2378
rect 189 -2432 193 -2421
rect 170 -2436 193 -2432
rect 196 -2408 200 -2371
rect 170 -2439 174 -2436
rect 196 -2439 200 -2412
rect 187 -2447 191 -2443
rect 179 -2522 183 -2518
rect 205 -2522 209 -2518
rect 222 -2522 226 -2518
rect 262 -2522 266 -2518
rect 283 -2522 287 -2518
rect 300 -2522 304 -2518
rect 340 -2522 344 -2518
rect 364 -2522 368 -2518
rect 401 -2522 405 -2518
rect 170 -2547 174 -2530
rect 170 -2598 174 -2551
rect 188 -2540 192 -2530
rect 188 -2598 192 -2544
rect 196 -2569 200 -2530
rect 214 -2562 218 -2530
rect 196 -2598 200 -2573
rect 214 -2598 218 -2566
rect 240 -2554 244 -2530
rect 240 -2591 244 -2558
rect 274 -2591 278 -2530
rect 292 -2547 296 -2530
rect 222 -2598 226 -2595
rect 230 -2595 244 -2591
rect 230 -2598 234 -2595
rect 258 -2598 262 -2595
rect 266 -2595 285 -2591
rect 266 -2598 270 -2595
rect 292 -2598 296 -2551
rect 318 -2562 322 -2530
rect 318 -2591 322 -2566
rect 352 -2584 356 -2530
rect 352 -2588 369 -2584
rect 300 -2598 304 -2595
rect 309 -2595 322 -2591
rect 309 -2598 313 -2595
rect 336 -2598 340 -2595
rect 360 -2598 364 -2588
rect 376 -2591 380 -2530
rect 384 -2584 388 -2530
rect 410 -2554 414 -2530
rect 384 -2588 403 -2584
rect 368 -2595 385 -2591
rect 368 -2598 372 -2595
rect 392 -2598 396 -2588
rect 410 -2598 414 -2558
rect 179 -2606 183 -2602
rect 205 -2606 209 -2602
rect 248 -2606 252 -2602
rect 283 -2606 287 -2602
rect 327 -2606 331 -2602
rect 344 -2606 348 -2602
rect 380 -2606 384 -2602
rect 401 -2606 405 -2602
rect 418 -2613 422 -2566
rect 435 -2569 439 -2412
rect 449 -2554 453 -2326
rect 464 -2387 468 -2100
rect 497 -2126 501 -2087
rect 497 -2141 501 -2130
rect 478 -2145 501 -2141
rect 504 -2117 508 -2080
rect 478 -2148 482 -2145
rect 504 -2148 508 -2121
rect 495 -2156 499 -2152
rect 487 -2231 491 -2227
rect 513 -2231 517 -2227
rect 530 -2231 534 -2227
rect 570 -2231 574 -2227
rect 591 -2231 595 -2227
rect 608 -2231 612 -2227
rect 648 -2231 652 -2227
rect 672 -2231 676 -2227
rect 709 -2231 713 -2227
rect 478 -2256 482 -2239
rect 478 -2307 482 -2260
rect 496 -2249 500 -2239
rect 496 -2307 500 -2253
rect 504 -2278 508 -2239
rect 522 -2271 526 -2239
rect 504 -2307 508 -2282
rect 522 -2307 526 -2275
rect 548 -2263 552 -2239
rect 548 -2300 552 -2267
rect 582 -2300 586 -2239
rect 600 -2256 604 -2239
rect 530 -2307 534 -2304
rect 538 -2304 552 -2300
rect 538 -2307 542 -2304
rect 566 -2307 570 -2304
rect 574 -2304 593 -2300
rect 574 -2307 578 -2304
rect 600 -2307 604 -2260
rect 626 -2271 630 -2239
rect 626 -2300 630 -2275
rect 660 -2293 664 -2239
rect 660 -2297 677 -2293
rect 608 -2307 612 -2304
rect 617 -2304 630 -2300
rect 617 -2307 621 -2304
rect 644 -2307 648 -2304
rect 668 -2307 672 -2297
rect 684 -2300 688 -2239
rect 692 -2293 696 -2239
rect 718 -2261 722 -2239
rect 692 -2297 711 -2293
rect 676 -2304 693 -2300
rect 676 -2307 680 -2304
rect 700 -2307 704 -2297
rect 718 -2307 722 -2265
rect 742 -2263 746 -2121
rect 487 -2315 491 -2311
rect 513 -2315 517 -2311
rect 556 -2315 560 -2311
rect 591 -2315 595 -2311
rect 635 -2315 639 -2311
rect 652 -2315 656 -2311
rect 688 -2315 692 -2311
rect 709 -2315 713 -2311
rect 726 -2329 730 -2275
rect 759 -2278 763 -2011
rect 772 -2096 776 -1778
rect 805 -1804 809 -1765
rect 805 -1819 809 -1808
rect 786 -1823 809 -1819
rect 812 -1795 816 -1758
rect 786 -1826 790 -1823
rect 812 -1826 816 -1799
rect 803 -1834 807 -1830
rect 795 -1909 799 -1905
rect 821 -1909 825 -1905
rect 838 -1909 842 -1905
rect 878 -1909 882 -1905
rect 899 -1909 903 -1905
rect 916 -1909 920 -1905
rect 956 -1909 960 -1905
rect 980 -1909 984 -1905
rect 1017 -1909 1021 -1905
rect 786 -1934 790 -1917
rect 786 -1985 790 -1938
rect 804 -1927 808 -1917
rect 804 -1985 808 -1931
rect 812 -1956 816 -1917
rect 830 -1949 834 -1917
rect 812 -1985 816 -1960
rect 830 -1985 834 -1953
rect 856 -1941 860 -1917
rect 856 -1978 860 -1945
rect 890 -1978 894 -1917
rect 908 -1934 912 -1917
rect 838 -1985 842 -1982
rect 846 -1982 860 -1978
rect 846 -1985 850 -1982
rect 874 -1985 878 -1982
rect 882 -1982 901 -1978
rect 882 -1985 886 -1982
rect 908 -1985 912 -1938
rect 934 -1949 938 -1917
rect 934 -1978 938 -1953
rect 968 -1971 972 -1917
rect 968 -1975 985 -1971
rect 916 -1985 920 -1982
rect 925 -1982 938 -1978
rect 925 -1985 929 -1982
rect 952 -1985 956 -1982
rect 976 -1985 980 -1975
rect 992 -1978 996 -1917
rect 1000 -1971 1004 -1917
rect 1000 -1975 1019 -1971
rect 984 -1982 1001 -1978
rect 984 -1985 988 -1982
rect 1008 -1985 1012 -1975
rect 1026 -1985 1030 -1917
rect 795 -1993 799 -1989
rect 821 -1993 825 -1989
rect 864 -1993 868 -1989
rect 899 -1993 903 -1989
rect 943 -1993 947 -1989
rect 960 -1993 964 -1989
rect 996 -1993 1000 -1989
rect 1017 -1993 1021 -1989
rect 1026 -2007 1030 -1989
rect 1042 -2000 1046 -1953
rect 786 -2072 790 -2068
rect 803 -2072 807 -2068
rect 794 -2083 798 -2080
rect 794 -2087 809 -2083
rect 772 -2100 787 -2096
rect 478 -2363 482 -2359
rect 495 -2363 499 -2359
rect 486 -2374 490 -2371
rect 486 -2378 501 -2374
rect 464 -2391 479 -2387
rect 170 -2654 174 -2650
rect 187 -2654 191 -2650
rect 178 -2665 182 -2662
rect 178 -2669 193 -2665
rect 156 -2682 171 -2678
rect -138 -2945 -134 -2941
rect -121 -2945 -117 -2941
rect -130 -2956 -126 -2953
rect -130 -2960 -115 -2956
rect -152 -2973 -137 -2969
rect -119 -2999 -115 -2960
rect -119 -3014 -115 -3003
rect -138 -3018 -115 -3014
rect -112 -2990 -108 -2953
rect -138 -3021 -134 -3018
rect -112 -3021 -108 -2994
rect -121 -3029 -117 -3025
rect -437 -3188 -433 -3184
rect -411 -3188 -407 -3184
rect -368 -3188 -364 -3184
rect -333 -3188 -329 -3184
rect -289 -3188 -285 -3184
rect -272 -3188 -268 -3184
rect -236 -3188 -232 -3184
rect -215 -3188 -211 -3184
rect -152 -3192 -148 -3096
rect -129 -3104 -125 -3100
rect -103 -3104 -99 -3100
rect -86 -3104 -82 -3100
rect -46 -3104 -42 -3100
rect -25 -3104 -21 -3100
rect -8 -3104 -4 -3100
rect 32 -3104 36 -3100
rect 56 -3104 60 -3100
rect 93 -3104 97 -3100
rect -138 -3129 -134 -3112
rect -138 -3180 -134 -3133
rect -120 -3122 -116 -3112
rect -120 -3180 -116 -3126
rect -112 -3151 -108 -3112
rect -94 -3144 -90 -3112
rect -112 -3180 -108 -3155
rect -94 -3180 -90 -3148
rect -68 -3136 -64 -3112
rect -68 -3173 -64 -3140
rect -34 -3173 -30 -3112
rect -16 -3129 -12 -3112
rect -86 -3180 -82 -3177
rect -78 -3177 -64 -3173
rect -78 -3180 -74 -3177
rect -50 -3180 -46 -3177
rect -42 -3177 -23 -3173
rect -42 -3180 -38 -3177
rect -16 -3180 -12 -3133
rect 10 -3144 14 -3112
rect 10 -3173 14 -3148
rect 44 -3166 48 -3112
rect 44 -3170 61 -3166
rect -8 -3180 -4 -3177
rect 1 -3177 14 -3173
rect 1 -3180 5 -3177
rect 28 -3180 32 -3177
rect 52 -3180 56 -3170
rect 68 -3173 72 -3112
rect 76 -3166 80 -3112
rect 102 -3136 106 -3112
rect 76 -3170 95 -3166
rect 60 -3177 77 -3173
rect 60 -3180 64 -3177
rect 84 -3180 88 -3170
rect 102 -3180 106 -3140
rect 126 -3151 130 -2994
rect 139 -3136 143 -2915
rect 156 -2969 160 -2682
rect 189 -2708 193 -2669
rect 189 -2723 193 -2712
rect 170 -2727 193 -2723
rect 196 -2699 200 -2662
rect 170 -2730 174 -2727
rect 196 -2730 200 -2703
rect 187 -2738 191 -2734
rect 179 -2813 183 -2809
rect 205 -2813 209 -2809
rect 222 -2813 226 -2809
rect 262 -2813 266 -2809
rect 283 -2813 287 -2809
rect 300 -2813 304 -2809
rect 340 -2813 344 -2809
rect 364 -2813 368 -2809
rect 401 -2813 405 -2809
rect 170 -2838 174 -2821
rect 170 -2889 174 -2842
rect 188 -2831 192 -2821
rect 188 -2889 192 -2835
rect 196 -2860 200 -2821
rect 214 -2853 218 -2821
rect 196 -2889 200 -2864
rect 214 -2889 218 -2857
rect 240 -2845 244 -2821
rect 240 -2882 244 -2849
rect 274 -2882 278 -2821
rect 292 -2838 296 -2821
rect 222 -2889 226 -2886
rect 230 -2886 244 -2882
rect 230 -2889 234 -2886
rect 258 -2889 262 -2886
rect 266 -2886 285 -2882
rect 266 -2889 270 -2886
rect 292 -2889 296 -2842
rect 318 -2853 322 -2821
rect 318 -2882 322 -2857
rect 352 -2875 356 -2821
rect 352 -2879 369 -2875
rect 300 -2889 304 -2886
rect 309 -2886 322 -2882
rect 309 -2889 313 -2886
rect 336 -2889 340 -2886
rect 360 -2889 364 -2879
rect 376 -2882 380 -2821
rect 384 -2875 388 -2821
rect 410 -2845 414 -2821
rect 384 -2879 403 -2875
rect 368 -2886 385 -2882
rect 368 -2889 372 -2886
rect 392 -2889 396 -2879
rect 410 -2889 414 -2849
rect 179 -2897 183 -2893
rect 205 -2897 209 -2893
rect 248 -2897 252 -2893
rect 283 -2897 287 -2893
rect 327 -2897 331 -2893
rect 344 -2897 348 -2893
rect 380 -2897 384 -2893
rect 401 -2897 405 -2893
rect 418 -2904 422 -2857
rect 435 -2860 439 -2703
rect 449 -2845 453 -2617
rect 464 -2678 468 -2391
rect 497 -2417 501 -2378
rect 497 -2432 501 -2421
rect 478 -2436 501 -2432
rect 504 -2408 508 -2371
rect 478 -2439 482 -2436
rect 504 -2439 508 -2412
rect 495 -2447 499 -2443
rect 487 -2522 491 -2518
rect 513 -2522 517 -2518
rect 530 -2522 534 -2518
rect 570 -2522 574 -2518
rect 591 -2522 595 -2518
rect 608 -2522 612 -2518
rect 648 -2522 652 -2518
rect 672 -2522 676 -2518
rect 709 -2522 713 -2518
rect 478 -2547 482 -2530
rect 478 -2598 482 -2551
rect 496 -2540 500 -2530
rect 496 -2598 500 -2544
rect 504 -2569 508 -2530
rect 522 -2562 526 -2530
rect 504 -2598 508 -2573
rect 522 -2598 526 -2566
rect 548 -2554 552 -2530
rect 548 -2591 552 -2558
rect 582 -2591 586 -2530
rect 600 -2547 604 -2530
rect 530 -2598 534 -2595
rect 538 -2595 552 -2591
rect 538 -2598 542 -2595
rect 566 -2598 570 -2595
rect 574 -2595 593 -2591
rect 574 -2598 578 -2595
rect 600 -2598 604 -2551
rect 626 -2562 630 -2530
rect 626 -2591 630 -2566
rect 660 -2584 664 -2530
rect 660 -2588 677 -2584
rect 608 -2598 612 -2595
rect 617 -2595 630 -2591
rect 617 -2598 621 -2595
rect 644 -2598 648 -2595
rect 668 -2598 672 -2588
rect 684 -2591 688 -2530
rect 692 -2584 696 -2530
rect 718 -2552 722 -2530
rect 692 -2588 711 -2584
rect 676 -2595 693 -2591
rect 676 -2598 680 -2595
rect 700 -2598 704 -2588
rect 718 -2598 722 -2556
rect 742 -2554 746 -2412
rect 487 -2606 491 -2602
rect 513 -2606 517 -2602
rect 556 -2606 560 -2602
rect 591 -2606 595 -2602
rect 635 -2606 639 -2602
rect 652 -2606 656 -2602
rect 688 -2606 692 -2602
rect 709 -2606 713 -2602
rect 726 -2620 730 -2566
rect 759 -2569 763 -2333
rect 772 -2387 776 -2100
rect 805 -2126 809 -2087
rect 805 -2141 809 -2130
rect 786 -2145 809 -2141
rect 812 -2117 816 -2080
rect 786 -2148 790 -2145
rect 812 -2148 816 -2121
rect 803 -2156 807 -2152
rect 795 -2231 799 -2227
rect 821 -2231 825 -2227
rect 838 -2231 842 -2227
rect 878 -2231 882 -2227
rect 899 -2231 903 -2227
rect 916 -2231 920 -2227
rect 956 -2231 960 -2227
rect 980 -2231 984 -2227
rect 1017 -2231 1021 -2227
rect 786 -2256 790 -2239
rect 786 -2307 790 -2260
rect 804 -2249 808 -2239
rect 804 -2307 808 -2253
rect 812 -2278 816 -2239
rect 830 -2271 834 -2239
rect 812 -2307 816 -2282
rect 830 -2307 834 -2275
rect 856 -2263 860 -2239
rect 856 -2300 860 -2267
rect 890 -2300 894 -2239
rect 908 -2256 912 -2239
rect 838 -2307 842 -2304
rect 846 -2304 860 -2300
rect 846 -2307 850 -2304
rect 874 -2307 878 -2304
rect 882 -2304 901 -2300
rect 882 -2307 886 -2304
rect 908 -2307 912 -2260
rect 934 -2271 938 -2239
rect 934 -2300 938 -2275
rect 968 -2293 972 -2239
rect 968 -2297 985 -2293
rect 916 -2307 920 -2304
rect 925 -2304 938 -2300
rect 925 -2307 929 -2304
rect 952 -2307 956 -2304
rect 976 -2307 980 -2297
rect 992 -2300 996 -2239
rect 1000 -2293 1004 -2239
rect 1000 -2297 1019 -2293
rect 984 -2304 1001 -2300
rect 984 -2307 988 -2304
rect 1008 -2307 1012 -2297
rect 1026 -2307 1030 -2239
rect 795 -2315 799 -2311
rect 821 -2315 825 -2311
rect 864 -2315 868 -2311
rect 899 -2315 903 -2311
rect 943 -2315 947 -2311
rect 960 -2315 964 -2311
rect 996 -2315 1000 -2311
rect 1017 -2315 1021 -2311
rect 1026 -2329 1030 -2311
rect 1039 -2322 1043 -2275
rect 786 -2363 790 -2359
rect 803 -2363 807 -2359
rect 794 -2374 798 -2371
rect 794 -2378 809 -2374
rect 772 -2391 787 -2387
rect 478 -2654 482 -2650
rect 495 -2654 499 -2650
rect 486 -2665 490 -2662
rect 486 -2669 501 -2665
rect 464 -2682 479 -2678
rect 170 -2945 174 -2941
rect 187 -2945 191 -2941
rect 178 -2956 182 -2953
rect 178 -2960 193 -2956
rect 156 -2973 171 -2969
rect 189 -2999 193 -2960
rect 189 -3014 193 -3003
rect 170 -3018 193 -3014
rect 196 -2990 200 -2953
rect 170 -3021 174 -3018
rect 196 -3021 200 -2994
rect 187 -3029 191 -3025
rect 179 -3104 183 -3100
rect 205 -3104 209 -3100
rect 222 -3104 226 -3100
rect 262 -3104 266 -3100
rect 283 -3104 287 -3100
rect 300 -3104 304 -3100
rect 340 -3104 344 -3100
rect 364 -3104 368 -3100
rect 401 -3104 405 -3100
rect 170 -3129 174 -3112
rect 170 -3180 174 -3133
rect 188 -3122 192 -3112
rect 188 -3180 192 -3126
rect 196 -3151 200 -3112
rect 214 -3144 218 -3112
rect 196 -3180 200 -3155
rect 214 -3180 218 -3148
rect 240 -3136 244 -3112
rect 240 -3173 244 -3140
rect 274 -3173 278 -3112
rect 292 -3129 296 -3112
rect 222 -3180 226 -3177
rect 230 -3177 244 -3173
rect 230 -3180 234 -3177
rect 258 -3180 262 -3177
rect 266 -3177 285 -3173
rect 266 -3180 270 -3177
rect 292 -3180 296 -3133
rect 318 -3144 322 -3112
rect 318 -3173 322 -3148
rect 352 -3166 356 -3112
rect 352 -3170 369 -3166
rect 300 -3180 304 -3177
rect 309 -3177 322 -3173
rect 309 -3180 313 -3177
rect 336 -3180 340 -3177
rect 360 -3180 364 -3170
rect 376 -3173 380 -3112
rect 384 -3166 388 -3112
rect 410 -3136 414 -3112
rect 384 -3170 403 -3166
rect 368 -3177 385 -3173
rect 368 -3180 372 -3177
rect 392 -3180 396 -3170
rect 410 -3180 414 -3140
rect 435 -3151 439 -2994
rect 447 -3136 451 -2908
rect 464 -2969 468 -2682
rect 497 -2708 501 -2669
rect 497 -2723 501 -2712
rect 478 -2727 501 -2723
rect 504 -2699 508 -2662
rect 478 -2730 482 -2727
rect 504 -2730 508 -2703
rect 495 -2738 499 -2734
rect 487 -2813 491 -2809
rect 513 -2813 517 -2809
rect 530 -2813 534 -2809
rect 570 -2813 574 -2809
rect 591 -2813 595 -2809
rect 608 -2813 612 -2809
rect 648 -2813 652 -2809
rect 672 -2813 676 -2809
rect 709 -2813 713 -2809
rect 478 -2838 482 -2821
rect 478 -2889 482 -2842
rect 496 -2831 500 -2821
rect 496 -2889 500 -2835
rect 504 -2860 508 -2821
rect 522 -2853 526 -2821
rect 504 -2889 508 -2864
rect 522 -2889 526 -2857
rect 548 -2845 552 -2821
rect 548 -2882 552 -2849
rect 582 -2882 586 -2821
rect 600 -2838 604 -2821
rect 530 -2889 534 -2886
rect 538 -2886 552 -2882
rect 538 -2889 542 -2886
rect 566 -2889 570 -2886
rect 574 -2886 593 -2882
rect 574 -2889 578 -2886
rect 600 -2889 604 -2842
rect 626 -2853 630 -2821
rect 626 -2882 630 -2857
rect 660 -2875 664 -2821
rect 660 -2879 677 -2875
rect 608 -2889 612 -2886
rect 617 -2886 630 -2882
rect 617 -2889 621 -2886
rect 644 -2889 648 -2886
rect 668 -2889 672 -2879
rect 684 -2882 688 -2821
rect 692 -2875 696 -2821
rect 718 -2843 722 -2821
rect 692 -2879 711 -2875
rect 676 -2886 693 -2882
rect 676 -2889 680 -2886
rect 700 -2889 704 -2879
rect 718 -2889 722 -2847
rect 742 -2845 746 -2703
rect 487 -2897 491 -2893
rect 513 -2897 517 -2893
rect 556 -2897 560 -2893
rect 591 -2897 595 -2893
rect 635 -2897 639 -2893
rect 652 -2897 656 -2893
rect 688 -2897 692 -2893
rect 709 -2897 713 -2893
rect 726 -2911 730 -2857
rect 759 -2860 763 -2624
rect 772 -2678 776 -2391
rect 805 -2417 809 -2378
rect 805 -2432 809 -2421
rect 786 -2436 809 -2432
rect 812 -2408 816 -2371
rect 786 -2439 790 -2436
rect 812 -2439 816 -2412
rect 803 -2447 807 -2443
rect 795 -2522 799 -2518
rect 821 -2522 825 -2518
rect 838 -2522 842 -2518
rect 878 -2522 882 -2518
rect 899 -2522 903 -2518
rect 916 -2522 920 -2518
rect 956 -2522 960 -2518
rect 980 -2522 984 -2518
rect 1017 -2522 1021 -2518
rect 786 -2547 790 -2530
rect 786 -2598 790 -2551
rect 804 -2540 808 -2530
rect 804 -2598 808 -2544
rect 812 -2569 816 -2530
rect 830 -2562 834 -2530
rect 812 -2598 816 -2573
rect 830 -2598 834 -2566
rect 856 -2554 860 -2530
rect 856 -2591 860 -2558
rect 890 -2591 894 -2530
rect 908 -2547 912 -2530
rect 838 -2598 842 -2595
rect 846 -2595 860 -2591
rect 846 -2598 850 -2595
rect 874 -2598 878 -2595
rect 882 -2595 901 -2591
rect 882 -2598 886 -2595
rect 908 -2598 912 -2551
rect 934 -2562 938 -2530
rect 934 -2591 938 -2566
rect 968 -2584 972 -2530
rect 968 -2588 985 -2584
rect 916 -2598 920 -2595
rect 925 -2595 938 -2591
rect 925 -2598 929 -2595
rect 952 -2598 956 -2595
rect 976 -2598 980 -2588
rect 992 -2591 996 -2530
rect 1000 -2584 1004 -2530
rect 1000 -2588 1019 -2584
rect 984 -2595 1001 -2591
rect 984 -2598 988 -2595
rect 1008 -2598 1012 -2588
rect 1026 -2598 1030 -2530
rect 795 -2606 799 -2602
rect 821 -2606 825 -2602
rect 864 -2606 868 -2602
rect 899 -2606 903 -2602
rect 943 -2606 947 -2602
rect 960 -2606 964 -2602
rect 996 -2606 1000 -2602
rect 1017 -2606 1021 -2602
rect 1026 -2620 1030 -2602
rect 1039 -2613 1043 -2566
rect 786 -2654 790 -2650
rect 803 -2654 807 -2650
rect 794 -2665 798 -2662
rect 794 -2669 809 -2665
rect 772 -2682 787 -2678
rect 478 -2945 482 -2941
rect 495 -2945 499 -2941
rect 486 -2956 490 -2953
rect 486 -2960 501 -2956
rect 464 -2973 479 -2969
rect 497 -2999 501 -2960
rect 497 -3014 501 -3003
rect 478 -3018 501 -3014
rect 504 -2990 508 -2953
rect 478 -3021 482 -3018
rect 504 -3021 508 -2994
rect 495 -3029 499 -3025
rect 487 -3104 491 -3100
rect 513 -3104 517 -3100
rect 530 -3104 534 -3100
rect 570 -3104 574 -3100
rect 591 -3104 595 -3100
rect 608 -3104 612 -3100
rect 648 -3104 652 -3100
rect 672 -3104 676 -3100
rect 709 -3104 713 -3100
rect 478 -3129 482 -3112
rect 478 -3180 482 -3133
rect 496 -3122 500 -3112
rect 496 -3180 500 -3126
rect 504 -3151 508 -3112
rect 522 -3144 526 -3112
rect 504 -3180 508 -3155
rect 522 -3180 526 -3148
rect 548 -3136 552 -3112
rect 548 -3173 552 -3140
rect 582 -3173 586 -3112
rect 600 -3129 604 -3112
rect 530 -3180 534 -3177
rect 538 -3177 552 -3173
rect 538 -3180 542 -3177
rect 566 -3180 570 -3177
rect 574 -3177 593 -3173
rect 574 -3180 578 -3177
rect 600 -3180 604 -3133
rect 626 -3144 630 -3112
rect 626 -3173 630 -3148
rect 660 -3166 664 -3112
rect 660 -3170 677 -3166
rect 608 -3180 612 -3177
rect 617 -3177 630 -3173
rect 617 -3180 621 -3177
rect 644 -3180 648 -3177
rect 668 -3180 672 -3170
rect 684 -3173 688 -3112
rect 692 -3166 696 -3112
rect 718 -3134 722 -3112
rect 692 -3170 711 -3166
rect 676 -3177 693 -3173
rect 676 -3180 680 -3177
rect 700 -3180 704 -3170
rect 718 -3180 722 -3138
rect 742 -3136 746 -2994
rect 752 -3151 756 -2915
rect 772 -2969 776 -2682
rect 805 -2708 809 -2669
rect 805 -2723 809 -2712
rect 786 -2727 809 -2723
rect 812 -2699 816 -2662
rect 786 -2730 790 -2727
rect 812 -2730 816 -2703
rect 803 -2738 807 -2734
rect 795 -2813 799 -2809
rect 821 -2813 825 -2809
rect 838 -2813 842 -2809
rect 878 -2813 882 -2809
rect 899 -2813 903 -2809
rect 916 -2813 920 -2809
rect 956 -2813 960 -2809
rect 980 -2813 984 -2809
rect 1017 -2813 1021 -2809
rect 786 -2838 790 -2821
rect 786 -2889 790 -2842
rect 804 -2831 808 -2821
rect 804 -2889 808 -2835
rect 812 -2860 816 -2821
rect 830 -2853 834 -2821
rect 812 -2889 816 -2864
rect 830 -2889 834 -2857
rect 856 -2845 860 -2821
rect 856 -2882 860 -2849
rect 890 -2882 894 -2821
rect 908 -2838 912 -2821
rect 838 -2889 842 -2886
rect 846 -2886 860 -2882
rect 846 -2889 850 -2886
rect 874 -2889 878 -2886
rect 882 -2886 901 -2882
rect 882 -2889 886 -2886
rect 908 -2889 912 -2842
rect 934 -2853 938 -2821
rect 934 -2882 938 -2857
rect 968 -2875 972 -2821
rect 968 -2879 985 -2875
rect 916 -2889 920 -2886
rect 925 -2886 938 -2882
rect 925 -2889 929 -2886
rect 952 -2889 956 -2886
rect 976 -2889 980 -2879
rect 992 -2882 996 -2821
rect 1000 -2875 1004 -2821
rect 1000 -2879 1019 -2875
rect 984 -2886 1001 -2882
rect 984 -2889 988 -2886
rect 1008 -2889 1012 -2879
rect 1026 -2889 1030 -2821
rect 795 -2897 799 -2893
rect 821 -2897 825 -2893
rect 864 -2897 868 -2893
rect 899 -2897 903 -2893
rect 943 -2897 947 -2893
rect 960 -2897 964 -2893
rect 996 -2897 1000 -2893
rect 1017 -2897 1021 -2893
rect 1026 -2911 1030 -2893
rect 1039 -2904 1043 -2857
rect 786 -2945 790 -2941
rect 803 -2945 807 -2941
rect 794 -2956 798 -2953
rect 794 -2960 809 -2956
rect 772 -2973 787 -2969
rect 805 -2999 809 -2960
rect 805 -3014 809 -3003
rect 786 -3018 809 -3014
rect 812 -2990 816 -2953
rect 786 -3021 790 -3018
rect 812 -3021 816 -2994
rect 803 -3029 807 -3025
rect 795 -3104 799 -3100
rect 821 -3104 825 -3100
rect 838 -3104 842 -3100
rect 878 -3104 882 -3100
rect 899 -3104 903 -3100
rect 916 -3104 920 -3100
rect 956 -3104 960 -3100
rect 980 -3104 984 -3100
rect 1017 -3104 1021 -3100
rect 786 -3129 790 -3112
rect 786 -3180 790 -3133
rect 804 -3122 808 -3112
rect 804 -3180 808 -3126
rect 812 -3151 816 -3112
rect 830 -3144 834 -3112
rect 812 -3180 816 -3155
rect 830 -3180 834 -3148
rect 856 -3136 860 -3112
rect 856 -3173 860 -3140
rect 890 -3173 894 -3112
rect 908 -3129 912 -3112
rect 838 -3180 842 -3177
rect 846 -3177 860 -3173
rect 846 -3180 850 -3177
rect 874 -3180 878 -3177
rect 882 -3177 901 -3173
rect 882 -3180 886 -3177
rect 908 -3180 912 -3133
rect 934 -3144 938 -3112
rect 934 -3173 938 -3148
rect 968 -3166 972 -3112
rect 968 -3170 985 -3166
rect 916 -3180 920 -3177
rect 925 -3177 938 -3173
rect 925 -3180 929 -3177
rect 952 -3180 956 -3177
rect 976 -3180 980 -3170
rect 992 -3173 996 -3112
rect 1000 -3166 1004 -3112
rect 1026 -3137 1030 -3112
rect 1026 -3141 1034 -3137
rect 1000 -3170 1019 -3166
rect 984 -3177 1001 -3173
rect 984 -3180 988 -3177
rect 1008 -3180 1012 -3170
rect 1026 -3180 1030 -3141
rect -129 -3188 -125 -3184
rect -103 -3188 -99 -3184
rect -60 -3188 -56 -3184
rect -25 -3188 -21 -3184
rect 19 -3188 23 -3184
rect 36 -3188 40 -3184
rect 72 -3188 76 -3184
rect 93 -3188 97 -3184
rect 179 -3188 183 -3184
rect 205 -3188 209 -3184
rect 248 -3188 252 -3184
rect 283 -3188 287 -3184
rect 327 -3188 331 -3184
rect 344 -3188 348 -3184
rect 380 -3188 384 -3184
rect 401 -3188 405 -3184
rect 487 -3188 491 -3184
rect 513 -3188 517 -3184
rect 556 -3188 560 -3184
rect 591 -3188 595 -3184
rect 635 -3188 639 -3184
rect 652 -3188 656 -3184
rect 688 -3188 692 -3184
rect 709 -3188 713 -3184
rect 795 -3188 799 -3184
rect 821 -3188 825 -3184
rect 864 -3188 868 -3184
rect 899 -3188 903 -3184
rect 943 -3188 947 -3184
rect 960 -3188 964 -3184
rect 996 -3188 1000 -3184
rect 1017 -3188 1021 -3184
<< metal2 >>
rect -1454 -984 -1307 -980
rect -1303 -984 -1290 -980
rect -1286 -984 -1063 -980
rect -1059 -984 -1046 -980
rect -1042 -984 -754 -980
rect -750 -984 -737 -980
rect -733 -984 -446 -980
rect -442 -984 -429 -980
rect -425 -984 -139 -980
rect -135 -984 -122 -980
rect -118 -984 170 -980
rect 174 -984 187 -980
rect 191 -984 478 -980
rect 482 -984 495 -980
rect 499 -984 786 -980
rect 790 -984 803 -980
rect 807 -984 1164 -980
rect -1454 -1130 -1427 -984
rect -1411 -1024 -1295 -1020
rect -1291 -1024 -1051 -1020
rect -1047 -1024 -742 -1020
rect -738 -1024 -434 -1020
rect -430 -1024 -127 -1020
rect -123 -1024 182 -1020
rect 186 -1024 490 -1020
rect 494 -1024 798 -1020
rect 802 -1024 1164 -1020
rect -1087 -1032 -728 -1028
rect -467 -1032 -113 -1028
rect 149 -1032 504 -1028
rect -1247 -1040 -1037 -1036
rect -778 -1040 -420 -1036
rect -166 -1040 196 -1036
rect 450 -1040 812 -1036
rect -1411 -1076 -1290 -1072
rect -1286 -1076 -1046 -1072
rect -1042 -1076 -737 -1072
rect -733 -1076 -429 -1072
rect -425 -1076 -122 -1072
rect -118 -1076 187 -1072
rect 191 -1076 495 -1072
rect 499 -1076 803 -1072
rect 807 -1076 1206 -1072
rect -1454 -1134 -1309 -1130
rect -1305 -1134 -1292 -1130
rect -1288 -1134 -1062 -1130
rect -1058 -1134 -1045 -1130
rect -1041 -1134 -754 -1130
rect -750 -1134 -737 -1130
rect -733 -1134 -446 -1130
rect -442 -1134 -429 -1130
rect -425 -1134 -138 -1130
rect -134 -1134 -121 -1130
rect -117 -1134 170 -1130
rect 174 -1134 187 -1130
rect 191 -1134 478 -1130
rect 482 -1134 495 -1130
rect 499 -1134 786 -1130
rect 790 -1134 803 -1130
rect 807 -1134 1164 -1130
rect -1454 -1294 -1427 -1134
rect -1411 -1174 -1297 -1170
rect -1293 -1174 -1050 -1170
rect -1046 -1174 -742 -1170
rect -738 -1174 -434 -1170
rect -430 -1174 -126 -1170
rect -122 -1174 182 -1170
rect 186 -1174 490 -1170
rect 494 -1174 798 -1170
rect 802 -1174 1164 -1170
rect -1099 -1187 -1036 -1183
rect -791 -1187 -728 -1183
rect -490 -1187 -420 -1183
rect -182 -1187 -112 -1183
rect 126 -1187 196 -1183
rect 434 -1187 504 -1183
rect 742 -1187 812 -1183
rect 1179 -1222 1206 -1076
rect -1411 -1226 -1292 -1222
rect -1288 -1226 -1045 -1222
rect -1041 -1226 -737 -1222
rect -733 -1226 -429 -1222
rect -425 -1226 -121 -1222
rect -117 -1226 187 -1222
rect 191 -1226 495 -1222
rect 499 -1226 803 -1222
rect 807 -1226 1206 -1222
rect -1454 -1298 -1221 -1294
rect -1217 -1298 -1204 -1294
rect -1200 -1298 -1164 -1294
rect -1160 -1298 -1143 -1294
rect -1139 -1298 -1053 -1294
rect -1049 -1298 -1027 -1294
rect -1023 -1298 -1010 -1294
rect -1006 -1298 -970 -1294
rect -966 -1298 -949 -1294
rect -945 -1298 -932 -1294
rect -928 -1298 -892 -1294
rect -888 -1298 -868 -1294
rect -864 -1298 -831 -1294
rect -827 -1298 -745 -1294
rect -741 -1298 -719 -1294
rect -715 -1298 -702 -1294
rect -698 -1298 -662 -1294
rect -658 -1298 -641 -1294
rect -637 -1298 -624 -1294
rect -620 -1298 -584 -1294
rect -580 -1298 -560 -1294
rect -556 -1298 -523 -1294
rect -519 -1298 -437 -1294
rect -433 -1298 -411 -1294
rect -407 -1298 -394 -1294
rect -390 -1298 -354 -1294
rect -350 -1298 -333 -1294
rect -329 -1298 -316 -1294
rect -312 -1298 -276 -1294
rect -272 -1298 -252 -1294
rect -248 -1298 -215 -1294
rect -211 -1298 -129 -1294
rect -125 -1298 -103 -1294
rect -99 -1298 -86 -1294
rect -82 -1298 -46 -1294
rect -42 -1298 -25 -1294
rect -21 -1298 -8 -1294
rect -4 -1298 32 -1294
rect 36 -1298 56 -1294
rect 60 -1298 93 -1294
rect 97 -1298 179 -1294
rect 183 -1298 205 -1294
rect 209 -1298 222 -1294
rect 226 -1298 262 -1294
rect 266 -1298 283 -1294
rect 287 -1298 300 -1294
rect 304 -1298 340 -1294
rect 344 -1298 364 -1294
rect 368 -1298 401 -1294
rect 405 -1298 487 -1294
rect 491 -1298 513 -1294
rect 517 -1298 530 -1294
rect 534 -1298 570 -1294
rect 574 -1298 591 -1294
rect 595 -1298 608 -1294
rect 612 -1298 648 -1294
rect 652 -1298 672 -1294
rect 676 -1298 709 -1294
rect 713 -1298 793 -1294
rect 797 -1298 810 -1294
rect 814 -1298 850 -1294
rect 854 -1298 871 -1294
rect 875 -1298 1164 -1294
rect -1454 -1451 -1427 -1298
rect -437 -1302 -433 -1298
rect -411 -1302 -407 -1298
rect -394 -1302 -390 -1298
rect -354 -1302 -350 -1298
rect -333 -1302 -329 -1298
rect -316 -1302 -312 -1298
rect -276 -1302 -272 -1298
rect -252 -1302 -248 -1298
rect -215 -1302 -211 -1298
rect -129 -1302 -125 -1298
rect -103 -1302 -99 -1298
rect -86 -1302 -82 -1298
rect -46 -1302 -42 -1298
rect -25 -1302 -21 -1298
rect -8 -1302 -4 -1298
rect 32 -1302 36 -1298
rect 56 -1302 60 -1298
rect 93 -1302 97 -1298
rect 179 -1302 183 -1298
rect 205 -1302 209 -1298
rect 222 -1302 226 -1298
rect 262 -1302 266 -1298
rect 283 -1302 287 -1298
rect 300 -1302 304 -1298
rect 340 -1302 344 -1298
rect 364 -1302 368 -1298
rect 401 -1302 405 -1298
rect 487 -1302 491 -1298
rect 513 -1302 517 -1298
rect 530 -1302 534 -1298
rect 570 -1302 574 -1298
rect 591 -1302 595 -1298
rect 608 -1302 612 -1298
rect 648 -1302 652 -1298
rect 672 -1302 676 -1298
rect 709 -1302 713 -1298
rect -1047 -1317 -985 -1313
rect -981 -1317 -951 -1313
rect -903 -1317 -873 -1313
rect -739 -1317 -677 -1313
rect -673 -1317 -643 -1313
rect -595 -1317 -565 -1313
rect -431 -1317 -369 -1313
rect -365 -1317 -335 -1313
rect -287 -1317 -257 -1313
rect -123 -1317 -61 -1313
rect -57 -1317 -27 -1313
rect 21 -1317 51 -1313
rect 185 -1317 247 -1313
rect 251 -1317 281 -1313
rect 329 -1317 359 -1313
rect 493 -1317 555 -1313
rect 559 -1317 589 -1313
rect 637 -1317 667 -1313
rect -1040 -1324 -1009 -1320
rect -732 -1324 -701 -1320
rect -424 -1324 -393 -1320
rect -116 -1324 -85 -1320
rect 192 -1324 223 -1320
rect 500 -1324 531 -1320
rect -1058 -1331 -975 -1327
rect -936 -1331 -833 -1327
rect -750 -1331 -667 -1327
rect -628 -1331 -525 -1327
rect -442 -1331 -359 -1327
rect -320 -1331 -217 -1327
rect -134 -1331 -51 -1327
rect -12 -1331 91 -1327
rect 174 -1331 257 -1327
rect 296 -1331 399 -1327
rect 482 -1331 565 -1327
rect 604 -1331 707 -1327
rect -1087 -1338 -1055 -1334
rect -1021 -1338 -992 -1334
rect -988 -1338 -907 -1334
rect -818 -1338 -791 -1334
rect -778 -1338 -747 -1334
rect -713 -1338 -684 -1334
rect -680 -1338 -599 -1334
rect -510 -1338 -490 -1334
rect -467 -1338 -439 -1334
rect -405 -1338 -376 -1334
rect -372 -1338 -291 -1334
rect -202 -1338 -182 -1334
rect -166 -1338 -131 -1334
rect -97 -1338 -68 -1334
rect -64 -1338 17 -1334
rect 106 -1338 126 -1334
rect 149 -1338 177 -1334
rect 211 -1338 240 -1334
rect 244 -1338 325 -1334
rect 414 -1338 434 -1334
rect 450 -1338 485 -1334
rect 519 -1338 548 -1334
rect 552 -1338 633 -1334
rect -795 -1342 -791 -1338
rect -494 -1342 -490 -1338
rect -186 -1342 -182 -1338
rect 122 -1342 126 -1338
rect 430 -1342 434 -1338
rect -1226 -1347 -1169 -1343
rect -1130 -1346 -1029 -1342
rect -1014 -1346 -931 -1342
rect -910 -1346 -815 -1342
rect -795 -1346 -721 -1342
rect -706 -1346 -623 -1342
rect -602 -1346 -505 -1342
rect -494 -1346 -413 -1342
rect -398 -1346 -315 -1342
rect -294 -1346 -198 -1342
rect -186 -1346 -105 -1342
rect -90 -1346 -7 -1342
rect 14 -1346 109 -1342
rect 122 -1346 203 -1342
rect 218 -1346 301 -1342
rect 322 -1346 417 -1342
rect 430 -1346 511 -1342
rect 526 -1346 609 -1342
rect 630 -1346 725 -1342
rect 788 -1347 845 -1343
rect -1247 -1354 -1219 -1350
rect -1215 -1354 -1179 -1350
rect -1175 -1354 -1159 -1350
rect -1099 -1353 -1051 -1349
rect -1032 -1353 -903 -1349
rect -791 -1353 -743 -1349
rect -724 -1353 -595 -1349
rect -490 -1353 -435 -1349
rect -416 -1353 -287 -1349
rect -182 -1353 -127 -1349
rect -108 -1353 21 -1349
rect 126 -1353 181 -1349
rect 200 -1353 329 -1349
rect 434 -1353 489 -1349
rect 508 -1353 637 -1349
rect 722 -1354 795 -1350
rect 799 -1354 835 -1350
rect 839 -1354 855 -1350
rect -1279 -1361 -1223 -1357
rect -1219 -1361 -1193 -1357
rect -1189 -1361 -1145 -1357
rect -1025 -1360 -921 -1356
rect -917 -1360 -887 -1356
rect -717 -1360 -613 -1356
rect -609 -1360 -579 -1356
rect -409 -1360 -305 -1356
rect -301 -1360 -271 -1356
rect -101 -1360 3 -1356
rect 7 -1360 37 -1356
rect 207 -1360 311 -1356
rect 315 -1360 345 -1356
rect 515 -1360 619 -1356
rect 623 -1360 653 -1356
rect 742 -1361 791 -1357
rect 795 -1361 821 -1357
rect 825 -1361 869 -1357
rect -1182 -1368 -1119 -1364
rect -1051 -1367 -999 -1363
rect -995 -1367 -965 -1363
rect -743 -1367 -691 -1363
rect -687 -1367 -657 -1363
rect -435 -1367 -383 -1363
rect -379 -1367 -349 -1363
rect -127 -1367 -75 -1363
rect -71 -1367 -41 -1363
rect 181 -1367 233 -1363
rect 237 -1367 267 -1363
rect 489 -1367 541 -1363
rect 545 -1367 575 -1363
rect 832 -1368 897 -1364
rect -1200 -1375 -1168 -1371
rect -1006 -1375 -974 -1371
rect -928 -1375 -896 -1371
rect -698 -1375 -666 -1371
rect -620 -1375 -588 -1371
rect -390 -1375 -358 -1371
rect -394 -1378 -390 -1375
rect -358 -1378 -354 -1375
rect -312 -1375 -280 -1371
rect -316 -1378 -312 -1375
rect -280 -1378 -276 -1375
rect -82 -1375 -50 -1371
rect -86 -1378 -82 -1375
rect -50 -1378 -46 -1375
rect -4 -1375 28 -1371
rect -8 -1378 -4 -1375
rect 28 -1378 32 -1375
rect 226 -1375 258 -1371
rect 222 -1378 226 -1375
rect 258 -1378 262 -1375
rect 304 -1375 336 -1371
rect 300 -1378 304 -1375
rect 336 -1378 340 -1375
rect 534 -1375 566 -1371
rect 530 -1378 534 -1375
rect 566 -1378 570 -1375
rect 612 -1375 644 -1371
rect 814 -1375 846 -1371
rect 608 -1378 612 -1375
rect 644 -1378 648 -1375
rect -437 -1386 -433 -1382
rect -411 -1386 -407 -1382
rect -368 -1386 -364 -1382
rect -333 -1386 -329 -1382
rect -289 -1386 -285 -1382
rect -272 -1386 -268 -1382
rect -236 -1386 -232 -1382
rect -215 -1386 -211 -1382
rect -129 -1386 -125 -1382
rect -103 -1386 -99 -1382
rect -60 -1386 -56 -1382
rect -25 -1386 -21 -1382
rect 19 -1386 23 -1382
rect 36 -1386 40 -1382
rect 72 -1386 76 -1382
rect 93 -1386 97 -1382
rect 179 -1386 183 -1382
rect 205 -1386 209 -1382
rect 248 -1386 252 -1382
rect 283 -1386 287 -1382
rect 327 -1386 331 -1382
rect 344 -1386 348 -1382
rect 380 -1386 384 -1382
rect 401 -1386 405 -1382
rect 487 -1386 491 -1382
rect 513 -1386 517 -1382
rect 556 -1386 560 -1382
rect 591 -1386 595 -1382
rect 635 -1386 639 -1382
rect 652 -1386 656 -1382
rect 688 -1386 692 -1382
rect 709 -1386 713 -1382
rect 1179 -1386 1206 -1226
rect -1411 -1390 -1221 -1386
rect -1217 -1390 -1177 -1386
rect -1173 -1390 -1143 -1386
rect -1139 -1390 -1053 -1386
rect -1049 -1390 -1027 -1386
rect -1023 -1390 -984 -1386
rect -980 -1390 -949 -1386
rect -945 -1390 -905 -1386
rect -901 -1390 -888 -1386
rect -884 -1390 -852 -1386
rect -848 -1390 -831 -1386
rect -827 -1390 -745 -1386
rect -741 -1390 -719 -1386
rect -715 -1390 -676 -1386
rect -672 -1390 -641 -1386
rect -637 -1390 -597 -1386
rect -593 -1390 -580 -1386
rect -576 -1390 -544 -1386
rect -540 -1390 -523 -1386
rect -519 -1390 -437 -1386
rect -433 -1390 -411 -1386
rect -407 -1390 -368 -1386
rect -364 -1390 -333 -1386
rect -329 -1390 -289 -1386
rect -285 -1390 -272 -1386
rect -268 -1390 -236 -1386
rect -232 -1390 -215 -1386
rect -211 -1390 -129 -1386
rect -125 -1390 -103 -1386
rect -99 -1390 -60 -1386
rect -56 -1390 -25 -1386
rect -21 -1390 19 -1386
rect 23 -1390 36 -1386
rect 40 -1390 72 -1386
rect 76 -1390 93 -1386
rect 97 -1390 179 -1386
rect 183 -1390 205 -1386
rect 209 -1390 248 -1386
rect 252 -1390 283 -1386
rect 287 -1390 327 -1386
rect 331 -1390 344 -1386
rect 348 -1390 380 -1386
rect 384 -1390 401 -1386
rect 405 -1390 487 -1386
rect 491 -1390 513 -1386
rect 517 -1390 556 -1386
rect 560 -1390 591 -1386
rect 595 -1390 635 -1386
rect 639 -1390 652 -1386
rect 656 -1390 688 -1386
rect 692 -1390 709 -1386
rect 713 -1390 793 -1386
rect 797 -1390 837 -1386
rect 841 -1390 871 -1386
rect 875 -1390 1206 -1386
rect -1253 -1397 -815 -1393
rect -1109 -1404 -505 -1400
rect -467 -1404 109 -1400
rect 149 -1404 725 -1400
rect 763 -1404 904 -1400
rect -778 -1411 -198 -1407
rect -166 -1411 417 -1407
rect 452 -1411 897 -1407
rect -1454 -1455 -1309 -1451
rect -1305 -1455 -1292 -1451
rect -1288 -1455 -1062 -1451
rect -1058 -1455 -1045 -1451
rect -1041 -1455 -754 -1451
rect -750 -1455 -737 -1451
rect -733 -1455 -446 -1451
rect -442 -1455 -429 -1451
rect -425 -1455 -138 -1451
rect -134 -1455 -121 -1451
rect -117 -1455 170 -1451
rect 174 -1455 187 -1451
rect 191 -1455 478 -1451
rect 482 -1455 495 -1451
rect 499 -1455 786 -1451
rect 790 -1455 803 -1451
rect 807 -1455 1164 -1451
rect -1454 -1610 -1427 -1455
rect -1411 -1495 -1297 -1491
rect -1293 -1495 -1050 -1491
rect -1046 -1495 -742 -1491
rect -738 -1495 -434 -1491
rect -430 -1495 -126 -1491
rect -122 -1495 182 -1491
rect 186 -1495 490 -1491
rect 494 -1495 798 -1491
rect 802 -1495 1164 -1491
rect -1091 -1508 -1036 -1504
rect -791 -1508 -728 -1504
rect -485 -1508 -420 -1504
rect -180 -1508 -112 -1504
rect 130 -1508 196 -1504
rect 438 -1508 504 -1504
rect 746 -1508 812 -1504
rect 1179 -1543 1206 -1390
rect -1411 -1547 -1292 -1543
rect -1288 -1547 -1045 -1543
rect -1041 -1547 -737 -1543
rect -733 -1547 -429 -1543
rect -425 -1547 -121 -1543
rect -117 -1547 187 -1543
rect 191 -1547 495 -1543
rect 499 -1547 803 -1543
rect 807 -1547 1206 -1543
rect -1454 -1614 -1225 -1610
rect -1221 -1614 -1208 -1610
rect -1204 -1614 -1168 -1610
rect -1164 -1614 -1147 -1610
rect -1143 -1614 -1053 -1610
rect -1049 -1614 -1027 -1610
rect -1023 -1614 -1010 -1610
rect -1006 -1614 -970 -1610
rect -966 -1614 -949 -1610
rect -945 -1614 -932 -1610
rect -928 -1614 -892 -1610
rect -888 -1614 -868 -1610
rect -864 -1614 -831 -1610
rect -827 -1614 -745 -1610
rect -741 -1614 -719 -1610
rect -715 -1614 -702 -1610
rect -698 -1614 -662 -1610
rect -658 -1614 -641 -1610
rect -637 -1614 -624 -1610
rect -620 -1614 -584 -1610
rect -580 -1614 -560 -1610
rect -556 -1614 -523 -1610
rect -519 -1614 -437 -1610
rect -433 -1614 -411 -1610
rect -407 -1614 -394 -1610
rect -390 -1614 -354 -1610
rect -350 -1614 -333 -1610
rect -329 -1614 -316 -1610
rect -312 -1614 -276 -1610
rect -272 -1614 -252 -1610
rect -248 -1614 -215 -1610
rect -211 -1614 -129 -1610
rect -125 -1614 -103 -1610
rect -99 -1614 -86 -1610
rect -82 -1614 -46 -1610
rect -42 -1614 -25 -1610
rect -21 -1614 -8 -1610
rect -4 -1614 32 -1610
rect 36 -1614 56 -1610
rect 60 -1614 93 -1610
rect 97 -1614 179 -1610
rect 183 -1614 205 -1610
rect 209 -1614 222 -1610
rect 226 -1614 262 -1610
rect 266 -1614 283 -1610
rect 287 -1614 300 -1610
rect 304 -1614 340 -1610
rect 344 -1614 364 -1610
rect 368 -1614 401 -1610
rect 405 -1614 487 -1610
rect 491 -1614 513 -1610
rect 517 -1614 530 -1610
rect 534 -1614 570 -1610
rect 574 -1614 591 -1610
rect 595 -1614 608 -1610
rect 612 -1614 648 -1610
rect 652 -1614 672 -1610
rect 676 -1614 709 -1610
rect 713 -1614 795 -1610
rect 799 -1614 821 -1610
rect 825 -1614 838 -1610
rect 842 -1614 878 -1610
rect 882 -1614 899 -1610
rect 903 -1614 916 -1610
rect 920 -1614 956 -1610
rect 960 -1614 980 -1610
rect 984 -1614 1017 -1610
rect 1021 -1614 1164 -1610
rect -1454 -1742 -1427 -1614
rect -1053 -1618 -1049 -1614
rect -1027 -1618 -1023 -1614
rect -1010 -1618 -1006 -1614
rect -970 -1618 -966 -1614
rect -949 -1618 -945 -1614
rect -932 -1618 -928 -1614
rect -892 -1618 -888 -1614
rect -868 -1618 -864 -1614
rect -831 -1618 -827 -1614
rect -745 -1618 -741 -1614
rect -719 -1618 -715 -1614
rect -702 -1618 -698 -1614
rect -662 -1618 -658 -1614
rect -641 -1618 -637 -1614
rect -624 -1618 -620 -1614
rect -584 -1618 -580 -1614
rect -560 -1618 -556 -1614
rect -523 -1618 -519 -1614
rect -437 -1618 -433 -1614
rect -411 -1618 -407 -1614
rect -394 -1618 -390 -1614
rect -354 -1618 -350 -1614
rect -333 -1618 -329 -1614
rect -316 -1618 -312 -1614
rect -276 -1618 -272 -1614
rect -252 -1618 -248 -1614
rect -215 -1618 -211 -1614
rect -129 -1618 -125 -1614
rect -103 -1618 -99 -1614
rect -86 -1618 -82 -1614
rect -46 -1618 -42 -1614
rect -25 -1618 -21 -1614
rect -8 -1618 -4 -1614
rect 32 -1618 36 -1614
rect 56 -1618 60 -1614
rect 93 -1618 97 -1614
rect 179 -1618 183 -1614
rect 205 -1618 209 -1614
rect 222 -1618 226 -1614
rect 262 -1618 266 -1614
rect 283 -1618 287 -1614
rect 300 -1618 304 -1614
rect 340 -1618 344 -1614
rect 364 -1618 368 -1614
rect 401 -1618 405 -1614
rect 487 -1618 491 -1614
rect 513 -1618 517 -1614
rect 530 -1618 534 -1614
rect 570 -1618 574 -1614
rect 591 -1618 595 -1614
rect 608 -1618 612 -1614
rect 648 -1618 652 -1614
rect 672 -1618 676 -1614
rect 709 -1618 713 -1614
rect 795 -1618 799 -1614
rect 821 -1618 825 -1614
rect 838 -1618 842 -1614
rect 878 -1618 882 -1614
rect 899 -1618 903 -1614
rect 916 -1618 920 -1614
rect 956 -1618 960 -1614
rect 980 -1618 984 -1614
rect 1017 -1618 1021 -1614
rect -1047 -1633 -985 -1629
rect -981 -1633 -951 -1629
rect -903 -1633 -873 -1629
rect -739 -1633 -677 -1629
rect -673 -1633 -643 -1629
rect -595 -1633 -565 -1629
rect -431 -1633 -369 -1629
rect -365 -1633 -335 -1629
rect -287 -1633 -257 -1629
rect -123 -1633 -61 -1629
rect -57 -1633 -27 -1629
rect 21 -1633 51 -1629
rect 185 -1633 247 -1629
rect 251 -1633 281 -1629
rect 329 -1633 359 -1629
rect 493 -1633 555 -1629
rect 559 -1633 589 -1629
rect 637 -1633 667 -1629
rect 801 -1633 863 -1629
rect 867 -1633 897 -1629
rect 945 -1633 975 -1629
rect -1040 -1640 -1009 -1636
rect -732 -1640 -701 -1636
rect -424 -1640 -393 -1636
rect -116 -1640 -85 -1636
rect 192 -1640 223 -1636
rect 500 -1640 531 -1636
rect 808 -1640 839 -1636
rect -1058 -1647 -975 -1643
rect -936 -1647 -833 -1643
rect -750 -1647 -667 -1643
rect -628 -1647 -525 -1643
rect -442 -1647 -359 -1643
rect -320 -1647 -217 -1643
rect -134 -1647 -51 -1643
rect -12 -1647 91 -1643
rect 174 -1647 257 -1643
rect 296 -1647 399 -1643
rect 482 -1647 565 -1643
rect 604 -1647 707 -1643
rect 790 -1647 873 -1643
rect 912 -1647 1015 -1643
rect -1109 -1654 -1055 -1650
rect -1021 -1654 -992 -1650
rect -988 -1654 -907 -1650
rect -818 -1654 -791 -1650
rect -778 -1654 -747 -1650
rect -713 -1654 -684 -1650
rect -680 -1654 -599 -1650
rect -510 -1651 -485 -1647
rect -795 -1658 -791 -1654
rect -489 -1658 -485 -1651
rect -467 -1654 -439 -1650
rect -405 -1654 -376 -1650
rect -372 -1654 -291 -1650
rect -202 -1654 -180 -1650
rect -166 -1654 -131 -1650
rect -97 -1654 -68 -1650
rect -64 -1654 17 -1650
rect 106 -1654 130 -1650
rect 149 -1654 177 -1650
rect 211 -1654 240 -1650
rect 244 -1654 325 -1650
rect 414 -1654 438 -1650
rect 452 -1654 485 -1650
rect 519 -1654 548 -1650
rect 552 -1654 633 -1650
rect 722 -1652 737 -1648
rect -184 -1658 -180 -1654
rect 126 -1658 130 -1654
rect 434 -1658 438 -1654
rect 733 -1658 737 -1652
rect 746 -1654 793 -1650
rect 827 -1654 856 -1650
rect 860 -1654 941 -1650
rect -1230 -1663 -1173 -1659
rect -1134 -1662 -1029 -1658
rect -1014 -1662 -931 -1658
rect -910 -1662 -814 -1658
rect -795 -1662 -721 -1658
rect -706 -1662 -623 -1658
rect -602 -1662 -505 -1658
rect -489 -1662 -413 -1658
rect -398 -1662 -315 -1658
rect -294 -1662 -198 -1658
rect -184 -1662 -105 -1658
rect -90 -1662 -7 -1658
rect 14 -1662 111 -1658
rect 126 -1662 203 -1658
rect 218 -1662 301 -1658
rect 322 -1662 418 -1658
rect 434 -1662 511 -1658
rect 526 -1662 609 -1658
rect 630 -1662 726 -1658
rect 733 -1662 819 -1658
rect 834 -1662 917 -1658
rect 938 -1662 1041 -1658
rect -1253 -1670 -1223 -1666
rect -1219 -1670 -1183 -1666
rect -1179 -1670 -1163 -1666
rect -1091 -1669 -1051 -1665
rect -1032 -1669 -903 -1665
rect -791 -1669 -743 -1665
rect -724 -1669 -595 -1665
rect -485 -1669 -435 -1665
rect -416 -1669 -287 -1665
rect -180 -1669 -127 -1665
rect -108 -1669 21 -1665
rect 130 -1669 181 -1665
rect 200 -1669 329 -1665
rect 438 -1669 489 -1665
rect 508 -1669 637 -1665
rect 763 -1669 797 -1665
rect 816 -1669 945 -1665
rect -1279 -1677 -1227 -1673
rect -1223 -1677 -1197 -1673
rect -1193 -1677 -1149 -1673
rect -1025 -1676 -921 -1672
rect -917 -1676 -887 -1672
rect -717 -1676 -613 -1672
rect -609 -1676 -579 -1672
rect -409 -1676 -305 -1672
rect -301 -1676 -271 -1672
rect -101 -1676 3 -1672
rect 7 -1676 37 -1672
rect 207 -1676 311 -1672
rect 315 -1676 345 -1672
rect 515 -1676 619 -1672
rect 623 -1676 653 -1672
rect 823 -1676 927 -1672
rect 931 -1676 961 -1672
rect -1186 -1684 -1122 -1680
rect -1051 -1683 -999 -1679
rect -995 -1683 -965 -1679
rect -743 -1683 -691 -1679
rect -687 -1683 -657 -1679
rect -435 -1683 -383 -1679
rect -379 -1683 -349 -1679
rect -127 -1683 -75 -1679
rect -71 -1683 -41 -1679
rect 181 -1683 233 -1679
rect 237 -1683 267 -1679
rect 489 -1683 541 -1679
rect 545 -1683 575 -1679
rect 797 -1683 849 -1679
rect 853 -1683 883 -1679
rect -1204 -1691 -1172 -1687
rect -1006 -1691 -974 -1687
rect -1010 -1694 -1006 -1691
rect -974 -1694 -970 -1691
rect -928 -1691 -896 -1687
rect -932 -1694 -928 -1691
rect -896 -1694 -892 -1691
rect -698 -1691 -666 -1687
rect -702 -1694 -698 -1691
rect -666 -1694 -662 -1691
rect -620 -1691 -588 -1687
rect -624 -1694 -620 -1691
rect -588 -1694 -584 -1691
rect -390 -1691 -358 -1687
rect -394 -1694 -390 -1691
rect -358 -1694 -354 -1691
rect -312 -1691 -280 -1687
rect -316 -1694 -312 -1691
rect -280 -1694 -276 -1691
rect -82 -1691 -50 -1687
rect -86 -1694 -82 -1691
rect -50 -1694 -46 -1691
rect -4 -1691 28 -1687
rect -8 -1694 -4 -1691
rect 28 -1694 32 -1691
rect 226 -1691 258 -1687
rect 222 -1694 226 -1691
rect 258 -1694 262 -1691
rect 304 -1691 336 -1687
rect 300 -1694 304 -1691
rect 336 -1694 340 -1691
rect 534 -1691 566 -1687
rect 530 -1694 534 -1691
rect 566 -1694 570 -1691
rect 612 -1691 644 -1687
rect 608 -1694 612 -1691
rect 644 -1694 648 -1691
rect 842 -1691 874 -1687
rect 838 -1694 842 -1691
rect 874 -1694 878 -1691
rect 920 -1691 952 -1687
rect 916 -1694 920 -1691
rect 952 -1694 956 -1691
rect -1053 -1702 -1049 -1698
rect -1027 -1702 -1023 -1698
rect -984 -1702 -980 -1698
rect -949 -1702 -945 -1698
rect -905 -1702 -901 -1698
rect -888 -1702 -884 -1698
rect -852 -1702 -848 -1698
rect -831 -1702 -827 -1698
rect -745 -1702 -741 -1698
rect -719 -1702 -715 -1698
rect -676 -1702 -672 -1698
rect -641 -1702 -637 -1698
rect -597 -1702 -593 -1698
rect -580 -1702 -576 -1698
rect -544 -1702 -540 -1698
rect -523 -1702 -519 -1698
rect -437 -1702 -433 -1698
rect -411 -1702 -407 -1698
rect -368 -1702 -364 -1698
rect -333 -1702 -329 -1698
rect -289 -1702 -285 -1698
rect -272 -1702 -268 -1698
rect -236 -1702 -232 -1698
rect -215 -1702 -211 -1698
rect -129 -1702 -125 -1698
rect -103 -1702 -99 -1698
rect -60 -1702 -56 -1698
rect -25 -1702 -21 -1698
rect 19 -1702 23 -1698
rect 36 -1702 40 -1698
rect 72 -1702 76 -1698
rect 93 -1702 97 -1698
rect 179 -1702 183 -1698
rect 205 -1702 209 -1698
rect 248 -1702 252 -1698
rect 283 -1702 287 -1698
rect 327 -1702 331 -1698
rect 344 -1702 348 -1698
rect 380 -1702 384 -1698
rect 401 -1702 405 -1698
rect 487 -1702 491 -1698
rect 513 -1702 517 -1698
rect 556 -1702 560 -1698
rect 591 -1702 595 -1698
rect 635 -1702 639 -1698
rect 652 -1702 656 -1698
rect 688 -1702 692 -1698
rect 709 -1702 713 -1698
rect 795 -1702 799 -1698
rect 821 -1702 825 -1698
rect 864 -1702 868 -1698
rect 899 -1702 903 -1698
rect 943 -1702 947 -1698
rect 960 -1702 964 -1698
rect 996 -1702 1000 -1698
rect 1017 -1702 1021 -1698
rect 1179 -1702 1206 -1547
rect -1411 -1706 -1225 -1702
rect -1221 -1706 -1181 -1702
rect -1177 -1706 -1147 -1702
rect -1143 -1706 -1053 -1702
rect -1049 -1706 -1027 -1702
rect -1023 -1706 -984 -1702
rect -980 -1706 -949 -1702
rect -945 -1706 -905 -1702
rect -901 -1706 -888 -1702
rect -884 -1706 -852 -1702
rect -848 -1706 -831 -1702
rect -827 -1706 -745 -1702
rect -741 -1706 -719 -1702
rect -715 -1706 -676 -1702
rect -672 -1706 -641 -1702
rect -637 -1706 -597 -1702
rect -593 -1706 -580 -1702
rect -576 -1706 -544 -1702
rect -540 -1706 -523 -1702
rect -519 -1706 -437 -1702
rect -433 -1706 -411 -1702
rect -407 -1706 -368 -1702
rect -364 -1706 -333 -1702
rect -329 -1706 -289 -1702
rect -285 -1706 -272 -1702
rect -268 -1706 -236 -1702
rect -232 -1706 -215 -1702
rect -211 -1706 -129 -1702
rect -125 -1706 -103 -1702
rect -99 -1706 -60 -1702
rect -56 -1706 -25 -1702
rect -21 -1706 19 -1702
rect 23 -1706 36 -1702
rect 40 -1706 72 -1702
rect 76 -1706 93 -1702
rect 97 -1706 179 -1702
rect 183 -1706 205 -1702
rect 209 -1706 248 -1702
rect 252 -1706 283 -1702
rect 287 -1706 327 -1702
rect 331 -1706 344 -1702
rect 348 -1706 380 -1702
rect 384 -1706 401 -1702
rect 405 -1706 487 -1702
rect 491 -1706 513 -1702
rect 517 -1706 556 -1702
rect 560 -1706 591 -1702
rect 595 -1706 635 -1702
rect 639 -1706 652 -1702
rect 656 -1706 688 -1702
rect 692 -1706 709 -1702
rect 713 -1706 795 -1702
rect 799 -1706 821 -1702
rect 825 -1706 864 -1702
rect 868 -1706 899 -1702
rect 903 -1706 943 -1702
rect 947 -1706 960 -1702
rect 964 -1706 996 -1702
rect 1000 -1706 1017 -1702
rect 1021 -1706 1206 -1702
rect -1253 -1713 -814 -1709
rect -776 -1713 -198 -1709
rect -162 -1713 418 -1709
rect 453 -1713 1041 -1709
rect -1086 -1720 -505 -1716
rect -472 -1720 111 -1716
rect 144 -1720 726 -1716
rect 763 -1720 1026 -1716
rect -1454 -1746 -1309 -1742
rect -1305 -1746 -1292 -1742
rect -1288 -1746 -1062 -1742
rect -1058 -1746 -1045 -1742
rect -1041 -1746 -754 -1742
rect -750 -1746 -737 -1742
rect -733 -1746 -446 -1742
rect -442 -1746 -429 -1742
rect -425 -1746 -138 -1742
rect -134 -1746 -121 -1742
rect -117 -1746 170 -1742
rect 174 -1746 187 -1742
rect 191 -1746 478 -1742
rect 482 -1746 495 -1742
rect 499 -1746 786 -1742
rect 790 -1746 803 -1742
rect 807 -1746 1164 -1742
rect -1454 -1901 -1427 -1746
rect -1411 -1786 -1297 -1782
rect -1293 -1786 -1050 -1782
rect -1046 -1786 -742 -1782
rect -738 -1786 -434 -1782
rect -430 -1786 -126 -1782
rect -122 -1786 182 -1782
rect 186 -1786 490 -1782
rect 494 -1786 798 -1782
rect 802 -1786 1164 -1782
rect -1102 -1799 -1036 -1795
rect -789 -1799 -728 -1795
rect -486 -1799 -420 -1795
rect -176 -1799 -112 -1795
rect 130 -1799 196 -1795
rect 439 -1799 504 -1795
rect 746 -1799 812 -1795
rect 1179 -1834 1206 -1706
rect -1411 -1838 -1292 -1834
rect -1288 -1838 -1045 -1834
rect -1041 -1838 -737 -1834
rect -733 -1838 -429 -1834
rect -425 -1838 -121 -1834
rect -117 -1838 187 -1834
rect 191 -1838 495 -1834
rect 499 -1838 803 -1834
rect 807 -1838 1206 -1834
rect -1454 -1905 -1225 -1901
rect -1221 -1905 -1208 -1901
rect -1204 -1905 -1168 -1901
rect -1164 -1905 -1147 -1901
rect -1143 -1905 -1053 -1901
rect -1049 -1905 -1027 -1901
rect -1023 -1905 -1010 -1901
rect -1006 -1905 -970 -1901
rect -966 -1905 -949 -1901
rect -945 -1905 -932 -1901
rect -928 -1905 -892 -1901
rect -888 -1905 -868 -1901
rect -864 -1905 -831 -1901
rect -827 -1905 -745 -1901
rect -741 -1905 -719 -1901
rect -715 -1905 -702 -1901
rect -698 -1905 -662 -1901
rect -658 -1905 -641 -1901
rect -637 -1905 -624 -1901
rect -620 -1905 -584 -1901
rect -580 -1905 -560 -1901
rect -556 -1905 -523 -1901
rect -519 -1905 -437 -1901
rect -433 -1905 -411 -1901
rect -407 -1905 -394 -1901
rect -390 -1905 -354 -1901
rect -350 -1905 -333 -1901
rect -329 -1905 -316 -1901
rect -312 -1905 -276 -1901
rect -272 -1905 -252 -1901
rect -248 -1905 -215 -1901
rect -211 -1905 -129 -1901
rect -125 -1905 -103 -1901
rect -99 -1905 -86 -1901
rect -82 -1905 -46 -1901
rect -42 -1905 -25 -1901
rect -21 -1905 -8 -1901
rect -4 -1905 32 -1901
rect 36 -1905 56 -1901
rect 60 -1905 93 -1901
rect 97 -1905 179 -1901
rect 183 -1905 205 -1901
rect 209 -1905 222 -1901
rect 226 -1905 262 -1901
rect 266 -1905 283 -1901
rect 287 -1905 300 -1901
rect 304 -1905 340 -1901
rect 344 -1905 364 -1901
rect 368 -1905 401 -1901
rect 405 -1905 487 -1901
rect 491 -1905 513 -1901
rect 517 -1905 530 -1901
rect 534 -1905 570 -1901
rect 574 -1905 591 -1901
rect 595 -1905 608 -1901
rect 612 -1905 648 -1901
rect 652 -1905 672 -1901
rect 676 -1905 709 -1901
rect 713 -1905 795 -1901
rect 799 -1905 821 -1901
rect 825 -1905 838 -1901
rect 842 -1905 878 -1901
rect 882 -1905 899 -1901
rect 903 -1905 916 -1901
rect 920 -1905 956 -1901
rect 960 -1905 980 -1901
rect 984 -1905 1017 -1901
rect 1021 -1905 1164 -1901
rect -1454 -2064 -1427 -1905
rect -1053 -1909 -1049 -1905
rect -1027 -1909 -1023 -1905
rect -1010 -1909 -1006 -1905
rect -970 -1909 -966 -1905
rect -949 -1909 -945 -1905
rect -932 -1909 -928 -1905
rect -892 -1909 -888 -1905
rect -868 -1909 -864 -1905
rect -831 -1909 -827 -1905
rect -745 -1909 -741 -1905
rect -719 -1909 -715 -1905
rect -702 -1909 -698 -1905
rect -662 -1909 -658 -1905
rect -641 -1909 -637 -1905
rect -624 -1909 -620 -1905
rect -584 -1909 -580 -1905
rect -560 -1909 -556 -1905
rect -523 -1909 -519 -1905
rect -437 -1909 -433 -1905
rect -411 -1909 -407 -1905
rect -394 -1909 -390 -1905
rect -354 -1909 -350 -1905
rect -333 -1909 -329 -1905
rect -316 -1909 -312 -1905
rect -276 -1909 -272 -1905
rect -252 -1909 -248 -1905
rect -215 -1909 -211 -1905
rect -129 -1909 -125 -1905
rect -103 -1909 -99 -1905
rect -86 -1909 -82 -1905
rect -46 -1909 -42 -1905
rect -25 -1909 -21 -1905
rect -8 -1909 -4 -1905
rect 32 -1909 36 -1905
rect 56 -1909 60 -1905
rect 93 -1909 97 -1905
rect 179 -1909 183 -1905
rect 205 -1909 209 -1905
rect 222 -1909 226 -1905
rect 262 -1909 266 -1905
rect 283 -1909 287 -1905
rect 300 -1909 304 -1905
rect 340 -1909 344 -1905
rect 364 -1909 368 -1905
rect 401 -1909 405 -1905
rect 487 -1909 491 -1905
rect 513 -1909 517 -1905
rect 530 -1909 534 -1905
rect 570 -1909 574 -1905
rect 591 -1909 595 -1905
rect 608 -1909 612 -1905
rect 648 -1909 652 -1905
rect 672 -1909 676 -1905
rect 709 -1909 713 -1905
rect 795 -1909 799 -1905
rect 821 -1909 825 -1905
rect 838 -1909 842 -1905
rect 878 -1909 882 -1905
rect 899 -1909 903 -1905
rect 916 -1909 920 -1905
rect 956 -1909 960 -1905
rect 980 -1909 984 -1905
rect 1017 -1909 1021 -1905
rect -1047 -1924 -985 -1920
rect -981 -1924 -951 -1920
rect -903 -1924 -873 -1920
rect -739 -1924 -677 -1920
rect -673 -1924 -643 -1920
rect -595 -1924 -565 -1920
rect -431 -1924 -369 -1920
rect -365 -1924 -335 -1920
rect -287 -1924 -257 -1920
rect -123 -1924 -61 -1920
rect -57 -1924 -27 -1920
rect 21 -1924 51 -1920
rect 185 -1924 247 -1920
rect 251 -1924 281 -1920
rect 329 -1924 359 -1920
rect 493 -1924 555 -1920
rect 559 -1924 589 -1920
rect 637 -1924 667 -1920
rect 801 -1924 863 -1920
rect 867 -1924 897 -1920
rect 945 -1924 975 -1920
rect -1040 -1931 -1009 -1927
rect -732 -1931 -701 -1927
rect -424 -1931 -393 -1927
rect -116 -1931 -85 -1927
rect 192 -1931 223 -1927
rect 500 -1931 531 -1927
rect 808 -1931 839 -1927
rect -1058 -1938 -975 -1934
rect -936 -1938 -833 -1934
rect -750 -1938 -667 -1934
rect -628 -1938 -525 -1934
rect -442 -1938 -359 -1934
rect -320 -1938 -217 -1934
rect -134 -1938 -51 -1934
rect -12 -1938 91 -1934
rect 174 -1938 257 -1934
rect 296 -1938 399 -1934
rect 482 -1938 565 -1934
rect 604 -1938 707 -1934
rect 790 -1938 873 -1934
rect 912 -1938 1015 -1934
rect -1102 -1945 -1055 -1941
rect -1021 -1945 -992 -1941
rect -988 -1945 -907 -1941
rect -818 -1945 -789 -1941
rect -776 -1945 -747 -1941
rect -713 -1945 -684 -1941
rect -680 -1945 -599 -1941
rect -510 -1944 -486 -1940
rect -793 -1949 -789 -1945
rect -490 -1949 -486 -1944
rect -472 -1945 -439 -1941
rect -405 -1945 -376 -1941
rect -372 -1945 -291 -1941
rect -202 -1945 -176 -1941
rect -162 -1945 -131 -1941
rect -97 -1945 -68 -1941
rect -64 -1945 17 -1941
rect 106 -1945 130 -1941
rect 144 -1945 177 -1941
rect 211 -1945 240 -1941
rect 244 -1945 325 -1941
rect 414 -1945 439 -1941
rect 453 -1945 485 -1941
rect 519 -1945 548 -1941
rect 552 -1945 633 -1941
rect 722 -1943 739 -1939
rect -180 -1949 -176 -1945
rect 126 -1949 130 -1945
rect 435 -1949 439 -1945
rect 735 -1949 739 -1943
rect 746 -1945 793 -1941
rect 827 -1945 856 -1941
rect 860 -1945 941 -1941
rect -1230 -1954 -1173 -1950
rect -1134 -1953 -1029 -1949
rect -1014 -1953 -931 -1949
rect -910 -1953 -815 -1949
rect -793 -1953 -721 -1949
rect -706 -1953 -623 -1949
rect -602 -1953 -506 -1949
rect -490 -1953 -413 -1949
rect -398 -1953 -315 -1949
rect -294 -1953 -199 -1949
rect -180 -1953 -105 -1949
rect -90 -1953 -7 -1949
rect 14 -1953 112 -1949
rect 126 -1953 203 -1949
rect 218 -1953 301 -1949
rect 322 -1953 417 -1949
rect 435 -1953 511 -1949
rect 526 -1953 609 -1949
rect 630 -1953 728 -1949
rect 735 -1953 819 -1949
rect 834 -1953 917 -1949
rect 938 -1953 1042 -1949
rect -1253 -1961 -1223 -1957
rect -1219 -1961 -1183 -1957
rect -1179 -1961 -1163 -1957
rect -1086 -1960 -1051 -1956
rect -1032 -1960 -903 -1956
rect -789 -1960 -743 -1956
rect -724 -1960 -595 -1956
rect -486 -1960 -435 -1956
rect -416 -1960 -287 -1956
rect -176 -1960 -127 -1956
rect -108 -1960 21 -1956
rect 130 -1960 181 -1956
rect 200 -1960 329 -1956
rect 439 -1960 489 -1956
rect 508 -1960 637 -1956
rect 763 -1960 797 -1956
rect 816 -1960 945 -1956
rect -1279 -1968 -1227 -1964
rect -1223 -1968 -1197 -1964
rect -1193 -1968 -1149 -1964
rect -1025 -1967 -921 -1963
rect -917 -1967 -887 -1963
rect -717 -1967 -613 -1963
rect -609 -1967 -579 -1963
rect -409 -1967 -305 -1963
rect -301 -1967 -271 -1963
rect -101 -1967 3 -1963
rect 7 -1967 37 -1963
rect 207 -1967 311 -1963
rect 315 -1967 345 -1963
rect 515 -1967 619 -1963
rect 623 -1967 653 -1963
rect 823 -1967 927 -1963
rect 931 -1967 961 -1963
rect -1186 -1975 -1122 -1971
rect -1051 -1974 -999 -1970
rect -995 -1974 -965 -1970
rect -743 -1974 -691 -1970
rect -687 -1974 -657 -1970
rect -435 -1974 -383 -1970
rect -379 -1974 -349 -1970
rect -127 -1974 -75 -1970
rect -71 -1974 -41 -1970
rect 181 -1974 233 -1970
rect 237 -1974 267 -1970
rect 489 -1974 541 -1970
rect 545 -1974 575 -1970
rect 797 -1974 849 -1970
rect 853 -1974 883 -1970
rect -1204 -1982 -1172 -1978
rect -1006 -1982 -974 -1978
rect -1010 -1985 -1006 -1982
rect -974 -1985 -970 -1982
rect -928 -1982 -896 -1978
rect -932 -1985 -928 -1982
rect -896 -1985 -892 -1982
rect -698 -1982 -666 -1978
rect -702 -1985 -698 -1982
rect -666 -1985 -662 -1982
rect -620 -1982 -588 -1978
rect -624 -1985 -620 -1982
rect -588 -1985 -584 -1982
rect -390 -1982 -358 -1978
rect -394 -1985 -390 -1982
rect -358 -1985 -354 -1982
rect -312 -1982 -280 -1978
rect -316 -1985 -312 -1982
rect -280 -1985 -276 -1982
rect -82 -1982 -50 -1978
rect -86 -1985 -82 -1982
rect -50 -1985 -46 -1982
rect -4 -1982 28 -1978
rect -8 -1985 -4 -1982
rect 28 -1985 32 -1982
rect 226 -1982 258 -1978
rect 222 -1985 226 -1982
rect 258 -1985 262 -1982
rect 304 -1982 336 -1978
rect 300 -1985 304 -1982
rect 336 -1985 340 -1982
rect 534 -1982 566 -1978
rect 530 -1985 534 -1982
rect 566 -1985 570 -1982
rect 612 -1982 644 -1978
rect 608 -1985 612 -1982
rect 644 -1985 648 -1982
rect 842 -1982 874 -1978
rect 838 -1985 842 -1982
rect 874 -1985 878 -1982
rect 920 -1982 952 -1978
rect 916 -1985 920 -1982
rect 952 -1985 956 -1982
rect -1053 -1993 -1049 -1989
rect -1027 -1993 -1023 -1989
rect -984 -1993 -980 -1989
rect -949 -1993 -945 -1989
rect -905 -1993 -901 -1989
rect -888 -1993 -884 -1989
rect -852 -1993 -848 -1989
rect -831 -1993 -827 -1989
rect -745 -1993 -741 -1989
rect -719 -1993 -715 -1989
rect -676 -1993 -672 -1989
rect -641 -1993 -637 -1989
rect -597 -1993 -593 -1989
rect -580 -1993 -576 -1989
rect -544 -1993 -540 -1989
rect -523 -1993 -519 -1989
rect -437 -1993 -433 -1989
rect -411 -1993 -407 -1989
rect -368 -1993 -364 -1989
rect -333 -1993 -329 -1989
rect -289 -1993 -285 -1989
rect -272 -1993 -268 -1989
rect -236 -1993 -232 -1989
rect -215 -1993 -211 -1989
rect -129 -1993 -125 -1989
rect -103 -1993 -99 -1989
rect -60 -1993 -56 -1989
rect -25 -1993 -21 -1989
rect 19 -1993 23 -1989
rect 36 -1993 40 -1989
rect 72 -1993 76 -1989
rect 93 -1993 97 -1989
rect 179 -1993 183 -1989
rect 205 -1993 209 -1989
rect 248 -1993 252 -1989
rect 283 -1993 287 -1989
rect 327 -1993 331 -1989
rect 344 -1993 348 -1989
rect 380 -1993 384 -1989
rect 401 -1993 405 -1989
rect 487 -1993 491 -1989
rect 513 -1993 517 -1989
rect 556 -1993 560 -1989
rect 591 -1993 595 -1989
rect 635 -1993 639 -1989
rect 652 -1993 656 -1989
rect 688 -1993 692 -1989
rect 709 -1993 713 -1989
rect 795 -1993 799 -1989
rect 821 -1993 825 -1989
rect 864 -1993 868 -1989
rect 899 -1993 903 -1989
rect 943 -1993 947 -1989
rect 960 -1993 964 -1989
rect 996 -1993 1000 -1989
rect 1017 -1993 1021 -1989
rect 1179 -1993 1206 -1838
rect -1411 -1997 -1225 -1993
rect -1221 -1997 -1181 -1993
rect -1177 -1997 -1147 -1993
rect -1143 -1997 -1053 -1993
rect -1049 -1997 -1027 -1993
rect -1023 -1997 -984 -1993
rect -980 -1997 -949 -1993
rect -945 -1997 -905 -1993
rect -901 -1997 -888 -1993
rect -884 -1997 -852 -1993
rect -848 -1997 -831 -1993
rect -827 -1997 -745 -1993
rect -741 -1997 -719 -1993
rect -715 -1997 -676 -1993
rect -672 -1997 -641 -1993
rect -637 -1997 -597 -1993
rect -593 -1997 -580 -1993
rect -576 -1997 -544 -1993
rect -540 -1997 -523 -1993
rect -519 -1997 -437 -1993
rect -433 -1997 -411 -1993
rect -407 -1997 -368 -1993
rect -364 -1997 -333 -1993
rect -329 -1997 -289 -1993
rect -285 -1997 -272 -1993
rect -268 -1997 -236 -1993
rect -232 -1997 -215 -1993
rect -211 -1997 -129 -1993
rect -125 -1997 -103 -1993
rect -99 -1997 -60 -1993
rect -56 -1997 -25 -1993
rect -21 -1997 19 -1993
rect 23 -1997 36 -1993
rect 40 -1997 72 -1993
rect 76 -1997 93 -1993
rect 97 -1997 179 -1993
rect 183 -1997 205 -1993
rect 209 -1997 248 -1993
rect 252 -1997 283 -1993
rect 287 -1997 327 -1993
rect 331 -1997 344 -1993
rect 348 -1997 380 -1993
rect 384 -1997 401 -1993
rect 405 -1997 487 -1993
rect 491 -1997 513 -1993
rect 517 -1997 556 -1993
rect 560 -1997 591 -1993
rect 595 -1997 635 -1993
rect 639 -1997 652 -1993
rect 656 -1997 688 -1993
rect 692 -1997 709 -1993
rect 713 -1997 795 -1993
rect 799 -1997 821 -1993
rect 825 -1997 864 -1993
rect 868 -1997 899 -1993
rect 903 -1997 943 -1993
rect 947 -1997 960 -1993
rect 964 -1997 996 -1993
rect 1000 -1997 1017 -1993
rect 1021 -1997 1206 -1993
rect -1253 -2004 -815 -2000
rect -776 -2004 -199 -2000
rect -162 -2004 417 -2000
rect 452 -2004 1042 -2000
rect -1086 -2011 -506 -2007
rect -472 -2011 112 -2007
rect 144 -2011 728 -2007
rect 763 -2011 1026 -2007
rect -1454 -2068 -1309 -2064
rect -1305 -2068 -1292 -2064
rect -1288 -2068 -1062 -2064
rect -1058 -2068 -1045 -2064
rect -1041 -2068 -754 -2064
rect -750 -2068 -737 -2064
rect -733 -2068 -446 -2064
rect -442 -2068 -429 -2064
rect -425 -2068 -138 -2064
rect -134 -2068 -121 -2064
rect -117 -2068 170 -2064
rect 174 -2068 187 -2064
rect 191 -2068 478 -2064
rect 482 -2068 495 -2064
rect 499 -2068 786 -2064
rect 790 -2068 803 -2064
rect 807 -2068 1164 -2064
rect -1454 -2223 -1427 -2068
rect -1411 -2108 -1297 -2104
rect -1293 -2108 -1050 -2104
rect -1046 -2108 -742 -2104
rect -738 -2108 -434 -2104
rect -430 -2108 -126 -2104
rect -122 -2108 182 -2104
rect 186 -2108 490 -2104
rect 494 -2108 798 -2104
rect 802 -2108 1164 -2104
rect -1102 -2121 -1036 -2117
rect -789 -2121 -728 -2117
rect -486 -2121 -420 -2117
rect -176 -2121 -112 -2117
rect 130 -2121 196 -2117
rect 438 -2121 504 -2117
rect 746 -2121 812 -2117
rect 1179 -2156 1206 -1997
rect -1411 -2160 -1292 -2156
rect -1288 -2160 -1045 -2156
rect -1041 -2160 -737 -2156
rect -733 -2160 -429 -2156
rect -425 -2160 -121 -2156
rect -117 -2160 187 -2156
rect 191 -2160 495 -2156
rect 499 -2160 803 -2156
rect 807 -2160 1206 -2156
rect -1454 -2227 -1225 -2223
rect -1221 -2227 -1208 -2223
rect -1204 -2227 -1168 -2223
rect -1164 -2227 -1147 -2223
rect -1143 -2227 -1053 -2223
rect -1049 -2227 -1027 -2223
rect -1023 -2227 -1010 -2223
rect -1006 -2227 -970 -2223
rect -966 -2227 -949 -2223
rect -945 -2227 -932 -2223
rect -928 -2227 -892 -2223
rect -888 -2227 -868 -2223
rect -864 -2227 -831 -2223
rect -827 -2227 -745 -2223
rect -741 -2227 -719 -2223
rect -715 -2227 -702 -2223
rect -698 -2227 -662 -2223
rect -658 -2227 -641 -2223
rect -637 -2227 -624 -2223
rect -620 -2227 -584 -2223
rect -580 -2227 -560 -2223
rect -556 -2227 -523 -2223
rect -519 -2227 -437 -2223
rect -433 -2227 -411 -2223
rect -407 -2227 -394 -2223
rect -390 -2227 -354 -2223
rect -350 -2227 -333 -2223
rect -329 -2227 -316 -2223
rect -312 -2227 -276 -2223
rect -272 -2227 -252 -2223
rect -248 -2227 -215 -2223
rect -211 -2227 -129 -2223
rect -125 -2227 -103 -2223
rect -99 -2227 -86 -2223
rect -82 -2227 -46 -2223
rect -42 -2227 -25 -2223
rect -21 -2227 -8 -2223
rect -4 -2227 32 -2223
rect 36 -2227 56 -2223
rect 60 -2227 93 -2223
rect 97 -2227 179 -2223
rect 183 -2227 205 -2223
rect 209 -2227 222 -2223
rect 226 -2227 262 -2223
rect 266 -2227 283 -2223
rect 287 -2227 300 -2223
rect 304 -2227 340 -2223
rect 344 -2227 364 -2223
rect 368 -2227 401 -2223
rect 405 -2227 487 -2223
rect 491 -2227 513 -2223
rect 517 -2227 530 -2223
rect 534 -2227 570 -2223
rect 574 -2227 591 -2223
rect 595 -2227 608 -2223
rect 612 -2227 648 -2223
rect 652 -2227 672 -2223
rect 676 -2227 709 -2223
rect 713 -2227 795 -2223
rect 799 -2227 821 -2223
rect 825 -2227 838 -2223
rect 842 -2227 878 -2223
rect 882 -2227 899 -2223
rect 903 -2227 916 -2223
rect 920 -2227 956 -2223
rect 960 -2227 980 -2223
rect 984 -2227 1017 -2223
rect 1021 -2227 1164 -2223
rect -1454 -2355 -1427 -2227
rect -1053 -2231 -1049 -2227
rect -1027 -2231 -1023 -2227
rect -1010 -2231 -1006 -2227
rect -970 -2231 -966 -2227
rect -949 -2231 -945 -2227
rect -932 -2231 -928 -2227
rect -892 -2231 -888 -2227
rect -868 -2231 -864 -2227
rect -831 -2231 -827 -2227
rect -745 -2231 -741 -2227
rect -719 -2231 -715 -2227
rect -702 -2231 -698 -2227
rect -662 -2231 -658 -2227
rect -641 -2231 -637 -2227
rect -624 -2231 -620 -2227
rect -584 -2231 -580 -2227
rect -560 -2231 -556 -2227
rect -523 -2231 -519 -2227
rect -437 -2231 -433 -2227
rect -411 -2231 -407 -2227
rect -394 -2231 -390 -2227
rect -354 -2231 -350 -2227
rect -333 -2231 -329 -2227
rect -316 -2231 -312 -2227
rect -276 -2231 -272 -2227
rect -252 -2231 -248 -2227
rect -215 -2231 -211 -2227
rect -129 -2231 -125 -2227
rect -103 -2231 -99 -2227
rect -86 -2231 -82 -2227
rect -46 -2231 -42 -2227
rect -25 -2231 -21 -2227
rect -8 -2231 -4 -2227
rect 32 -2231 36 -2227
rect 56 -2231 60 -2227
rect 93 -2231 97 -2227
rect 179 -2231 183 -2227
rect 205 -2231 209 -2227
rect 222 -2231 226 -2227
rect 262 -2231 266 -2227
rect 283 -2231 287 -2227
rect 300 -2231 304 -2227
rect 340 -2231 344 -2227
rect 364 -2231 368 -2227
rect 401 -2231 405 -2227
rect 487 -2231 491 -2227
rect 513 -2231 517 -2227
rect 530 -2231 534 -2227
rect 570 -2231 574 -2227
rect 591 -2231 595 -2227
rect 608 -2231 612 -2227
rect 648 -2231 652 -2227
rect 672 -2231 676 -2227
rect 709 -2231 713 -2227
rect 795 -2231 799 -2227
rect 821 -2231 825 -2227
rect 838 -2231 842 -2227
rect 878 -2231 882 -2227
rect 899 -2231 903 -2227
rect 916 -2231 920 -2227
rect 956 -2231 960 -2227
rect 980 -2231 984 -2227
rect 1017 -2231 1021 -2227
rect -1047 -2246 -985 -2242
rect -981 -2246 -951 -2242
rect -903 -2246 -873 -2242
rect -739 -2246 -677 -2242
rect -673 -2246 -643 -2242
rect -595 -2246 -565 -2242
rect -431 -2246 -369 -2242
rect -365 -2246 -335 -2242
rect -287 -2246 -257 -2242
rect -123 -2246 -61 -2242
rect -57 -2246 -27 -2242
rect 21 -2246 51 -2242
rect 185 -2246 247 -2242
rect 251 -2246 281 -2242
rect 329 -2246 359 -2242
rect 493 -2246 555 -2242
rect 559 -2246 589 -2242
rect 637 -2246 667 -2242
rect 801 -2246 863 -2242
rect 867 -2246 897 -2242
rect 945 -2246 975 -2242
rect -1040 -2253 -1009 -2249
rect -732 -2253 -701 -2249
rect -424 -2253 -393 -2249
rect -116 -2253 -85 -2249
rect 192 -2253 223 -2249
rect 500 -2253 531 -2249
rect 808 -2253 839 -2249
rect -1058 -2260 -975 -2256
rect -936 -2260 -833 -2256
rect -750 -2260 -667 -2256
rect -628 -2260 -525 -2256
rect -442 -2260 -359 -2256
rect -320 -2260 -217 -2256
rect -134 -2260 -51 -2256
rect -12 -2260 91 -2256
rect 174 -2260 257 -2256
rect 296 -2260 399 -2256
rect 482 -2260 565 -2256
rect 604 -2260 707 -2256
rect 790 -2260 873 -2256
rect 912 -2260 1015 -2256
rect -1102 -2267 -1055 -2263
rect -1021 -2267 -992 -2263
rect -988 -2267 -907 -2263
rect -818 -2267 -789 -2263
rect -776 -2267 -747 -2263
rect -713 -2267 -684 -2263
rect -680 -2267 -599 -2263
rect -510 -2266 -486 -2262
rect -793 -2271 -789 -2267
rect -490 -2271 -486 -2266
rect -472 -2267 -439 -2263
rect -405 -2267 -376 -2263
rect -372 -2267 -291 -2263
rect -202 -2267 -176 -2263
rect -162 -2267 -131 -2263
rect -97 -2267 -68 -2263
rect -64 -2267 17 -2263
rect 106 -2267 130 -2263
rect 144 -2267 177 -2263
rect 211 -2267 240 -2263
rect 244 -2267 325 -2263
rect 414 -2267 439 -2263
rect 453 -2267 485 -2263
rect 519 -2267 548 -2263
rect 552 -2267 633 -2263
rect 722 -2265 739 -2261
rect -180 -2271 -176 -2267
rect 126 -2271 130 -2267
rect 435 -2271 439 -2267
rect 735 -2271 739 -2265
rect 746 -2267 793 -2263
rect 827 -2267 856 -2263
rect 860 -2267 941 -2263
rect -1230 -2276 -1173 -2272
rect -1134 -2275 -1029 -2271
rect -1014 -2275 -931 -2271
rect -910 -2275 -814 -2271
rect -793 -2275 -721 -2271
rect -706 -2275 -623 -2271
rect -602 -2275 -505 -2271
rect -490 -2275 -413 -2271
rect -398 -2275 -315 -2271
rect -294 -2275 -198 -2271
rect -180 -2275 -105 -2271
rect -90 -2275 -7 -2271
rect 14 -2275 111 -2271
rect 126 -2275 203 -2271
rect 218 -2275 301 -2271
rect 322 -2275 418 -2271
rect 435 -2275 511 -2271
rect 526 -2275 609 -2271
rect 630 -2275 726 -2271
rect 735 -2275 819 -2271
rect 834 -2275 917 -2271
rect 938 -2275 1039 -2271
rect -1253 -2283 -1223 -2279
rect -1219 -2283 -1183 -2279
rect -1179 -2283 -1163 -2279
rect -1086 -2282 -1051 -2278
rect -1032 -2282 -903 -2278
rect -789 -2282 -743 -2278
rect -724 -2282 -595 -2278
rect -486 -2282 -435 -2278
rect -416 -2282 -287 -2278
rect -176 -2282 -127 -2278
rect -108 -2282 21 -2278
rect 130 -2282 181 -2278
rect 200 -2282 329 -2278
rect 439 -2282 489 -2278
rect 508 -2282 637 -2278
rect 763 -2282 797 -2278
rect 816 -2282 945 -2278
rect -1279 -2290 -1227 -2286
rect -1223 -2290 -1197 -2286
rect -1193 -2290 -1149 -2286
rect -1025 -2289 -921 -2285
rect -917 -2289 -887 -2285
rect -717 -2289 -613 -2285
rect -609 -2289 -579 -2285
rect -409 -2289 -305 -2285
rect -301 -2289 -271 -2285
rect -101 -2289 3 -2285
rect 7 -2289 37 -2285
rect 207 -2289 311 -2285
rect 315 -2289 345 -2285
rect 515 -2289 619 -2285
rect 623 -2289 653 -2285
rect 823 -2289 927 -2285
rect 931 -2289 961 -2285
rect -1186 -2297 -1122 -2293
rect -1051 -2296 -999 -2292
rect -995 -2296 -965 -2292
rect -743 -2296 -691 -2292
rect -687 -2296 -657 -2292
rect -435 -2296 -383 -2292
rect -379 -2296 -349 -2292
rect -127 -2296 -75 -2292
rect -71 -2296 -41 -2292
rect 181 -2296 233 -2292
rect 237 -2296 267 -2292
rect 489 -2296 541 -2292
rect 545 -2296 575 -2292
rect 797 -2296 849 -2292
rect 853 -2296 883 -2292
rect -1204 -2304 -1172 -2300
rect -1006 -2304 -974 -2300
rect -1010 -2307 -1006 -2304
rect -974 -2307 -970 -2304
rect -928 -2304 -896 -2300
rect -932 -2307 -928 -2304
rect -896 -2307 -892 -2304
rect -698 -2304 -666 -2300
rect -702 -2307 -698 -2304
rect -666 -2307 -662 -2304
rect -620 -2304 -588 -2300
rect -624 -2307 -620 -2304
rect -588 -2307 -584 -2304
rect -390 -2304 -358 -2300
rect -394 -2307 -390 -2304
rect -358 -2307 -354 -2304
rect -312 -2304 -280 -2300
rect -316 -2307 -312 -2304
rect -280 -2307 -276 -2304
rect -82 -2304 -50 -2300
rect -86 -2307 -82 -2304
rect -50 -2307 -46 -2304
rect -4 -2304 28 -2300
rect -8 -2307 -4 -2304
rect 28 -2307 32 -2304
rect 226 -2304 258 -2300
rect 222 -2307 226 -2304
rect 258 -2307 262 -2304
rect 304 -2304 336 -2300
rect 300 -2307 304 -2304
rect 336 -2307 340 -2304
rect 534 -2304 566 -2300
rect 530 -2307 534 -2304
rect 566 -2307 570 -2304
rect 612 -2304 644 -2300
rect 608 -2307 612 -2304
rect 644 -2307 648 -2304
rect 842 -2304 874 -2300
rect 838 -2307 842 -2304
rect 874 -2307 878 -2304
rect 920 -2304 952 -2300
rect 916 -2307 920 -2304
rect 952 -2307 956 -2304
rect -1053 -2315 -1049 -2311
rect -1027 -2315 -1023 -2311
rect -984 -2315 -980 -2311
rect -949 -2315 -945 -2311
rect -905 -2315 -901 -2311
rect -888 -2315 -884 -2311
rect -852 -2315 -848 -2311
rect -831 -2315 -827 -2311
rect -745 -2315 -741 -2311
rect -719 -2315 -715 -2311
rect -676 -2315 -672 -2311
rect -641 -2315 -637 -2311
rect -597 -2315 -593 -2311
rect -580 -2315 -576 -2311
rect -544 -2315 -540 -2311
rect -523 -2315 -519 -2311
rect -437 -2315 -433 -2311
rect -411 -2315 -407 -2311
rect -368 -2315 -364 -2311
rect -333 -2315 -329 -2311
rect -289 -2315 -285 -2311
rect -272 -2315 -268 -2311
rect -236 -2315 -232 -2311
rect -215 -2315 -211 -2311
rect -129 -2315 -125 -2311
rect -103 -2315 -99 -2311
rect -60 -2315 -56 -2311
rect -25 -2315 -21 -2311
rect 19 -2315 23 -2311
rect 36 -2315 40 -2311
rect 72 -2315 76 -2311
rect 93 -2315 97 -2311
rect 179 -2315 183 -2311
rect 205 -2315 209 -2311
rect 248 -2315 252 -2311
rect 283 -2315 287 -2311
rect 327 -2315 331 -2311
rect 344 -2315 348 -2311
rect 380 -2315 384 -2311
rect 401 -2315 405 -2311
rect 487 -2315 491 -2311
rect 513 -2315 517 -2311
rect 556 -2315 560 -2311
rect 591 -2315 595 -2311
rect 635 -2315 639 -2311
rect 652 -2315 656 -2311
rect 688 -2315 692 -2311
rect 709 -2315 713 -2311
rect 795 -2315 799 -2311
rect 821 -2315 825 -2311
rect 864 -2315 868 -2311
rect 899 -2315 903 -2311
rect 943 -2315 947 -2311
rect 960 -2315 964 -2311
rect 996 -2315 1000 -2311
rect 1017 -2315 1021 -2311
rect 1179 -2315 1206 -2160
rect -1411 -2319 -1225 -2315
rect -1221 -2319 -1181 -2315
rect -1177 -2319 -1147 -2315
rect -1143 -2319 -1053 -2315
rect -1049 -2319 -1027 -2315
rect -1023 -2319 -984 -2315
rect -980 -2319 -949 -2315
rect -945 -2319 -905 -2315
rect -901 -2319 -888 -2315
rect -884 -2319 -852 -2315
rect -848 -2319 -831 -2315
rect -827 -2319 -745 -2315
rect -741 -2319 -719 -2315
rect -715 -2319 -676 -2315
rect -672 -2319 -641 -2315
rect -637 -2319 -597 -2315
rect -593 -2319 -580 -2315
rect -576 -2319 -544 -2315
rect -540 -2319 -523 -2315
rect -519 -2319 -437 -2315
rect -433 -2319 -411 -2315
rect -407 -2319 -368 -2315
rect -364 -2319 -333 -2315
rect -329 -2319 -289 -2315
rect -285 -2319 -272 -2315
rect -268 -2319 -236 -2315
rect -232 -2319 -215 -2315
rect -211 -2319 -129 -2315
rect -125 -2319 -103 -2315
rect -99 -2319 -60 -2315
rect -56 -2319 -25 -2315
rect -21 -2319 19 -2315
rect 23 -2319 36 -2315
rect 40 -2319 72 -2315
rect 76 -2319 93 -2315
rect 97 -2319 179 -2315
rect 183 -2319 205 -2315
rect 209 -2319 248 -2315
rect 252 -2319 283 -2315
rect 287 -2319 327 -2315
rect 331 -2319 344 -2315
rect 348 -2319 380 -2315
rect 384 -2319 401 -2315
rect 405 -2319 487 -2315
rect 491 -2319 513 -2315
rect 517 -2319 556 -2315
rect 560 -2319 591 -2315
rect 595 -2319 635 -2315
rect 639 -2319 652 -2315
rect 656 -2319 688 -2315
rect 692 -2319 709 -2315
rect 713 -2319 795 -2315
rect 799 -2319 821 -2315
rect 825 -2319 864 -2315
rect 868 -2319 899 -2315
rect 903 -2319 943 -2315
rect 947 -2319 960 -2315
rect 964 -2319 996 -2315
rect 1000 -2319 1017 -2315
rect 1021 -2319 1206 -2315
rect -1253 -2326 -814 -2322
rect -776 -2326 -198 -2322
rect -162 -2326 418 -2322
rect 453 -2326 1039 -2322
rect -1086 -2333 -505 -2329
rect -472 -2333 111 -2329
rect 144 -2333 726 -2329
rect 763 -2333 1026 -2329
rect -1454 -2359 -1309 -2355
rect -1305 -2359 -1292 -2355
rect -1288 -2359 -1062 -2355
rect -1058 -2359 -1045 -2355
rect -1041 -2359 -754 -2355
rect -750 -2359 -737 -2355
rect -733 -2359 -446 -2355
rect -442 -2359 -429 -2355
rect -425 -2359 -138 -2355
rect -134 -2359 -121 -2355
rect -117 -2359 170 -2355
rect 174 -2359 187 -2355
rect 191 -2359 478 -2355
rect 482 -2359 495 -2355
rect 499 -2359 786 -2355
rect 790 -2359 803 -2355
rect 807 -2359 1164 -2355
rect -1454 -2514 -1427 -2359
rect -1411 -2399 -1297 -2395
rect -1293 -2399 -1050 -2395
rect -1046 -2399 -742 -2395
rect -738 -2399 -434 -2395
rect -430 -2399 -126 -2395
rect -122 -2399 182 -2395
rect 186 -2399 490 -2395
rect 494 -2399 798 -2395
rect 802 -2399 1164 -2395
rect -1102 -2412 -1036 -2408
rect -789 -2412 -728 -2408
rect -486 -2412 -420 -2408
rect -176 -2412 -112 -2408
rect 130 -2412 196 -2408
rect 439 -2412 504 -2408
rect 746 -2412 812 -2408
rect 1179 -2447 1206 -2319
rect -1411 -2451 -1292 -2447
rect -1288 -2451 -1045 -2447
rect -1041 -2451 -737 -2447
rect -733 -2451 -429 -2447
rect -425 -2451 -121 -2447
rect -117 -2451 187 -2447
rect 191 -2451 495 -2447
rect 499 -2451 803 -2447
rect 807 -2451 1206 -2447
rect -1454 -2518 -1225 -2514
rect -1221 -2518 -1208 -2514
rect -1204 -2518 -1168 -2514
rect -1164 -2518 -1147 -2514
rect -1143 -2518 -1053 -2514
rect -1049 -2518 -1027 -2514
rect -1023 -2518 -1010 -2514
rect -1006 -2518 -970 -2514
rect -966 -2518 -949 -2514
rect -945 -2518 -932 -2514
rect -928 -2518 -892 -2514
rect -888 -2518 -868 -2514
rect -864 -2518 -831 -2514
rect -827 -2518 -745 -2514
rect -741 -2518 -719 -2514
rect -715 -2518 -702 -2514
rect -698 -2518 -662 -2514
rect -658 -2518 -641 -2514
rect -637 -2518 -624 -2514
rect -620 -2518 -584 -2514
rect -580 -2518 -560 -2514
rect -556 -2518 -523 -2514
rect -519 -2518 -437 -2514
rect -433 -2518 -411 -2514
rect -407 -2518 -394 -2514
rect -390 -2518 -354 -2514
rect -350 -2518 -333 -2514
rect -329 -2518 -316 -2514
rect -312 -2518 -276 -2514
rect -272 -2518 -252 -2514
rect -248 -2518 -215 -2514
rect -211 -2518 -129 -2514
rect -125 -2518 -103 -2514
rect -99 -2518 -86 -2514
rect -82 -2518 -46 -2514
rect -42 -2518 -25 -2514
rect -21 -2518 -8 -2514
rect -4 -2518 32 -2514
rect 36 -2518 56 -2514
rect 60 -2518 93 -2514
rect 97 -2518 179 -2514
rect 183 -2518 205 -2514
rect 209 -2518 222 -2514
rect 226 -2518 262 -2514
rect 266 -2518 283 -2514
rect 287 -2518 300 -2514
rect 304 -2518 340 -2514
rect 344 -2518 364 -2514
rect 368 -2518 401 -2514
rect 405 -2518 487 -2514
rect 491 -2518 513 -2514
rect 517 -2518 530 -2514
rect 534 -2518 570 -2514
rect 574 -2518 591 -2514
rect 595 -2518 608 -2514
rect 612 -2518 648 -2514
rect 652 -2518 672 -2514
rect 676 -2518 709 -2514
rect 713 -2518 795 -2514
rect 799 -2518 821 -2514
rect 825 -2518 838 -2514
rect 842 -2518 878 -2514
rect 882 -2518 899 -2514
rect 903 -2518 916 -2514
rect 920 -2518 956 -2514
rect 960 -2518 980 -2514
rect 984 -2518 1017 -2514
rect 1021 -2518 1164 -2514
rect -1454 -2646 -1427 -2518
rect -1053 -2522 -1049 -2518
rect -1027 -2522 -1023 -2518
rect -1010 -2522 -1006 -2518
rect -970 -2522 -966 -2518
rect -949 -2522 -945 -2518
rect -932 -2522 -928 -2518
rect -892 -2522 -888 -2518
rect -868 -2522 -864 -2518
rect -831 -2522 -827 -2518
rect -745 -2522 -741 -2518
rect -719 -2522 -715 -2518
rect -702 -2522 -698 -2518
rect -662 -2522 -658 -2518
rect -641 -2522 -637 -2518
rect -624 -2522 -620 -2518
rect -584 -2522 -580 -2518
rect -560 -2522 -556 -2518
rect -523 -2522 -519 -2518
rect -437 -2522 -433 -2518
rect -411 -2522 -407 -2518
rect -394 -2522 -390 -2518
rect -354 -2522 -350 -2518
rect -333 -2522 -329 -2518
rect -316 -2522 -312 -2518
rect -276 -2522 -272 -2518
rect -252 -2522 -248 -2518
rect -215 -2522 -211 -2518
rect -129 -2522 -125 -2518
rect -103 -2522 -99 -2518
rect -86 -2522 -82 -2518
rect -46 -2522 -42 -2518
rect -25 -2522 -21 -2518
rect -8 -2522 -4 -2518
rect 32 -2522 36 -2518
rect 56 -2522 60 -2518
rect 93 -2522 97 -2518
rect 179 -2522 183 -2518
rect 205 -2522 209 -2518
rect 222 -2522 226 -2518
rect 262 -2522 266 -2518
rect 283 -2522 287 -2518
rect 300 -2522 304 -2518
rect 340 -2522 344 -2518
rect 364 -2522 368 -2518
rect 401 -2522 405 -2518
rect 487 -2522 491 -2518
rect 513 -2522 517 -2518
rect 530 -2522 534 -2518
rect 570 -2522 574 -2518
rect 591 -2522 595 -2518
rect 608 -2522 612 -2518
rect 648 -2522 652 -2518
rect 672 -2522 676 -2518
rect 709 -2522 713 -2518
rect 795 -2522 799 -2518
rect 821 -2522 825 -2518
rect 838 -2522 842 -2518
rect 878 -2522 882 -2518
rect 899 -2522 903 -2518
rect 916 -2522 920 -2518
rect 956 -2522 960 -2518
rect 980 -2522 984 -2518
rect 1017 -2522 1021 -2518
rect -1047 -2537 -985 -2533
rect -981 -2537 -951 -2533
rect -903 -2537 -873 -2533
rect -739 -2537 -677 -2533
rect -673 -2537 -643 -2533
rect -595 -2537 -565 -2533
rect -431 -2537 -369 -2533
rect -365 -2537 -335 -2533
rect -287 -2537 -257 -2533
rect -123 -2537 -61 -2533
rect -57 -2537 -27 -2533
rect 21 -2537 51 -2533
rect 185 -2537 247 -2533
rect 251 -2537 281 -2533
rect 329 -2537 359 -2533
rect 493 -2537 555 -2533
rect 559 -2537 589 -2533
rect 637 -2537 667 -2533
rect 801 -2537 863 -2533
rect 867 -2537 897 -2533
rect 945 -2537 975 -2533
rect -1040 -2544 -1009 -2540
rect -732 -2544 -701 -2540
rect -424 -2544 -393 -2540
rect -116 -2544 -85 -2540
rect 192 -2544 223 -2540
rect 500 -2544 531 -2540
rect 808 -2544 839 -2540
rect -1058 -2551 -975 -2547
rect -936 -2551 -833 -2547
rect -750 -2551 -667 -2547
rect -628 -2551 -525 -2547
rect -442 -2551 -359 -2547
rect -320 -2551 -217 -2547
rect -134 -2551 -51 -2547
rect -12 -2551 91 -2547
rect 174 -2551 257 -2547
rect 296 -2551 399 -2547
rect 482 -2551 565 -2547
rect 604 -2551 707 -2547
rect 790 -2551 873 -2547
rect 912 -2551 1015 -2547
rect -1102 -2558 -1055 -2554
rect -1021 -2558 -992 -2554
rect -988 -2558 -907 -2554
rect -818 -2558 -789 -2554
rect -776 -2558 -747 -2554
rect -713 -2558 -684 -2554
rect -680 -2558 -599 -2554
rect -510 -2557 -486 -2553
rect -793 -2562 -789 -2558
rect -490 -2562 -486 -2557
rect -472 -2558 -439 -2554
rect -405 -2558 -376 -2554
rect -372 -2558 -291 -2554
rect -202 -2558 -176 -2554
rect -162 -2558 -131 -2554
rect -97 -2558 -68 -2554
rect -64 -2558 17 -2554
rect 106 -2558 130 -2554
rect 144 -2558 177 -2554
rect 211 -2558 240 -2554
rect 244 -2558 325 -2554
rect 414 -2558 439 -2554
rect 453 -2558 485 -2554
rect 519 -2558 548 -2554
rect 552 -2558 633 -2554
rect 722 -2556 739 -2552
rect -180 -2562 -176 -2558
rect 126 -2562 130 -2558
rect 435 -2562 439 -2558
rect 735 -2562 739 -2556
rect 746 -2558 793 -2554
rect 827 -2558 856 -2554
rect 860 -2558 941 -2554
rect -1230 -2567 -1173 -2563
rect -1134 -2566 -1029 -2562
rect -1014 -2566 -931 -2562
rect -910 -2566 -814 -2562
rect -793 -2566 -721 -2562
rect -706 -2566 -623 -2562
rect -602 -2566 -505 -2562
rect -490 -2566 -413 -2562
rect -398 -2566 -315 -2562
rect -294 -2566 -198 -2562
rect -180 -2566 -105 -2562
rect -90 -2566 -7 -2562
rect 14 -2566 111 -2562
rect 126 -2566 203 -2562
rect 218 -2566 301 -2562
rect 322 -2566 418 -2562
rect 435 -2566 511 -2562
rect 526 -2566 609 -2562
rect 630 -2566 726 -2562
rect 735 -2566 819 -2562
rect 834 -2566 917 -2562
rect 938 -2566 1039 -2562
rect -1253 -2574 -1223 -2570
rect -1219 -2574 -1183 -2570
rect -1179 -2574 -1163 -2570
rect -1086 -2573 -1051 -2569
rect -1032 -2573 -903 -2569
rect -789 -2573 -743 -2569
rect -724 -2573 -595 -2569
rect -486 -2573 -435 -2569
rect -416 -2573 -287 -2569
rect -176 -2573 -127 -2569
rect -108 -2573 21 -2569
rect 130 -2573 181 -2569
rect 200 -2573 329 -2569
rect 439 -2573 489 -2569
rect 508 -2573 637 -2569
rect 763 -2573 797 -2569
rect 816 -2573 945 -2569
rect -1279 -2581 -1227 -2577
rect -1223 -2581 -1197 -2577
rect -1193 -2581 -1149 -2577
rect -1025 -2580 -921 -2576
rect -917 -2580 -887 -2576
rect -717 -2580 -613 -2576
rect -609 -2580 -579 -2576
rect -409 -2580 -305 -2576
rect -301 -2580 -271 -2576
rect -101 -2580 3 -2576
rect 7 -2580 37 -2576
rect 207 -2580 311 -2576
rect 315 -2580 345 -2576
rect 515 -2580 619 -2576
rect 623 -2580 653 -2576
rect 823 -2580 927 -2576
rect 931 -2580 961 -2576
rect -1186 -2588 -1122 -2584
rect -1051 -2587 -999 -2583
rect -995 -2587 -965 -2583
rect -743 -2587 -691 -2583
rect -687 -2587 -657 -2583
rect -435 -2587 -383 -2583
rect -379 -2587 -349 -2583
rect -127 -2587 -75 -2583
rect -71 -2587 -41 -2583
rect 181 -2587 233 -2583
rect 237 -2587 267 -2583
rect 489 -2587 541 -2583
rect 545 -2587 575 -2583
rect 797 -2587 849 -2583
rect 853 -2587 883 -2583
rect -1204 -2595 -1172 -2591
rect -1006 -2595 -974 -2591
rect -1010 -2598 -1006 -2595
rect -974 -2598 -970 -2595
rect -928 -2595 -896 -2591
rect -932 -2598 -928 -2595
rect -896 -2598 -892 -2595
rect -698 -2595 -666 -2591
rect -702 -2598 -698 -2595
rect -666 -2598 -662 -2595
rect -620 -2595 -588 -2591
rect -624 -2598 -620 -2595
rect -588 -2598 -584 -2595
rect -390 -2595 -358 -2591
rect -394 -2598 -390 -2595
rect -358 -2598 -354 -2595
rect -312 -2595 -280 -2591
rect -316 -2598 -312 -2595
rect -280 -2598 -276 -2595
rect -82 -2595 -50 -2591
rect -86 -2598 -82 -2595
rect -50 -2598 -46 -2595
rect -4 -2595 28 -2591
rect -8 -2598 -4 -2595
rect 28 -2598 32 -2595
rect 226 -2595 258 -2591
rect 222 -2598 226 -2595
rect 258 -2598 262 -2595
rect 304 -2595 336 -2591
rect 300 -2598 304 -2595
rect 336 -2598 340 -2595
rect 534 -2595 566 -2591
rect 530 -2598 534 -2595
rect 566 -2598 570 -2595
rect 612 -2595 644 -2591
rect 608 -2598 612 -2595
rect 644 -2598 648 -2595
rect 842 -2595 874 -2591
rect 838 -2598 842 -2595
rect 874 -2598 878 -2595
rect 920 -2595 952 -2591
rect 916 -2598 920 -2595
rect 952 -2598 956 -2595
rect -1053 -2606 -1049 -2602
rect -1027 -2606 -1023 -2602
rect -984 -2606 -980 -2602
rect -949 -2606 -945 -2602
rect -905 -2606 -901 -2602
rect -888 -2606 -884 -2602
rect -852 -2606 -848 -2602
rect -831 -2606 -827 -2602
rect -745 -2606 -741 -2602
rect -719 -2606 -715 -2602
rect -676 -2606 -672 -2602
rect -641 -2606 -637 -2602
rect -597 -2606 -593 -2602
rect -580 -2606 -576 -2602
rect -544 -2606 -540 -2602
rect -523 -2606 -519 -2602
rect -437 -2606 -433 -2602
rect -411 -2606 -407 -2602
rect -368 -2606 -364 -2602
rect -333 -2606 -329 -2602
rect -289 -2606 -285 -2602
rect -272 -2606 -268 -2602
rect -236 -2606 -232 -2602
rect -215 -2606 -211 -2602
rect -129 -2606 -125 -2602
rect -103 -2606 -99 -2602
rect -60 -2606 -56 -2602
rect -25 -2606 -21 -2602
rect 19 -2606 23 -2602
rect 36 -2606 40 -2602
rect 72 -2606 76 -2602
rect 93 -2606 97 -2602
rect 179 -2606 183 -2602
rect 205 -2606 209 -2602
rect 248 -2606 252 -2602
rect 283 -2606 287 -2602
rect 327 -2606 331 -2602
rect 344 -2606 348 -2602
rect 380 -2606 384 -2602
rect 401 -2606 405 -2602
rect 487 -2606 491 -2602
rect 513 -2606 517 -2602
rect 556 -2606 560 -2602
rect 591 -2606 595 -2602
rect 635 -2606 639 -2602
rect 652 -2606 656 -2602
rect 688 -2606 692 -2602
rect 709 -2606 713 -2602
rect 795 -2606 799 -2602
rect 821 -2606 825 -2602
rect 864 -2606 868 -2602
rect 899 -2606 903 -2602
rect 943 -2606 947 -2602
rect 960 -2606 964 -2602
rect 996 -2606 1000 -2602
rect 1017 -2606 1021 -2602
rect 1179 -2606 1206 -2451
rect -1411 -2610 -1225 -2606
rect -1221 -2610 -1181 -2606
rect -1177 -2610 -1147 -2606
rect -1143 -2610 -1053 -2606
rect -1049 -2610 -1027 -2606
rect -1023 -2610 -984 -2606
rect -980 -2610 -949 -2606
rect -945 -2610 -905 -2606
rect -901 -2610 -888 -2606
rect -884 -2610 -852 -2606
rect -848 -2610 -831 -2606
rect -827 -2610 -745 -2606
rect -741 -2610 -719 -2606
rect -715 -2610 -676 -2606
rect -672 -2610 -641 -2606
rect -637 -2610 -597 -2606
rect -593 -2610 -580 -2606
rect -576 -2610 -544 -2606
rect -540 -2610 -523 -2606
rect -519 -2610 -437 -2606
rect -433 -2610 -411 -2606
rect -407 -2610 -368 -2606
rect -364 -2610 -333 -2606
rect -329 -2610 -289 -2606
rect -285 -2610 -272 -2606
rect -268 -2610 -236 -2606
rect -232 -2610 -215 -2606
rect -211 -2610 -129 -2606
rect -125 -2610 -103 -2606
rect -99 -2610 -60 -2606
rect -56 -2610 -25 -2606
rect -21 -2610 19 -2606
rect 23 -2610 36 -2606
rect 40 -2610 72 -2606
rect 76 -2610 93 -2606
rect 97 -2610 179 -2606
rect 183 -2610 205 -2606
rect 209 -2610 248 -2606
rect 252 -2610 283 -2606
rect 287 -2610 327 -2606
rect 331 -2610 344 -2606
rect 348 -2610 380 -2606
rect 384 -2610 401 -2606
rect 405 -2610 487 -2606
rect 491 -2610 513 -2606
rect 517 -2610 556 -2606
rect 560 -2610 591 -2606
rect 595 -2610 635 -2606
rect 639 -2610 652 -2606
rect 656 -2610 688 -2606
rect 692 -2610 709 -2606
rect 713 -2610 795 -2606
rect 799 -2610 821 -2606
rect 825 -2610 864 -2606
rect 868 -2610 899 -2606
rect 903 -2610 943 -2606
rect 947 -2610 960 -2606
rect 964 -2610 996 -2606
rect 1000 -2610 1017 -2606
rect 1021 -2610 1206 -2606
rect -1253 -2617 -814 -2613
rect -776 -2617 -198 -2613
rect -162 -2617 418 -2613
rect 453 -2617 1039 -2613
rect -1086 -2624 -505 -2620
rect -472 -2624 111 -2620
rect 144 -2624 726 -2620
rect 763 -2624 1026 -2620
rect -1454 -2650 -1309 -2646
rect -1305 -2650 -1292 -2646
rect -1288 -2650 -1062 -2646
rect -1058 -2650 -1045 -2646
rect -1041 -2650 -754 -2646
rect -750 -2650 -737 -2646
rect -733 -2650 -446 -2646
rect -442 -2650 -429 -2646
rect -425 -2650 -138 -2646
rect -134 -2650 -121 -2646
rect -117 -2650 170 -2646
rect 174 -2650 187 -2646
rect 191 -2650 478 -2646
rect 482 -2650 495 -2646
rect 499 -2650 786 -2646
rect 790 -2650 803 -2646
rect 807 -2650 1164 -2646
rect -1454 -2805 -1427 -2650
rect -1411 -2690 -1297 -2686
rect -1293 -2690 -1050 -2686
rect -1046 -2690 -742 -2686
rect -738 -2690 -434 -2686
rect -430 -2690 -126 -2686
rect -122 -2690 182 -2686
rect 186 -2690 490 -2686
rect 494 -2690 798 -2686
rect 802 -2690 1164 -2686
rect -1102 -2703 -1036 -2699
rect -789 -2703 -728 -2699
rect -486 -2703 -420 -2699
rect -176 -2703 -112 -2699
rect 130 -2703 196 -2699
rect 439 -2703 504 -2699
rect 746 -2703 812 -2699
rect 1179 -2738 1206 -2610
rect -1411 -2742 -1292 -2738
rect -1288 -2742 -1045 -2738
rect -1041 -2742 -737 -2738
rect -733 -2742 -429 -2738
rect -425 -2742 -121 -2738
rect -117 -2742 187 -2738
rect 191 -2742 495 -2738
rect 499 -2742 803 -2738
rect 807 -2742 1206 -2738
rect -1454 -2809 -1225 -2805
rect -1221 -2809 -1208 -2805
rect -1204 -2809 -1168 -2805
rect -1164 -2809 -1147 -2805
rect -1143 -2809 -1053 -2805
rect -1049 -2809 -1027 -2805
rect -1023 -2809 -1010 -2805
rect -1006 -2809 -970 -2805
rect -966 -2809 -949 -2805
rect -945 -2809 -932 -2805
rect -928 -2809 -892 -2805
rect -888 -2809 -868 -2805
rect -864 -2809 -831 -2805
rect -827 -2809 -745 -2805
rect -741 -2809 -719 -2805
rect -715 -2809 -702 -2805
rect -698 -2809 -662 -2805
rect -658 -2809 -641 -2805
rect -637 -2809 -624 -2805
rect -620 -2809 -584 -2805
rect -580 -2809 -560 -2805
rect -556 -2809 -523 -2805
rect -519 -2809 -437 -2805
rect -433 -2809 -411 -2805
rect -407 -2809 -394 -2805
rect -390 -2809 -354 -2805
rect -350 -2809 -333 -2805
rect -329 -2809 -316 -2805
rect -312 -2809 -276 -2805
rect -272 -2809 -252 -2805
rect -248 -2809 -215 -2805
rect -211 -2809 -129 -2805
rect -125 -2809 -103 -2805
rect -99 -2809 -86 -2805
rect -82 -2809 -46 -2805
rect -42 -2809 -25 -2805
rect -21 -2809 -8 -2805
rect -4 -2809 32 -2805
rect 36 -2809 56 -2805
rect 60 -2809 93 -2805
rect 97 -2809 179 -2805
rect 183 -2809 205 -2805
rect 209 -2809 222 -2805
rect 226 -2809 262 -2805
rect 266 -2809 283 -2805
rect 287 -2809 300 -2805
rect 304 -2809 340 -2805
rect 344 -2809 364 -2805
rect 368 -2809 401 -2805
rect 405 -2809 487 -2805
rect 491 -2809 513 -2805
rect 517 -2809 530 -2805
rect 534 -2809 570 -2805
rect 574 -2809 591 -2805
rect 595 -2809 608 -2805
rect 612 -2809 648 -2805
rect 652 -2809 672 -2805
rect 676 -2809 709 -2805
rect 713 -2809 795 -2805
rect 799 -2809 821 -2805
rect 825 -2809 838 -2805
rect 842 -2809 878 -2805
rect 882 -2809 899 -2805
rect 903 -2809 916 -2805
rect 920 -2809 956 -2805
rect 960 -2809 980 -2805
rect 984 -2809 1017 -2805
rect 1021 -2809 1164 -2805
rect -1454 -2937 -1427 -2809
rect -1053 -2813 -1049 -2809
rect -1027 -2813 -1023 -2809
rect -1010 -2813 -1006 -2809
rect -970 -2813 -966 -2809
rect -949 -2813 -945 -2809
rect -932 -2813 -928 -2809
rect -892 -2813 -888 -2809
rect -868 -2813 -864 -2809
rect -831 -2813 -827 -2809
rect -745 -2813 -741 -2809
rect -719 -2813 -715 -2809
rect -702 -2813 -698 -2809
rect -662 -2813 -658 -2809
rect -641 -2813 -637 -2809
rect -624 -2813 -620 -2809
rect -584 -2813 -580 -2809
rect -560 -2813 -556 -2809
rect -523 -2813 -519 -2809
rect -437 -2813 -433 -2809
rect -411 -2813 -407 -2809
rect -394 -2813 -390 -2809
rect -354 -2813 -350 -2809
rect -333 -2813 -329 -2809
rect -316 -2813 -312 -2809
rect -276 -2813 -272 -2809
rect -252 -2813 -248 -2809
rect -215 -2813 -211 -2809
rect -129 -2813 -125 -2809
rect -103 -2813 -99 -2809
rect -86 -2813 -82 -2809
rect -46 -2813 -42 -2809
rect -25 -2813 -21 -2809
rect -8 -2813 -4 -2809
rect 32 -2813 36 -2809
rect 56 -2813 60 -2809
rect 93 -2813 97 -2809
rect 179 -2813 183 -2809
rect 205 -2813 209 -2809
rect 222 -2813 226 -2809
rect 262 -2813 266 -2809
rect 283 -2813 287 -2809
rect 300 -2813 304 -2809
rect 340 -2813 344 -2809
rect 364 -2813 368 -2809
rect 401 -2813 405 -2809
rect 487 -2813 491 -2809
rect 513 -2813 517 -2809
rect 530 -2813 534 -2809
rect 570 -2813 574 -2809
rect 591 -2813 595 -2809
rect 608 -2813 612 -2809
rect 648 -2813 652 -2809
rect 672 -2813 676 -2809
rect 709 -2813 713 -2809
rect 795 -2813 799 -2809
rect 821 -2813 825 -2809
rect 838 -2813 842 -2809
rect 878 -2813 882 -2809
rect 899 -2813 903 -2809
rect 916 -2813 920 -2809
rect 956 -2813 960 -2809
rect 980 -2813 984 -2809
rect 1017 -2813 1021 -2809
rect -1047 -2828 -985 -2824
rect -981 -2828 -951 -2824
rect -903 -2828 -873 -2824
rect -739 -2828 -677 -2824
rect -673 -2828 -643 -2824
rect -595 -2828 -565 -2824
rect -431 -2828 -369 -2824
rect -365 -2828 -335 -2824
rect -287 -2828 -257 -2824
rect -123 -2828 -61 -2824
rect -57 -2828 -27 -2824
rect 21 -2828 51 -2824
rect 185 -2828 247 -2824
rect 251 -2828 281 -2824
rect 329 -2828 359 -2824
rect 493 -2828 555 -2824
rect 559 -2828 589 -2824
rect 637 -2828 667 -2824
rect 801 -2828 863 -2824
rect 867 -2828 897 -2824
rect 945 -2828 975 -2824
rect -1040 -2835 -1009 -2831
rect -732 -2835 -701 -2831
rect -424 -2835 -393 -2831
rect -116 -2835 -85 -2831
rect 192 -2835 223 -2831
rect 500 -2835 531 -2831
rect 808 -2835 839 -2831
rect -1058 -2842 -975 -2838
rect -936 -2842 -833 -2838
rect -750 -2842 -667 -2838
rect -628 -2842 -525 -2838
rect -442 -2842 -359 -2838
rect -320 -2842 -217 -2838
rect -134 -2842 -51 -2838
rect -12 -2842 91 -2838
rect 174 -2842 257 -2838
rect 296 -2842 399 -2838
rect 482 -2842 565 -2838
rect 604 -2842 707 -2838
rect 790 -2842 873 -2838
rect 912 -2842 1015 -2838
rect -1102 -2849 -1055 -2845
rect -1021 -2849 -992 -2845
rect -988 -2849 -907 -2845
rect -818 -2849 -789 -2845
rect -776 -2849 -747 -2845
rect -713 -2849 -684 -2845
rect -680 -2849 -599 -2845
rect -510 -2848 -486 -2844
rect -793 -2853 -789 -2849
rect -490 -2853 -486 -2848
rect -472 -2849 -439 -2845
rect -405 -2849 -376 -2845
rect -372 -2849 -291 -2845
rect -202 -2849 -176 -2845
rect -162 -2849 -131 -2845
rect -97 -2849 -68 -2845
rect -64 -2849 17 -2845
rect 106 -2849 130 -2845
rect 144 -2849 177 -2845
rect 211 -2849 240 -2845
rect 244 -2849 325 -2845
rect 414 -2849 439 -2845
rect 453 -2849 485 -2845
rect 519 -2849 548 -2845
rect 552 -2849 633 -2845
rect 722 -2847 739 -2843
rect -180 -2853 -176 -2849
rect 126 -2853 130 -2849
rect 435 -2853 439 -2849
rect 735 -2853 739 -2847
rect 746 -2849 793 -2845
rect 827 -2849 856 -2845
rect 860 -2849 941 -2845
rect -1230 -2858 -1173 -2854
rect -1134 -2857 -1029 -2853
rect -1014 -2857 -931 -2853
rect -910 -2857 -814 -2853
rect -793 -2857 -721 -2853
rect -706 -2857 -623 -2853
rect -602 -2857 -505 -2853
rect -490 -2857 -413 -2853
rect -398 -2857 -315 -2853
rect -294 -2857 -198 -2853
rect -180 -2857 -105 -2853
rect -90 -2857 -7 -2853
rect 14 -2857 111 -2853
rect 126 -2857 203 -2853
rect 218 -2857 301 -2853
rect 322 -2857 418 -2853
rect 435 -2857 511 -2853
rect 526 -2857 609 -2853
rect 630 -2857 726 -2853
rect 735 -2857 819 -2853
rect 834 -2857 917 -2853
rect 938 -2857 1039 -2853
rect -1253 -2865 -1223 -2861
rect -1219 -2865 -1183 -2861
rect -1179 -2865 -1163 -2861
rect -1086 -2864 -1051 -2860
rect -1032 -2864 -903 -2860
rect -789 -2864 -743 -2860
rect -724 -2864 -595 -2860
rect -486 -2864 -435 -2860
rect -416 -2864 -287 -2860
rect -176 -2864 -127 -2860
rect -108 -2864 21 -2860
rect 130 -2864 181 -2860
rect 200 -2864 329 -2860
rect 439 -2864 489 -2860
rect 508 -2864 637 -2860
rect 763 -2864 797 -2860
rect 816 -2864 945 -2860
rect -1279 -2872 -1227 -2868
rect -1223 -2872 -1197 -2868
rect -1193 -2872 -1149 -2868
rect -1025 -2871 -921 -2867
rect -917 -2871 -887 -2867
rect -717 -2871 -613 -2867
rect -609 -2871 -579 -2867
rect -409 -2871 -305 -2867
rect -301 -2871 -271 -2867
rect -101 -2871 3 -2867
rect 7 -2871 37 -2867
rect 207 -2871 311 -2867
rect 315 -2871 345 -2867
rect 515 -2871 619 -2867
rect 623 -2871 653 -2867
rect 823 -2871 927 -2867
rect 931 -2871 961 -2867
rect -1186 -2879 -1122 -2875
rect -1051 -2878 -999 -2874
rect -995 -2878 -965 -2874
rect -743 -2878 -691 -2874
rect -687 -2878 -657 -2874
rect -435 -2878 -383 -2874
rect -379 -2878 -349 -2874
rect -127 -2878 -75 -2874
rect -71 -2878 -41 -2874
rect 181 -2878 233 -2874
rect 237 -2878 267 -2874
rect 489 -2878 541 -2874
rect 545 -2878 575 -2874
rect 797 -2878 849 -2874
rect 853 -2878 883 -2874
rect -1204 -2886 -1172 -2882
rect -1006 -2886 -974 -2882
rect -1010 -2889 -1006 -2886
rect -974 -2889 -970 -2886
rect -928 -2886 -896 -2882
rect -932 -2889 -928 -2886
rect -896 -2889 -892 -2886
rect -698 -2886 -666 -2882
rect -702 -2889 -698 -2886
rect -666 -2889 -662 -2886
rect -620 -2886 -588 -2882
rect -624 -2889 -620 -2886
rect -588 -2889 -584 -2886
rect -390 -2886 -358 -2882
rect -394 -2889 -390 -2886
rect -358 -2889 -354 -2886
rect -312 -2886 -280 -2882
rect -316 -2889 -312 -2886
rect -280 -2889 -276 -2886
rect -82 -2886 -50 -2882
rect -86 -2889 -82 -2886
rect -50 -2889 -46 -2886
rect -4 -2886 28 -2882
rect -8 -2889 -4 -2886
rect 28 -2889 32 -2886
rect 226 -2886 258 -2882
rect 222 -2889 226 -2886
rect 258 -2889 262 -2886
rect 304 -2886 336 -2882
rect 300 -2889 304 -2886
rect 336 -2889 340 -2886
rect 534 -2886 566 -2882
rect 530 -2889 534 -2886
rect 566 -2889 570 -2886
rect 612 -2886 644 -2882
rect 608 -2889 612 -2886
rect 644 -2889 648 -2886
rect 842 -2886 874 -2882
rect 838 -2889 842 -2886
rect 874 -2889 878 -2886
rect 920 -2886 952 -2882
rect 916 -2889 920 -2886
rect 952 -2889 956 -2886
rect -1053 -2897 -1049 -2893
rect -1027 -2897 -1023 -2893
rect -984 -2897 -980 -2893
rect -949 -2897 -945 -2893
rect -905 -2897 -901 -2893
rect -888 -2897 -884 -2893
rect -852 -2897 -848 -2893
rect -831 -2897 -827 -2893
rect -745 -2897 -741 -2893
rect -719 -2897 -715 -2893
rect -676 -2897 -672 -2893
rect -641 -2897 -637 -2893
rect -597 -2897 -593 -2893
rect -580 -2897 -576 -2893
rect -544 -2897 -540 -2893
rect -523 -2897 -519 -2893
rect -437 -2897 -433 -2893
rect -411 -2897 -407 -2893
rect -368 -2897 -364 -2893
rect -333 -2897 -329 -2893
rect -289 -2897 -285 -2893
rect -272 -2897 -268 -2893
rect -236 -2897 -232 -2893
rect -215 -2897 -211 -2893
rect -129 -2897 -125 -2893
rect -103 -2897 -99 -2893
rect -60 -2897 -56 -2893
rect -25 -2897 -21 -2893
rect 19 -2897 23 -2893
rect 36 -2897 40 -2893
rect 72 -2897 76 -2893
rect 93 -2897 97 -2893
rect 179 -2897 183 -2893
rect 205 -2897 209 -2893
rect 248 -2897 252 -2893
rect 283 -2897 287 -2893
rect 327 -2897 331 -2893
rect 344 -2897 348 -2893
rect 380 -2897 384 -2893
rect 401 -2897 405 -2893
rect 487 -2897 491 -2893
rect 513 -2897 517 -2893
rect 556 -2897 560 -2893
rect 591 -2897 595 -2893
rect 635 -2897 639 -2893
rect 652 -2897 656 -2893
rect 688 -2897 692 -2893
rect 709 -2897 713 -2893
rect 795 -2897 799 -2893
rect 821 -2897 825 -2893
rect 864 -2897 868 -2893
rect 899 -2897 903 -2893
rect 943 -2897 947 -2893
rect 960 -2897 964 -2893
rect 996 -2897 1000 -2893
rect 1017 -2897 1021 -2893
rect 1179 -2897 1206 -2742
rect -1411 -2901 -1225 -2897
rect -1221 -2901 -1181 -2897
rect -1177 -2901 -1147 -2897
rect -1143 -2901 -1053 -2897
rect -1049 -2901 -1027 -2897
rect -1023 -2901 -984 -2897
rect -980 -2901 -949 -2897
rect -945 -2901 -905 -2897
rect -901 -2901 -888 -2897
rect -884 -2901 -852 -2897
rect -848 -2901 -831 -2897
rect -827 -2901 -745 -2897
rect -741 -2901 -719 -2897
rect -715 -2901 -676 -2897
rect -672 -2901 -641 -2897
rect -637 -2901 -597 -2897
rect -593 -2901 -580 -2897
rect -576 -2901 -544 -2897
rect -540 -2901 -523 -2897
rect -519 -2901 -437 -2897
rect -433 -2901 -411 -2897
rect -407 -2901 -368 -2897
rect -364 -2901 -333 -2897
rect -329 -2901 -289 -2897
rect -285 -2901 -272 -2897
rect -268 -2901 -236 -2897
rect -232 -2901 -215 -2897
rect -211 -2901 -129 -2897
rect -125 -2901 -103 -2897
rect -99 -2901 -60 -2897
rect -56 -2901 -25 -2897
rect -21 -2901 19 -2897
rect 23 -2901 36 -2897
rect 40 -2901 72 -2897
rect 76 -2901 93 -2897
rect 97 -2901 179 -2897
rect 183 -2901 205 -2897
rect 209 -2901 248 -2897
rect 252 -2901 283 -2897
rect 287 -2901 327 -2897
rect 331 -2901 344 -2897
rect 348 -2901 380 -2897
rect 384 -2901 401 -2897
rect 405 -2901 487 -2897
rect 491 -2901 513 -2897
rect 517 -2901 556 -2897
rect 560 -2901 591 -2897
rect 595 -2901 635 -2897
rect 639 -2901 652 -2897
rect 656 -2901 688 -2897
rect 692 -2901 709 -2897
rect 713 -2901 795 -2897
rect 799 -2901 821 -2897
rect 825 -2901 864 -2897
rect 868 -2901 899 -2897
rect 903 -2901 943 -2897
rect 947 -2901 960 -2897
rect 964 -2901 996 -2897
rect 1000 -2901 1017 -2897
rect 1021 -2901 1206 -2897
rect -1253 -2908 -814 -2904
rect -776 -2908 -198 -2904
rect -165 -2908 418 -2904
rect 451 -2908 1039 -2904
rect -1086 -2915 -505 -2911
rect -472 -2915 111 -2911
rect 143 -2915 726 -2911
rect 756 -2915 1026 -2911
rect -1454 -2941 -1309 -2937
rect -1305 -2941 -1292 -2937
rect -1288 -2941 -1062 -2937
rect -1058 -2941 -1045 -2937
rect -1041 -2941 -754 -2937
rect -750 -2941 -737 -2937
rect -733 -2941 -446 -2937
rect -442 -2941 -429 -2937
rect -425 -2941 -138 -2937
rect -134 -2941 -121 -2937
rect -117 -2941 170 -2937
rect 174 -2941 187 -2937
rect 191 -2941 478 -2937
rect 482 -2941 495 -2937
rect 499 -2941 786 -2937
rect 790 -2941 803 -2937
rect 807 -2941 1164 -2937
rect -1454 -3096 -1427 -2941
rect -1411 -2981 -1297 -2977
rect -1293 -2981 -1050 -2977
rect -1046 -2981 -742 -2977
rect -738 -2981 -434 -2977
rect -430 -2981 -126 -2977
rect -122 -2981 182 -2977
rect 186 -2981 490 -2977
rect 494 -2981 798 -2977
rect 802 -2981 1164 -2977
rect -1102 -2994 -1036 -2990
rect -789 -2994 -728 -2990
rect -486 -2994 -420 -2990
rect -176 -2994 -112 -2990
rect 130 -2994 196 -2990
rect 439 -2994 504 -2990
rect 746 -2994 812 -2990
rect 1179 -3029 1206 -2901
rect -1411 -3033 -1292 -3029
rect -1288 -3033 -1045 -3029
rect -1041 -3033 -737 -3029
rect -733 -3033 -429 -3029
rect -425 -3033 -121 -3029
rect -117 -3033 187 -3029
rect 191 -3033 495 -3029
rect 499 -3033 803 -3029
rect 807 -3033 1206 -3029
rect -1454 -3100 -1225 -3096
rect -1221 -3100 -1208 -3096
rect -1204 -3100 -1168 -3096
rect -1164 -3100 -1147 -3096
rect -1143 -3100 -1053 -3096
rect -1049 -3100 -1027 -3096
rect -1023 -3100 -1010 -3096
rect -1006 -3100 -970 -3096
rect -966 -3100 -949 -3096
rect -945 -3100 -932 -3096
rect -928 -3100 -892 -3096
rect -888 -3100 -868 -3096
rect -864 -3100 -831 -3096
rect -827 -3100 -745 -3096
rect -741 -3100 -719 -3096
rect -715 -3100 -702 -3096
rect -698 -3100 -662 -3096
rect -658 -3100 -641 -3096
rect -637 -3100 -624 -3096
rect -620 -3100 -584 -3096
rect -580 -3100 -560 -3096
rect -556 -3100 -523 -3096
rect -519 -3100 -437 -3096
rect -433 -3100 -411 -3096
rect -407 -3100 -394 -3096
rect -390 -3100 -354 -3096
rect -350 -3100 -333 -3096
rect -329 -3100 -316 -3096
rect -312 -3100 -276 -3096
rect -272 -3100 -252 -3096
rect -248 -3100 -215 -3096
rect -211 -3100 -129 -3096
rect -125 -3100 -103 -3096
rect -99 -3100 -86 -3096
rect -82 -3100 -46 -3096
rect -42 -3100 -25 -3096
rect -21 -3100 -8 -3096
rect -4 -3100 32 -3096
rect 36 -3100 56 -3096
rect 60 -3100 93 -3096
rect 97 -3100 179 -3096
rect 183 -3100 205 -3096
rect 209 -3100 222 -3096
rect 226 -3100 262 -3096
rect 266 -3100 283 -3096
rect 287 -3100 300 -3096
rect 304 -3100 340 -3096
rect 344 -3100 364 -3096
rect 368 -3100 401 -3096
rect 405 -3100 487 -3096
rect 491 -3100 513 -3096
rect 517 -3100 530 -3096
rect 534 -3100 570 -3096
rect 574 -3100 591 -3096
rect 595 -3100 608 -3096
rect 612 -3100 648 -3096
rect 652 -3100 672 -3096
rect 676 -3100 709 -3096
rect 713 -3100 795 -3096
rect 799 -3100 821 -3096
rect 825 -3100 838 -3096
rect 842 -3100 878 -3096
rect 882 -3100 899 -3096
rect 903 -3100 916 -3096
rect 920 -3100 956 -3096
rect 960 -3100 980 -3096
rect 984 -3100 1017 -3096
rect 1021 -3100 1164 -3096
rect -1053 -3104 -1049 -3100
rect -1027 -3104 -1023 -3100
rect -1010 -3104 -1006 -3100
rect -970 -3104 -966 -3100
rect -949 -3104 -945 -3100
rect -932 -3104 -928 -3100
rect -892 -3104 -888 -3100
rect -868 -3104 -864 -3100
rect -831 -3104 -827 -3100
rect -745 -3104 -741 -3100
rect -719 -3104 -715 -3100
rect -702 -3104 -698 -3100
rect -662 -3104 -658 -3100
rect -641 -3104 -637 -3100
rect -624 -3104 -620 -3100
rect -584 -3104 -580 -3100
rect -560 -3104 -556 -3100
rect -523 -3104 -519 -3100
rect -437 -3104 -433 -3100
rect -411 -3104 -407 -3100
rect -394 -3104 -390 -3100
rect -354 -3104 -350 -3100
rect -333 -3104 -329 -3100
rect -316 -3104 -312 -3100
rect -276 -3104 -272 -3100
rect -252 -3104 -248 -3100
rect -215 -3104 -211 -3100
rect -129 -3104 -125 -3100
rect -103 -3104 -99 -3100
rect -86 -3104 -82 -3100
rect -46 -3104 -42 -3100
rect -25 -3104 -21 -3100
rect -8 -3104 -4 -3100
rect 32 -3104 36 -3100
rect 56 -3104 60 -3100
rect 93 -3104 97 -3100
rect 179 -3104 183 -3100
rect 205 -3104 209 -3100
rect 222 -3104 226 -3100
rect 262 -3104 266 -3100
rect 283 -3104 287 -3100
rect 300 -3104 304 -3100
rect 340 -3104 344 -3100
rect 364 -3104 368 -3100
rect 401 -3104 405 -3100
rect 487 -3104 491 -3100
rect 513 -3104 517 -3100
rect 530 -3104 534 -3100
rect 570 -3104 574 -3100
rect 591 -3104 595 -3100
rect 608 -3104 612 -3100
rect 648 -3104 652 -3100
rect 672 -3104 676 -3100
rect 709 -3104 713 -3100
rect 795 -3104 799 -3100
rect 821 -3104 825 -3100
rect 838 -3104 842 -3100
rect 878 -3104 882 -3100
rect 899 -3104 903 -3100
rect 916 -3104 920 -3100
rect 956 -3104 960 -3100
rect 980 -3104 984 -3100
rect 1017 -3104 1021 -3100
rect -1047 -3119 -985 -3115
rect -981 -3119 -951 -3115
rect -903 -3119 -873 -3115
rect -739 -3119 -677 -3115
rect -673 -3119 -643 -3115
rect -595 -3119 -565 -3115
rect -431 -3119 -369 -3115
rect -365 -3119 -335 -3115
rect -287 -3119 -257 -3115
rect -123 -3119 -61 -3115
rect -57 -3119 -27 -3115
rect 21 -3119 51 -3115
rect 185 -3119 247 -3115
rect 251 -3119 281 -3115
rect 329 -3119 359 -3115
rect 493 -3119 555 -3115
rect 559 -3119 589 -3115
rect 637 -3119 667 -3115
rect 801 -3119 863 -3115
rect 867 -3119 897 -3115
rect 945 -3119 975 -3115
rect -1040 -3126 -1009 -3122
rect -732 -3126 -701 -3122
rect -424 -3126 -393 -3122
rect -116 -3126 -85 -3122
rect 192 -3126 223 -3122
rect 500 -3126 531 -3122
rect 808 -3126 839 -3122
rect -1058 -3133 -975 -3129
rect -936 -3133 -833 -3129
rect -750 -3133 -667 -3129
rect -628 -3133 -525 -3129
rect -442 -3133 -359 -3129
rect -320 -3133 -217 -3129
rect -134 -3133 -51 -3129
rect -12 -3133 91 -3129
rect 174 -3133 257 -3129
rect 296 -3133 399 -3129
rect 482 -3133 565 -3129
rect 604 -3133 707 -3129
rect 790 -3133 873 -3129
rect 912 -3133 1015 -3129
rect -1102 -3140 -1055 -3136
rect -1021 -3140 -992 -3136
rect -988 -3140 -907 -3136
rect -818 -3140 -789 -3136
rect -776 -3140 -747 -3136
rect -713 -3140 -684 -3136
rect -680 -3140 -599 -3136
rect -510 -3139 -486 -3135
rect -793 -3144 -789 -3140
rect -490 -3144 -486 -3139
rect -472 -3140 -439 -3136
rect -405 -3140 -376 -3136
rect -372 -3140 -291 -3136
rect -202 -3140 -176 -3136
rect -165 -3140 -131 -3136
rect -97 -3140 -68 -3136
rect -64 -3140 17 -3136
rect 106 -3140 130 -3136
rect 143 -3140 177 -3136
rect 211 -3140 240 -3136
rect 244 -3140 325 -3136
rect 414 -3140 439 -3136
rect 451 -3140 485 -3136
rect 519 -3140 548 -3136
rect 552 -3140 633 -3136
rect 722 -3138 739 -3134
rect -180 -3144 -176 -3140
rect 126 -3144 130 -3140
rect 435 -3144 439 -3140
rect 735 -3144 739 -3138
rect 746 -3140 793 -3136
rect 827 -3140 856 -3136
rect 860 -3140 941 -3136
rect -1230 -3149 -1173 -3145
rect -1134 -3148 -1029 -3144
rect -1014 -3148 -931 -3144
rect -910 -3148 -814 -3144
rect -793 -3148 -721 -3144
rect -706 -3148 -623 -3144
rect -602 -3148 -505 -3144
rect -490 -3148 -413 -3144
rect -398 -3148 -315 -3144
rect -294 -3148 -198 -3144
rect -180 -3148 -105 -3144
rect -90 -3148 -7 -3144
rect 14 -3148 111 -3144
rect 126 -3148 203 -3144
rect 218 -3148 301 -3144
rect 322 -3148 418 -3144
rect 435 -3148 511 -3144
rect 526 -3148 609 -3144
rect 630 -3148 726 -3144
rect 735 -3148 819 -3144
rect 834 -3148 917 -3144
rect 938 -3148 1034 -3144
rect -1253 -3156 -1223 -3152
rect -1219 -3156 -1183 -3152
rect -1179 -3156 -1163 -3152
rect -1086 -3155 -1051 -3151
rect -1032 -3155 -903 -3151
rect -789 -3155 -743 -3151
rect -724 -3155 -595 -3151
rect -486 -3155 -435 -3151
rect -416 -3155 -287 -3151
rect -176 -3155 -127 -3151
rect -108 -3155 21 -3151
rect 130 -3155 181 -3151
rect 200 -3155 329 -3151
rect 439 -3155 489 -3151
rect 508 -3155 637 -3151
rect 756 -3155 797 -3151
rect 816 -3155 945 -3151
rect -1279 -3163 -1227 -3159
rect -1223 -3163 -1197 -3159
rect -1193 -3163 -1149 -3159
rect -1025 -3162 -921 -3158
rect -917 -3162 -887 -3158
rect -717 -3162 -613 -3158
rect -609 -3162 -579 -3158
rect -409 -3162 -305 -3158
rect -301 -3162 -271 -3158
rect -101 -3162 3 -3158
rect 7 -3162 37 -3158
rect 207 -3162 311 -3158
rect 315 -3162 345 -3158
rect 515 -3162 619 -3158
rect 623 -3162 653 -3158
rect 823 -3162 927 -3158
rect 931 -3162 961 -3158
rect -1186 -3170 -1122 -3166
rect -1051 -3169 -999 -3165
rect -995 -3169 -965 -3165
rect -743 -3169 -691 -3165
rect -687 -3169 -657 -3165
rect -435 -3169 -383 -3165
rect -379 -3169 -349 -3165
rect -127 -3169 -75 -3165
rect -71 -3169 -41 -3165
rect 181 -3169 233 -3165
rect 237 -3169 267 -3165
rect 489 -3169 541 -3165
rect 545 -3169 575 -3165
rect 797 -3169 849 -3165
rect 853 -3169 883 -3165
rect -1204 -3177 -1172 -3173
rect -1006 -3177 -974 -3173
rect -1010 -3180 -1006 -3177
rect -974 -3180 -970 -3177
rect -928 -3177 -896 -3173
rect -932 -3180 -928 -3177
rect -896 -3180 -892 -3177
rect -698 -3177 -666 -3173
rect -702 -3180 -698 -3177
rect -666 -3180 -662 -3177
rect -620 -3177 -588 -3173
rect -624 -3180 -620 -3177
rect -588 -3180 -584 -3177
rect -390 -3177 -358 -3173
rect -394 -3180 -390 -3177
rect -358 -3180 -354 -3177
rect -312 -3177 -280 -3173
rect -316 -3180 -312 -3177
rect -280 -3180 -276 -3177
rect -82 -3177 -50 -3173
rect -86 -3180 -82 -3177
rect -50 -3180 -46 -3177
rect -4 -3177 28 -3173
rect -8 -3180 -4 -3177
rect 28 -3180 32 -3177
rect 226 -3177 258 -3173
rect 222 -3180 226 -3177
rect 258 -3180 262 -3177
rect 304 -3177 336 -3173
rect 300 -3180 304 -3177
rect 336 -3180 340 -3177
rect 534 -3177 566 -3173
rect 530 -3180 534 -3177
rect 566 -3180 570 -3177
rect 612 -3177 644 -3173
rect 608 -3180 612 -3177
rect 644 -3180 648 -3177
rect 842 -3177 874 -3173
rect 838 -3180 842 -3177
rect 874 -3180 878 -3177
rect 920 -3177 952 -3173
rect 916 -3180 920 -3177
rect 952 -3180 956 -3177
rect -1053 -3188 -1049 -3184
rect -1027 -3188 -1023 -3184
rect -984 -3188 -980 -3184
rect -949 -3188 -945 -3184
rect -905 -3188 -901 -3184
rect -888 -3188 -884 -3184
rect -852 -3188 -848 -3184
rect -831 -3188 -827 -3184
rect -745 -3188 -741 -3184
rect -719 -3188 -715 -3184
rect -676 -3188 -672 -3184
rect -641 -3188 -637 -3184
rect -597 -3188 -593 -3184
rect -580 -3188 -576 -3184
rect -544 -3188 -540 -3184
rect -523 -3188 -519 -3184
rect -437 -3188 -433 -3184
rect -411 -3188 -407 -3184
rect -368 -3188 -364 -3184
rect -333 -3188 -329 -3184
rect -289 -3188 -285 -3184
rect -272 -3188 -268 -3184
rect -236 -3188 -232 -3184
rect -215 -3188 -211 -3184
rect -129 -3188 -125 -3184
rect -103 -3188 -99 -3184
rect -60 -3188 -56 -3184
rect -25 -3188 -21 -3184
rect 19 -3188 23 -3184
rect 36 -3188 40 -3184
rect 72 -3188 76 -3184
rect 93 -3188 97 -3184
rect 179 -3188 183 -3184
rect 205 -3188 209 -3184
rect 248 -3188 252 -3184
rect 283 -3188 287 -3184
rect 327 -3188 331 -3184
rect 344 -3188 348 -3184
rect 380 -3188 384 -3184
rect 401 -3188 405 -3184
rect 487 -3188 491 -3184
rect 513 -3188 517 -3184
rect 556 -3188 560 -3184
rect 591 -3188 595 -3184
rect 635 -3188 639 -3184
rect 652 -3188 656 -3184
rect 688 -3188 692 -3184
rect 709 -3188 713 -3184
rect 795 -3188 799 -3184
rect 821 -3188 825 -3184
rect 864 -3188 868 -3184
rect 899 -3188 903 -3184
rect 943 -3188 947 -3184
rect 960 -3188 964 -3184
rect 996 -3188 1000 -3184
rect 1017 -3188 1021 -3184
rect 1179 -3188 1206 -3033
rect -1411 -3192 -1225 -3188
rect -1221 -3192 -1181 -3188
rect -1177 -3192 -1147 -3188
rect -1143 -3192 -1053 -3188
rect -1049 -3192 -1027 -3188
rect -1023 -3192 -984 -3188
rect -980 -3192 -949 -3188
rect -945 -3192 -905 -3188
rect -901 -3192 -888 -3188
rect -884 -3192 -852 -3188
rect -848 -3192 -831 -3188
rect -827 -3192 -745 -3188
rect -741 -3192 -719 -3188
rect -715 -3192 -676 -3188
rect -672 -3192 -641 -3188
rect -637 -3192 -597 -3188
rect -593 -3192 -580 -3188
rect -576 -3192 -544 -3188
rect -540 -3192 -523 -3188
rect -519 -3192 -437 -3188
rect -433 -3192 -411 -3188
rect -407 -3192 -368 -3188
rect -364 -3192 -333 -3188
rect -329 -3192 -289 -3188
rect -285 -3192 -272 -3188
rect -268 -3192 -236 -3188
rect -232 -3192 -215 -3188
rect -211 -3192 -129 -3188
rect -125 -3192 -103 -3188
rect -99 -3192 -60 -3188
rect -56 -3192 -25 -3188
rect -21 -3192 19 -3188
rect 23 -3192 36 -3188
rect 40 -3192 72 -3188
rect 76 -3192 93 -3188
rect 97 -3192 179 -3188
rect 183 -3192 205 -3188
rect 209 -3192 248 -3188
rect 252 -3192 283 -3188
rect 287 -3192 327 -3188
rect 331 -3192 344 -3188
rect 348 -3192 380 -3188
rect 384 -3192 401 -3188
rect 405 -3192 487 -3188
rect 491 -3192 513 -3188
rect 517 -3192 556 -3188
rect 560 -3192 591 -3188
rect 595 -3192 635 -3188
rect 639 -3192 652 -3188
rect 656 -3192 688 -3188
rect 692 -3192 709 -3188
rect 713 -3192 795 -3188
rect 799 -3192 821 -3188
rect 825 -3192 864 -3188
rect 868 -3192 899 -3188
rect 903 -3192 943 -3188
rect 947 -3192 960 -3188
rect 964 -3192 996 -3188
rect 1000 -3192 1017 -3188
rect 1021 -3192 1206 -3188
<< ntransistor >>
rect -1302 -1068 -1300 -1064
rect -1294 -1068 -1292 -1064
rect -1284 -1068 -1282 -1064
rect -1058 -1068 -1056 -1064
rect -1050 -1068 -1048 -1064
rect -1040 -1068 -1038 -1064
rect -749 -1068 -747 -1064
rect -741 -1068 -739 -1064
rect -731 -1068 -729 -1064
rect -441 -1068 -439 -1064
rect -433 -1068 -431 -1064
rect -423 -1068 -421 -1064
rect -134 -1068 -132 -1064
rect -126 -1068 -124 -1064
rect -116 -1068 -114 -1064
rect 175 -1068 177 -1064
rect 183 -1068 185 -1064
rect 193 -1068 195 -1064
rect 483 -1068 485 -1064
rect 491 -1068 493 -1064
rect 501 -1068 503 -1064
rect 791 -1068 793 -1064
rect 799 -1068 801 -1064
rect 809 -1068 811 -1064
rect -1304 -1218 -1302 -1214
rect -1296 -1218 -1294 -1214
rect -1286 -1218 -1284 -1214
rect -1057 -1218 -1055 -1214
rect -1049 -1218 -1047 -1214
rect -1039 -1218 -1037 -1214
rect -749 -1218 -747 -1214
rect -741 -1218 -739 -1214
rect -731 -1218 -729 -1214
rect -441 -1218 -439 -1214
rect -433 -1218 -431 -1214
rect -423 -1218 -421 -1214
rect -133 -1218 -131 -1214
rect -125 -1218 -123 -1214
rect -115 -1218 -113 -1214
rect 175 -1218 177 -1214
rect 183 -1218 185 -1214
rect 193 -1218 195 -1214
rect 483 -1218 485 -1214
rect 491 -1218 493 -1214
rect 501 -1218 503 -1214
rect 791 -1218 793 -1214
rect 799 -1218 801 -1214
rect 809 -1218 811 -1214
rect -1225 -1382 -1223 -1378
rect -1215 -1382 -1213 -1378
rect -1199 -1382 -1197 -1378
rect -1189 -1382 -1187 -1378
rect -1181 -1382 -1179 -1378
rect -1171 -1382 -1169 -1378
rect -1155 -1382 -1153 -1378
rect -1147 -1382 -1145 -1378
rect -1137 -1382 -1135 -1378
rect -1057 -1382 -1055 -1378
rect -1047 -1382 -1045 -1378
rect -1031 -1382 -1029 -1378
rect -1021 -1382 -1019 -1378
rect -1005 -1382 -1003 -1378
rect -995 -1382 -993 -1378
rect -987 -1382 -985 -1378
rect -977 -1382 -975 -1378
rect -961 -1382 -959 -1378
rect -953 -1382 -951 -1378
rect -943 -1382 -941 -1378
rect -927 -1382 -925 -1378
rect -917 -1382 -915 -1378
rect -909 -1382 -907 -1378
rect -899 -1382 -897 -1378
rect -883 -1382 -881 -1378
rect -875 -1382 -873 -1378
rect -859 -1382 -857 -1378
rect -843 -1382 -841 -1378
rect -835 -1382 -833 -1378
rect -825 -1382 -823 -1378
rect -749 -1382 -747 -1378
rect -739 -1382 -737 -1378
rect -723 -1382 -721 -1378
rect -713 -1382 -711 -1378
rect -697 -1382 -695 -1378
rect -687 -1382 -685 -1378
rect -679 -1382 -677 -1378
rect -669 -1382 -667 -1378
rect -653 -1382 -651 -1378
rect -645 -1382 -643 -1378
rect -635 -1382 -633 -1378
rect -619 -1382 -617 -1378
rect -609 -1382 -607 -1378
rect -601 -1382 -599 -1378
rect -591 -1382 -589 -1378
rect -575 -1382 -573 -1378
rect -567 -1382 -565 -1378
rect -551 -1382 -549 -1378
rect -535 -1382 -533 -1378
rect -527 -1382 -525 -1378
rect -517 -1382 -515 -1378
rect -441 -1382 -439 -1378
rect -431 -1382 -429 -1378
rect -415 -1382 -413 -1378
rect -405 -1382 -403 -1378
rect -389 -1382 -387 -1378
rect -379 -1382 -377 -1378
rect -371 -1382 -369 -1378
rect -361 -1382 -359 -1378
rect -345 -1382 -343 -1378
rect -337 -1382 -335 -1378
rect -327 -1382 -325 -1378
rect -311 -1382 -309 -1378
rect -301 -1382 -299 -1378
rect -293 -1382 -291 -1378
rect -283 -1382 -281 -1378
rect -267 -1382 -265 -1378
rect -259 -1382 -257 -1378
rect -243 -1382 -241 -1378
rect -227 -1382 -225 -1378
rect -219 -1382 -217 -1378
rect -209 -1382 -207 -1378
rect -133 -1382 -131 -1378
rect -123 -1382 -121 -1378
rect -107 -1382 -105 -1378
rect -97 -1382 -95 -1378
rect -81 -1382 -79 -1378
rect -71 -1382 -69 -1378
rect -63 -1382 -61 -1378
rect -53 -1382 -51 -1378
rect -37 -1382 -35 -1378
rect -29 -1382 -27 -1378
rect -19 -1382 -17 -1378
rect -3 -1382 -1 -1378
rect 7 -1382 9 -1378
rect 15 -1382 17 -1378
rect 25 -1382 27 -1378
rect 41 -1382 43 -1378
rect 49 -1382 51 -1378
rect 65 -1382 67 -1378
rect 81 -1382 83 -1378
rect 89 -1382 91 -1378
rect 99 -1382 101 -1378
rect 175 -1382 177 -1378
rect 185 -1382 187 -1378
rect 201 -1382 203 -1378
rect 211 -1382 213 -1378
rect 227 -1382 229 -1378
rect 237 -1382 239 -1378
rect 245 -1382 247 -1378
rect 255 -1382 257 -1378
rect 271 -1382 273 -1378
rect 279 -1382 281 -1378
rect 289 -1382 291 -1378
rect 305 -1382 307 -1378
rect 315 -1382 317 -1378
rect 323 -1382 325 -1378
rect 333 -1382 335 -1378
rect 349 -1382 351 -1378
rect 357 -1382 359 -1378
rect 373 -1382 375 -1378
rect 389 -1382 391 -1378
rect 397 -1382 399 -1378
rect 407 -1382 409 -1378
rect 483 -1382 485 -1378
rect 493 -1382 495 -1378
rect 509 -1382 511 -1378
rect 519 -1382 521 -1378
rect 535 -1382 537 -1378
rect 545 -1382 547 -1378
rect 553 -1382 555 -1378
rect 563 -1382 565 -1378
rect 579 -1382 581 -1378
rect 587 -1382 589 -1378
rect 597 -1382 599 -1378
rect 613 -1382 615 -1378
rect 623 -1382 625 -1378
rect 631 -1382 633 -1378
rect 641 -1382 643 -1378
rect 657 -1382 659 -1378
rect 665 -1382 667 -1378
rect 681 -1382 683 -1378
rect 697 -1382 699 -1378
rect 705 -1382 707 -1378
rect 715 -1382 717 -1378
rect 789 -1382 791 -1378
rect 799 -1382 801 -1378
rect 815 -1382 817 -1378
rect 825 -1382 827 -1378
rect 833 -1382 835 -1378
rect 843 -1382 845 -1378
rect 859 -1382 861 -1378
rect 867 -1382 869 -1378
rect 877 -1382 879 -1378
rect -1304 -1539 -1302 -1535
rect -1296 -1539 -1294 -1535
rect -1286 -1539 -1284 -1535
rect -1057 -1539 -1055 -1535
rect -1049 -1539 -1047 -1535
rect -1039 -1539 -1037 -1535
rect -749 -1539 -747 -1535
rect -741 -1539 -739 -1535
rect -731 -1539 -729 -1535
rect -441 -1539 -439 -1535
rect -433 -1539 -431 -1535
rect -423 -1539 -421 -1535
rect -133 -1539 -131 -1535
rect -125 -1539 -123 -1535
rect -115 -1539 -113 -1535
rect 175 -1539 177 -1535
rect 183 -1539 185 -1535
rect 193 -1539 195 -1535
rect 483 -1539 485 -1535
rect 491 -1539 493 -1535
rect 501 -1539 503 -1535
rect 791 -1539 793 -1535
rect 799 -1539 801 -1535
rect 809 -1539 811 -1535
rect -1229 -1698 -1227 -1694
rect -1219 -1698 -1217 -1694
rect -1203 -1698 -1201 -1694
rect -1193 -1698 -1191 -1694
rect -1185 -1698 -1183 -1694
rect -1175 -1698 -1173 -1694
rect -1159 -1698 -1157 -1694
rect -1151 -1698 -1149 -1694
rect -1141 -1698 -1139 -1694
rect -1057 -1698 -1055 -1694
rect -1047 -1698 -1045 -1694
rect -1031 -1698 -1029 -1694
rect -1021 -1698 -1019 -1694
rect -1005 -1698 -1003 -1694
rect -995 -1698 -993 -1694
rect -987 -1698 -985 -1694
rect -977 -1698 -975 -1694
rect -961 -1698 -959 -1694
rect -953 -1698 -951 -1694
rect -943 -1698 -941 -1694
rect -927 -1698 -925 -1694
rect -917 -1698 -915 -1694
rect -909 -1698 -907 -1694
rect -899 -1698 -897 -1694
rect -883 -1698 -881 -1694
rect -875 -1698 -873 -1694
rect -859 -1698 -857 -1694
rect -843 -1698 -841 -1694
rect -835 -1698 -833 -1694
rect -825 -1698 -823 -1694
rect -749 -1698 -747 -1694
rect -739 -1698 -737 -1694
rect -723 -1698 -721 -1694
rect -713 -1698 -711 -1694
rect -697 -1698 -695 -1694
rect -687 -1698 -685 -1694
rect -679 -1698 -677 -1694
rect -669 -1698 -667 -1694
rect -653 -1698 -651 -1694
rect -645 -1698 -643 -1694
rect -635 -1698 -633 -1694
rect -619 -1698 -617 -1694
rect -609 -1698 -607 -1694
rect -601 -1698 -599 -1694
rect -591 -1698 -589 -1694
rect -575 -1698 -573 -1694
rect -567 -1698 -565 -1694
rect -551 -1698 -549 -1694
rect -535 -1698 -533 -1694
rect -527 -1698 -525 -1694
rect -517 -1698 -515 -1694
rect -441 -1698 -439 -1694
rect -431 -1698 -429 -1694
rect -415 -1698 -413 -1694
rect -405 -1698 -403 -1694
rect -389 -1698 -387 -1694
rect -379 -1698 -377 -1694
rect -371 -1698 -369 -1694
rect -361 -1698 -359 -1694
rect -345 -1698 -343 -1694
rect -337 -1698 -335 -1694
rect -327 -1698 -325 -1694
rect -311 -1698 -309 -1694
rect -301 -1698 -299 -1694
rect -293 -1698 -291 -1694
rect -283 -1698 -281 -1694
rect -267 -1698 -265 -1694
rect -259 -1698 -257 -1694
rect -243 -1698 -241 -1694
rect -227 -1698 -225 -1694
rect -219 -1698 -217 -1694
rect -209 -1698 -207 -1694
rect -133 -1698 -131 -1694
rect -123 -1698 -121 -1694
rect -107 -1698 -105 -1694
rect -97 -1698 -95 -1694
rect -81 -1698 -79 -1694
rect -71 -1698 -69 -1694
rect -63 -1698 -61 -1694
rect -53 -1698 -51 -1694
rect -37 -1698 -35 -1694
rect -29 -1698 -27 -1694
rect -19 -1698 -17 -1694
rect -3 -1698 -1 -1694
rect 7 -1698 9 -1694
rect 15 -1698 17 -1694
rect 25 -1698 27 -1694
rect 41 -1698 43 -1694
rect 49 -1698 51 -1694
rect 65 -1698 67 -1694
rect 81 -1698 83 -1694
rect 89 -1698 91 -1694
rect 99 -1698 101 -1694
rect 175 -1698 177 -1694
rect 185 -1698 187 -1694
rect 201 -1698 203 -1694
rect 211 -1698 213 -1694
rect 227 -1698 229 -1694
rect 237 -1698 239 -1694
rect 245 -1698 247 -1694
rect 255 -1698 257 -1694
rect 271 -1698 273 -1694
rect 279 -1698 281 -1694
rect 289 -1698 291 -1694
rect 305 -1698 307 -1694
rect 315 -1698 317 -1694
rect 323 -1698 325 -1694
rect 333 -1698 335 -1694
rect 349 -1698 351 -1694
rect 357 -1698 359 -1694
rect 373 -1698 375 -1694
rect 389 -1698 391 -1694
rect 397 -1698 399 -1694
rect 407 -1698 409 -1694
rect 483 -1698 485 -1694
rect 493 -1698 495 -1694
rect 509 -1698 511 -1694
rect 519 -1698 521 -1694
rect 535 -1698 537 -1694
rect 545 -1698 547 -1694
rect 553 -1698 555 -1694
rect 563 -1698 565 -1694
rect 579 -1698 581 -1694
rect 587 -1698 589 -1694
rect 597 -1698 599 -1694
rect 613 -1698 615 -1694
rect 623 -1698 625 -1694
rect 631 -1698 633 -1694
rect 641 -1698 643 -1694
rect 657 -1698 659 -1694
rect 665 -1698 667 -1694
rect 681 -1698 683 -1694
rect 697 -1698 699 -1694
rect 705 -1698 707 -1694
rect 715 -1698 717 -1694
rect 791 -1698 793 -1694
rect 801 -1698 803 -1694
rect 817 -1698 819 -1694
rect 827 -1698 829 -1694
rect 843 -1698 845 -1694
rect 853 -1698 855 -1694
rect 861 -1698 863 -1694
rect 871 -1698 873 -1694
rect 887 -1698 889 -1694
rect 895 -1698 897 -1694
rect 905 -1698 907 -1694
rect 921 -1698 923 -1694
rect 931 -1698 933 -1694
rect 939 -1698 941 -1694
rect 949 -1698 951 -1694
rect 965 -1698 967 -1694
rect 973 -1698 975 -1694
rect 989 -1698 991 -1694
rect 1005 -1698 1007 -1694
rect 1013 -1698 1015 -1694
rect 1023 -1698 1025 -1694
rect -1304 -1830 -1302 -1826
rect -1296 -1830 -1294 -1826
rect -1286 -1830 -1284 -1826
rect -1057 -1830 -1055 -1826
rect -1049 -1830 -1047 -1826
rect -1039 -1830 -1037 -1826
rect -749 -1830 -747 -1826
rect -741 -1830 -739 -1826
rect -731 -1830 -729 -1826
rect -441 -1830 -439 -1826
rect -433 -1830 -431 -1826
rect -423 -1830 -421 -1826
rect -133 -1830 -131 -1826
rect -125 -1830 -123 -1826
rect -115 -1830 -113 -1826
rect 175 -1830 177 -1826
rect 183 -1830 185 -1826
rect 193 -1830 195 -1826
rect 483 -1830 485 -1826
rect 491 -1830 493 -1826
rect 501 -1830 503 -1826
rect 791 -1830 793 -1826
rect 799 -1830 801 -1826
rect 809 -1830 811 -1826
rect -1229 -1989 -1227 -1985
rect -1219 -1989 -1217 -1985
rect -1203 -1989 -1201 -1985
rect -1193 -1989 -1191 -1985
rect -1185 -1989 -1183 -1985
rect -1175 -1989 -1173 -1985
rect -1159 -1989 -1157 -1985
rect -1151 -1989 -1149 -1985
rect -1141 -1989 -1139 -1985
rect -1057 -1989 -1055 -1985
rect -1047 -1989 -1045 -1985
rect -1031 -1989 -1029 -1985
rect -1021 -1989 -1019 -1985
rect -1005 -1989 -1003 -1985
rect -995 -1989 -993 -1985
rect -987 -1989 -985 -1985
rect -977 -1989 -975 -1985
rect -961 -1989 -959 -1985
rect -953 -1989 -951 -1985
rect -943 -1989 -941 -1985
rect -927 -1989 -925 -1985
rect -917 -1989 -915 -1985
rect -909 -1989 -907 -1985
rect -899 -1989 -897 -1985
rect -883 -1989 -881 -1985
rect -875 -1989 -873 -1985
rect -859 -1989 -857 -1985
rect -843 -1989 -841 -1985
rect -835 -1989 -833 -1985
rect -825 -1989 -823 -1985
rect -749 -1989 -747 -1985
rect -739 -1989 -737 -1985
rect -723 -1989 -721 -1985
rect -713 -1989 -711 -1985
rect -697 -1989 -695 -1985
rect -687 -1989 -685 -1985
rect -679 -1989 -677 -1985
rect -669 -1989 -667 -1985
rect -653 -1989 -651 -1985
rect -645 -1989 -643 -1985
rect -635 -1989 -633 -1985
rect -619 -1989 -617 -1985
rect -609 -1989 -607 -1985
rect -601 -1989 -599 -1985
rect -591 -1989 -589 -1985
rect -575 -1989 -573 -1985
rect -567 -1989 -565 -1985
rect -551 -1989 -549 -1985
rect -535 -1989 -533 -1985
rect -527 -1989 -525 -1985
rect -517 -1989 -515 -1985
rect -441 -1989 -439 -1985
rect -431 -1989 -429 -1985
rect -415 -1989 -413 -1985
rect -405 -1989 -403 -1985
rect -389 -1989 -387 -1985
rect -379 -1989 -377 -1985
rect -371 -1989 -369 -1985
rect -361 -1989 -359 -1985
rect -345 -1989 -343 -1985
rect -337 -1989 -335 -1985
rect -327 -1989 -325 -1985
rect -311 -1989 -309 -1985
rect -301 -1989 -299 -1985
rect -293 -1989 -291 -1985
rect -283 -1989 -281 -1985
rect -267 -1989 -265 -1985
rect -259 -1989 -257 -1985
rect -243 -1989 -241 -1985
rect -227 -1989 -225 -1985
rect -219 -1989 -217 -1985
rect -209 -1989 -207 -1985
rect -133 -1989 -131 -1985
rect -123 -1989 -121 -1985
rect -107 -1989 -105 -1985
rect -97 -1989 -95 -1985
rect -81 -1989 -79 -1985
rect -71 -1989 -69 -1985
rect -63 -1989 -61 -1985
rect -53 -1989 -51 -1985
rect -37 -1989 -35 -1985
rect -29 -1989 -27 -1985
rect -19 -1989 -17 -1985
rect -3 -1989 -1 -1985
rect 7 -1989 9 -1985
rect 15 -1989 17 -1985
rect 25 -1989 27 -1985
rect 41 -1989 43 -1985
rect 49 -1989 51 -1985
rect 65 -1989 67 -1985
rect 81 -1989 83 -1985
rect 89 -1989 91 -1985
rect 99 -1989 101 -1985
rect 175 -1989 177 -1985
rect 185 -1989 187 -1985
rect 201 -1989 203 -1985
rect 211 -1989 213 -1985
rect 227 -1989 229 -1985
rect 237 -1989 239 -1985
rect 245 -1989 247 -1985
rect 255 -1989 257 -1985
rect 271 -1989 273 -1985
rect 279 -1989 281 -1985
rect 289 -1989 291 -1985
rect 305 -1989 307 -1985
rect 315 -1989 317 -1985
rect 323 -1989 325 -1985
rect 333 -1989 335 -1985
rect 349 -1989 351 -1985
rect 357 -1989 359 -1985
rect 373 -1989 375 -1985
rect 389 -1989 391 -1985
rect 397 -1989 399 -1985
rect 407 -1989 409 -1985
rect 483 -1989 485 -1985
rect 493 -1989 495 -1985
rect 509 -1989 511 -1985
rect 519 -1989 521 -1985
rect 535 -1989 537 -1985
rect 545 -1989 547 -1985
rect 553 -1989 555 -1985
rect 563 -1989 565 -1985
rect 579 -1989 581 -1985
rect 587 -1989 589 -1985
rect 597 -1989 599 -1985
rect 613 -1989 615 -1985
rect 623 -1989 625 -1985
rect 631 -1989 633 -1985
rect 641 -1989 643 -1985
rect 657 -1989 659 -1985
rect 665 -1989 667 -1985
rect 681 -1989 683 -1985
rect 697 -1989 699 -1985
rect 705 -1989 707 -1985
rect 715 -1989 717 -1985
rect 791 -1989 793 -1985
rect 801 -1989 803 -1985
rect 817 -1989 819 -1985
rect 827 -1989 829 -1985
rect 843 -1989 845 -1985
rect 853 -1989 855 -1985
rect 861 -1989 863 -1985
rect 871 -1989 873 -1985
rect 887 -1989 889 -1985
rect 895 -1989 897 -1985
rect 905 -1989 907 -1985
rect 921 -1989 923 -1985
rect 931 -1989 933 -1985
rect 939 -1989 941 -1985
rect 949 -1989 951 -1985
rect 965 -1989 967 -1985
rect 973 -1989 975 -1985
rect 989 -1989 991 -1985
rect 1005 -1989 1007 -1985
rect 1013 -1989 1015 -1985
rect 1023 -1989 1025 -1985
rect -1304 -2152 -1302 -2148
rect -1296 -2152 -1294 -2148
rect -1286 -2152 -1284 -2148
rect -1057 -2152 -1055 -2148
rect -1049 -2152 -1047 -2148
rect -1039 -2152 -1037 -2148
rect -749 -2152 -747 -2148
rect -741 -2152 -739 -2148
rect -731 -2152 -729 -2148
rect -441 -2152 -439 -2148
rect -433 -2152 -431 -2148
rect -423 -2152 -421 -2148
rect -133 -2152 -131 -2148
rect -125 -2152 -123 -2148
rect -115 -2152 -113 -2148
rect 175 -2152 177 -2148
rect 183 -2152 185 -2148
rect 193 -2152 195 -2148
rect 483 -2152 485 -2148
rect 491 -2152 493 -2148
rect 501 -2152 503 -2148
rect 791 -2152 793 -2148
rect 799 -2152 801 -2148
rect 809 -2152 811 -2148
rect -1229 -2311 -1227 -2307
rect -1219 -2311 -1217 -2307
rect -1203 -2311 -1201 -2307
rect -1193 -2311 -1191 -2307
rect -1185 -2311 -1183 -2307
rect -1175 -2311 -1173 -2307
rect -1159 -2311 -1157 -2307
rect -1151 -2311 -1149 -2307
rect -1141 -2311 -1139 -2307
rect -1057 -2311 -1055 -2307
rect -1047 -2311 -1045 -2307
rect -1031 -2311 -1029 -2307
rect -1021 -2311 -1019 -2307
rect -1005 -2311 -1003 -2307
rect -995 -2311 -993 -2307
rect -987 -2311 -985 -2307
rect -977 -2311 -975 -2307
rect -961 -2311 -959 -2307
rect -953 -2311 -951 -2307
rect -943 -2311 -941 -2307
rect -927 -2311 -925 -2307
rect -917 -2311 -915 -2307
rect -909 -2311 -907 -2307
rect -899 -2311 -897 -2307
rect -883 -2311 -881 -2307
rect -875 -2311 -873 -2307
rect -859 -2311 -857 -2307
rect -843 -2311 -841 -2307
rect -835 -2311 -833 -2307
rect -825 -2311 -823 -2307
rect -749 -2311 -747 -2307
rect -739 -2311 -737 -2307
rect -723 -2311 -721 -2307
rect -713 -2311 -711 -2307
rect -697 -2311 -695 -2307
rect -687 -2311 -685 -2307
rect -679 -2311 -677 -2307
rect -669 -2311 -667 -2307
rect -653 -2311 -651 -2307
rect -645 -2311 -643 -2307
rect -635 -2311 -633 -2307
rect -619 -2311 -617 -2307
rect -609 -2311 -607 -2307
rect -601 -2311 -599 -2307
rect -591 -2311 -589 -2307
rect -575 -2311 -573 -2307
rect -567 -2311 -565 -2307
rect -551 -2311 -549 -2307
rect -535 -2311 -533 -2307
rect -527 -2311 -525 -2307
rect -517 -2311 -515 -2307
rect -441 -2311 -439 -2307
rect -431 -2311 -429 -2307
rect -415 -2311 -413 -2307
rect -405 -2311 -403 -2307
rect -389 -2311 -387 -2307
rect -379 -2311 -377 -2307
rect -371 -2311 -369 -2307
rect -361 -2311 -359 -2307
rect -345 -2311 -343 -2307
rect -337 -2311 -335 -2307
rect -327 -2311 -325 -2307
rect -311 -2311 -309 -2307
rect -301 -2311 -299 -2307
rect -293 -2311 -291 -2307
rect -283 -2311 -281 -2307
rect -267 -2311 -265 -2307
rect -259 -2311 -257 -2307
rect -243 -2311 -241 -2307
rect -227 -2311 -225 -2307
rect -219 -2311 -217 -2307
rect -209 -2311 -207 -2307
rect -133 -2311 -131 -2307
rect -123 -2311 -121 -2307
rect -107 -2311 -105 -2307
rect -97 -2311 -95 -2307
rect -81 -2311 -79 -2307
rect -71 -2311 -69 -2307
rect -63 -2311 -61 -2307
rect -53 -2311 -51 -2307
rect -37 -2311 -35 -2307
rect -29 -2311 -27 -2307
rect -19 -2311 -17 -2307
rect -3 -2311 -1 -2307
rect 7 -2311 9 -2307
rect 15 -2311 17 -2307
rect 25 -2311 27 -2307
rect 41 -2311 43 -2307
rect 49 -2311 51 -2307
rect 65 -2311 67 -2307
rect 81 -2311 83 -2307
rect 89 -2311 91 -2307
rect 99 -2311 101 -2307
rect 175 -2311 177 -2307
rect 185 -2311 187 -2307
rect 201 -2311 203 -2307
rect 211 -2311 213 -2307
rect 227 -2311 229 -2307
rect 237 -2311 239 -2307
rect 245 -2311 247 -2307
rect 255 -2311 257 -2307
rect 271 -2311 273 -2307
rect 279 -2311 281 -2307
rect 289 -2311 291 -2307
rect 305 -2311 307 -2307
rect 315 -2311 317 -2307
rect 323 -2311 325 -2307
rect 333 -2311 335 -2307
rect 349 -2311 351 -2307
rect 357 -2311 359 -2307
rect 373 -2311 375 -2307
rect 389 -2311 391 -2307
rect 397 -2311 399 -2307
rect 407 -2311 409 -2307
rect 483 -2311 485 -2307
rect 493 -2311 495 -2307
rect 509 -2311 511 -2307
rect 519 -2311 521 -2307
rect 535 -2311 537 -2307
rect 545 -2311 547 -2307
rect 553 -2311 555 -2307
rect 563 -2311 565 -2307
rect 579 -2311 581 -2307
rect 587 -2311 589 -2307
rect 597 -2311 599 -2307
rect 613 -2311 615 -2307
rect 623 -2311 625 -2307
rect 631 -2311 633 -2307
rect 641 -2311 643 -2307
rect 657 -2311 659 -2307
rect 665 -2311 667 -2307
rect 681 -2311 683 -2307
rect 697 -2311 699 -2307
rect 705 -2311 707 -2307
rect 715 -2311 717 -2307
rect 791 -2311 793 -2307
rect 801 -2311 803 -2307
rect 817 -2311 819 -2307
rect 827 -2311 829 -2307
rect 843 -2311 845 -2307
rect 853 -2311 855 -2307
rect 861 -2311 863 -2307
rect 871 -2311 873 -2307
rect 887 -2311 889 -2307
rect 895 -2311 897 -2307
rect 905 -2311 907 -2307
rect 921 -2311 923 -2307
rect 931 -2311 933 -2307
rect 939 -2311 941 -2307
rect 949 -2311 951 -2307
rect 965 -2311 967 -2307
rect 973 -2311 975 -2307
rect 989 -2311 991 -2307
rect 1005 -2311 1007 -2307
rect 1013 -2311 1015 -2307
rect 1023 -2311 1025 -2307
rect -1304 -2443 -1302 -2439
rect -1296 -2443 -1294 -2439
rect -1286 -2443 -1284 -2439
rect -1057 -2443 -1055 -2439
rect -1049 -2443 -1047 -2439
rect -1039 -2443 -1037 -2439
rect -749 -2443 -747 -2439
rect -741 -2443 -739 -2439
rect -731 -2443 -729 -2439
rect -441 -2443 -439 -2439
rect -433 -2443 -431 -2439
rect -423 -2443 -421 -2439
rect -133 -2443 -131 -2439
rect -125 -2443 -123 -2439
rect -115 -2443 -113 -2439
rect 175 -2443 177 -2439
rect 183 -2443 185 -2439
rect 193 -2443 195 -2439
rect 483 -2443 485 -2439
rect 491 -2443 493 -2439
rect 501 -2443 503 -2439
rect 791 -2443 793 -2439
rect 799 -2443 801 -2439
rect 809 -2443 811 -2439
rect -1229 -2602 -1227 -2598
rect -1219 -2602 -1217 -2598
rect -1203 -2602 -1201 -2598
rect -1193 -2602 -1191 -2598
rect -1185 -2602 -1183 -2598
rect -1175 -2602 -1173 -2598
rect -1159 -2602 -1157 -2598
rect -1151 -2602 -1149 -2598
rect -1141 -2602 -1139 -2598
rect -1057 -2602 -1055 -2598
rect -1047 -2602 -1045 -2598
rect -1031 -2602 -1029 -2598
rect -1021 -2602 -1019 -2598
rect -1005 -2602 -1003 -2598
rect -995 -2602 -993 -2598
rect -987 -2602 -985 -2598
rect -977 -2602 -975 -2598
rect -961 -2602 -959 -2598
rect -953 -2602 -951 -2598
rect -943 -2602 -941 -2598
rect -927 -2602 -925 -2598
rect -917 -2602 -915 -2598
rect -909 -2602 -907 -2598
rect -899 -2602 -897 -2598
rect -883 -2602 -881 -2598
rect -875 -2602 -873 -2598
rect -859 -2602 -857 -2598
rect -843 -2602 -841 -2598
rect -835 -2602 -833 -2598
rect -825 -2602 -823 -2598
rect -749 -2602 -747 -2598
rect -739 -2602 -737 -2598
rect -723 -2602 -721 -2598
rect -713 -2602 -711 -2598
rect -697 -2602 -695 -2598
rect -687 -2602 -685 -2598
rect -679 -2602 -677 -2598
rect -669 -2602 -667 -2598
rect -653 -2602 -651 -2598
rect -645 -2602 -643 -2598
rect -635 -2602 -633 -2598
rect -619 -2602 -617 -2598
rect -609 -2602 -607 -2598
rect -601 -2602 -599 -2598
rect -591 -2602 -589 -2598
rect -575 -2602 -573 -2598
rect -567 -2602 -565 -2598
rect -551 -2602 -549 -2598
rect -535 -2602 -533 -2598
rect -527 -2602 -525 -2598
rect -517 -2602 -515 -2598
rect -441 -2602 -439 -2598
rect -431 -2602 -429 -2598
rect -415 -2602 -413 -2598
rect -405 -2602 -403 -2598
rect -389 -2602 -387 -2598
rect -379 -2602 -377 -2598
rect -371 -2602 -369 -2598
rect -361 -2602 -359 -2598
rect -345 -2602 -343 -2598
rect -337 -2602 -335 -2598
rect -327 -2602 -325 -2598
rect -311 -2602 -309 -2598
rect -301 -2602 -299 -2598
rect -293 -2602 -291 -2598
rect -283 -2602 -281 -2598
rect -267 -2602 -265 -2598
rect -259 -2602 -257 -2598
rect -243 -2602 -241 -2598
rect -227 -2602 -225 -2598
rect -219 -2602 -217 -2598
rect -209 -2602 -207 -2598
rect -133 -2602 -131 -2598
rect -123 -2602 -121 -2598
rect -107 -2602 -105 -2598
rect -97 -2602 -95 -2598
rect -81 -2602 -79 -2598
rect -71 -2602 -69 -2598
rect -63 -2602 -61 -2598
rect -53 -2602 -51 -2598
rect -37 -2602 -35 -2598
rect -29 -2602 -27 -2598
rect -19 -2602 -17 -2598
rect -3 -2602 -1 -2598
rect 7 -2602 9 -2598
rect 15 -2602 17 -2598
rect 25 -2602 27 -2598
rect 41 -2602 43 -2598
rect 49 -2602 51 -2598
rect 65 -2602 67 -2598
rect 81 -2602 83 -2598
rect 89 -2602 91 -2598
rect 99 -2602 101 -2598
rect 175 -2602 177 -2598
rect 185 -2602 187 -2598
rect 201 -2602 203 -2598
rect 211 -2602 213 -2598
rect 227 -2602 229 -2598
rect 237 -2602 239 -2598
rect 245 -2602 247 -2598
rect 255 -2602 257 -2598
rect 271 -2602 273 -2598
rect 279 -2602 281 -2598
rect 289 -2602 291 -2598
rect 305 -2602 307 -2598
rect 315 -2602 317 -2598
rect 323 -2602 325 -2598
rect 333 -2602 335 -2598
rect 349 -2602 351 -2598
rect 357 -2602 359 -2598
rect 373 -2602 375 -2598
rect 389 -2602 391 -2598
rect 397 -2602 399 -2598
rect 407 -2602 409 -2598
rect 483 -2602 485 -2598
rect 493 -2602 495 -2598
rect 509 -2602 511 -2598
rect 519 -2602 521 -2598
rect 535 -2602 537 -2598
rect 545 -2602 547 -2598
rect 553 -2602 555 -2598
rect 563 -2602 565 -2598
rect 579 -2602 581 -2598
rect 587 -2602 589 -2598
rect 597 -2602 599 -2598
rect 613 -2602 615 -2598
rect 623 -2602 625 -2598
rect 631 -2602 633 -2598
rect 641 -2602 643 -2598
rect 657 -2602 659 -2598
rect 665 -2602 667 -2598
rect 681 -2602 683 -2598
rect 697 -2602 699 -2598
rect 705 -2602 707 -2598
rect 715 -2602 717 -2598
rect 791 -2602 793 -2598
rect 801 -2602 803 -2598
rect 817 -2602 819 -2598
rect 827 -2602 829 -2598
rect 843 -2602 845 -2598
rect 853 -2602 855 -2598
rect 861 -2602 863 -2598
rect 871 -2602 873 -2598
rect 887 -2602 889 -2598
rect 895 -2602 897 -2598
rect 905 -2602 907 -2598
rect 921 -2602 923 -2598
rect 931 -2602 933 -2598
rect 939 -2602 941 -2598
rect 949 -2602 951 -2598
rect 965 -2602 967 -2598
rect 973 -2602 975 -2598
rect 989 -2602 991 -2598
rect 1005 -2602 1007 -2598
rect 1013 -2602 1015 -2598
rect 1023 -2602 1025 -2598
rect -1304 -2734 -1302 -2730
rect -1296 -2734 -1294 -2730
rect -1286 -2734 -1284 -2730
rect -1057 -2734 -1055 -2730
rect -1049 -2734 -1047 -2730
rect -1039 -2734 -1037 -2730
rect -749 -2734 -747 -2730
rect -741 -2734 -739 -2730
rect -731 -2734 -729 -2730
rect -441 -2734 -439 -2730
rect -433 -2734 -431 -2730
rect -423 -2734 -421 -2730
rect -133 -2734 -131 -2730
rect -125 -2734 -123 -2730
rect -115 -2734 -113 -2730
rect 175 -2734 177 -2730
rect 183 -2734 185 -2730
rect 193 -2734 195 -2730
rect 483 -2734 485 -2730
rect 491 -2734 493 -2730
rect 501 -2734 503 -2730
rect 791 -2734 793 -2730
rect 799 -2734 801 -2730
rect 809 -2734 811 -2730
rect -1229 -2893 -1227 -2889
rect -1219 -2893 -1217 -2889
rect -1203 -2893 -1201 -2889
rect -1193 -2893 -1191 -2889
rect -1185 -2893 -1183 -2889
rect -1175 -2893 -1173 -2889
rect -1159 -2893 -1157 -2889
rect -1151 -2893 -1149 -2889
rect -1141 -2893 -1139 -2889
rect -1057 -2893 -1055 -2889
rect -1047 -2893 -1045 -2889
rect -1031 -2893 -1029 -2889
rect -1021 -2893 -1019 -2889
rect -1005 -2893 -1003 -2889
rect -995 -2893 -993 -2889
rect -987 -2893 -985 -2889
rect -977 -2893 -975 -2889
rect -961 -2893 -959 -2889
rect -953 -2893 -951 -2889
rect -943 -2893 -941 -2889
rect -927 -2893 -925 -2889
rect -917 -2893 -915 -2889
rect -909 -2893 -907 -2889
rect -899 -2893 -897 -2889
rect -883 -2893 -881 -2889
rect -875 -2893 -873 -2889
rect -859 -2893 -857 -2889
rect -843 -2893 -841 -2889
rect -835 -2893 -833 -2889
rect -825 -2893 -823 -2889
rect -749 -2893 -747 -2889
rect -739 -2893 -737 -2889
rect -723 -2893 -721 -2889
rect -713 -2893 -711 -2889
rect -697 -2893 -695 -2889
rect -687 -2893 -685 -2889
rect -679 -2893 -677 -2889
rect -669 -2893 -667 -2889
rect -653 -2893 -651 -2889
rect -645 -2893 -643 -2889
rect -635 -2893 -633 -2889
rect -619 -2893 -617 -2889
rect -609 -2893 -607 -2889
rect -601 -2893 -599 -2889
rect -591 -2893 -589 -2889
rect -575 -2893 -573 -2889
rect -567 -2893 -565 -2889
rect -551 -2893 -549 -2889
rect -535 -2893 -533 -2889
rect -527 -2893 -525 -2889
rect -517 -2893 -515 -2889
rect -441 -2893 -439 -2889
rect -431 -2893 -429 -2889
rect -415 -2893 -413 -2889
rect -405 -2893 -403 -2889
rect -389 -2893 -387 -2889
rect -379 -2893 -377 -2889
rect -371 -2893 -369 -2889
rect -361 -2893 -359 -2889
rect -345 -2893 -343 -2889
rect -337 -2893 -335 -2889
rect -327 -2893 -325 -2889
rect -311 -2893 -309 -2889
rect -301 -2893 -299 -2889
rect -293 -2893 -291 -2889
rect -283 -2893 -281 -2889
rect -267 -2893 -265 -2889
rect -259 -2893 -257 -2889
rect -243 -2893 -241 -2889
rect -227 -2893 -225 -2889
rect -219 -2893 -217 -2889
rect -209 -2893 -207 -2889
rect -133 -2893 -131 -2889
rect -123 -2893 -121 -2889
rect -107 -2893 -105 -2889
rect -97 -2893 -95 -2889
rect -81 -2893 -79 -2889
rect -71 -2893 -69 -2889
rect -63 -2893 -61 -2889
rect -53 -2893 -51 -2889
rect -37 -2893 -35 -2889
rect -29 -2893 -27 -2889
rect -19 -2893 -17 -2889
rect -3 -2893 -1 -2889
rect 7 -2893 9 -2889
rect 15 -2893 17 -2889
rect 25 -2893 27 -2889
rect 41 -2893 43 -2889
rect 49 -2893 51 -2889
rect 65 -2893 67 -2889
rect 81 -2893 83 -2889
rect 89 -2893 91 -2889
rect 99 -2893 101 -2889
rect 175 -2893 177 -2889
rect 185 -2893 187 -2889
rect 201 -2893 203 -2889
rect 211 -2893 213 -2889
rect 227 -2893 229 -2889
rect 237 -2893 239 -2889
rect 245 -2893 247 -2889
rect 255 -2893 257 -2889
rect 271 -2893 273 -2889
rect 279 -2893 281 -2889
rect 289 -2893 291 -2889
rect 305 -2893 307 -2889
rect 315 -2893 317 -2889
rect 323 -2893 325 -2889
rect 333 -2893 335 -2889
rect 349 -2893 351 -2889
rect 357 -2893 359 -2889
rect 373 -2893 375 -2889
rect 389 -2893 391 -2889
rect 397 -2893 399 -2889
rect 407 -2893 409 -2889
rect 483 -2893 485 -2889
rect 493 -2893 495 -2889
rect 509 -2893 511 -2889
rect 519 -2893 521 -2889
rect 535 -2893 537 -2889
rect 545 -2893 547 -2889
rect 553 -2893 555 -2889
rect 563 -2893 565 -2889
rect 579 -2893 581 -2889
rect 587 -2893 589 -2889
rect 597 -2893 599 -2889
rect 613 -2893 615 -2889
rect 623 -2893 625 -2889
rect 631 -2893 633 -2889
rect 641 -2893 643 -2889
rect 657 -2893 659 -2889
rect 665 -2893 667 -2889
rect 681 -2893 683 -2889
rect 697 -2893 699 -2889
rect 705 -2893 707 -2889
rect 715 -2893 717 -2889
rect 791 -2893 793 -2889
rect 801 -2893 803 -2889
rect 817 -2893 819 -2889
rect 827 -2893 829 -2889
rect 843 -2893 845 -2889
rect 853 -2893 855 -2889
rect 861 -2893 863 -2889
rect 871 -2893 873 -2889
rect 887 -2893 889 -2889
rect 895 -2893 897 -2889
rect 905 -2893 907 -2889
rect 921 -2893 923 -2889
rect 931 -2893 933 -2889
rect 939 -2893 941 -2889
rect 949 -2893 951 -2889
rect 965 -2893 967 -2889
rect 973 -2893 975 -2889
rect 989 -2893 991 -2889
rect 1005 -2893 1007 -2889
rect 1013 -2893 1015 -2889
rect 1023 -2893 1025 -2889
rect -1304 -3025 -1302 -3021
rect -1296 -3025 -1294 -3021
rect -1286 -3025 -1284 -3021
rect -1057 -3025 -1055 -3021
rect -1049 -3025 -1047 -3021
rect -1039 -3025 -1037 -3021
rect -749 -3025 -747 -3021
rect -741 -3025 -739 -3021
rect -731 -3025 -729 -3021
rect -441 -3025 -439 -3021
rect -433 -3025 -431 -3021
rect -423 -3025 -421 -3021
rect -133 -3025 -131 -3021
rect -125 -3025 -123 -3021
rect -115 -3025 -113 -3021
rect 175 -3025 177 -3021
rect 183 -3025 185 -3021
rect 193 -3025 195 -3021
rect 483 -3025 485 -3021
rect 491 -3025 493 -3021
rect 501 -3025 503 -3021
rect 791 -3025 793 -3021
rect 799 -3025 801 -3021
rect 809 -3025 811 -3021
rect -1229 -3184 -1227 -3180
rect -1219 -3184 -1217 -3180
rect -1203 -3184 -1201 -3180
rect -1193 -3184 -1191 -3180
rect -1185 -3184 -1183 -3180
rect -1175 -3184 -1173 -3180
rect -1159 -3184 -1157 -3180
rect -1151 -3184 -1149 -3180
rect -1141 -3184 -1139 -3180
rect -1057 -3184 -1055 -3180
rect -1047 -3184 -1045 -3180
rect -1031 -3184 -1029 -3180
rect -1021 -3184 -1019 -3180
rect -1005 -3184 -1003 -3180
rect -995 -3184 -993 -3180
rect -987 -3184 -985 -3180
rect -977 -3184 -975 -3180
rect -961 -3184 -959 -3180
rect -953 -3184 -951 -3180
rect -943 -3184 -941 -3180
rect -927 -3184 -925 -3180
rect -917 -3184 -915 -3180
rect -909 -3184 -907 -3180
rect -899 -3184 -897 -3180
rect -883 -3184 -881 -3180
rect -875 -3184 -873 -3180
rect -859 -3184 -857 -3180
rect -843 -3184 -841 -3180
rect -835 -3184 -833 -3180
rect -825 -3184 -823 -3180
rect -749 -3184 -747 -3180
rect -739 -3184 -737 -3180
rect -723 -3184 -721 -3180
rect -713 -3184 -711 -3180
rect -697 -3184 -695 -3180
rect -687 -3184 -685 -3180
rect -679 -3184 -677 -3180
rect -669 -3184 -667 -3180
rect -653 -3184 -651 -3180
rect -645 -3184 -643 -3180
rect -635 -3184 -633 -3180
rect -619 -3184 -617 -3180
rect -609 -3184 -607 -3180
rect -601 -3184 -599 -3180
rect -591 -3184 -589 -3180
rect -575 -3184 -573 -3180
rect -567 -3184 -565 -3180
rect -551 -3184 -549 -3180
rect -535 -3184 -533 -3180
rect -527 -3184 -525 -3180
rect -517 -3184 -515 -3180
rect -441 -3184 -439 -3180
rect -431 -3184 -429 -3180
rect -415 -3184 -413 -3180
rect -405 -3184 -403 -3180
rect -389 -3184 -387 -3180
rect -379 -3184 -377 -3180
rect -371 -3184 -369 -3180
rect -361 -3184 -359 -3180
rect -345 -3184 -343 -3180
rect -337 -3184 -335 -3180
rect -327 -3184 -325 -3180
rect -311 -3184 -309 -3180
rect -301 -3184 -299 -3180
rect -293 -3184 -291 -3180
rect -283 -3184 -281 -3180
rect -267 -3184 -265 -3180
rect -259 -3184 -257 -3180
rect -243 -3184 -241 -3180
rect -227 -3184 -225 -3180
rect -219 -3184 -217 -3180
rect -209 -3184 -207 -3180
rect -133 -3184 -131 -3180
rect -123 -3184 -121 -3180
rect -107 -3184 -105 -3180
rect -97 -3184 -95 -3180
rect -81 -3184 -79 -3180
rect -71 -3184 -69 -3180
rect -63 -3184 -61 -3180
rect -53 -3184 -51 -3180
rect -37 -3184 -35 -3180
rect -29 -3184 -27 -3180
rect -19 -3184 -17 -3180
rect -3 -3184 -1 -3180
rect 7 -3184 9 -3180
rect 15 -3184 17 -3180
rect 25 -3184 27 -3180
rect 41 -3184 43 -3180
rect 49 -3184 51 -3180
rect 65 -3184 67 -3180
rect 81 -3184 83 -3180
rect 89 -3184 91 -3180
rect 99 -3184 101 -3180
rect 175 -3184 177 -3180
rect 185 -3184 187 -3180
rect 201 -3184 203 -3180
rect 211 -3184 213 -3180
rect 227 -3184 229 -3180
rect 237 -3184 239 -3180
rect 245 -3184 247 -3180
rect 255 -3184 257 -3180
rect 271 -3184 273 -3180
rect 279 -3184 281 -3180
rect 289 -3184 291 -3180
rect 305 -3184 307 -3180
rect 315 -3184 317 -3180
rect 323 -3184 325 -3180
rect 333 -3184 335 -3180
rect 349 -3184 351 -3180
rect 357 -3184 359 -3180
rect 373 -3184 375 -3180
rect 389 -3184 391 -3180
rect 397 -3184 399 -3180
rect 407 -3184 409 -3180
rect 483 -3184 485 -3180
rect 493 -3184 495 -3180
rect 509 -3184 511 -3180
rect 519 -3184 521 -3180
rect 535 -3184 537 -3180
rect 545 -3184 547 -3180
rect 553 -3184 555 -3180
rect 563 -3184 565 -3180
rect 579 -3184 581 -3180
rect 587 -3184 589 -3180
rect 597 -3184 599 -3180
rect 613 -3184 615 -3180
rect 623 -3184 625 -3180
rect 631 -3184 633 -3180
rect 641 -3184 643 -3180
rect 657 -3184 659 -3180
rect 665 -3184 667 -3180
rect 681 -3184 683 -3180
rect 697 -3184 699 -3180
rect 705 -3184 707 -3180
rect 715 -3184 717 -3180
rect 791 -3184 793 -3180
rect 801 -3184 803 -3180
rect 817 -3184 819 -3180
rect 827 -3184 829 -3180
rect 843 -3184 845 -3180
rect 853 -3184 855 -3180
rect 861 -3184 863 -3180
rect 871 -3184 873 -3180
rect 887 -3184 889 -3180
rect 895 -3184 897 -3180
rect 905 -3184 907 -3180
rect 921 -3184 923 -3180
rect 931 -3184 933 -3180
rect 939 -3184 941 -3180
rect 949 -3184 951 -3180
rect 965 -3184 967 -3180
rect 973 -3184 975 -3180
rect 989 -3184 991 -3180
rect 1005 -3184 1007 -3180
rect 1013 -3184 1015 -3180
rect 1023 -3184 1025 -3180
<< ptransistor >>
rect -1302 -996 -1300 -988
rect -1294 -996 -1292 -988
rect -1284 -996 -1282 -988
rect -1058 -996 -1056 -988
rect -1050 -996 -1048 -988
rect -1040 -996 -1038 -988
rect -749 -996 -747 -988
rect -741 -996 -739 -988
rect -731 -996 -729 -988
rect -441 -996 -439 -988
rect -433 -996 -431 -988
rect -423 -996 -421 -988
rect -134 -996 -132 -988
rect -126 -996 -124 -988
rect -116 -996 -114 -988
rect 175 -996 177 -988
rect 183 -996 185 -988
rect 193 -996 195 -988
rect 483 -996 485 -988
rect 491 -996 493 -988
rect 501 -996 503 -988
rect 791 -996 793 -988
rect 799 -996 801 -988
rect 809 -996 811 -988
rect -1304 -1146 -1302 -1138
rect -1296 -1146 -1294 -1138
rect -1286 -1146 -1284 -1138
rect -1057 -1146 -1055 -1138
rect -1049 -1146 -1047 -1138
rect -1039 -1146 -1037 -1138
rect -749 -1146 -747 -1138
rect -741 -1146 -739 -1138
rect -731 -1146 -729 -1138
rect -441 -1146 -439 -1138
rect -433 -1146 -431 -1138
rect -423 -1146 -421 -1138
rect -133 -1146 -131 -1138
rect -125 -1146 -123 -1138
rect -115 -1146 -113 -1138
rect 175 -1146 177 -1138
rect 183 -1146 185 -1138
rect 193 -1146 195 -1138
rect 483 -1146 485 -1138
rect 491 -1146 493 -1138
rect 501 -1146 503 -1138
rect 791 -1146 793 -1138
rect 799 -1146 801 -1138
rect 809 -1146 811 -1138
rect -1225 -1310 -1223 -1302
rect -1215 -1310 -1213 -1302
rect -1199 -1310 -1197 -1302
rect -1189 -1310 -1187 -1302
rect -1181 -1310 -1179 -1302
rect -1171 -1310 -1169 -1302
rect -1155 -1310 -1153 -1302
rect -1147 -1310 -1145 -1302
rect -1137 -1310 -1135 -1302
rect -1057 -1310 -1055 -1302
rect -1047 -1310 -1045 -1302
rect -1031 -1310 -1029 -1302
rect -1021 -1310 -1019 -1302
rect -1005 -1310 -1003 -1302
rect -995 -1310 -993 -1302
rect -987 -1310 -985 -1302
rect -977 -1310 -975 -1302
rect -961 -1310 -959 -1302
rect -953 -1310 -951 -1302
rect -943 -1310 -941 -1302
rect -927 -1310 -925 -1302
rect -917 -1310 -915 -1302
rect -909 -1310 -907 -1302
rect -899 -1310 -897 -1302
rect -883 -1310 -881 -1302
rect -875 -1310 -873 -1302
rect -859 -1310 -857 -1302
rect -843 -1310 -841 -1302
rect -835 -1310 -833 -1302
rect -825 -1310 -823 -1302
rect -749 -1310 -747 -1302
rect -739 -1310 -737 -1302
rect -723 -1310 -721 -1302
rect -713 -1310 -711 -1302
rect -697 -1310 -695 -1302
rect -687 -1310 -685 -1302
rect -679 -1310 -677 -1302
rect -669 -1310 -667 -1302
rect -653 -1310 -651 -1302
rect -645 -1310 -643 -1302
rect -635 -1310 -633 -1302
rect -619 -1310 -617 -1302
rect -609 -1310 -607 -1302
rect -601 -1310 -599 -1302
rect -591 -1310 -589 -1302
rect -575 -1310 -573 -1302
rect -567 -1310 -565 -1302
rect -551 -1310 -549 -1302
rect -535 -1310 -533 -1302
rect -527 -1310 -525 -1302
rect -517 -1310 -515 -1302
rect -441 -1310 -439 -1302
rect -431 -1310 -429 -1302
rect -415 -1310 -413 -1302
rect -405 -1310 -403 -1302
rect -389 -1310 -387 -1302
rect -379 -1310 -377 -1302
rect -371 -1310 -369 -1302
rect -361 -1310 -359 -1302
rect -345 -1310 -343 -1302
rect -337 -1310 -335 -1302
rect -327 -1310 -325 -1302
rect -311 -1310 -309 -1302
rect -301 -1310 -299 -1302
rect -293 -1310 -291 -1302
rect -283 -1310 -281 -1302
rect -267 -1310 -265 -1302
rect -259 -1310 -257 -1302
rect -243 -1310 -241 -1302
rect -227 -1310 -225 -1302
rect -219 -1310 -217 -1302
rect -209 -1310 -207 -1302
rect -133 -1310 -131 -1302
rect -123 -1310 -121 -1302
rect -107 -1310 -105 -1302
rect -97 -1310 -95 -1302
rect -81 -1310 -79 -1302
rect -71 -1310 -69 -1302
rect -63 -1310 -61 -1302
rect -53 -1310 -51 -1302
rect -37 -1310 -35 -1302
rect -29 -1310 -27 -1302
rect -19 -1310 -17 -1302
rect -3 -1310 -1 -1302
rect 7 -1310 9 -1302
rect 15 -1310 17 -1302
rect 25 -1310 27 -1302
rect 41 -1310 43 -1302
rect 49 -1310 51 -1302
rect 65 -1310 67 -1302
rect 81 -1310 83 -1302
rect 89 -1310 91 -1302
rect 99 -1310 101 -1302
rect 175 -1310 177 -1302
rect 185 -1310 187 -1302
rect 201 -1310 203 -1302
rect 211 -1310 213 -1302
rect 227 -1310 229 -1302
rect 237 -1310 239 -1302
rect 245 -1310 247 -1302
rect 255 -1310 257 -1302
rect 271 -1310 273 -1302
rect 279 -1310 281 -1302
rect 289 -1310 291 -1302
rect 305 -1310 307 -1302
rect 315 -1310 317 -1302
rect 323 -1310 325 -1302
rect 333 -1310 335 -1302
rect 349 -1310 351 -1302
rect 357 -1310 359 -1302
rect 373 -1310 375 -1302
rect 389 -1310 391 -1302
rect 397 -1310 399 -1302
rect 407 -1310 409 -1302
rect 483 -1310 485 -1302
rect 493 -1310 495 -1302
rect 509 -1310 511 -1302
rect 519 -1310 521 -1302
rect 535 -1310 537 -1302
rect 545 -1310 547 -1302
rect 553 -1310 555 -1302
rect 563 -1310 565 -1302
rect 579 -1310 581 -1302
rect 587 -1310 589 -1302
rect 597 -1310 599 -1302
rect 613 -1310 615 -1302
rect 623 -1310 625 -1302
rect 631 -1310 633 -1302
rect 641 -1310 643 -1302
rect 657 -1310 659 -1302
rect 665 -1310 667 -1302
rect 681 -1310 683 -1302
rect 697 -1310 699 -1302
rect 705 -1310 707 -1302
rect 715 -1310 717 -1302
rect 789 -1310 791 -1302
rect 799 -1310 801 -1302
rect 815 -1310 817 -1302
rect 825 -1310 827 -1302
rect 833 -1310 835 -1302
rect 843 -1310 845 -1302
rect 859 -1310 861 -1302
rect 867 -1310 869 -1302
rect 877 -1310 879 -1302
rect -1304 -1467 -1302 -1459
rect -1296 -1467 -1294 -1459
rect -1286 -1467 -1284 -1459
rect -1057 -1467 -1055 -1459
rect -1049 -1467 -1047 -1459
rect -1039 -1467 -1037 -1459
rect -749 -1467 -747 -1459
rect -741 -1467 -739 -1459
rect -731 -1467 -729 -1459
rect -441 -1467 -439 -1459
rect -433 -1467 -431 -1459
rect -423 -1467 -421 -1459
rect -133 -1467 -131 -1459
rect -125 -1467 -123 -1459
rect -115 -1467 -113 -1459
rect 175 -1467 177 -1459
rect 183 -1467 185 -1459
rect 193 -1467 195 -1459
rect 483 -1467 485 -1459
rect 491 -1467 493 -1459
rect 501 -1467 503 -1459
rect 791 -1467 793 -1459
rect 799 -1467 801 -1459
rect 809 -1467 811 -1459
rect -1229 -1626 -1227 -1618
rect -1219 -1626 -1217 -1618
rect -1203 -1626 -1201 -1618
rect -1193 -1626 -1191 -1618
rect -1185 -1626 -1183 -1618
rect -1175 -1626 -1173 -1618
rect -1159 -1626 -1157 -1618
rect -1151 -1626 -1149 -1618
rect -1141 -1626 -1139 -1618
rect -1057 -1626 -1055 -1618
rect -1047 -1626 -1045 -1618
rect -1031 -1626 -1029 -1618
rect -1021 -1626 -1019 -1618
rect -1005 -1626 -1003 -1618
rect -995 -1626 -993 -1618
rect -987 -1626 -985 -1618
rect -977 -1626 -975 -1618
rect -961 -1626 -959 -1618
rect -953 -1626 -951 -1618
rect -943 -1626 -941 -1618
rect -927 -1626 -925 -1618
rect -917 -1626 -915 -1618
rect -909 -1626 -907 -1618
rect -899 -1626 -897 -1618
rect -883 -1626 -881 -1618
rect -875 -1626 -873 -1618
rect -859 -1626 -857 -1618
rect -843 -1626 -841 -1618
rect -835 -1626 -833 -1618
rect -825 -1626 -823 -1618
rect -749 -1626 -747 -1618
rect -739 -1626 -737 -1618
rect -723 -1626 -721 -1618
rect -713 -1626 -711 -1618
rect -697 -1626 -695 -1618
rect -687 -1626 -685 -1618
rect -679 -1626 -677 -1618
rect -669 -1626 -667 -1618
rect -653 -1626 -651 -1618
rect -645 -1626 -643 -1618
rect -635 -1626 -633 -1618
rect -619 -1626 -617 -1618
rect -609 -1626 -607 -1618
rect -601 -1626 -599 -1618
rect -591 -1626 -589 -1618
rect -575 -1626 -573 -1618
rect -567 -1626 -565 -1618
rect -551 -1626 -549 -1618
rect -535 -1626 -533 -1618
rect -527 -1626 -525 -1618
rect -517 -1626 -515 -1618
rect -441 -1626 -439 -1618
rect -431 -1626 -429 -1618
rect -415 -1626 -413 -1618
rect -405 -1626 -403 -1618
rect -389 -1626 -387 -1618
rect -379 -1626 -377 -1618
rect -371 -1626 -369 -1618
rect -361 -1626 -359 -1618
rect -345 -1626 -343 -1618
rect -337 -1626 -335 -1618
rect -327 -1626 -325 -1618
rect -311 -1626 -309 -1618
rect -301 -1626 -299 -1618
rect -293 -1626 -291 -1618
rect -283 -1626 -281 -1618
rect -267 -1626 -265 -1618
rect -259 -1626 -257 -1618
rect -243 -1626 -241 -1618
rect -227 -1626 -225 -1618
rect -219 -1626 -217 -1618
rect -209 -1626 -207 -1618
rect -133 -1626 -131 -1618
rect -123 -1626 -121 -1618
rect -107 -1626 -105 -1618
rect -97 -1626 -95 -1618
rect -81 -1626 -79 -1618
rect -71 -1626 -69 -1618
rect -63 -1626 -61 -1618
rect -53 -1626 -51 -1618
rect -37 -1626 -35 -1618
rect -29 -1626 -27 -1618
rect -19 -1626 -17 -1618
rect -3 -1626 -1 -1618
rect 7 -1626 9 -1618
rect 15 -1626 17 -1618
rect 25 -1626 27 -1618
rect 41 -1626 43 -1618
rect 49 -1626 51 -1618
rect 65 -1626 67 -1618
rect 81 -1626 83 -1618
rect 89 -1626 91 -1618
rect 99 -1626 101 -1618
rect 175 -1626 177 -1618
rect 185 -1626 187 -1618
rect 201 -1626 203 -1618
rect 211 -1626 213 -1618
rect 227 -1626 229 -1618
rect 237 -1626 239 -1618
rect 245 -1626 247 -1618
rect 255 -1626 257 -1618
rect 271 -1626 273 -1618
rect 279 -1626 281 -1618
rect 289 -1626 291 -1618
rect 305 -1626 307 -1618
rect 315 -1626 317 -1618
rect 323 -1626 325 -1618
rect 333 -1626 335 -1618
rect 349 -1626 351 -1618
rect 357 -1626 359 -1618
rect 373 -1626 375 -1618
rect 389 -1626 391 -1618
rect 397 -1626 399 -1618
rect 407 -1626 409 -1618
rect 483 -1626 485 -1618
rect 493 -1626 495 -1618
rect 509 -1626 511 -1618
rect 519 -1626 521 -1618
rect 535 -1626 537 -1618
rect 545 -1626 547 -1618
rect 553 -1626 555 -1618
rect 563 -1626 565 -1618
rect 579 -1626 581 -1618
rect 587 -1626 589 -1618
rect 597 -1626 599 -1618
rect 613 -1626 615 -1618
rect 623 -1626 625 -1618
rect 631 -1626 633 -1618
rect 641 -1626 643 -1618
rect 657 -1626 659 -1618
rect 665 -1626 667 -1618
rect 681 -1626 683 -1618
rect 697 -1626 699 -1618
rect 705 -1626 707 -1618
rect 715 -1626 717 -1618
rect 791 -1626 793 -1618
rect 801 -1626 803 -1618
rect 817 -1626 819 -1618
rect 827 -1626 829 -1618
rect 843 -1626 845 -1618
rect 853 -1626 855 -1618
rect 861 -1626 863 -1618
rect 871 -1626 873 -1618
rect 887 -1626 889 -1618
rect 895 -1626 897 -1618
rect 905 -1626 907 -1618
rect 921 -1626 923 -1618
rect 931 -1626 933 -1618
rect 939 -1626 941 -1618
rect 949 -1626 951 -1618
rect 965 -1626 967 -1618
rect 973 -1626 975 -1618
rect 989 -1626 991 -1618
rect 1005 -1626 1007 -1618
rect 1013 -1626 1015 -1618
rect 1023 -1626 1025 -1618
rect -1304 -1758 -1302 -1750
rect -1296 -1758 -1294 -1750
rect -1286 -1758 -1284 -1750
rect -1057 -1758 -1055 -1750
rect -1049 -1758 -1047 -1750
rect -1039 -1758 -1037 -1750
rect -749 -1758 -747 -1750
rect -741 -1758 -739 -1750
rect -731 -1758 -729 -1750
rect -441 -1758 -439 -1750
rect -433 -1758 -431 -1750
rect -423 -1758 -421 -1750
rect -133 -1758 -131 -1750
rect -125 -1758 -123 -1750
rect -115 -1758 -113 -1750
rect 175 -1758 177 -1750
rect 183 -1758 185 -1750
rect 193 -1758 195 -1750
rect 483 -1758 485 -1750
rect 491 -1758 493 -1750
rect 501 -1758 503 -1750
rect 791 -1758 793 -1750
rect 799 -1758 801 -1750
rect 809 -1758 811 -1750
rect -1229 -1917 -1227 -1909
rect -1219 -1917 -1217 -1909
rect -1203 -1917 -1201 -1909
rect -1193 -1917 -1191 -1909
rect -1185 -1917 -1183 -1909
rect -1175 -1917 -1173 -1909
rect -1159 -1917 -1157 -1909
rect -1151 -1917 -1149 -1909
rect -1141 -1917 -1139 -1909
rect -1057 -1917 -1055 -1909
rect -1047 -1917 -1045 -1909
rect -1031 -1917 -1029 -1909
rect -1021 -1917 -1019 -1909
rect -1005 -1917 -1003 -1909
rect -995 -1917 -993 -1909
rect -987 -1917 -985 -1909
rect -977 -1917 -975 -1909
rect -961 -1917 -959 -1909
rect -953 -1917 -951 -1909
rect -943 -1917 -941 -1909
rect -927 -1917 -925 -1909
rect -917 -1917 -915 -1909
rect -909 -1917 -907 -1909
rect -899 -1917 -897 -1909
rect -883 -1917 -881 -1909
rect -875 -1917 -873 -1909
rect -859 -1917 -857 -1909
rect -843 -1917 -841 -1909
rect -835 -1917 -833 -1909
rect -825 -1917 -823 -1909
rect -749 -1917 -747 -1909
rect -739 -1917 -737 -1909
rect -723 -1917 -721 -1909
rect -713 -1917 -711 -1909
rect -697 -1917 -695 -1909
rect -687 -1917 -685 -1909
rect -679 -1917 -677 -1909
rect -669 -1917 -667 -1909
rect -653 -1917 -651 -1909
rect -645 -1917 -643 -1909
rect -635 -1917 -633 -1909
rect -619 -1917 -617 -1909
rect -609 -1917 -607 -1909
rect -601 -1917 -599 -1909
rect -591 -1917 -589 -1909
rect -575 -1917 -573 -1909
rect -567 -1917 -565 -1909
rect -551 -1917 -549 -1909
rect -535 -1917 -533 -1909
rect -527 -1917 -525 -1909
rect -517 -1917 -515 -1909
rect -441 -1917 -439 -1909
rect -431 -1917 -429 -1909
rect -415 -1917 -413 -1909
rect -405 -1917 -403 -1909
rect -389 -1917 -387 -1909
rect -379 -1917 -377 -1909
rect -371 -1917 -369 -1909
rect -361 -1917 -359 -1909
rect -345 -1917 -343 -1909
rect -337 -1917 -335 -1909
rect -327 -1917 -325 -1909
rect -311 -1917 -309 -1909
rect -301 -1917 -299 -1909
rect -293 -1917 -291 -1909
rect -283 -1917 -281 -1909
rect -267 -1917 -265 -1909
rect -259 -1917 -257 -1909
rect -243 -1917 -241 -1909
rect -227 -1917 -225 -1909
rect -219 -1917 -217 -1909
rect -209 -1917 -207 -1909
rect -133 -1917 -131 -1909
rect -123 -1917 -121 -1909
rect -107 -1917 -105 -1909
rect -97 -1917 -95 -1909
rect -81 -1917 -79 -1909
rect -71 -1917 -69 -1909
rect -63 -1917 -61 -1909
rect -53 -1917 -51 -1909
rect -37 -1917 -35 -1909
rect -29 -1917 -27 -1909
rect -19 -1917 -17 -1909
rect -3 -1917 -1 -1909
rect 7 -1917 9 -1909
rect 15 -1917 17 -1909
rect 25 -1917 27 -1909
rect 41 -1917 43 -1909
rect 49 -1917 51 -1909
rect 65 -1917 67 -1909
rect 81 -1917 83 -1909
rect 89 -1917 91 -1909
rect 99 -1917 101 -1909
rect 175 -1917 177 -1909
rect 185 -1917 187 -1909
rect 201 -1917 203 -1909
rect 211 -1917 213 -1909
rect 227 -1917 229 -1909
rect 237 -1917 239 -1909
rect 245 -1917 247 -1909
rect 255 -1917 257 -1909
rect 271 -1917 273 -1909
rect 279 -1917 281 -1909
rect 289 -1917 291 -1909
rect 305 -1917 307 -1909
rect 315 -1917 317 -1909
rect 323 -1917 325 -1909
rect 333 -1917 335 -1909
rect 349 -1917 351 -1909
rect 357 -1917 359 -1909
rect 373 -1917 375 -1909
rect 389 -1917 391 -1909
rect 397 -1917 399 -1909
rect 407 -1917 409 -1909
rect 483 -1917 485 -1909
rect 493 -1917 495 -1909
rect 509 -1917 511 -1909
rect 519 -1917 521 -1909
rect 535 -1917 537 -1909
rect 545 -1917 547 -1909
rect 553 -1917 555 -1909
rect 563 -1917 565 -1909
rect 579 -1917 581 -1909
rect 587 -1917 589 -1909
rect 597 -1917 599 -1909
rect 613 -1917 615 -1909
rect 623 -1917 625 -1909
rect 631 -1917 633 -1909
rect 641 -1917 643 -1909
rect 657 -1917 659 -1909
rect 665 -1917 667 -1909
rect 681 -1917 683 -1909
rect 697 -1917 699 -1909
rect 705 -1917 707 -1909
rect 715 -1917 717 -1909
rect 791 -1917 793 -1909
rect 801 -1917 803 -1909
rect 817 -1917 819 -1909
rect 827 -1917 829 -1909
rect 843 -1917 845 -1909
rect 853 -1917 855 -1909
rect 861 -1917 863 -1909
rect 871 -1917 873 -1909
rect 887 -1917 889 -1909
rect 895 -1917 897 -1909
rect 905 -1917 907 -1909
rect 921 -1917 923 -1909
rect 931 -1917 933 -1909
rect 939 -1917 941 -1909
rect 949 -1917 951 -1909
rect 965 -1917 967 -1909
rect 973 -1917 975 -1909
rect 989 -1917 991 -1909
rect 1005 -1917 1007 -1909
rect 1013 -1917 1015 -1909
rect 1023 -1917 1025 -1909
rect -1304 -2080 -1302 -2072
rect -1296 -2080 -1294 -2072
rect -1286 -2080 -1284 -2072
rect -1057 -2080 -1055 -2072
rect -1049 -2080 -1047 -2072
rect -1039 -2080 -1037 -2072
rect -749 -2080 -747 -2072
rect -741 -2080 -739 -2072
rect -731 -2080 -729 -2072
rect -441 -2080 -439 -2072
rect -433 -2080 -431 -2072
rect -423 -2080 -421 -2072
rect -133 -2080 -131 -2072
rect -125 -2080 -123 -2072
rect -115 -2080 -113 -2072
rect 175 -2080 177 -2072
rect 183 -2080 185 -2072
rect 193 -2080 195 -2072
rect 483 -2080 485 -2072
rect 491 -2080 493 -2072
rect 501 -2080 503 -2072
rect 791 -2080 793 -2072
rect 799 -2080 801 -2072
rect 809 -2080 811 -2072
rect -1229 -2239 -1227 -2231
rect -1219 -2239 -1217 -2231
rect -1203 -2239 -1201 -2231
rect -1193 -2239 -1191 -2231
rect -1185 -2239 -1183 -2231
rect -1175 -2239 -1173 -2231
rect -1159 -2239 -1157 -2231
rect -1151 -2239 -1149 -2231
rect -1141 -2239 -1139 -2231
rect -1057 -2239 -1055 -2231
rect -1047 -2239 -1045 -2231
rect -1031 -2239 -1029 -2231
rect -1021 -2239 -1019 -2231
rect -1005 -2239 -1003 -2231
rect -995 -2239 -993 -2231
rect -987 -2239 -985 -2231
rect -977 -2239 -975 -2231
rect -961 -2239 -959 -2231
rect -953 -2239 -951 -2231
rect -943 -2239 -941 -2231
rect -927 -2239 -925 -2231
rect -917 -2239 -915 -2231
rect -909 -2239 -907 -2231
rect -899 -2239 -897 -2231
rect -883 -2239 -881 -2231
rect -875 -2239 -873 -2231
rect -859 -2239 -857 -2231
rect -843 -2239 -841 -2231
rect -835 -2239 -833 -2231
rect -825 -2239 -823 -2231
rect -749 -2239 -747 -2231
rect -739 -2239 -737 -2231
rect -723 -2239 -721 -2231
rect -713 -2239 -711 -2231
rect -697 -2239 -695 -2231
rect -687 -2239 -685 -2231
rect -679 -2239 -677 -2231
rect -669 -2239 -667 -2231
rect -653 -2239 -651 -2231
rect -645 -2239 -643 -2231
rect -635 -2239 -633 -2231
rect -619 -2239 -617 -2231
rect -609 -2239 -607 -2231
rect -601 -2239 -599 -2231
rect -591 -2239 -589 -2231
rect -575 -2239 -573 -2231
rect -567 -2239 -565 -2231
rect -551 -2239 -549 -2231
rect -535 -2239 -533 -2231
rect -527 -2239 -525 -2231
rect -517 -2239 -515 -2231
rect -441 -2239 -439 -2231
rect -431 -2239 -429 -2231
rect -415 -2239 -413 -2231
rect -405 -2239 -403 -2231
rect -389 -2239 -387 -2231
rect -379 -2239 -377 -2231
rect -371 -2239 -369 -2231
rect -361 -2239 -359 -2231
rect -345 -2239 -343 -2231
rect -337 -2239 -335 -2231
rect -327 -2239 -325 -2231
rect -311 -2239 -309 -2231
rect -301 -2239 -299 -2231
rect -293 -2239 -291 -2231
rect -283 -2239 -281 -2231
rect -267 -2239 -265 -2231
rect -259 -2239 -257 -2231
rect -243 -2239 -241 -2231
rect -227 -2239 -225 -2231
rect -219 -2239 -217 -2231
rect -209 -2239 -207 -2231
rect -133 -2239 -131 -2231
rect -123 -2239 -121 -2231
rect -107 -2239 -105 -2231
rect -97 -2239 -95 -2231
rect -81 -2239 -79 -2231
rect -71 -2239 -69 -2231
rect -63 -2239 -61 -2231
rect -53 -2239 -51 -2231
rect -37 -2239 -35 -2231
rect -29 -2239 -27 -2231
rect -19 -2239 -17 -2231
rect -3 -2239 -1 -2231
rect 7 -2239 9 -2231
rect 15 -2239 17 -2231
rect 25 -2239 27 -2231
rect 41 -2239 43 -2231
rect 49 -2239 51 -2231
rect 65 -2239 67 -2231
rect 81 -2239 83 -2231
rect 89 -2239 91 -2231
rect 99 -2239 101 -2231
rect 175 -2239 177 -2231
rect 185 -2239 187 -2231
rect 201 -2239 203 -2231
rect 211 -2239 213 -2231
rect 227 -2239 229 -2231
rect 237 -2239 239 -2231
rect 245 -2239 247 -2231
rect 255 -2239 257 -2231
rect 271 -2239 273 -2231
rect 279 -2239 281 -2231
rect 289 -2239 291 -2231
rect 305 -2239 307 -2231
rect 315 -2239 317 -2231
rect 323 -2239 325 -2231
rect 333 -2239 335 -2231
rect 349 -2239 351 -2231
rect 357 -2239 359 -2231
rect 373 -2239 375 -2231
rect 389 -2239 391 -2231
rect 397 -2239 399 -2231
rect 407 -2239 409 -2231
rect 483 -2239 485 -2231
rect 493 -2239 495 -2231
rect 509 -2239 511 -2231
rect 519 -2239 521 -2231
rect 535 -2239 537 -2231
rect 545 -2239 547 -2231
rect 553 -2239 555 -2231
rect 563 -2239 565 -2231
rect 579 -2239 581 -2231
rect 587 -2239 589 -2231
rect 597 -2239 599 -2231
rect 613 -2239 615 -2231
rect 623 -2239 625 -2231
rect 631 -2239 633 -2231
rect 641 -2239 643 -2231
rect 657 -2239 659 -2231
rect 665 -2239 667 -2231
rect 681 -2239 683 -2231
rect 697 -2239 699 -2231
rect 705 -2239 707 -2231
rect 715 -2239 717 -2231
rect 791 -2239 793 -2231
rect 801 -2239 803 -2231
rect 817 -2239 819 -2231
rect 827 -2239 829 -2231
rect 843 -2239 845 -2231
rect 853 -2239 855 -2231
rect 861 -2239 863 -2231
rect 871 -2239 873 -2231
rect 887 -2239 889 -2231
rect 895 -2239 897 -2231
rect 905 -2239 907 -2231
rect 921 -2239 923 -2231
rect 931 -2239 933 -2231
rect 939 -2239 941 -2231
rect 949 -2239 951 -2231
rect 965 -2239 967 -2231
rect 973 -2239 975 -2231
rect 989 -2239 991 -2231
rect 1005 -2239 1007 -2231
rect 1013 -2239 1015 -2231
rect 1023 -2239 1025 -2231
rect -1304 -2371 -1302 -2363
rect -1296 -2371 -1294 -2363
rect -1286 -2371 -1284 -2363
rect -1057 -2371 -1055 -2363
rect -1049 -2371 -1047 -2363
rect -1039 -2371 -1037 -2363
rect -749 -2371 -747 -2363
rect -741 -2371 -739 -2363
rect -731 -2371 -729 -2363
rect -441 -2371 -439 -2363
rect -433 -2371 -431 -2363
rect -423 -2371 -421 -2363
rect -133 -2371 -131 -2363
rect -125 -2371 -123 -2363
rect -115 -2371 -113 -2363
rect 175 -2371 177 -2363
rect 183 -2371 185 -2363
rect 193 -2371 195 -2363
rect 483 -2371 485 -2363
rect 491 -2371 493 -2363
rect 501 -2371 503 -2363
rect 791 -2371 793 -2363
rect 799 -2371 801 -2363
rect 809 -2371 811 -2363
rect -1229 -2530 -1227 -2522
rect -1219 -2530 -1217 -2522
rect -1203 -2530 -1201 -2522
rect -1193 -2530 -1191 -2522
rect -1185 -2530 -1183 -2522
rect -1175 -2530 -1173 -2522
rect -1159 -2530 -1157 -2522
rect -1151 -2530 -1149 -2522
rect -1141 -2530 -1139 -2522
rect -1057 -2530 -1055 -2522
rect -1047 -2530 -1045 -2522
rect -1031 -2530 -1029 -2522
rect -1021 -2530 -1019 -2522
rect -1005 -2530 -1003 -2522
rect -995 -2530 -993 -2522
rect -987 -2530 -985 -2522
rect -977 -2530 -975 -2522
rect -961 -2530 -959 -2522
rect -953 -2530 -951 -2522
rect -943 -2530 -941 -2522
rect -927 -2530 -925 -2522
rect -917 -2530 -915 -2522
rect -909 -2530 -907 -2522
rect -899 -2530 -897 -2522
rect -883 -2530 -881 -2522
rect -875 -2530 -873 -2522
rect -859 -2530 -857 -2522
rect -843 -2530 -841 -2522
rect -835 -2530 -833 -2522
rect -825 -2530 -823 -2522
rect -749 -2530 -747 -2522
rect -739 -2530 -737 -2522
rect -723 -2530 -721 -2522
rect -713 -2530 -711 -2522
rect -697 -2530 -695 -2522
rect -687 -2530 -685 -2522
rect -679 -2530 -677 -2522
rect -669 -2530 -667 -2522
rect -653 -2530 -651 -2522
rect -645 -2530 -643 -2522
rect -635 -2530 -633 -2522
rect -619 -2530 -617 -2522
rect -609 -2530 -607 -2522
rect -601 -2530 -599 -2522
rect -591 -2530 -589 -2522
rect -575 -2530 -573 -2522
rect -567 -2530 -565 -2522
rect -551 -2530 -549 -2522
rect -535 -2530 -533 -2522
rect -527 -2530 -525 -2522
rect -517 -2530 -515 -2522
rect -441 -2530 -439 -2522
rect -431 -2530 -429 -2522
rect -415 -2530 -413 -2522
rect -405 -2530 -403 -2522
rect -389 -2530 -387 -2522
rect -379 -2530 -377 -2522
rect -371 -2530 -369 -2522
rect -361 -2530 -359 -2522
rect -345 -2530 -343 -2522
rect -337 -2530 -335 -2522
rect -327 -2530 -325 -2522
rect -311 -2530 -309 -2522
rect -301 -2530 -299 -2522
rect -293 -2530 -291 -2522
rect -283 -2530 -281 -2522
rect -267 -2530 -265 -2522
rect -259 -2530 -257 -2522
rect -243 -2530 -241 -2522
rect -227 -2530 -225 -2522
rect -219 -2530 -217 -2522
rect -209 -2530 -207 -2522
rect -133 -2530 -131 -2522
rect -123 -2530 -121 -2522
rect -107 -2530 -105 -2522
rect -97 -2530 -95 -2522
rect -81 -2530 -79 -2522
rect -71 -2530 -69 -2522
rect -63 -2530 -61 -2522
rect -53 -2530 -51 -2522
rect -37 -2530 -35 -2522
rect -29 -2530 -27 -2522
rect -19 -2530 -17 -2522
rect -3 -2530 -1 -2522
rect 7 -2530 9 -2522
rect 15 -2530 17 -2522
rect 25 -2530 27 -2522
rect 41 -2530 43 -2522
rect 49 -2530 51 -2522
rect 65 -2530 67 -2522
rect 81 -2530 83 -2522
rect 89 -2530 91 -2522
rect 99 -2530 101 -2522
rect 175 -2530 177 -2522
rect 185 -2530 187 -2522
rect 201 -2530 203 -2522
rect 211 -2530 213 -2522
rect 227 -2530 229 -2522
rect 237 -2530 239 -2522
rect 245 -2530 247 -2522
rect 255 -2530 257 -2522
rect 271 -2530 273 -2522
rect 279 -2530 281 -2522
rect 289 -2530 291 -2522
rect 305 -2530 307 -2522
rect 315 -2530 317 -2522
rect 323 -2530 325 -2522
rect 333 -2530 335 -2522
rect 349 -2530 351 -2522
rect 357 -2530 359 -2522
rect 373 -2530 375 -2522
rect 389 -2530 391 -2522
rect 397 -2530 399 -2522
rect 407 -2530 409 -2522
rect 483 -2530 485 -2522
rect 493 -2530 495 -2522
rect 509 -2530 511 -2522
rect 519 -2530 521 -2522
rect 535 -2530 537 -2522
rect 545 -2530 547 -2522
rect 553 -2530 555 -2522
rect 563 -2530 565 -2522
rect 579 -2530 581 -2522
rect 587 -2530 589 -2522
rect 597 -2530 599 -2522
rect 613 -2530 615 -2522
rect 623 -2530 625 -2522
rect 631 -2530 633 -2522
rect 641 -2530 643 -2522
rect 657 -2530 659 -2522
rect 665 -2530 667 -2522
rect 681 -2530 683 -2522
rect 697 -2530 699 -2522
rect 705 -2530 707 -2522
rect 715 -2530 717 -2522
rect 791 -2530 793 -2522
rect 801 -2530 803 -2522
rect 817 -2530 819 -2522
rect 827 -2530 829 -2522
rect 843 -2530 845 -2522
rect 853 -2530 855 -2522
rect 861 -2530 863 -2522
rect 871 -2530 873 -2522
rect 887 -2530 889 -2522
rect 895 -2530 897 -2522
rect 905 -2530 907 -2522
rect 921 -2530 923 -2522
rect 931 -2530 933 -2522
rect 939 -2530 941 -2522
rect 949 -2530 951 -2522
rect 965 -2530 967 -2522
rect 973 -2530 975 -2522
rect 989 -2530 991 -2522
rect 1005 -2530 1007 -2522
rect 1013 -2530 1015 -2522
rect 1023 -2530 1025 -2522
rect -1304 -2662 -1302 -2654
rect -1296 -2662 -1294 -2654
rect -1286 -2662 -1284 -2654
rect -1057 -2662 -1055 -2654
rect -1049 -2662 -1047 -2654
rect -1039 -2662 -1037 -2654
rect -749 -2662 -747 -2654
rect -741 -2662 -739 -2654
rect -731 -2662 -729 -2654
rect -441 -2662 -439 -2654
rect -433 -2662 -431 -2654
rect -423 -2662 -421 -2654
rect -133 -2662 -131 -2654
rect -125 -2662 -123 -2654
rect -115 -2662 -113 -2654
rect 175 -2662 177 -2654
rect 183 -2662 185 -2654
rect 193 -2662 195 -2654
rect 483 -2662 485 -2654
rect 491 -2662 493 -2654
rect 501 -2662 503 -2654
rect 791 -2662 793 -2654
rect 799 -2662 801 -2654
rect 809 -2662 811 -2654
rect -1229 -2821 -1227 -2813
rect -1219 -2821 -1217 -2813
rect -1203 -2821 -1201 -2813
rect -1193 -2821 -1191 -2813
rect -1185 -2821 -1183 -2813
rect -1175 -2821 -1173 -2813
rect -1159 -2821 -1157 -2813
rect -1151 -2821 -1149 -2813
rect -1141 -2821 -1139 -2813
rect -1057 -2821 -1055 -2813
rect -1047 -2821 -1045 -2813
rect -1031 -2821 -1029 -2813
rect -1021 -2821 -1019 -2813
rect -1005 -2821 -1003 -2813
rect -995 -2821 -993 -2813
rect -987 -2821 -985 -2813
rect -977 -2821 -975 -2813
rect -961 -2821 -959 -2813
rect -953 -2821 -951 -2813
rect -943 -2821 -941 -2813
rect -927 -2821 -925 -2813
rect -917 -2821 -915 -2813
rect -909 -2821 -907 -2813
rect -899 -2821 -897 -2813
rect -883 -2821 -881 -2813
rect -875 -2821 -873 -2813
rect -859 -2821 -857 -2813
rect -843 -2821 -841 -2813
rect -835 -2821 -833 -2813
rect -825 -2821 -823 -2813
rect -749 -2821 -747 -2813
rect -739 -2821 -737 -2813
rect -723 -2821 -721 -2813
rect -713 -2821 -711 -2813
rect -697 -2821 -695 -2813
rect -687 -2821 -685 -2813
rect -679 -2821 -677 -2813
rect -669 -2821 -667 -2813
rect -653 -2821 -651 -2813
rect -645 -2821 -643 -2813
rect -635 -2821 -633 -2813
rect -619 -2821 -617 -2813
rect -609 -2821 -607 -2813
rect -601 -2821 -599 -2813
rect -591 -2821 -589 -2813
rect -575 -2821 -573 -2813
rect -567 -2821 -565 -2813
rect -551 -2821 -549 -2813
rect -535 -2821 -533 -2813
rect -527 -2821 -525 -2813
rect -517 -2821 -515 -2813
rect -441 -2821 -439 -2813
rect -431 -2821 -429 -2813
rect -415 -2821 -413 -2813
rect -405 -2821 -403 -2813
rect -389 -2821 -387 -2813
rect -379 -2821 -377 -2813
rect -371 -2821 -369 -2813
rect -361 -2821 -359 -2813
rect -345 -2821 -343 -2813
rect -337 -2821 -335 -2813
rect -327 -2821 -325 -2813
rect -311 -2821 -309 -2813
rect -301 -2821 -299 -2813
rect -293 -2821 -291 -2813
rect -283 -2821 -281 -2813
rect -267 -2821 -265 -2813
rect -259 -2821 -257 -2813
rect -243 -2821 -241 -2813
rect -227 -2821 -225 -2813
rect -219 -2821 -217 -2813
rect -209 -2821 -207 -2813
rect -133 -2821 -131 -2813
rect -123 -2821 -121 -2813
rect -107 -2821 -105 -2813
rect -97 -2821 -95 -2813
rect -81 -2821 -79 -2813
rect -71 -2821 -69 -2813
rect -63 -2821 -61 -2813
rect -53 -2821 -51 -2813
rect -37 -2821 -35 -2813
rect -29 -2821 -27 -2813
rect -19 -2821 -17 -2813
rect -3 -2821 -1 -2813
rect 7 -2821 9 -2813
rect 15 -2821 17 -2813
rect 25 -2821 27 -2813
rect 41 -2821 43 -2813
rect 49 -2821 51 -2813
rect 65 -2821 67 -2813
rect 81 -2821 83 -2813
rect 89 -2821 91 -2813
rect 99 -2821 101 -2813
rect 175 -2821 177 -2813
rect 185 -2821 187 -2813
rect 201 -2821 203 -2813
rect 211 -2821 213 -2813
rect 227 -2821 229 -2813
rect 237 -2821 239 -2813
rect 245 -2821 247 -2813
rect 255 -2821 257 -2813
rect 271 -2821 273 -2813
rect 279 -2821 281 -2813
rect 289 -2821 291 -2813
rect 305 -2821 307 -2813
rect 315 -2821 317 -2813
rect 323 -2821 325 -2813
rect 333 -2821 335 -2813
rect 349 -2821 351 -2813
rect 357 -2821 359 -2813
rect 373 -2821 375 -2813
rect 389 -2821 391 -2813
rect 397 -2821 399 -2813
rect 407 -2821 409 -2813
rect 483 -2821 485 -2813
rect 493 -2821 495 -2813
rect 509 -2821 511 -2813
rect 519 -2821 521 -2813
rect 535 -2821 537 -2813
rect 545 -2821 547 -2813
rect 553 -2821 555 -2813
rect 563 -2821 565 -2813
rect 579 -2821 581 -2813
rect 587 -2821 589 -2813
rect 597 -2821 599 -2813
rect 613 -2821 615 -2813
rect 623 -2821 625 -2813
rect 631 -2821 633 -2813
rect 641 -2821 643 -2813
rect 657 -2821 659 -2813
rect 665 -2821 667 -2813
rect 681 -2821 683 -2813
rect 697 -2821 699 -2813
rect 705 -2821 707 -2813
rect 715 -2821 717 -2813
rect 791 -2821 793 -2813
rect 801 -2821 803 -2813
rect 817 -2821 819 -2813
rect 827 -2821 829 -2813
rect 843 -2821 845 -2813
rect 853 -2821 855 -2813
rect 861 -2821 863 -2813
rect 871 -2821 873 -2813
rect 887 -2821 889 -2813
rect 895 -2821 897 -2813
rect 905 -2821 907 -2813
rect 921 -2821 923 -2813
rect 931 -2821 933 -2813
rect 939 -2821 941 -2813
rect 949 -2821 951 -2813
rect 965 -2821 967 -2813
rect 973 -2821 975 -2813
rect 989 -2821 991 -2813
rect 1005 -2821 1007 -2813
rect 1013 -2821 1015 -2813
rect 1023 -2821 1025 -2813
rect -1304 -2953 -1302 -2945
rect -1296 -2953 -1294 -2945
rect -1286 -2953 -1284 -2945
rect -1057 -2953 -1055 -2945
rect -1049 -2953 -1047 -2945
rect -1039 -2953 -1037 -2945
rect -749 -2953 -747 -2945
rect -741 -2953 -739 -2945
rect -731 -2953 -729 -2945
rect -441 -2953 -439 -2945
rect -433 -2953 -431 -2945
rect -423 -2953 -421 -2945
rect -133 -2953 -131 -2945
rect -125 -2953 -123 -2945
rect -115 -2953 -113 -2945
rect 175 -2953 177 -2945
rect 183 -2953 185 -2945
rect 193 -2953 195 -2945
rect 483 -2953 485 -2945
rect 491 -2953 493 -2945
rect 501 -2953 503 -2945
rect 791 -2953 793 -2945
rect 799 -2953 801 -2945
rect 809 -2953 811 -2945
rect -1229 -3112 -1227 -3104
rect -1219 -3112 -1217 -3104
rect -1203 -3112 -1201 -3104
rect -1193 -3112 -1191 -3104
rect -1185 -3112 -1183 -3104
rect -1175 -3112 -1173 -3104
rect -1159 -3112 -1157 -3104
rect -1151 -3112 -1149 -3104
rect -1141 -3112 -1139 -3104
rect -1057 -3112 -1055 -3104
rect -1047 -3112 -1045 -3104
rect -1031 -3112 -1029 -3104
rect -1021 -3112 -1019 -3104
rect -1005 -3112 -1003 -3104
rect -995 -3112 -993 -3104
rect -987 -3112 -985 -3104
rect -977 -3112 -975 -3104
rect -961 -3112 -959 -3104
rect -953 -3112 -951 -3104
rect -943 -3112 -941 -3104
rect -927 -3112 -925 -3104
rect -917 -3112 -915 -3104
rect -909 -3112 -907 -3104
rect -899 -3112 -897 -3104
rect -883 -3112 -881 -3104
rect -875 -3112 -873 -3104
rect -859 -3112 -857 -3104
rect -843 -3112 -841 -3104
rect -835 -3112 -833 -3104
rect -825 -3112 -823 -3104
rect -749 -3112 -747 -3104
rect -739 -3112 -737 -3104
rect -723 -3112 -721 -3104
rect -713 -3112 -711 -3104
rect -697 -3112 -695 -3104
rect -687 -3112 -685 -3104
rect -679 -3112 -677 -3104
rect -669 -3112 -667 -3104
rect -653 -3112 -651 -3104
rect -645 -3112 -643 -3104
rect -635 -3112 -633 -3104
rect -619 -3112 -617 -3104
rect -609 -3112 -607 -3104
rect -601 -3112 -599 -3104
rect -591 -3112 -589 -3104
rect -575 -3112 -573 -3104
rect -567 -3112 -565 -3104
rect -551 -3112 -549 -3104
rect -535 -3112 -533 -3104
rect -527 -3112 -525 -3104
rect -517 -3112 -515 -3104
rect -441 -3112 -439 -3104
rect -431 -3112 -429 -3104
rect -415 -3112 -413 -3104
rect -405 -3112 -403 -3104
rect -389 -3112 -387 -3104
rect -379 -3112 -377 -3104
rect -371 -3112 -369 -3104
rect -361 -3112 -359 -3104
rect -345 -3112 -343 -3104
rect -337 -3112 -335 -3104
rect -327 -3112 -325 -3104
rect -311 -3112 -309 -3104
rect -301 -3112 -299 -3104
rect -293 -3112 -291 -3104
rect -283 -3112 -281 -3104
rect -267 -3112 -265 -3104
rect -259 -3112 -257 -3104
rect -243 -3112 -241 -3104
rect -227 -3112 -225 -3104
rect -219 -3112 -217 -3104
rect -209 -3112 -207 -3104
rect -133 -3112 -131 -3104
rect -123 -3112 -121 -3104
rect -107 -3112 -105 -3104
rect -97 -3112 -95 -3104
rect -81 -3112 -79 -3104
rect -71 -3112 -69 -3104
rect -63 -3112 -61 -3104
rect -53 -3112 -51 -3104
rect -37 -3112 -35 -3104
rect -29 -3112 -27 -3104
rect -19 -3112 -17 -3104
rect -3 -3112 -1 -3104
rect 7 -3112 9 -3104
rect 15 -3112 17 -3104
rect 25 -3112 27 -3104
rect 41 -3112 43 -3104
rect 49 -3112 51 -3104
rect 65 -3112 67 -3104
rect 81 -3112 83 -3104
rect 89 -3112 91 -3104
rect 99 -3112 101 -3104
rect 175 -3112 177 -3104
rect 185 -3112 187 -3104
rect 201 -3112 203 -3104
rect 211 -3112 213 -3104
rect 227 -3112 229 -3104
rect 237 -3112 239 -3104
rect 245 -3112 247 -3104
rect 255 -3112 257 -3104
rect 271 -3112 273 -3104
rect 279 -3112 281 -3104
rect 289 -3112 291 -3104
rect 305 -3112 307 -3104
rect 315 -3112 317 -3104
rect 323 -3112 325 -3104
rect 333 -3112 335 -3104
rect 349 -3112 351 -3104
rect 357 -3112 359 -3104
rect 373 -3112 375 -3104
rect 389 -3112 391 -3104
rect 397 -3112 399 -3104
rect 407 -3112 409 -3104
rect 483 -3112 485 -3104
rect 493 -3112 495 -3104
rect 509 -3112 511 -3104
rect 519 -3112 521 -3104
rect 535 -3112 537 -3104
rect 545 -3112 547 -3104
rect 553 -3112 555 -3104
rect 563 -3112 565 -3104
rect 579 -3112 581 -3104
rect 587 -3112 589 -3104
rect 597 -3112 599 -3104
rect 613 -3112 615 -3104
rect 623 -3112 625 -3104
rect 631 -3112 633 -3104
rect 641 -3112 643 -3104
rect 657 -3112 659 -3104
rect 665 -3112 667 -3104
rect 681 -3112 683 -3104
rect 697 -3112 699 -3104
rect 705 -3112 707 -3104
rect 715 -3112 717 -3104
rect 791 -3112 793 -3104
rect 801 -3112 803 -3104
rect 817 -3112 819 -3104
rect 827 -3112 829 -3104
rect 843 -3112 845 -3104
rect 853 -3112 855 -3104
rect 861 -3112 863 -3104
rect 871 -3112 873 -3104
rect 887 -3112 889 -3104
rect 895 -3112 897 -3104
rect 905 -3112 907 -3104
rect 921 -3112 923 -3104
rect 931 -3112 933 -3104
rect 939 -3112 941 -3104
rect 949 -3112 951 -3104
rect 965 -3112 967 -3104
rect 973 -3112 975 -3104
rect 989 -3112 991 -3104
rect 1005 -3112 1007 -3104
rect 1013 -3112 1015 -3104
rect 1023 -3112 1025 -3104
<< polycontact >>
rect -1306 -1016 -1302 -1012
rect -1295 -1024 -1291 -1020
rect -1288 -1046 -1284 -1042
rect -1062 -1016 -1058 -1012
rect -1051 -1024 -1047 -1020
rect -1044 -1048 -1040 -1044
rect -753 -1016 -749 -1012
rect -742 -1024 -738 -1020
rect -735 -1048 -731 -1044
rect -445 -1016 -441 -1012
rect -434 -1024 -430 -1020
rect -427 -1048 -423 -1044
rect -138 -1016 -134 -1012
rect -127 -1024 -123 -1020
rect -120 -1061 -116 -1057
rect 171 -1016 175 -1012
rect 182 -1024 186 -1020
rect 189 -1061 193 -1057
rect 479 -1016 483 -1012
rect 490 -1024 494 -1020
rect 497 -1061 501 -1057
rect 787 -1016 791 -1012
rect 798 -1024 802 -1020
rect 805 -1061 809 -1057
rect -1308 -1166 -1304 -1162
rect -1297 -1174 -1293 -1170
rect -1290 -1196 -1286 -1192
rect -1061 -1166 -1057 -1162
rect -1050 -1174 -1046 -1170
rect -1043 -1196 -1039 -1192
rect -753 -1166 -749 -1162
rect -742 -1174 -738 -1170
rect -735 -1196 -731 -1192
rect -445 -1166 -441 -1162
rect -434 -1174 -430 -1170
rect -427 -1196 -423 -1192
rect -137 -1166 -133 -1162
rect -126 -1174 -122 -1170
rect -119 -1196 -115 -1192
rect 171 -1166 175 -1162
rect 182 -1174 186 -1170
rect 189 -1196 193 -1192
rect 479 -1166 483 -1162
rect 490 -1174 494 -1170
rect 497 -1196 501 -1192
rect 787 -1166 791 -1162
rect 798 -1174 802 -1170
rect 805 -1196 809 -1192
rect -1219 -1354 -1215 -1350
rect -1223 -1361 -1219 -1357
rect -1203 -1341 -1199 -1337
rect -1193 -1361 -1189 -1357
rect -1179 -1354 -1175 -1350
rect -1169 -1347 -1165 -1343
rect -1159 -1354 -1155 -1350
rect -1145 -1361 -1141 -1357
rect -1141 -1375 -1137 -1371
rect -1051 -1317 -1047 -1313
rect -1055 -1338 -1051 -1334
rect -1051 -1353 -1047 -1349
rect -1055 -1367 -1051 -1363
rect -1025 -1338 -1021 -1334
rect -1029 -1346 -1025 -1342
rect -1029 -1360 -1025 -1356
rect -1009 -1324 -1005 -1320
rect -999 -1367 -995 -1363
rect -985 -1317 -981 -1313
rect -975 -1331 -971 -1327
rect -965 -1367 -961 -1363
rect -951 -1317 -947 -1313
rect -947 -1375 -943 -1371
rect -931 -1346 -927 -1342
rect -921 -1360 -917 -1356
rect -907 -1317 -903 -1313
rect -907 -1338 -903 -1334
rect -903 -1353 -899 -1349
rect -887 -1360 -883 -1356
rect -873 -1317 -869 -1313
rect -863 -1368 -859 -1364
rect -847 -1375 -843 -1371
rect -833 -1331 -829 -1327
rect -829 -1368 -825 -1364
rect -743 -1317 -739 -1313
rect -747 -1338 -743 -1334
rect -743 -1353 -739 -1349
rect -747 -1367 -743 -1363
rect -717 -1338 -713 -1334
rect -721 -1346 -717 -1342
rect -721 -1360 -717 -1356
rect -701 -1324 -697 -1320
rect -691 -1367 -687 -1363
rect -677 -1317 -673 -1313
rect -667 -1331 -663 -1327
rect -657 -1367 -653 -1363
rect -643 -1317 -639 -1313
rect -639 -1375 -635 -1371
rect -623 -1346 -619 -1342
rect -613 -1360 -609 -1356
rect -599 -1317 -595 -1313
rect -599 -1338 -595 -1334
rect -595 -1353 -591 -1349
rect -579 -1360 -575 -1356
rect -565 -1317 -561 -1313
rect -555 -1368 -551 -1364
rect -539 -1375 -535 -1371
rect -525 -1331 -521 -1327
rect -521 -1368 -517 -1364
rect -435 -1317 -431 -1313
rect -439 -1338 -435 -1334
rect -435 -1353 -431 -1349
rect -439 -1367 -435 -1363
rect -409 -1338 -405 -1334
rect -413 -1346 -409 -1342
rect -413 -1360 -409 -1356
rect -393 -1324 -389 -1320
rect -383 -1367 -379 -1363
rect -369 -1317 -365 -1313
rect -359 -1331 -355 -1327
rect -349 -1367 -345 -1363
rect -335 -1317 -331 -1313
rect -331 -1375 -327 -1371
rect -315 -1346 -311 -1342
rect -305 -1360 -301 -1356
rect -291 -1317 -287 -1313
rect -291 -1338 -287 -1334
rect -287 -1353 -283 -1349
rect -271 -1360 -267 -1356
rect -257 -1317 -253 -1313
rect -247 -1368 -243 -1364
rect -231 -1375 -227 -1371
rect -217 -1331 -213 -1327
rect -213 -1368 -209 -1364
rect -127 -1317 -123 -1313
rect -131 -1338 -127 -1334
rect -127 -1353 -123 -1349
rect -131 -1367 -127 -1363
rect -101 -1338 -97 -1334
rect -105 -1346 -101 -1342
rect -105 -1360 -101 -1356
rect -85 -1324 -81 -1320
rect -75 -1367 -71 -1363
rect -61 -1317 -57 -1313
rect -51 -1331 -47 -1327
rect -41 -1367 -37 -1363
rect -27 -1317 -23 -1313
rect -23 -1375 -19 -1371
rect -7 -1346 -3 -1342
rect 3 -1360 7 -1356
rect 17 -1317 21 -1313
rect 17 -1338 21 -1334
rect 21 -1353 25 -1349
rect 37 -1360 41 -1356
rect 51 -1317 55 -1313
rect 61 -1368 65 -1364
rect 77 -1375 81 -1371
rect 91 -1331 95 -1327
rect 95 -1368 99 -1364
rect 181 -1317 185 -1313
rect 177 -1338 181 -1334
rect 181 -1353 185 -1349
rect 177 -1367 181 -1363
rect 207 -1338 211 -1334
rect 203 -1346 207 -1342
rect 203 -1360 207 -1356
rect 223 -1324 227 -1320
rect 233 -1367 237 -1363
rect 247 -1317 251 -1313
rect 257 -1331 261 -1327
rect 267 -1367 271 -1363
rect 281 -1317 285 -1313
rect 285 -1375 289 -1371
rect 301 -1346 305 -1342
rect 311 -1360 315 -1356
rect 325 -1317 329 -1313
rect 325 -1338 329 -1334
rect 329 -1353 333 -1349
rect 345 -1360 349 -1356
rect 359 -1317 363 -1313
rect 369 -1368 373 -1364
rect 385 -1375 389 -1371
rect 399 -1331 403 -1327
rect 403 -1368 407 -1364
rect 489 -1317 493 -1313
rect 485 -1338 489 -1334
rect 489 -1353 493 -1349
rect 485 -1367 489 -1363
rect 515 -1338 519 -1334
rect 511 -1346 515 -1342
rect 511 -1360 515 -1356
rect 531 -1324 535 -1320
rect 541 -1367 545 -1363
rect 555 -1317 559 -1313
rect 565 -1331 569 -1327
rect 575 -1367 579 -1363
rect 589 -1317 593 -1313
rect 593 -1375 597 -1371
rect 609 -1346 613 -1342
rect 619 -1360 623 -1356
rect 633 -1317 637 -1313
rect 633 -1338 637 -1334
rect 637 -1353 641 -1349
rect 653 -1360 657 -1356
rect 667 -1317 671 -1313
rect 677 -1368 681 -1364
rect 693 -1375 697 -1371
rect 707 -1331 711 -1327
rect 711 -1368 715 -1364
rect 795 -1354 799 -1350
rect 791 -1361 795 -1357
rect 811 -1341 815 -1337
rect 821 -1361 825 -1357
rect 835 -1354 839 -1350
rect 845 -1347 849 -1343
rect 855 -1354 859 -1350
rect 869 -1361 873 -1357
rect 873 -1375 877 -1371
rect -1308 -1487 -1304 -1483
rect -1297 -1495 -1293 -1491
rect -1290 -1517 -1286 -1513
rect -1061 -1487 -1057 -1483
rect -1050 -1495 -1046 -1491
rect -1043 -1517 -1039 -1513
rect -753 -1487 -749 -1483
rect -742 -1495 -738 -1491
rect -735 -1517 -731 -1513
rect -445 -1487 -441 -1483
rect -434 -1495 -430 -1491
rect -427 -1517 -423 -1513
rect -137 -1487 -133 -1483
rect -126 -1495 -122 -1491
rect -119 -1517 -115 -1513
rect 171 -1487 175 -1483
rect 182 -1495 186 -1491
rect 189 -1517 193 -1513
rect 479 -1487 483 -1483
rect 490 -1495 494 -1491
rect 497 -1517 501 -1513
rect 787 -1487 791 -1483
rect 798 -1495 802 -1491
rect 805 -1517 809 -1513
rect -1223 -1670 -1219 -1666
rect -1227 -1677 -1223 -1673
rect -1207 -1657 -1203 -1653
rect -1197 -1677 -1193 -1673
rect -1183 -1670 -1179 -1666
rect -1173 -1663 -1169 -1659
rect -1163 -1670 -1159 -1666
rect -1149 -1677 -1145 -1673
rect -1145 -1691 -1141 -1687
rect -1051 -1633 -1047 -1629
rect -1055 -1654 -1051 -1650
rect -1051 -1669 -1047 -1665
rect -1055 -1683 -1051 -1679
rect -1025 -1654 -1021 -1650
rect -1029 -1662 -1025 -1658
rect -1029 -1676 -1025 -1672
rect -1009 -1640 -1005 -1636
rect -999 -1683 -995 -1679
rect -985 -1633 -981 -1629
rect -975 -1647 -971 -1643
rect -965 -1683 -961 -1679
rect -951 -1633 -947 -1629
rect -947 -1691 -943 -1687
rect -931 -1662 -927 -1658
rect -921 -1676 -917 -1672
rect -907 -1633 -903 -1629
rect -907 -1654 -903 -1650
rect -903 -1669 -899 -1665
rect -887 -1676 -883 -1672
rect -873 -1633 -869 -1629
rect -863 -1684 -859 -1680
rect -847 -1691 -843 -1687
rect -833 -1647 -829 -1643
rect -829 -1684 -825 -1680
rect -743 -1633 -739 -1629
rect -747 -1654 -743 -1650
rect -743 -1669 -739 -1665
rect -747 -1683 -743 -1679
rect -717 -1654 -713 -1650
rect -721 -1662 -717 -1658
rect -721 -1676 -717 -1672
rect -701 -1640 -697 -1636
rect -691 -1683 -687 -1679
rect -677 -1633 -673 -1629
rect -667 -1647 -663 -1643
rect -657 -1683 -653 -1679
rect -643 -1633 -639 -1629
rect -639 -1691 -635 -1687
rect -623 -1662 -619 -1658
rect -613 -1676 -609 -1672
rect -599 -1633 -595 -1629
rect -599 -1654 -595 -1650
rect -595 -1669 -591 -1665
rect -579 -1676 -575 -1672
rect -565 -1633 -561 -1629
rect -555 -1684 -551 -1680
rect -539 -1691 -535 -1687
rect -525 -1647 -521 -1643
rect -521 -1684 -517 -1680
rect -435 -1633 -431 -1629
rect -439 -1654 -435 -1650
rect -435 -1669 -431 -1665
rect -439 -1683 -435 -1679
rect -409 -1654 -405 -1650
rect -413 -1662 -409 -1658
rect -413 -1676 -409 -1672
rect -393 -1640 -389 -1636
rect -383 -1683 -379 -1679
rect -369 -1633 -365 -1629
rect -359 -1647 -355 -1643
rect -349 -1683 -345 -1679
rect -335 -1633 -331 -1629
rect -331 -1691 -327 -1687
rect -315 -1662 -311 -1658
rect -305 -1676 -301 -1672
rect -291 -1633 -287 -1629
rect -291 -1654 -287 -1650
rect -287 -1669 -283 -1665
rect -271 -1676 -267 -1672
rect -257 -1633 -253 -1629
rect -247 -1684 -243 -1680
rect -231 -1691 -227 -1687
rect -217 -1647 -213 -1643
rect -213 -1684 -209 -1680
rect -127 -1633 -123 -1629
rect -131 -1654 -127 -1650
rect -127 -1669 -123 -1665
rect -131 -1683 -127 -1679
rect -101 -1654 -97 -1650
rect -105 -1662 -101 -1658
rect -105 -1676 -101 -1672
rect -85 -1640 -81 -1636
rect -75 -1683 -71 -1679
rect -61 -1633 -57 -1629
rect -51 -1647 -47 -1643
rect -41 -1683 -37 -1679
rect -27 -1633 -23 -1629
rect -23 -1691 -19 -1687
rect -7 -1662 -3 -1658
rect 3 -1676 7 -1672
rect 17 -1633 21 -1629
rect 17 -1654 21 -1650
rect 21 -1669 25 -1665
rect 37 -1676 41 -1672
rect 51 -1633 55 -1629
rect 61 -1684 65 -1680
rect 77 -1691 81 -1687
rect 91 -1647 95 -1643
rect 95 -1684 99 -1680
rect 181 -1633 185 -1629
rect 177 -1654 181 -1650
rect 181 -1669 185 -1665
rect 177 -1683 181 -1679
rect 207 -1654 211 -1650
rect 203 -1662 207 -1658
rect 203 -1676 207 -1672
rect 223 -1640 227 -1636
rect 233 -1683 237 -1679
rect 247 -1633 251 -1629
rect 257 -1647 261 -1643
rect 267 -1683 271 -1679
rect 281 -1633 285 -1629
rect 285 -1691 289 -1687
rect 301 -1662 305 -1658
rect 311 -1676 315 -1672
rect 325 -1633 329 -1629
rect 325 -1654 329 -1650
rect 329 -1669 333 -1665
rect 345 -1676 349 -1672
rect 359 -1633 363 -1629
rect 369 -1684 373 -1680
rect 385 -1691 389 -1687
rect 399 -1647 403 -1643
rect 403 -1684 407 -1680
rect 489 -1633 493 -1629
rect 485 -1654 489 -1650
rect 489 -1669 493 -1665
rect 485 -1683 489 -1679
rect 515 -1654 519 -1650
rect 511 -1662 515 -1658
rect 511 -1676 515 -1672
rect 531 -1640 535 -1636
rect 541 -1683 545 -1679
rect 555 -1633 559 -1629
rect 565 -1647 569 -1643
rect 575 -1683 579 -1679
rect 589 -1633 593 -1629
rect 593 -1691 597 -1687
rect 609 -1662 613 -1658
rect 619 -1676 623 -1672
rect 633 -1633 637 -1629
rect 633 -1654 637 -1650
rect 637 -1669 641 -1665
rect 653 -1676 657 -1672
rect 667 -1633 671 -1629
rect 677 -1684 681 -1680
rect 693 -1691 697 -1687
rect 707 -1647 711 -1643
rect 711 -1684 715 -1680
rect 797 -1633 801 -1629
rect 793 -1654 797 -1650
rect 797 -1669 801 -1665
rect 793 -1683 797 -1679
rect 823 -1654 827 -1650
rect 819 -1662 823 -1658
rect 819 -1676 823 -1672
rect 839 -1640 843 -1636
rect 849 -1683 853 -1679
rect 863 -1633 867 -1629
rect 873 -1647 877 -1643
rect 883 -1683 887 -1679
rect 897 -1633 901 -1629
rect 901 -1691 905 -1687
rect 917 -1662 921 -1658
rect 927 -1676 931 -1672
rect 941 -1633 945 -1629
rect 941 -1654 945 -1650
rect 945 -1669 949 -1665
rect 961 -1676 965 -1672
rect 975 -1633 979 -1629
rect 985 -1684 989 -1680
rect 1001 -1691 1005 -1687
rect 1015 -1647 1019 -1643
rect 1019 -1684 1023 -1680
rect -1308 -1778 -1304 -1774
rect -1297 -1786 -1293 -1782
rect -1290 -1808 -1286 -1804
rect -1061 -1778 -1057 -1774
rect -1050 -1786 -1046 -1782
rect -1043 -1808 -1039 -1804
rect -753 -1778 -749 -1774
rect -742 -1786 -738 -1782
rect -735 -1808 -731 -1804
rect -445 -1778 -441 -1774
rect -434 -1786 -430 -1782
rect -427 -1808 -423 -1804
rect -137 -1778 -133 -1774
rect -126 -1786 -122 -1782
rect -119 -1808 -115 -1804
rect 171 -1778 175 -1774
rect 182 -1786 186 -1782
rect 189 -1808 193 -1804
rect 479 -1778 483 -1774
rect 490 -1786 494 -1782
rect 497 -1808 501 -1804
rect 787 -1778 791 -1774
rect 798 -1786 802 -1782
rect 805 -1808 809 -1804
rect -1223 -1961 -1219 -1957
rect -1227 -1968 -1223 -1964
rect -1207 -1948 -1203 -1944
rect -1197 -1968 -1193 -1964
rect -1183 -1961 -1179 -1957
rect -1173 -1954 -1169 -1950
rect -1163 -1961 -1159 -1957
rect -1149 -1968 -1145 -1964
rect -1145 -1982 -1141 -1978
rect -1051 -1924 -1047 -1920
rect -1055 -1945 -1051 -1941
rect -1051 -1960 -1047 -1956
rect -1055 -1974 -1051 -1970
rect -1025 -1945 -1021 -1941
rect -1029 -1953 -1025 -1949
rect -1029 -1967 -1025 -1963
rect -1009 -1931 -1005 -1927
rect -999 -1974 -995 -1970
rect -985 -1924 -981 -1920
rect -975 -1938 -971 -1934
rect -965 -1974 -961 -1970
rect -951 -1924 -947 -1920
rect -947 -1982 -943 -1978
rect -931 -1953 -927 -1949
rect -921 -1967 -917 -1963
rect -907 -1924 -903 -1920
rect -907 -1945 -903 -1941
rect -903 -1960 -899 -1956
rect -887 -1967 -883 -1963
rect -873 -1924 -869 -1920
rect -863 -1975 -859 -1971
rect -847 -1982 -843 -1978
rect -833 -1938 -829 -1934
rect -829 -1975 -825 -1971
rect -743 -1924 -739 -1920
rect -747 -1945 -743 -1941
rect -743 -1960 -739 -1956
rect -747 -1974 -743 -1970
rect -717 -1945 -713 -1941
rect -721 -1953 -717 -1949
rect -721 -1967 -717 -1963
rect -701 -1931 -697 -1927
rect -691 -1974 -687 -1970
rect -677 -1924 -673 -1920
rect -667 -1938 -663 -1934
rect -657 -1974 -653 -1970
rect -643 -1924 -639 -1920
rect -639 -1982 -635 -1978
rect -623 -1953 -619 -1949
rect -613 -1967 -609 -1963
rect -599 -1924 -595 -1920
rect -599 -1945 -595 -1941
rect -595 -1960 -591 -1956
rect -579 -1967 -575 -1963
rect -565 -1924 -561 -1920
rect -555 -1975 -551 -1971
rect -539 -1982 -535 -1978
rect -525 -1938 -521 -1934
rect -521 -1975 -517 -1971
rect -435 -1924 -431 -1920
rect -439 -1945 -435 -1941
rect -435 -1960 -431 -1956
rect -439 -1974 -435 -1970
rect -409 -1945 -405 -1941
rect -413 -1953 -409 -1949
rect -413 -1967 -409 -1963
rect -393 -1931 -389 -1927
rect -383 -1974 -379 -1970
rect -369 -1924 -365 -1920
rect -359 -1938 -355 -1934
rect -349 -1974 -345 -1970
rect -335 -1924 -331 -1920
rect -331 -1982 -327 -1978
rect -315 -1953 -311 -1949
rect -305 -1967 -301 -1963
rect -291 -1924 -287 -1920
rect -291 -1945 -287 -1941
rect -287 -1960 -283 -1956
rect -271 -1967 -267 -1963
rect -257 -1924 -253 -1920
rect -247 -1975 -243 -1971
rect -231 -1982 -227 -1978
rect -217 -1938 -213 -1934
rect -213 -1975 -209 -1971
rect -127 -1924 -123 -1920
rect -131 -1945 -127 -1941
rect -127 -1960 -123 -1956
rect -131 -1974 -127 -1970
rect -101 -1945 -97 -1941
rect -105 -1953 -101 -1949
rect -105 -1967 -101 -1963
rect -85 -1931 -81 -1927
rect -75 -1974 -71 -1970
rect -61 -1924 -57 -1920
rect -51 -1938 -47 -1934
rect -41 -1974 -37 -1970
rect -27 -1924 -23 -1920
rect -23 -1982 -19 -1978
rect -7 -1953 -3 -1949
rect 3 -1967 7 -1963
rect 17 -1924 21 -1920
rect 17 -1945 21 -1941
rect 21 -1960 25 -1956
rect 37 -1967 41 -1963
rect 51 -1924 55 -1920
rect 61 -1975 65 -1971
rect 77 -1982 81 -1978
rect 91 -1938 95 -1934
rect 95 -1975 99 -1971
rect 181 -1924 185 -1920
rect 177 -1945 181 -1941
rect 181 -1960 185 -1956
rect 177 -1974 181 -1970
rect 207 -1945 211 -1941
rect 203 -1953 207 -1949
rect 203 -1967 207 -1963
rect 223 -1931 227 -1927
rect 233 -1974 237 -1970
rect 247 -1924 251 -1920
rect 257 -1938 261 -1934
rect 267 -1974 271 -1970
rect 281 -1924 285 -1920
rect 285 -1982 289 -1978
rect 301 -1953 305 -1949
rect 311 -1967 315 -1963
rect 325 -1924 329 -1920
rect 325 -1945 329 -1941
rect 329 -1960 333 -1956
rect 345 -1967 349 -1963
rect 359 -1924 363 -1920
rect 369 -1975 373 -1971
rect 385 -1982 389 -1978
rect 399 -1938 403 -1934
rect 403 -1975 407 -1971
rect 489 -1924 493 -1920
rect 485 -1945 489 -1941
rect 489 -1960 493 -1956
rect 485 -1974 489 -1970
rect 515 -1945 519 -1941
rect 511 -1953 515 -1949
rect 511 -1967 515 -1963
rect 531 -1931 535 -1927
rect 541 -1974 545 -1970
rect 555 -1924 559 -1920
rect 565 -1938 569 -1934
rect 575 -1974 579 -1970
rect 589 -1924 593 -1920
rect 593 -1982 597 -1978
rect 609 -1953 613 -1949
rect 619 -1967 623 -1963
rect 633 -1924 637 -1920
rect 633 -1945 637 -1941
rect 637 -1960 641 -1956
rect 653 -1967 657 -1963
rect 667 -1924 671 -1920
rect 677 -1975 681 -1971
rect 693 -1982 697 -1978
rect 707 -1938 711 -1934
rect 711 -1975 715 -1971
rect 797 -1924 801 -1920
rect 793 -1945 797 -1941
rect 797 -1960 801 -1956
rect 793 -1974 797 -1970
rect 823 -1945 827 -1941
rect 819 -1953 823 -1949
rect 819 -1967 823 -1963
rect 839 -1931 843 -1927
rect 849 -1974 853 -1970
rect 863 -1924 867 -1920
rect 873 -1938 877 -1934
rect 883 -1974 887 -1970
rect 897 -1924 901 -1920
rect 901 -1982 905 -1978
rect 917 -1953 921 -1949
rect 927 -1967 931 -1963
rect 941 -1924 945 -1920
rect 941 -1945 945 -1941
rect 945 -1960 949 -1956
rect 961 -1967 965 -1963
rect 975 -1924 979 -1920
rect 985 -1975 989 -1971
rect 1001 -1982 1005 -1978
rect 1015 -1938 1019 -1934
rect 1019 -1975 1023 -1971
rect -1308 -2100 -1304 -2096
rect -1297 -2108 -1293 -2104
rect -1290 -2130 -1286 -2126
rect -1061 -2100 -1057 -2096
rect -1050 -2108 -1046 -2104
rect -1043 -2130 -1039 -2126
rect -753 -2100 -749 -2096
rect -742 -2108 -738 -2104
rect -735 -2130 -731 -2126
rect -445 -2100 -441 -2096
rect -434 -2108 -430 -2104
rect -427 -2130 -423 -2126
rect -137 -2100 -133 -2096
rect -126 -2108 -122 -2104
rect -119 -2130 -115 -2126
rect 171 -2100 175 -2096
rect 182 -2108 186 -2104
rect 189 -2130 193 -2126
rect 479 -2100 483 -2096
rect 490 -2108 494 -2104
rect 497 -2130 501 -2126
rect 787 -2100 791 -2096
rect 798 -2108 802 -2104
rect 805 -2130 809 -2126
rect -1223 -2283 -1219 -2279
rect -1227 -2290 -1223 -2286
rect -1207 -2270 -1203 -2266
rect -1197 -2290 -1193 -2286
rect -1183 -2283 -1179 -2279
rect -1173 -2276 -1169 -2272
rect -1163 -2283 -1159 -2279
rect -1149 -2290 -1145 -2286
rect -1145 -2304 -1141 -2300
rect -1051 -2246 -1047 -2242
rect -1055 -2267 -1051 -2263
rect -1051 -2282 -1047 -2278
rect -1055 -2296 -1051 -2292
rect -1025 -2267 -1021 -2263
rect -1029 -2275 -1025 -2271
rect -1029 -2289 -1025 -2285
rect -1009 -2253 -1005 -2249
rect -999 -2296 -995 -2292
rect -985 -2246 -981 -2242
rect -975 -2260 -971 -2256
rect -965 -2296 -961 -2292
rect -951 -2246 -947 -2242
rect -947 -2304 -943 -2300
rect -931 -2275 -927 -2271
rect -921 -2289 -917 -2285
rect -907 -2246 -903 -2242
rect -907 -2267 -903 -2263
rect -903 -2282 -899 -2278
rect -887 -2289 -883 -2285
rect -873 -2246 -869 -2242
rect -863 -2297 -859 -2293
rect -847 -2304 -843 -2300
rect -833 -2260 -829 -2256
rect -829 -2297 -825 -2293
rect -743 -2246 -739 -2242
rect -747 -2267 -743 -2263
rect -743 -2282 -739 -2278
rect -747 -2296 -743 -2292
rect -717 -2267 -713 -2263
rect -721 -2275 -717 -2271
rect -721 -2289 -717 -2285
rect -701 -2253 -697 -2249
rect -691 -2296 -687 -2292
rect -677 -2246 -673 -2242
rect -667 -2260 -663 -2256
rect -657 -2296 -653 -2292
rect -643 -2246 -639 -2242
rect -639 -2304 -635 -2300
rect -623 -2275 -619 -2271
rect -613 -2289 -609 -2285
rect -599 -2246 -595 -2242
rect -599 -2267 -595 -2263
rect -595 -2282 -591 -2278
rect -579 -2289 -575 -2285
rect -565 -2246 -561 -2242
rect -555 -2297 -551 -2293
rect -539 -2304 -535 -2300
rect -525 -2260 -521 -2256
rect -521 -2297 -517 -2293
rect -435 -2246 -431 -2242
rect -439 -2267 -435 -2263
rect -435 -2282 -431 -2278
rect -439 -2296 -435 -2292
rect -409 -2267 -405 -2263
rect -413 -2275 -409 -2271
rect -413 -2289 -409 -2285
rect -393 -2253 -389 -2249
rect -383 -2296 -379 -2292
rect -369 -2246 -365 -2242
rect -359 -2260 -355 -2256
rect -349 -2296 -345 -2292
rect -335 -2246 -331 -2242
rect -331 -2304 -327 -2300
rect -315 -2275 -311 -2271
rect -305 -2289 -301 -2285
rect -291 -2246 -287 -2242
rect -291 -2267 -287 -2263
rect -287 -2282 -283 -2278
rect -271 -2289 -267 -2285
rect -257 -2246 -253 -2242
rect -247 -2297 -243 -2293
rect -231 -2304 -227 -2300
rect -217 -2260 -213 -2256
rect -213 -2297 -209 -2293
rect -127 -2246 -123 -2242
rect -131 -2267 -127 -2263
rect -127 -2282 -123 -2278
rect -131 -2296 -127 -2292
rect -101 -2267 -97 -2263
rect -105 -2275 -101 -2271
rect -105 -2289 -101 -2285
rect -85 -2253 -81 -2249
rect -75 -2296 -71 -2292
rect -61 -2246 -57 -2242
rect -51 -2260 -47 -2256
rect -41 -2296 -37 -2292
rect -27 -2246 -23 -2242
rect -23 -2304 -19 -2300
rect -7 -2275 -3 -2271
rect 3 -2289 7 -2285
rect 17 -2246 21 -2242
rect 17 -2267 21 -2263
rect 21 -2282 25 -2278
rect 37 -2289 41 -2285
rect 51 -2246 55 -2242
rect 61 -2297 65 -2293
rect 77 -2304 81 -2300
rect 91 -2260 95 -2256
rect 95 -2297 99 -2293
rect 181 -2246 185 -2242
rect 177 -2267 181 -2263
rect 181 -2282 185 -2278
rect 177 -2296 181 -2292
rect 207 -2267 211 -2263
rect 203 -2275 207 -2271
rect 203 -2289 207 -2285
rect 223 -2253 227 -2249
rect 233 -2296 237 -2292
rect 247 -2246 251 -2242
rect 257 -2260 261 -2256
rect 267 -2296 271 -2292
rect 281 -2246 285 -2242
rect 285 -2304 289 -2300
rect 301 -2275 305 -2271
rect 311 -2289 315 -2285
rect 325 -2246 329 -2242
rect 325 -2267 329 -2263
rect 329 -2282 333 -2278
rect 345 -2289 349 -2285
rect 359 -2246 363 -2242
rect 369 -2297 373 -2293
rect 385 -2304 389 -2300
rect 399 -2260 403 -2256
rect 403 -2297 407 -2293
rect 489 -2246 493 -2242
rect 485 -2267 489 -2263
rect 489 -2282 493 -2278
rect 485 -2296 489 -2292
rect 515 -2267 519 -2263
rect 511 -2275 515 -2271
rect 511 -2289 515 -2285
rect 531 -2253 535 -2249
rect 541 -2296 545 -2292
rect 555 -2246 559 -2242
rect 565 -2260 569 -2256
rect 575 -2296 579 -2292
rect 589 -2246 593 -2242
rect 593 -2304 597 -2300
rect 609 -2275 613 -2271
rect 619 -2289 623 -2285
rect 633 -2246 637 -2242
rect 633 -2267 637 -2263
rect 637 -2282 641 -2278
rect 653 -2289 657 -2285
rect 667 -2246 671 -2242
rect 677 -2297 681 -2293
rect 693 -2304 697 -2300
rect 707 -2260 711 -2256
rect 711 -2297 715 -2293
rect 797 -2246 801 -2242
rect 793 -2267 797 -2263
rect 797 -2282 801 -2278
rect 793 -2296 797 -2292
rect 823 -2267 827 -2263
rect 819 -2275 823 -2271
rect 819 -2289 823 -2285
rect 839 -2253 843 -2249
rect 849 -2296 853 -2292
rect 863 -2246 867 -2242
rect 873 -2260 877 -2256
rect 883 -2296 887 -2292
rect 897 -2246 901 -2242
rect 901 -2304 905 -2300
rect 917 -2275 921 -2271
rect 927 -2289 931 -2285
rect 941 -2246 945 -2242
rect 941 -2267 945 -2263
rect 945 -2282 949 -2278
rect 961 -2289 965 -2285
rect 975 -2246 979 -2242
rect 985 -2297 989 -2293
rect 1001 -2304 1005 -2300
rect 1015 -2260 1019 -2256
rect 1019 -2297 1023 -2293
rect -1308 -2391 -1304 -2387
rect -1297 -2399 -1293 -2395
rect -1290 -2421 -1286 -2417
rect -1061 -2391 -1057 -2387
rect -1050 -2399 -1046 -2395
rect -1043 -2421 -1039 -2417
rect -753 -2391 -749 -2387
rect -742 -2399 -738 -2395
rect -735 -2421 -731 -2417
rect -445 -2391 -441 -2387
rect -434 -2399 -430 -2395
rect -427 -2421 -423 -2417
rect -137 -2391 -133 -2387
rect -126 -2399 -122 -2395
rect -119 -2421 -115 -2417
rect 171 -2391 175 -2387
rect 182 -2399 186 -2395
rect 189 -2421 193 -2417
rect 479 -2391 483 -2387
rect 490 -2399 494 -2395
rect 497 -2421 501 -2417
rect 787 -2391 791 -2387
rect 798 -2399 802 -2395
rect 805 -2421 809 -2417
rect -1223 -2574 -1219 -2570
rect -1227 -2581 -1223 -2577
rect -1207 -2561 -1203 -2557
rect -1197 -2581 -1193 -2577
rect -1183 -2574 -1179 -2570
rect -1173 -2567 -1169 -2563
rect -1163 -2574 -1159 -2570
rect -1149 -2581 -1145 -2577
rect -1145 -2595 -1141 -2591
rect -1051 -2537 -1047 -2533
rect -1055 -2558 -1051 -2554
rect -1051 -2573 -1047 -2569
rect -1055 -2587 -1051 -2583
rect -1025 -2558 -1021 -2554
rect -1029 -2566 -1025 -2562
rect -1029 -2580 -1025 -2576
rect -1009 -2544 -1005 -2540
rect -999 -2587 -995 -2583
rect -985 -2537 -981 -2533
rect -975 -2551 -971 -2547
rect -965 -2587 -961 -2583
rect -951 -2537 -947 -2533
rect -947 -2595 -943 -2591
rect -931 -2566 -927 -2562
rect -921 -2580 -917 -2576
rect -907 -2537 -903 -2533
rect -907 -2558 -903 -2554
rect -903 -2573 -899 -2569
rect -887 -2580 -883 -2576
rect -873 -2537 -869 -2533
rect -863 -2588 -859 -2584
rect -847 -2595 -843 -2591
rect -833 -2551 -829 -2547
rect -829 -2588 -825 -2584
rect -743 -2537 -739 -2533
rect -747 -2558 -743 -2554
rect -743 -2573 -739 -2569
rect -747 -2587 -743 -2583
rect -717 -2558 -713 -2554
rect -721 -2566 -717 -2562
rect -721 -2580 -717 -2576
rect -701 -2544 -697 -2540
rect -691 -2587 -687 -2583
rect -677 -2537 -673 -2533
rect -667 -2551 -663 -2547
rect -657 -2587 -653 -2583
rect -643 -2537 -639 -2533
rect -639 -2595 -635 -2591
rect -623 -2566 -619 -2562
rect -613 -2580 -609 -2576
rect -599 -2537 -595 -2533
rect -599 -2558 -595 -2554
rect -595 -2573 -591 -2569
rect -579 -2580 -575 -2576
rect -565 -2537 -561 -2533
rect -555 -2588 -551 -2584
rect -539 -2595 -535 -2591
rect -525 -2551 -521 -2547
rect -521 -2588 -517 -2584
rect -435 -2537 -431 -2533
rect -439 -2558 -435 -2554
rect -435 -2573 -431 -2569
rect -439 -2587 -435 -2583
rect -409 -2558 -405 -2554
rect -413 -2566 -409 -2562
rect -413 -2580 -409 -2576
rect -393 -2544 -389 -2540
rect -383 -2587 -379 -2583
rect -369 -2537 -365 -2533
rect -359 -2551 -355 -2547
rect -349 -2587 -345 -2583
rect -335 -2537 -331 -2533
rect -331 -2595 -327 -2591
rect -315 -2566 -311 -2562
rect -305 -2580 -301 -2576
rect -291 -2537 -287 -2533
rect -291 -2558 -287 -2554
rect -287 -2573 -283 -2569
rect -271 -2580 -267 -2576
rect -257 -2537 -253 -2533
rect -247 -2588 -243 -2584
rect -231 -2595 -227 -2591
rect -217 -2551 -213 -2547
rect -213 -2588 -209 -2584
rect -127 -2537 -123 -2533
rect -131 -2558 -127 -2554
rect -127 -2573 -123 -2569
rect -131 -2587 -127 -2583
rect -101 -2558 -97 -2554
rect -105 -2566 -101 -2562
rect -105 -2580 -101 -2576
rect -85 -2544 -81 -2540
rect -75 -2587 -71 -2583
rect -61 -2537 -57 -2533
rect -51 -2551 -47 -2547
rect -41 -2587 -37 -2583
rect -27 -2537 -23 -2533
rect -23 -2595 -19 -2591
rect -7 -2566 -3 -2562
rect 3 -2580 7 -2576
rect 17 -2537 21 -2533
rect 17 -2558 21 -2554
rect 21 -2573 25 -2569
rect 37 -2580 41 -2576
rect 51 -2537 55 -2533
rect 61 -2588 65 -2584
rect 77 -2595 81 -2591
rect 91 -2551 95 -2547
rect 95 -2588 99 -2584
rect 181 -2537 185 -2533
rect 177 -2558 181 -2554
rect 181 -2573 185 -2569
rect 177 -2587 181 -2583
rect 207 -2558 211 -2554
rect 203 -2566 207 -2562
rect 203 -2580 207 -2576
rect 223 -2544 227 -2540
rect 233 -2587 237 -2583
rect 247 -2537 251 -2533
rect 257 -2551 261 -2547
rect 267 -2587 271 -2583
rect 281 -2537 285 -2533
rect 285 -2595 289 -2591
rect 301 -2566 305 -2562
rect 311 -2580 315 -2576
rect 325 -2537 329 -2533
rect 325 -2558 329 -2554
rect 329 -2573 333 -2569
rect 345 -2580 349 -2576
rect 359 -2537 363 -2533
rect 369 -2588 373 -2584
rect 385 -2595 389 -2591
rect 399 -2551 403 -2547
rect 403 -2588 407 -2584
rect 489 -2537 493 -2533
rect 485 -2558 489 -2554
rect 489 -2573 493 -2569
rect 485 -2587 489 -2583
rect 515 -2558 519 -2554
rect 511 -2566 515 -2562
rect 511 -2580 515 -2576
rect 531 -2544 535 -2540
rect 541 -2587 545 -2583
rect 555 -2537 559 -2533
rect 565 -2551 569 -2547
rect 575 -2587 579 -2583
rect 589 -2537 593 -2533
rect 593 -2595 597 -2591
rect 609 -2566 613 -2562
rect 619 -2580 623 -2576
rect 633 -2537 637 -2533
rect 633 -2558 637 -2554
rect 637 -2573 641 -2569
rect 653 -2580 657 -2576
rect 667 -2537 671 -2533
rect 677 -2588 681 -2584
rect 693 -2595 697 -2591
rect 707 -2551 711 -2547
rect 711 -2588 715 -2584
rect 797 -2537 801 -2533
rect 793 -2558 797 -2554
rect 797 -2573 801 -2569
rect 793 -2587 797 -2583
rect 823 -2558 827 -2554
rect 819 -2566 823 -2562
rect 819 -2580 823 -2576
rect 839 -2544 843 -2540
rect 849 -2587 853 -2583
rect 863 -2537 867 -2533
rect 873 -2551 877 -2547
rect 883 -2587 887 -2583
rect 897 -2537 901 -2533
rect 901 -2595 905 -2591
rect 917 -2566 921 -2562
rect 927 -2580 931 -2576
rect 941 -2537 945 -2533
rect 941 -2558 945 -2554
rect 945 -2573 949 -2569
rect 961 -2580 965 -2576
rect 975 -2537 979 -2533
rect 985 -2588 989 -2584
rect 1001 -2595 1005 -2591
rect 1015 -2551 1019 -2547
rect 1019 -2588 1023 -2584
rect -1308 -2682 -1304 -2678
rect -1297 -2690 -1293 -2686
rect -1290 -2712 -1286 -2708
rect -1061 -2682 -1057 -2678
rect -1050 -2690 -1046 -2686
rect -1043 -2712 -1039 -2708
rect -753 -2682 -749 -2678
rect -742 -2690 -738 -2686
rect -735 -2712 -731 -2708
rect -445 -2682 -441 -2678
rect -434 -2690 -430 -2686
rect -427 -2712 -423 -2708
rect -137 -2682 -133 -2678
rect -126 -2690 -122 -2686
rect -119 -2712 -115 -2708
rect 171 -2682 175 -2678
rect 182 -2690 186 -2686
rect 189 -2712 193 -2708
rect 479 -2682 483 -2678
rect 490 -2690 494 -2686
rect 497 -2712 501 -2708
rect 787 -2682 791 -2678
rect 798 -2690 802 -2686
rect 805 -2712 809 -2708
rect -1223 -2865 -1219 -2861
rect -1227 -2872 -1223 -2868
rect -1207 -2852 -1203 -2848
rect -1197 -2872 -1193 -2868
rect -1183 -2865 -1179 -2861
rect -1173 -2858 -1169 -2854
rect -1163 -2865 -1159 -2861
rect -1149 -2872 -1145 -2868
rect -1145 -2886 -1141 -2882
rect -1051 -2828 -1047 -2824
rect -1055 -2849 -1051 -2845
rect -1051 -2864 -1047 -2860
rect -1055 -2878 -1051 -2874
rect -1025 -2849 -1021 -2845
rect -1029 -2857 -1025 -2853
rect -1029 -2871 -1025 -2867
rect -1009 -2835 -1005 -2831
rect -999 -2878 -995 -2874
rect -985 -2828 -981 -2824
rect -975 -2842 -971 -2838
rect -965 -2878 -961 -2874
rect -951 -2828 -947 -2824
rect -947 -2886 -943 -2882
rect -931 -2857 -927 -2853
rect -921 -2871 -917 -2867
rect -907 -2828 -903 -2824
rect -907 -2849 -903 -2845
rect -903 -2864 -899 -2860
rect -887 -2871 -883 -2867
rect -873 -2828 -869 -2824
rect -863 -2879 -859 -2875
rect -847 -2886 -843 -2882
rect -833 -2842 -829 -2838
rect -829 -2879 -825 -2875
rect -743 -2828 -739 -2824
rect -747 -2849 -743 -2845
rect -743 -2864 -739 -2860
rect -747 -2878 -743 -2874
rect -717 -2849 -713 -2845
rect -721 -2857 -717 -2853
rect -721 -2871 -717 -2867
rect -701 -2835 -697 -2831
rect -691 -2878 -687 -2874
rect -677 -2828 -673 -2824
rect -667 -2842 -663 -2838
rect -657 -2878 -653 -2874
rect -643 -2828 -639 -2824
rect -639 -2886 -635 -2882
rect -623 -2857 -619 -2853
rect -613 -2871 -609 -2867
rect -599 -2828 -595 -2824
rect -599 -2849 -595 -2845
rect -595 -2864 -591 -2860
rect -579 -2871 -575 -2867
rect -565 -2828 -561 -2824
rect -555 -2879 -551 -2875
rect -539 -2886 -535 -2882
rect -525 -2842 -521 -2838
rect -521 -2879 -517 -2875
rect -435 -2828 -431 -2824
rect -439 -2849 -435 -2845
rect -435 -2864 -431 -2860
rect -439 -2878 -435 -2874
rect -409 -2849 -405 -2845
rect -413 -2857 -409 -2853
rect -413 -2871 -409 -2867
rect -393 -2835 -389 -2831
rect -383 -2878 -379 -2874
rect -369 -2828 -365 -2824
rect -359 -2842 -355 -2838
rect -349 -2878 -345 -2874
rect -335 -2828 -331 -2824
rect -331 -2886 -327 -2882
rect -315 -2857 -311 -2853
rect -305 -2871 -301 -2867
rect -291 -2828 -287 -2824
rect -291 -2849 -287 -2845
rect -287 -2864 -283 -2860
rect -271 -2871 -267 -2867
rect -257 -2828 -253 -2824
rect -247 -2879 -243 -2875
rect -231 -2886 -227 -2882
rect -217 -2842 -213 -2838
rect -213 -2879 -209 -2875
rect -127 -2828 -123 -2824
rect -131 -2849 -127 -2845
rect -127 -2864 -123 -2860
rect -131 -2878 -127 -2874
rect -101 -2849 -97 -2845
rect -105 -2857 -101 -2853
rect -105 -2871 -101 -2867
rect -85 -2835 -81 -2831
rect -75 -2878 -71 -2874
rect -61 -2828 -57 -2824
rect -51 -2842 -47 -2838
rect -41 -2878 -37 -2874
rect -27 -2828 -23 -2824
rect -23 -2886 -19 -2882
rect -7 -2857 -3 -2853
rect 3 -2871 7 -2867
rect 17 -2828 21 -2824
rect 17 -2849 21 -2845
rect 21 -2864 25 -2860
rect 37 -2871 41 -2867
rect 51 -2828 55 -2824
rect 61 -2879 65 -2875
rect 77 -2886 81 -2882
rect 91 -2842 95 -2838
rect 95 -2879 99 -2875
rect 181 -2828 185 -2824
rect 177 -2849 181 -2845
rect 181 -2864 185 -2860
rect 177 -2878 181 -2874
rect 207 -2849 211 -2845
rect 203 -2857 207 -2853
rect 203 -2871 207 -2867
rect 223 -2835 227 -2831
rect 233 -2878 237 -2874
rect 247 -2828 251 -2824
rect 257 -2842 261 -2838
rect 267 -2878 271 -2874
rect 281 -2828 285 -2824
rect 285 -2886 289 -2882
rect 301 -2857 305 -2853
rect 311 -2871 315 -2867
rect 325 -2828 329 -2824
rect 325 -2849 329 -2845
rect 329 -2864 333 -2860
rect 345 -2871 349 -2867
rect 359 -2828 363 -2824
rect 369 -2879 373 -2875
rect 385 -2886 389 -2882
rect 399 -2842 403 -2838
rect 403 -2879 407 -2875
rect 489 -2828 493 -2824
rect 485 -2849 489 -2845
rect 489 -2864 493 -2860
rect 485 -2878 489 -2874
rect 515 -2849 519 -2845
rect 511 -2857 515 -2853
rect 511 -2871 515 -2867
rect 531 -2835 535 -2831
rect 541 -2878 545 -2874
rect 555 -2828 559 -2824
rect 565 -2842 569 -2838
rect 575 -2878 579 -2874
rect 589 -2828 593 -2824
rect 593 -2886 597 -2882
rect 609 -2857 613 -2853
rect 619 -2871 623 -2867
rect 633 -2828 637 -2824
rect 633 -2849 637 -2845
rect 637 -2864 641 -2860
rect 653 -2871 657 -2867
rect 667 -2828 671 -2824
rect 677 -2879 681 -2875
rect 693 -2886 697 -2882
rect 707 -2842 711 -2838
rect 711 -2879 715 -2875
rect 797 -2828 801 -2824
rect 793 -2849 797 -2845
rect 797 -2864 801 -2860
rect 793 -2878 797 -2874
rect 823 -2849 827 -2845
rect 819 -2857 823 -2853
rect 819 -2871 823 -2867
rect 839 -2835 843 -2831
rect 849 -2878 853 -2874
rect 863 -2828 867 -2824
rect 873 -2842 877 -2838
rect 883 -2878 887 -2874
rect 897 -2828 901 -2824
rect 901 -2886 905 -2882
rect 917 -2857 921 -2853
rect 927 -2871 931 -2867
rect 941 -2828 945 -2824
rect 941 -2849 945 -2845
rect 945 -2864 949 -2860
rect 961 -2871 965 -2867
rect 975 -2828 979 -2824
rect 985 -2879 989 -2875
rect 1001 -2886 1005 -2882
rect 1015 -2842 1019 -2838
rect 1019 -2879 1023 -2875
rect -1308 -2973 -1304 -2969
rect -1297 -2981 -1293 -2977
rect -1290 -3003 -1286 -2999
rect -1061 -2973 -1057 -2969
rect -1050 -2981 -1046 -2977
rect -1043 -3003 -1039 -2999
rect -753 -2973 -749 -2969
rect -742 -2981 -738 -2977
rect -735 -3003 -731 -2999
rect -445 -2973 -441 -2969
rect -434 -2981 -430 -2977
rect -427 -3003 -423 -2999
rect -137 -2973 -133 -2969
rect -126 -2981 -122 -2977
rect -119 -3003 -115 -2999
rect 171 -2973 175 -2969
rect 182 -2981 186 -2977
rect 189 -3003 193 -2999
rect 479 -2973 483 -2969
rect 490 -2981 494 -2977
rect 497 -3003 501 -2999
rect 787 -2973 791 -2969
rect 798 -2981 802 -2977
rect 805 -3003 809 -2999
rect -1223 -3156 -1219 -3152
rect -1227 -3163 -1223 -3159
rect -1207 -3143 -1203 -3139
rect -1197 -3163 -1193 -3159
rect -1183 -3156 -1179 -3152
rect -1173 -3149 -1169 -3145
rect -1163 -3156 -1159 -3152
rect -1149 -3163 -1145 -3159
rect -1145 -3177 -1141 -3173
rect -1051 -3119 -1047 -3115
rect -1055 -3140 -1051 -3136
rect -1051 -3155 -1047 -3151
rect -1055 -3169 -1051 -3165
rect -1025 -3140 -1021 -3136
rect -1029 -3148 -1025 -3144
rect -1029 -3162 -1025 -3158
rect -1009 -3126 -1005 -3122
rect -999 -3169 -995 -3165
rect -985 -3119 -981 -3115
rect -975 -3133 -971 -3129
rect -965 -3169 -961 -3165
rect -951 -3119 -947 -3115
rect -947 -3177 -943 -3173
rect -931 -3148 -927 -3144
rect -921 -3162 -917 -3158
rect -907 -3119 -903 -3115
rect -907 -3140 -903 -3136
rect -903 -3155 -899 -3151
rect -887 -3162 -883 -3158
rect -873 -3119 -869 -3115
rect -863 -3170 -859 -3166
rect -847 -3177 -843 -3173
rect -833 -3133 -829 -3129
rect -829 -3170 -825 -3166
rect -743 -3119 -739 -3115
rect -747 -3140 -743 -3136
rect -743 -3155 -739 -3151
rect -747 -3169 -743 -3165
rect -717 -3140 -713 -3136
rect -721 -3148 -717 -3144
rect -721 -3162 -717 -3158
rect -701 -3126 -697 -3122
rect -691 -3169 -687 -3165
rect -677 -3119 -673 -3115
rect -667 -3133 -663 -3129
rect -657 -3169 -653 -3165
rect -643 -3119 -639 -3115
rect -639 -3177 -635 -3173
rect -623 -3148 -619 -3144
rect -613 -3162 -609 -3158
rect -599 -3119 -595 -3115
rect -599 -3140 -595 -3136
rect -595 -3155 -591 -3151
rect -579 -3162 -575 -3158
rect -565 -3119 -561 -3115
rect -555 -3170 -551 -3166
rect -539 -3177 -535 -3173
rect -525 -3133 -521 -3129
rect -521 -3170 -517 -3166
rect -435 -3119 -431 -3115
rect -439 -3140 -435 -3136
rect -435 -3155 -431 -3151
rect -439 -3169 -435 -3165
rect -409 -3140 -405 -3136
rect -413 -3148 -409 -3144
rect -413 -3162 -409 -3158
rect -393 -3126 -389 -3122
rect -383 -3169 -379 -3165
rect -369 -3119 -365 -3115
rect -359 -3133 -355 -3129
rect -349 -3169 -345 -3165
rect -335 -3119 -331 -3115
rect -331 -3177 -327 -3173
rect -315 -3148 -311 -3144
rect -305 -3162 -301 -3158
rect -291 -3119 -287 -3115
rect -291 -3140 -287 -3136
rect -287 -3155 -283 -3151
rect -271 -3162 -267 -3158
rect -257 -3119 -253 -3115
rect -247 -3170 -243 -3166
rect -231 -3177 -227 -3173
rect -217 -3133 -213 -3129
rect -213 -3170 -209 -3166
rect -127 -3119 -123 -3115
rect -131 -3140 -127 -3136
rect -127 -3155 -123 -3151
rect -131 -3169 -127 -3165
rect -101 -3140 -97 -3136
rect -105 -3148 -101 -3144
rect -105 -3162 -101 -3158
rect -85 -3126 -81 -3122
rect -75 -3169 -71 -3165
rect -61 -3119 -57 -3115
rect -51 -3133 -47 -3129
rect -41 -3169 -37 -3165
rect -27 -3119 -23 -3115
rect -23 -3177 -19 -3173
rect -7 -3148 -3 -3144
rect 3 -3162 7 -3158
rect 17 -3119 21 -3115
rect 17 -3140 21 -3136
rect 21 -3155 25 -3151
rect 37 -3162 41 -3158
rect 51 -3119 55 -3115
rect 61 -3170 65 -3166
rect 77 -3177 81 -3173
rect 91 -3133 95 -3129
rect 95 -3170 99 -3166
rect 181 -3119 185 -3115
rect 177 -3140 181 -3136
rect 181 -3155 185 -3151
rect 177 -3169 181 -3165
rect 207 -3140 211 -3136
rect 203 -3148 207 -3144
rect 203 -3162 207 -3158
rect 223 -3126 227 -3122
rect 233 -3169 237 -3165
rect 247 -3119 251 -3115
rect 257 -3133 261 -3129
rect 267 -3169 271 -3165
rect 281 -3119 285 -3115
rect 285 -3177 289 -3173
rect 301 -3148 305 -3144
rect 311 -3162 315 -3158
rect 325 -3119 329 -3115
rect 325 -3140 329 -3136
rect 329 -3155 333 -3151
rect 345 -3162 349 -3158
rect 359 -3119 363 -3115
rect 369 -3170 373 -3166
rect 385 -3177 389 -3173
rect 399 -3133 403 -3129
rect 403 -3170 407 -3166
rect 489 -3119 493 -3115
rect 485 -3140 489 -3136
rect 489 -3155 493 -3151
rect 485 -3169 489 -3165
rect 515 -3140 519 -3136
rect 511 -3148 515 -3144
rect 511 -3162 515 -3158
rect 531 -3126 535 -3122
rect 541 -3169 545 -3165
rect 555 -3119 559 -3115
rect 565 -3133 569 -3129
rect 575 -3169 579 -3165
rect 589 -3119 593 -3115
rect 593 -3177 597 -3173
rect 609 -3148 613 -3144
rect 619 -3162 623 -3158
rect 633 -3119 637 -3115
rect 633 -3140 637 -3136
rect 637 -3155 641 -3151
rect 653 -3162 657 -3158
rect 667 -3119 671 -3115
rect 677 -3170 681 -3166
rect 693 -3177 697 -3173
rect 707 -3133 711 -3129
rect 711 -3170 715 -3166
rect 797 -3119 801 -3115
rect 793 -3140 797 -3136
rect 797 -3155 801 -3151
rect 793 -3169 797 -3165
rect 823 -3140 827 -3136
rect 819 -3148 823 -3144
rect 819 -3162 823 -3158
rect 839 -3126 843 -3122
rect 849 -3169 853 -3165
rect 863 -3119 867 -3115
rect 873 -3133 877 -3129
rect 883 -3169 887 -3165
rect 897 -3119 901 -3115
rect 901 -3177 905 -3173
rect 917 -3148 921 -3144
rect 927 -3162 931 -3158
rect 941 -3119 945 -3115
rect 941 -3140 945 -3136
rect 945 -3155 949 -3151
rect 961 -3162 965 -3158
rect 975 -3119 979 -3115
rect 985 -3170 989 -3166
rect 1001 -3177 1005 -3173
rect 1015 -3133 1019 -3129
rect 1019 -3170 1023 -3166
<< ndcontact >>
rect -1307 -1068 -1303 -1064
rect -1290 -1068 -1286 -1064
rect -1281 -1068 -1277 -1064
rect -1063 -1068 -1059 -1064
rect -1046 -1068 -1042 -1064
rect -1037 -1068 -1033 -1064
rect -754 -1068 -750 -1064
rect -737 -1068 -733 -1064
rect -728 -1068 -724 -1064
rect -446 -1068 -442 -1064
rect -429 -1068 -425 -1064
rect -420 -1068 -416 -1064
rect -139 -1068 -135 -1064
rect -122 -1068 -118 -1064
rect -113 -1068 -109 -1064
rect 170 -1068 174 -1064
rect 187 -1068 191 -1064
rect 196 -1068 200 -1064
rect 478 -1068 482 -1064
rect 495 -1068 499 -1064
rect 504 -1068 508 -1064
rect 786 -1068 790 -1064
rect 803 -1068 807 -1064
rect 812 -1068 816 -1064
rect -1309 -1218 -1305 -1214
rect -1292 -1218 -1288 -1214
rect -1283 -1218 -1279 -1214
rect -1062 -1218 -1058 -1214
rect -1045 -1218 -1041 -1214
rect -1036 -1218 -1032 -1214
rect -754 -1218 -750 -1214
rect -737 -1218 -733 -1214
rect -728 -1218 -724 -1214
rect -446 -1218 -442 -1214
rect -429 -1218 -425 -1214
rect -420 -1218 -416 -1214
rect -138 -1218 -134 -1214
rect -121 -1218 -117 -1214
rect -112 -1218 -108 -1214
rect 170 -1218 174 -1214
rect 187 -1218 191 -1214
rect 196 -1218 200 -1214
rect 478 -1218 482 -1214
rect 495 -1218 499 -1214
rect 504 -1218 508 -1214
rect 786 -1218 790 -1214
rect 803 -1218 807 -1214
rect 812 -1218 816 -1214
rect -1230 -1382 -1226 -1378
rect -1221 -1382 -1217 -1378
rect -1212 -1382 -1208 -1378
rect -1204 -1382 -1200 -1378
rect -1195 -1382 -1191 -1378
rect -1177 -1382 -1173 -1378
rect -1168 -1382 -1164 -1378
rect -1160 -1382 -1156 -1378
rect -1143 -1382 -1139 -1378
rect -1134 -1382 -1130 -1378
rect -1062 -1382 -1058 -1378
rect -1053 -1382 -1049 -1378
rect -1044 -1382 -1040 -1378
rect -1036 -1382 -1032 -1378
rect -1027 -1382 -1023 -1378
rect -1018 -1382 -1014 -1378
rect -1010 -1382 -1006 -1378
rect -1002 -1382 -998 -1378
rect -984 -1382 -980 -1378
rect -974 -1382 -970 -1378
rect -966 -1382 -962 -1378
rect -949 -1382 -945 -1378
rect -940 -1382 -936 -1378
rect -932 -1382 -928 -1378
rect -923 -1382 -919 -1378
rect -905 -1382 -901 -1378
rect -896 -1382 -892 -1378
rect -888 -1382 -884 -1378
rect -872 -1382 -868 -1378
rect -864 -1382 -860 -1378
rect -852 -1382 -848 -1378
rect -840 -1382 -836 -1378
rect -831 -1382 -827 -1378
rect -822 -1382 -818 -1378
rect -754 -1382 -750 -1378
rect -745 -1382 -741 -1378
rect -736 -1382 -732 -1378
rect -728 -1382 -724 -1378
rect -719 -1382 -715 -1378
rect -710 -1382 -706 -1378
rect -702 -1382 -698 -1378
rect -694 -1382 -690 -1378
rect -676 -1382 -672 -1378
rect -666 -1382 -662 -1378
rect -658 -1382 -654 -1378
rect -641 -1382 -637 -1378
rect -632 -1382 -628 -1378
rect -624 -1382 -620 -1378
rect -615 -1382 -611 -1378
rect -597 -1382 -593 -1378
rect -588 -1382 -584 -1378
rect -580 -1382 -576 -1378
rect -564 -1382 -560 -1378
rect -556 -1382 -552 -1378
rect -544 -1382 -540 -1378
rect -532 -1382 -528 -1378
rect -523 -1382 -519 -1378
rect -514 -1382 -510 -1378
rect -446 -1382 -442 -1378
rect -437 -1382 -433 -1378
rect -428 -1382 -424 -1378
rect -420 -1382 -416 -1378
rect -411 -1382 -407 -1378
rect -402 -1382 -398 -1378
rect -394 -1382 -390 -1378
rect -386 -1382 -382 -1378
rect -368 -1382 -364 -1378
rect -358 -1382 -354 -1378
rect -350 -1382 -346 -1378
rect -333 -1382 -329 -1378
rect -324 -1382 -320 -1378
rect -316 -1382 -312 -1378
rect -307 -1382 -303 -1378
rect -289 -1382 -285 -1378
rect -280 -1382 -276 -1378
rect -272 -1382 -268 -1378
rect -256 -1382 -252 -1378
rect -248 -1382 -244 -1378
rect -236 -1382 -232 -1378
rect -224 -1382 -220 -1378
rect -215 -1382 -211 -1378
rect -206 -1382 -202 -1378
rect -138 -1382 -134 -1378
rect -129 -1382 -125 -1378
rect -120 -1382 -116 -1378
rect -112 -1382 -108 -1378
rect -103 -1382 -99 -1378
rect -94 -1382 -90 -1378
rect -86 -1382 -82 -1378
rect -78 -1382 -74 -1378
rect -60 -1382 -56 -1378
rect -50 -1382 -46 -1378
rect -42 -1382 -38 -1378
rect -25 -1382 -21 -1378
rect -16 -1382 -12 -1378
rect -8 -1382 -4 -1378
rect 1 -1382 5 -1378
rect 19 -1382 23 -1378
rect 28 -1382 32 -1378
rect 36 -1382 40 -1378
rect 52 -1382 56 -1378
rect 60 -1382 64 -1378
rect 72 -1382 76 -1378
rect 84 -1382 88 -1378
rect 93 -1382 97 -1378
rect 102 -1382 106 -1378
rect 170 -1382 174 -1378
rect 179 -1382 183 -1378
rect 188 -1382 192 -1378
rect 196 -1382 200 -1378
rect 205 -1382 209 -1378
rect 214 -1382 218 -1378
rect 222 -1382 226 -1378
rect 230 -1382 234 -1378
rect 248 -1382 252 -1378
rect 258 -1382 262 -1378
rect 266 -1382 270 -1378
rect 283 -1382 287 -1378
rect 292 -1382 296 -1378
rect 300 -1382 304 -1378
rect 309 -1382 313 -1378
rect 327 -1382 331 -1378
rect 336 -1382 340 -1378
rect 344 -1382 348 -1378
rect 360 -1382 364 -1378
rect 368 -1382 372 -1378
rect 380 -1382 384 -1378
rect 392 -1382 396 -1378
rect 401 -1382 405 -1378
rect 410 -1382 414 -1378
rect 478 -1382 482 -1378
rect 487 -1382 491 -1378
rect 496 -1382 500 -1378
rect 504 -1382 508 -1378
rect 513 -1382 517 -1378
rect 522 -1382 526 -1378
rect 530 -1382 534 -1378
rect 538 -1382 542 -1378
rect 556 -1382 560 -1378
rect 566 -1382 570 -1378
rect 574 -1382 578 -1378
rect 591 -1382 595 -1378
rect 600 -1382 604 -1378
rect 608 -1382 612 -1378
rect 617 -1382 621 -1378
rect 635 -1382 639 -1378
rect 644 -1382 648 -1378
rect 652 -1382 656 -1378
rect 668 -1382 672 -1378
rect 676 -1382 680 -1378
rect 688 -1382 692 -1378
rect 700 -1382 704 -1378
rect 709 -1382 713 -1378
rect 718 -1382 722 -1378
rect 784 -1382 788 -1378
rect 793 -1382 797 -1378
rect 802 -1382 806 -1378
rect 810 -1382 814 -1378
rect 819 -1382 823 -1378
rect 837 -1382 841 -1378
rect 846 -1382 850 -1378
rect 854 -1382 858 -1378
rect 871 -1382 875 -1378
rect 880 -1382 884 -1378
rect -1309 -1539 -1305 -1535
rect -1292 -1539 -1288 -1535
rect -1283 -1539 -1279 -1535
rect -1062 -1539 -1058 -1535
rect -1045 -1539 -1041 -1535
rect -1036 -1539 -1032 -1535
rect -754 -1539 -750 -1535
rect -737 -1539 -733 -1535
rect -728 -1539 -724 -1535
rect -446 -1539 -442 -1535
rect -429 -1539 -425 -1535
rect -420 -1539 -416 -1535
rect -138 -1539 -134 -1535
rect -121 -1539 -117 -1535
rect -112 -1539 -108 -1535
rect 170 -1539 174 -1535
rect 187 -1539 191 -1535
rect 196 -1539 200 -1535
rect 478 -1539 482 -1535
rect 495 -1539 499 -1535
rect 504 -1539 508 -1535
rect 786 -1539 790 -1535
rect 803 -1539 807 -1535
rect 812 -1539 816 -1535
rect -1234 -1698 -1230 -1694
rect -1225 -1698 -1221 -1694
rect -1216 -1698 -1212 -1694
rect -1208 -1698 -1204 -1694
rect -1199 -1698 -1195 -1694
rect -1181 -1698 -1177 -1694
rect -1172 -1698 -1168 -1694
rect -1164 -1698 -1160 -1694
rect -1147 -1698 -1143 -1694
rect -1138 -1698 -1134 -1694
rect -1062 -1698 -1058 -1694
rect -1053 -1698 -1049 -1694
rect -1044 -1698 -1040 -1694
rect -1036 -1698 -1032 -1694
rect -1027 -1698 -1023 -1694
rect -1018 -1698 -1014 -1694
rect -1010 -1698 -1006 -1694
rect -1002 -1698 -998 -1694
rect -984 -1698 -980 -1694
rect -974 -1698 -970 -1694
rect -966 -1698 -962 -1694
rect -949 -1698 -945 -1694
rect -940 -1698 -936 -1694
rect -932 -1698 -928 -1694
rect -923 -1698 -919 -1694
rect -905 -1698 -901 -1694
rect -896 -1698 -892 -1694
rect -888 -1698 -884 -1694
rect -872 -1698 -868 -1694
rect -864 -1698 -860 -1694
rect -852 -1698 -848 -1694
rect -840 -1698 -836 -1694
rect -831 -1698 -827 -1694
rect -822 -1698 -818 -1694
rect -754 -1698 -750 -1694
rect -745 -1698 -741 -1694
rect -736 -1698 -732 -1694
rect -728 -1698 -724 -1694
rect -719 -1698 -715 -1694
rect -710 -1698 -706 -1694
rect -702 -1698 -698 -1694
rect -694 -1698 -690 -1694
rect -676 -1698 -672 -1694
rect -666 -1698 -662 -1694
rect -658 -1698 -654 -1694
rect -641 -1698 -637 -1694
rect -632 -1698 -628 -1694
rect -624 -1698 -620 -1694
rect -615 -1698 -611 -1694
rect -597 -1698 -593 -1694
rect -588 -1698 -584 -1694
rect -580 -1698 -576 -1694
rect -564 -1698 -560 -1694
rect -556 -1698 -552 -1694
rect -544 -1698 -540 -1694
rect -532 -1698 -528 -1694
rect -523 -1698 -519 -1694
rect -514 -1698 -510 -1694
rect -446 -1698 -442 -1694
rect -437 -1698 -433 -1694
rect -428 -1698 -424 -1694
rect -420 -1698 -416 -1694
rect -411 -1698 -407 -1694
rect -402 -1698 -398 -1694
rect -394 -1698 -390 -1694
rect -386 -1698 -382 -1694
rect -368 -1698 -364 -1694
rect -358 -1698 -354 -1694
rect -350 -1698 -346 -1694
rect -333 -1698 -329 -1694
rect -324 -1698 -320 -1694
rect -316 -1698 -312 -1694
rect -307 -1698 -303 -1694
rect -289 -1698 -285 -1694
rect -280 -1698 -276 -1694
rect -272 -1698 -268 -1694
rect -256 -1698 -252 -1694
rect -248 -1698 -244 -1694
rect -236 -1698 -232 -1694
rect -224 -1698 -220 -1694
rect -215 -1698 -211 -1694
rect -206 -1698 -202 -1694
rect -138 -1698 -134 -1694
rect -129 -1698 -125 -1694
rect -120 -1698 -116 -1694
rect -112 -1698 -108 -1694
rect -103 -1698 -99 -1694
rect -94 -1698 -90 -1694
rect -86 -1698 -82 -1694
rect -78 -1698 -74 -1694
rect -60 -1698 -56 -1694
rect -50 -1698 -46 -1694
rect -42 -1698 -38 -1694
rect -25 -1698 -21 -1694
rect -16 -1698 -12 -1694
rect -8 -1698 -4 -1694
rect 1 -1698 5 -1694
rect 19 -1698 23 -1694
rect 28 -1698 32 -1694
rect 36 -1698 40 -1694
rect 52 -1698 56 -1694
rect 60 -1698 64 -1694
rect 72 -1698 76 -1694
rect 84 -1698 88 -1694
rect 93 -1698 97 -1694
rect 102 -1698 106 -1694
rect 170 -1698 174 -1694
rect 179 -1698 183 -1694
rect 188 -1698 192 -1694
rect 196 -1698 200 -1694
rect 205 -1698 209 -1694
rect 214 -1698 218 -1694
rect 222 -1698 226 -1694
rect 230 -1698 234 -1694
rect 248 -1698 252 -1694
rect 258 -1698 262 -1694
rect 266 -1698 270 -1694
rect 283 -1698 287 -1694
rect 292 -1698 296 -1694
rect 300 -1698 304 -1694
rect 309 -1698 313 -1694
rect 327 -1698 331 -1694
rect 336 -1698 340 -1694
rect 344 -1698 348 -1694
rect 360 -1698 364 -1694
rect 368 -1698 372 -1694
rect 380 -1698 384 -1694
rect 392 -1698 396 -1694
rect 401 -1698 405 -1694
rect 410 -1698 414 -1694
rect 478 -1698 482 -1694
rect 487 -1698 491 -1694
rect 496 -1698 500 -1694
rect 504 -1698 508 -1694
rect 513 -1698 517 -1694
rect 522 -1698 526 -1694
rect 530 -1698 534 -1694
rect 538 -1698 542 -1694
rect 556 -1698 560 -1694
rect 566 -1698 570 -1694
rect 574 -1698 578 -1694
rect 591 -1698 595 -1694
rect 600 -1698 604 -1694
rect 608 -1698 612 -1694
rect 617 -1698 621 -1694
rect 635 -1698 639 -1694
rect 644 -1698 648 -1694
rect 652 -1698 656 -1694
rect 668 -1698 672 -1694
rect 676 -1698 680 -1694
rect 688 -1698 692 -1694
rect 700 -1698 704 -1694
rect 709 -1698 713 -1694
rect 718 -1698 722 -1694
rect 786 -1698 790 -1694
rect 795 -1698 799 -1694
rect 804 -1698 808 -1694
rect 812 -1698 816 -1694
rect 821 -1698 825 -1694
rect 830 -1698 834 -1694
rect 838 -1698 842 -1694
rect 846 -1698 850 -1694
rect 864 -1698 868 -1694
rect 874 -1698 878 -1694
rect 882 -1698 886 -1694
rect 899 -1698 903 -1694
rect 908 -1698 912 -1694
rect 916 -1698 920 -1694
rect 925 -1698 929 -1694
rect 943 -1698 947 -1694
rect 952 -1698 956 -1694
rect 960 -1698 964 -1694
rect 976 -1698 980 -1694
rect 984 -1698 988 -1694
rect 996 -1698 1000 -1694
rect 1008 -1698 1012 -1694
rect 1017 -1698 1021 -1694
rect 1026 -1698 1030 -1694
rect -1309 -1830 -1305 -1826
rect -1292 -1830 -1288 -1826
rect -1283 -1830 -1279 -1826
rect -1062 -1830 -1058 -1826
rect -1045 -1830 -1041 -1826
rect -1036 -1830 -1032 -1826
rect -754 -1830 -750 -1826
rect -737 -1830 -733 -1826
rect -728 -1830 -724 -1826
rect -446 -1830 -442 -1826
rect -429 -1830 -425 -1826
rect -420 -1830 -416 -1826
rect -138 -1830 -134 -1826
rect -121 -1830 -117 -1826
rect -112 -1830 -108 -1826
rect 170 -1830 174 -1826
rect 187 -1830 191 -1826
rect 196 -1830 200 -1826
rect 478 -1830 482 -1826
rect 495 -1830 499 -1826
rect 504 -1830 508 -1826
rect 786 -1830 790 -1826
rect 803 -1830 807 -1826
rect 812 -1830 816 -1826
rect -1234 -1989 -1230 -1985
rect -1225 -1989 -1221 -1985
rect -1216 -1989 -1212 -1985
rect -1208 -1989 -1204 -1985
rect -1199 -1989 -1195 -1985
rect -1181 -1989 -1177 -1985
rect -1172 -1989 -1168 -1985
rect -1164 -1989 -1160 -1985
rect -1147 -1989 -1143 -1985
rect -1138 -1989 -1134 -1985
rect -1062 -1989 -1058 -1985
rect -1053 -1989 -1049 -1985
rect -1044 -1989 -1040 -1985
rect -1036 -1989 -1032 -1985
rect -1027 -1989 -1023 -1985
rect -1018 -1989 -1014 -1985
rect -1010 -1989 -1006 -1985
rect -1002 -1989 -998 -1985
rect -984 -1989 -980 -1985
rect -974 -1989 -970 -1985
rect -966 -1989 -962 -1985
rect -949 -1989 -945 -1985
rect -940 -1989 -936 -1985
rect -932 -1989 -928 -1985
rect -923 -1989 -919 -1985
rect -905 -1989 -901 -1985
rect -896 -1989 -892 -1985
rect -888 -1989 -884 -1985
rect -872 -1989 -868 -1985
rect -864 -1989 -860 -1985
rect -852 -1989 -848 -1985
rect -840 -1989 -836 -1985
rect -831 -1989 -827 -1985
rect -822 -1989 -818 -1985
rect -754 -1989 -750 -1985
rect -745 -1989 -741 -1985
rect -736 -1989 -732 -1985
rect -728 -1989 -724 -1985
rect -719 -1989 -715 -1985
rect -710 -1989 -706 -1985
rect -702 -1989 -698 -1985
rect -694 -1989 -690 -1985
rect -676 -1989 -672 -1985
rect -666 -1989 -662 -1985
rect -658 -1989 -654 -1985
rect -641 -1989 -637 -1985
rect -632 -1989 -628 -1985
rect -624 -1989 -620 -1985
rect -615 -1989 -611 -1985
rect -597 -1989 -593 -1985
rect -588 -1989 -584 -1985
rect -580 -1989 -576 -1985
rect -564 -1989 -560 -1985
rect -556 -1989 -552 -1985
rect -544 -1989 -540 -1985
rect -532 -1989 -528 -1985
rect -523 -1989 -519 -1985
rect -514 -1989 -510 -1985
rect -446 -1989 -442 -1985
rect -437 -1989 -433 -1985
rect -428 -1989 -424 -1985
rect -420 -1989 -416 -1985
rect -411 -1989 -407 -1985
rect -402 -1989 -398 -1985
rect -394 -1989 -390 -1985
rect -386 -1989 -382 -1985
rect -368 -1989 -364 -1985
rect -358 -1989 -354 -1985
rect -350 -1989 -346 -1985
rect -333 -1989 -329 -1985
rect -324 -1989 -320 -1985
rect -316 -1989 -312 -1985
rect -307 -1989 -303 -1985
rect -289 -1989 -285 -1985
rect -280 -1989 -276 -1985
rect -272 -1989 -268 -1985
rect -256 -1989 -252 -1985
rect -248 -1989 -244 -1985
rect -236 -1989 -232 -1985
rect -224 -1989 -220 -1985
rect -215 -1989 -211 -1985
rect -206 -1989 -202 -1985
rect -138 -1989 -134 -1985
rect -129 -1989 -125 -1985
rect -120 -1989 -116 -1985
rect -112 -1989 -108 -1985
rect -103 -1989 -99 -1985
rect -94 -1989 -90 -1985
rect -86 -1989 -82 -1985
rect -78 -1989 -74 -1985
rect -60 -1989 -56 -1985
rect -50 -1989 -46 -1985
rect -42 -1989 -38 -1985
rect -25 -1989 -21 -1985
rect -16 -1989 -12 -1985
rect -8 -1989 -4 -1985
rect 1 -1989 5 -1985
rect 19 -1989 23 -1985
rect 28 -1989 32 -1985
rect 36 -1989 40 -1985
rect 52 -1989 56 -1985
rect 60 -1989 64 -1985
rect 72 -1989 76 -1985
rect 84 -1989 88 -1985
rect 93 -1989 97 -1985
rect 102 -1989 106 -1985
rect 170 -1989 174 -1985
rect 179 -1989 183 -1985
rect 188 -1989 192 -1985
rect 196 -1989 200 -1985
rect 205 -1989 209 -1985
rect 214 -1989 218 -1985
rect 222 -1989 226 -1985
rect 230 -1989 234 -1985
rect 248 -1989 252 -1985
rect 258 -1989 262 -1985
rect 266 -1989 270 -1985
rect 283 -1989 287 -1985
rect 292 -1989 296 -1985
rect 300 -1989 304 -1985
rect 309 -1989 313 -1985
rect 327 -1989 331 -1985
rect 336 -1989 340 -1985
rect 344 -1989 348 -1985
rect 360 -1989 364 -1985
rect 368 -1989 372 -1985
rect 380 -1989 384 -1985
rect 392 -1989 396 -1985
rect 401 -1989 405 -1985
rect 410 -1989 414 -1985
rect 478 -1989 482 -1985
rect 487 -1989 491 -1985
rect 496 -1989 500 -1985
rect 504 -1989 508 -1985
rect 513 -1989 517 -1985
rect 522 -1989 526 -1985
rect 530 -1989 534 -1985
rect 538 -1989 542 -1985
rect 556 -1989 560 -1985
rect 566 -1989 570 -1985
rect 574 -1989 578 -1985
rect 591 -1989 595 -1985
rect 600 -1989 604 -1985
rect 608 -1989 612 -1985
rect 617 -1989 621 -1985
rect 635 -1989 639 -1985
rect 644 -1989 648 -1985
rect 652 -1989 656 -1985
rect 668 -1989 672 -1985
rect 676 -1989 680 -1985
rect 688 -1989 692 -1985
rect 700 -1989 704 -1985
rect 709 -1989 713 -1985
rect 718 -1989 722 -1985
rect 786 -1989 790 -1985
rect 795 -1989 799 -1985
rect 804 -1989 808 -1985
rect 812 -1989 816 -1985
rect 821 -1989 825 -1985
rect 830 -1989 834 -1985
rect 838 -1989 842 -1985
rect 846 -1989 850 -1985
rect 864 -1989 868 -1985
rect 874 -1989 878 -1985
rect 882 -1989 886 -1985
rect 899 -1989 903 -1985
rect 908 -1989 912 -1985
rect 916 -1989 920 -1985
rect 925 -1989 929 -1985
rect 943 -1989 947 -1985
rect 952 -1989 956 -1985
rect 960 -1989 964 -1985
rect 976 -1989 980 -1985
rect 984 -1989 988 -1985
rect 996 -1989 1000 -1985
rect 1008 -1989 1012 -1985
rect 1017 -1989 1021 -1985
rect 1026 -1989 1030 -1985
rect -1309 -2152 -1305 -2148
rect -1292 -2152 -1288 -2148
rect -1283 -2152 -1279 -2148
rect -1062 -2152 -1058 -2148
rect -1045 -2152 -1041 -2148
rect -1036 -2152 -1032 -2148
rect -754 -2152 -750 -2148
rect -737 -2152 -733 -2148
rect -728 -2152 -724 -2148
rect -446 -2152 -442 -2148
rect -429 -2152 -425 -2148
rect -420 -2152 -416 -2148
rect -138 -2152 -134 -2148
rect -121 -2152 -117 -2148
rect -112 -2152 -108 -2148
rect 170 -2152 174 -2148
rect 187 -2152 191 -2148
rect 196 -2152 200 -2148
rect 478 -2152 482 -2148
rect 495 -2152 499 -2148
rect 504 -2152 508 -2148
rect 786 -2152 790 -2148
rect 803 -2152 807 -2148
rect 812 -2152 816 -2148
rect -1234 -2311 -1230 -2307
rect -1225 -2311 -1221 -2307
rect -1216 -2311 -1212 -2307
rect -1208 -2311 -1204 -2307
rect -1199 -2311 -1195 -2307
rect -1181 -2311 -1177 -2307
rect -1172 -2311 -1168 -2307
rect -1164 -2311 -1160 -2307
rect -1147 -2311 -1143 -2307
rect -1138 -2311 -1134 -2307
rect -1062 -2311 -1058 -2307
rect -1053 -2311 -1049 -2307
rect -1044 -2311 -1040 -2307
rect -1036 -2311 -1032 -2307
rect -1027 -2311 -1023 -2307
rect -1018 -2311 -1014 -2307
rect -1010 -2311 -1006 -2307
rect -1002 -2311 -998 -2307
rect -984 -2311 -980 -2307
rect -974 -2311 -970 -2307
rect -966 -2311 -962 -2307
rect -949 -2311 -945 -2307
rect -940 -2311 -936 -2307
rect -932 -2311 -928 -2307
rect -923 -2311 -919 -2307
rect -905 -2311 -901 -2307
rect -896 -2311 -892 -2307
rect -888 -2311 -884 -2307
rect -872 -2311 -868 -2307
rect -864 -2311 -860 -2307
rect -852 -2311 -848 -2307
rect -840 -2311 -836 -2307
rect -831 -2311 -827 -2307
rect -822 -2311 -818 -2307
rect -754 -2311 -750 -2307
rect -745 -2311 -741 -2307
rect -736 -2311 -732 -2307
rect -728 -2311 -724 -2307
rect -719 -2311 -715 -2307
rect -710 -2311 -706 -2307
rect -702 -2311 -698 -2307
rect -694 -2311 -690 -2307
rect -676 -2311 -672 -2307
rect -666 -2311 -662 -2307
rect -658 -2311 -654 -2307
rect -641 -2311 -637 -2307
rect -632 -2311 -628 -2307
rect -624 -2311 -620 -2307
rect -615 -2311 -611 -2307
rect -597 -2311 -593 -2307
rect -588 -2311 -584 -2307
rect -580 -2311 -576 -2307
rect -564 -2311 -560 -2307
rect -556 -2311 -552 -2307
rect -544 -2311 -540 -2307
rect -532 -2311 -528 -2307
rect -523 -2311 -519 -2307
rect -514 -2311 -510 -2307
rect -446 -2311 -442 -2307
rect -437 -2311 -433 -2307
rect -428 -2311 -424 -2307
rect -420 -2311 -416 -2307
rect -411 -2311 -407 -2307
rect -402 -2311 -398 -2307
rect -394 -2311 -390 -2307
rect -386 -2311 -382 -2307
rect -368 -2311 -364 -2307
rect -358 -2311 -354 -2307
rect -350 -2311 -346 -2307
rect -333 -2311 -329 -2307
rect -324 -2311 -320 -2307
rect -316 -2311 -312 -2307
rect -307 -2311 -303 -2307
rect -289 -2311 -285 -2307
rect -280 -2311 -276 -2307
rect -272 -2311 -268 -2307
rect -256 -2311 -252 -2307
rect -248 -2311 -244 -2307
rect -236 -2311 -232 -2307
rect -224 -2311 -220 -2307
rect -215 -2311 -211 -2307
rect -206 -2311 -202 -2307
rect -138 -2311 -134 -2307
rect -129 -2311 -125 -2307
rect -120 -2311 -116 -2307
rect -112 -2311 -108 -2307
rect -103 -2311 -99 -2307
rect -94 -2311 -90 -2307
rect -86 -2311 -82 -2307
rect -78 -2311 -74 -2307
rect -60 -2311 -56 -2307
rect -50 -2311 -46 -2307
rect -42 -2311 -38 -2307
rect -25 -2311 -21 -2307
rect -16 -2311 -12 -2307
rect -8 -2311 -4 -2307
rect 1 -2311 5 -2307
rect 19 -2311 23 -2307
rect 28 -2311 32 -2307
rect 36 -2311 40 -2307
rect 52 -2311 56 -2307
rect 60 -2311 64 -2307
rect 72 -2311 76 -2307
rect 84 -2311 88 -2307
rect 93 -2311 97 -2307
rect 102 -2311 106 -2307
rect 170 -2311 174 -2307
rect 179 -2311 183 -2307
rect 188 -2311 192 -2307
rect 196 -2311 200 -2307
rect 205 -2311 209 -2307
rect 214 -2311 218 -2307
rect 222 -2311 226 -2307
rect 230 -2311 234 -2307
rect 248 -2311 252 -2307
rect 258 -2311 262 -2307
rect 266 -2311 270 -2307
rect 283 -2311 287 -2307
rect 292 -2311 296 -2307
rect 300 -2311 304 -2307
rect 309 -2311 313 -2307
rect 327 -2311 331 -2307
rect 336 -2311 340 -2307
rect 344 -2311 348 -2307
rect 360 -2311 364 -2307
rect 368 -2311 372 -2307
rect 380 -2311 384 -2307
rect 392 -2311 396 -2307
rect 401 -2311 405 -2307
rect 410 -2311 414 -2307
rect 478 -2311 482 -2307
rect 487 -2311 491 -2307
rect 496 -2311 500 -2307
rect 504 -2311 508 -2307
rect 513 -2311 517 -2307
rect 522 -2311 526 -2307
rect 530 -2311 534 -2307
rect 538 -2311 542 -2307
rect 556 -2311 560 -2307
rect 566 -2311 570 -2307
rect 574 -2311 578 -2307
rect 591 -2311 595 -2307
rect 600 -2311 604 -2307
rect 608 -2311 612 -2307
rect 617 -2311 621 -2307
rect 635 -2311 639 -2307
rect 644 -2311 648 -2307
rect 652 -2311 656 -2307
rect 668 -2311 672 -2307
rect 676 -2311 680 -2307
rect 688 -2311 692 -2307
rect 700 -2311 704 -2307
rect 709 -2311 713 -2307
rect 718 -2311 722 -2307
rect 786 -2311 790 -2307
rect 795 -2311 799 -2307
rect 804 -2311 808 -2307
rect 812 -2311 816 -2307
rect 821 -2311 825 -2307
rect 830 -2311 834 -2307
rect 838 -2311 842 -2307
rect 846 -2311 850 -2307
rect 864 -2311 868 -2307
rect 874 -2311 878 -2307
rect 882 -2311 886 -2307
rect 899 -2311 903 -2307
rect 908 -2311 912 -2307
rect 916 -2311 920 -2307
rect 925 -2311 929 -2307
rect 943 -2311 947 -2307
rect 952 -2311 956 -2307
rect 960 -2311 964 -2307
rect 976 -2311 980 -2307
rect 984 -2311 988 -2307
rect 996 -2311 1000 -2307
rect 1008 -2311 1012 -2307
rect 1017 -2311 1021 -2307
rect 1026 -2311 1030 -2307
rect -1309 -2443 -1305 -2439
rect -1292 -2443 -1288 -2439
rect -1283 -2443 -1279 -2439
rect -1062 -2443 -1058 -2439
rect -1045 -2443 -1041 -2439
rect -1036 -2443 -1032 -2439
rect -754 -2443 -750 -2439
rect -737 -2443 -733 -2439
rect -728 -2443 -724 -2439
rect -446 -2443 -442 -2439
rect -429 -2443 -425 -2439
rect -420 -2443 -416 -2439
rect -138 -2443 -134 -2439
rect -121 -2443 -117 -2439
rect -112 -2443 -108 -2439
rect 170 -2443 174 -2439
rect 187 -2443 191 -2439
rect 196 -2443 200 -2439
rect 478 -2443 482 -2439
rect 495 -2443 499 -2439
rect 504 -2443 508 -2439
rect 786 -2443 790 -2439
rect 803 -2443 807 -2439
rect 812 -2443 816 -2439
rect -1234 -2602 -1230 -2598
rect -1225 -2602 -1221 -2598
rect -1216 -2602 -1212 -2598
rect -1208 -2602 -1204 -2598
rect -1199 -2602 -1195 -2598
rect -1181 -2602 -1177 -2598
rect -1172 -2602 -1168 -2598
rect -1164 -2602 -1160 -2598
rect -1147 -2602 -1143 -2598
rect -1138 -2602 -1134 -2598
rect -1062 -2602 -1058 -2598
rect -1053 -2602 -1049 -2598
rect -1044 -2602 -1040 -2598
rect -1036 -2602 -1032 -2598
rect -1027 -2602 -1023 -2598
rect -1018 -2602 -1014 -2598
rect -1010 -2602 -1006 -2598
rect -1002 -2602 -998 -2598
rect -984 -2602 -980 -2598
rect -974 -2602 -970 -2598
rect -966 -2602 -962 -2598
rect -949 -2602 -945 -2598
rect -940 -2602 -936 -2598
rect -932 -2602 -928 -2598
rect -923 -2602 -919 -2598
rect -905 -2602 -901 -2598
rect -896 -2602 -892 -2598
rect -888 -2602 -884 -2598
rect -872 -2602 -868 -2598
rect -864 -2602 -860 -2598
rect -852 -2602 -848 -2598
rect -840 -2602 -836 -2598
rect -831 -2602 -827 -2598
rect -822 -2602 -818 -2598
rect -754 -2602 -750 -2598
rect -745 -2602 -741 -2598
rect -736 -2602 -732 -2598
rect -728 -2602 -724 -2598
rect -719 -2602 -715 -2598
rect -710 -2602 -706 -2598
rect -702 -2602 -698 -2598
rect -694 -2602 -690 -2598
rect -676 -2602 -672 -2598
rect -666 -2602 -662 -2598
rect -658 -2602 -654 -2598
rect -641 -2602 -637 -2598
rect -632 -2602 -628 -2598
rect -624 -2602 -620 -2598
rect -615 -2602 -611 -2598
rect -597 -2602 -593 -2598
rect -588 -2602 -584 -2598
rect -580 -2602 -576 -2598
rect -564 -2602 -560 -2598
rect -556 -2602 -552 -2598
rect -544 -2602 -540 -2598
rect -532 -2602 -528 -2598
rect -523 -2602 -519 -2598
rect -514 -2602 -510 -2598
rect -446 -2602 -442 -2598
rect -437 -2602 -433 -2598
rect -428 -2602 -424 -2598
rect -420 -2602 -416 -2598
rect -411 -2602 -407 -2598
rect -402 -2602 -398 -2598
rect -394 -2602 -390 -2598
rect -386 -2602 -382 -2598
rect -368 -2602 -364 -2598
rect -358 -2602 -354 -2598
rect -350 -2602 -346 -2598
rect -333 -2602 -329 -2598
rect -324 -2602 -320 -2598
rect -316 -2602 -312 -2598
rect -307 -2602 -303 -2598
rect -289 -2602 -285 -2598
rect -280 -2602 -276 -2598
rect -272 -2602 -268 -2598
rect -256 -2602 -252 -2598
rect -248 -2602 -244 -2598
rect -236 -2602 -232 -2598
rect -224 -2602 -220 -2598
rect -215 -2602 -211 -2598
rect -206 -2602 -202 -2598
rect -138 -2602 -134 -2598
rect -129 -2602 -125 -2598
rect -120 -2602 -116 -2598
rect -112 -2602 -108 -2598
rect -103 -2602 -99 -2598
rect -94 -2602 -90 -2598
rect -86 -2602 -82 -2598
rect -78 -2602 -74 -2598
rect -60 -2602 -56 -2598
rect -50 -2602 -46 -2598
rect -42 -2602 -38 -2598
rect -25 -2602 -21 -2598
rect -16 -2602 -12 -2598
rect -8 -2602 -4 -2598
rect 1 -2602 5 -2598
rect 19 -2602 23 -2598
rect 28 -2602 32 -2598
rect 36 -2602 40 -2598
rect 52 -2602 56 -2598
rect 60 -2602 64 -2598
rect 72 -2602 76 -2598
rect 84 -2602 88 -2598
rect 93 -2602 97 -2598
rect 102 -2602 106 -2598
rect 170 -2602 174 -2598
rect 179 -2602 183 -2598
rect 188 -2602 192 -2598
rect 196 -2602 200 -2598
rect 205 -2602 209 -2598
rect 214 -2602 218 -2598
rect 222 -2602 226 -2598
rect 230 -2602 234 -2598
rect 248 -2602 252 -2598
rect 258 -2602 262 -2598
rect 266 -2602 270 -2598
rect 283 -2602 287 -2598
rect 292 -2602 296 -2598
rect 300 -2602 304 -2598
rect 309 -2602 313 -2598
rect 327 -2602 331 -2598
rect 336 -2602 340 -2598
rect 344 -2602 348 -2598
rect 360 -2602 364 -2598
rect 368 -2602 372 -2598
rect 380 -2602 384 -2598
rect 392 -2602 396 -2598
rect 401 -2602 405 -2598
rect 410 -2602 414 -2598
rect 478 -2602 482 -2598
rect 487 -2602 491 -2598
rect 496 -2602 500 -2598
rect 504 -2602 508 -2598
rect 513 -2602 517 -2598
rect 522 -2602 526 -2598
rect 530 -2602 534 -2598
rect 538 -2602 542 -2598
rect 556 -2602 560 -2598
rect 566 -2602 570 -2598
rect 574 -2602 578 -2598
rect 591 -2602 595 -2598
rect 600 -2602 604 -2598
rect 608 -2602 612 -2598
rect 617 -2602 621 -2598
rect 635 -2602 639 -2598
rect 644 -2602 648 -2598
rect 652 -2602 656 -2598
rect 668 -2602 672 -2598
rect 676 -2602 680 -2598
rect 688 -2602 692 -2598
rect 700 -2602 704 -2598
rect 709 -2602 713 -2598
rect 718 -2602 722 -2598
rect 786 -2602 790 -2598
rect 795 -2602 799 -2598
rect 804 -2602 808 -2598
rect 812 -2602 816 -2598
rect 821 -2602 825 -2598
rect 830 -2602 834 -2598
rect 838 -2602 842 -2598
rect 846 -2602 850 -2598
rect 864 -2602 868 -2598
rect 874 -2602 878 -2598
rect 882 -2602 886 -2598
rect 899 -2602 903 -2598
rect 908 -2602 912 -2598
rect 916 -2602 920 -2598
rect 925 -2602 929 -2598
rect 943 -2602 947 -2598
rect 952 -2602 956 -2598
rect 960 -2602 964 -2598
rect 976 -2602 980 -2598
rect 984 -2602 988 -2598
rect 996 -2602 1000 -2598
rect 1008 -2602 1012 -2598
rect 1017 -2602 1021 -2598
rect 1026 -2602 1030 -2598
rect -1309 -2734 -1305 -2730
rect -1292 -2734 -1288 -2730
rect -1283 -2734 -1279 -2730
rect -1062 -2734 -1058 -2730
rect -1045 -2734 -1041 -2730
rect -1036 -2734 -1032 -2730
rect -754 -2734 -750 -2730
rect -737 -2734 -733 -2730
rect -728 -2734 -724 -2730
rect -446 -2734 -442 -2730
rect -429 -2734 -425 -2730
rect -420 -2734 -416 -2730
rect -138 -2734 -134 -2730
rect -121 -2734 -117 -2730
rect -112 -2734 -108 -2730
rect 170 -2734 174 -2730
rect 187 -2734 191 -2730
rect 196 -2734 200 -2730
rect 478 -2734 482 -2730
rect 495 -2734 499 -2730
rect 504 -2734 508 -2730
rect 786 -2734 790 -2730
rect 803 -2734 807 -2730
rect 812 -2734 816 -2730
rect -1234 -2893 -1230 -2889
rect -1225 -2893 -1221 -2889
rect -1216 -2893 -1212 -2889
rect -1208 -2893 -1204 -2889
rect -1199 -2893 -1195 -2889
rect -1181 -2893 -1177 -2889
rect -1172 -2893 -1168 -2889
rect -1164 -2893 -1160 -2889
rect -1147 -2893 -1143 -2889
rect -1138 -2893 -1134 -2889
rect -1062 -2893 -1058 -2889
rect -1053 -2893 -1049 -2889
rect -1044 -2893 -1040 -2889
rect -1036 -2893 -1032 -2889
rect -1027 -2893 -1023 -2889
rect -1018 -2893 -1014 -2889
rect -1010 -2893 -1006 -2889
rect -1002 -2893 -998 -2889
rect -984 -2893 -980 -2889
rect -974 -2893 -970 -2889
rect -966 -2893 -962 -2889
rect -949 -2893 -945 -2889
rect -940 -2893 -936 -2889
rect -932 -2893 -928 -2889
rect -923 -2893 -919 -2889
rect -905 -2893 -901 -2889
rect -896 -2893 -892 -2889
rect -888 -2893 -884 -2889
rect -872 -2893 -868 -2889
rect -864 -2893 -860 -2889
rect -852 -2893 -848 -2889
rect -840 -2893 -836 -2889
rect -831 -2893 -827 -2889
rect -822 -2893 -818 -2889
rect -754 -2893 -750 -2889
rect -745 -2893 -741 -2889
rect -736 -2893 -732 -2889
rect -728 -2893 -724 -2889
rect -719 -2893 -715 -2889
rect -710 -2893 -706 -2889
rect -702 -2893 -698 -2889
rect -694 -2893 -690 -2889
rect -676 -2893 -672 -2889
rect -666 -2893 -662 -2889
rect -658 -2893 -654 -2889
rect -641 -2893 -637 -2889
rect -632 -2893 -628 -2889
rect -624 -2893 -620 -2889
rect -615 -2893 -611 -2889
rect -597 -2893 -593 -2889
rect -588 -2893 -584 -2889
rect -580 -2893 -576 -2889
rect -564 -2893 -560 -2889
rect -556 -2893 -552 -2889
rect -544 -2893 -540 -2889
rect -532 -2893 -528 -2889
rect -523 -2893 -519 -2889
rect -514 -2893 -510 -2889
rect -446 -2893 -442 -2889
rect -437 -2893 -433 -2889
rect -428 -2893 -424 -2889
rect -420 -2893 -416 -2889
rect -411 -2893 -407 -2889
rect -402 -2893 -398 -2889
rect -394 -2893 -390 -2889
rect -386 -2893 -382 -2889
rect -368 -2893 -364 -2889
rect -358 -2893 -354 -2889
rect -350 -2893 -346 -2889
rect -333 -2893 -329 -2889
rect -324 -2893 -320 -2889
rect -316 -2893 -312 -2889
rect -307 -2893 -303 -2889
rect -289 -2893 -285 -2889
rect -280 -2893 -276 -2889
rect -272 -2893 -268 -2889
rect -256 -2893 -252 -2889
rect -248 -2893 -244 -2889
rect -236 -2893 -232 -2889
rect -224 -2893 -220 -2889
rect -215 -2893 -211 -2889
rect -206 -2893 -202 -2889
rect -138 -2893 -134 -2889
rect -129 -2893 -125 -2889
rect -120 -2893 -116 -2889
rect -112 -2893 -108 -2889
rect -103 -2893 -99 -2889
rect -94 -2893 -90 -2889
rect -86 -2893 -82 -2889
rect -78 -2893 -74 -2889
rect -60 -2893 -56 -2889
rect -50 -2893 -46 -2889
rect -42 -2893 -38 -2889
rect -25 -2893 -21 -2889
rect -16 -2893 -12 -2889
rect -8 -2893 -4 -2889
rect 1 -2893 5 -2889
rect 19 -2893 23 -2889
rect 28 -2893 32 -2889
rect 36 -2893 40 -2889
rect 52 -2893 56 -2889
rect 60 -2893 64 -2889
rect 72 -2893 76 -2889
rect 84 -2893 88 -2889
rect 93 -2893 97 -2889
rect 102 -2893 106 -2889
rect 170 -2893 174 -2889
rect 179 -2893 183 -2889
rect 188 -2893 192 -2889
rect 196 -2893 200 -2889
rect 205 -2893 209 -2889
rect 214 -2893 218 -2889
rect 222 -2893 226 -2889
rect 230 -2893 234 -2889
rect 248 -2893 252 -2889
rect 258 -2893 262 -2889
rect 266 -2893 270 -2889
rect 283 -2893 287 -2889
rect 292 -2893 296 -2889
rect 300 -2893 304 -2889
rect 309 -2893 313 -2889
rect 327 -2893 331 -2889
rect 336 -2893 340 -2889
rect 344 -2893 348 -2889
rect 360 -2893 364 -2889
rect 368 -2893 372 -2889
rect 380 -2893 384 -2889
rect 392 -2893 396 -2889
rect 401 -2893 405 -2889
rect 410 -2893 414 -2889
rect 478 -2893 482 -2889
rect 487 -2893 491 -2889
rect 496 -2893 500 -2889
rect 504 -2893 508 -2889
rect 513 -2893 517 -2889
rect 522 -2893 526 -2889
rect 530 -2893 534 -2889
rect 538 -2893 542 -2889
rect 556 -2893 560 -2889
rect 566 -2893 570 -2889
rect 574 -2893 578 -2889
rect 591 -2893 595 -2889
rect 600 -2893 604 -2889
rect 608 -2893 612 -2889
rect 617 -2893 621 -2889
rect 635 -2893 639 -2889
rect 644 -2893 648 -2889
rect 652 -2893 656 -2889
rect 668 -2893 672 -2889
rect 676 -2893 680 -2889
rect 688 -2893 692 -2889
rect 700 -2893 704 -2889
rect 709 -2893 713 -2889
rect 718 -2893 722 -2889
rect 786 -2893 790 -2889
rect 795 -2893 799 -2889
rect 804 -2893 808 -2889
rect 812 -2893 816 -2889
rect 821 -2893 825 -2889
rect 830 -2893 834 -2889
rect 838 -2893 842 -2889
rect 846 -2893 850 -2889
rect 864 -2893 868 -2889
rect 874 -2893 878 -2889
rect 882 -2893 886 -2889
rect 899 -2893 903 -2889
rect 908 -2893 912 -2889
rect 916 -2893 920 -2889
rect 925 -2893 929 -2889
rect 943 -2893 947 -2889
rect 952 -2893 956 -2889
rect 960 -2893 964 -2889
rect 976 -2893 980 -2889
rect 984 -2893 988 -2889
rect 996 -2893 1000 -2889
rect 1008 -2893 1012 -2889
rect 1017 -2893 1021 -2889
rect 1026 -2893 1030 -2889
rect -1309 -3025 -1305 -3021
rect -1292 -3025 -1288 -3021
rect -1283 -3025 -1279 -3021
rect -1062 -3025 -1058 -3021
rect -1045 -3025 -1041 -3021
rect -1036 -3025 -1032 -3021
rect -754 -3025 -750 -3021
rect -737 -3025 -733 -3021
rect -728 -3025 -724 -3021
rect -446 -3025 -442 -3021
rect -429 -3025 -425 -3021
rect -420 -3025 -416 -3021
rect -138 -3025 -134 -3021
rect -121 -3025 -117 -3021
rect -112 -3025 -108 -3021
rect 170 -3025 174 -3021
rect 187 -3025 191 -3021
rect 196 -3025 200 -3021
rect 478 -3025 482 -3021
rect 495 -3025 499 -3021
rect 504 -3025 508 -3021
rect 786 -3025 790 -3021
rect 803 -3025 807 -3021
rect 812 -3025 816 -3021
rect -1234 -3184 -1230 -3180
rect -1225 -3184 -1221 -3180
rect -1216 -3184 -1212 -3180
rect -1208 -3184 -1204 -3180
rect -1199 -3184 -1195 -3180
rect -1181 -3184 -1177 -3180
rect -1172 -3184 -1168 -3180
rect -1164 -3184 -1160 -3180
rect -1147 -3184 -1143 -3180
rect -1138 -3184 -1134 -3180
rect -1062 -3184 -1058 -3180
rect -1053 -3184 -1049 -3180
rect -1044 -3184 -1040 -3180
rect -1036 -3184 -1032 -3180
rect -1027 -3184 -1023 -3180
rect -1018 -3184 -1014 -3180
rect -1010 -3184 -1006 -3180
rect -1002 -3184 -998 -3180
rect -984 -3184 -980 -3180
rect -974 -3184 -970 -3180
rect -966 -3184 -962 -3180
rect -949 -3184 -945 -3180
rect -940 -3184 -936 -3180
rect -932 -3184 -928 -3180
rect -923 -3184 -919 -3180
rect -905 -3184 -901 -3180
rect -896 -3184 -892 -3180
rect -888 -3184 -884 -3180
rect -872 -3184 -868 -3180
rect -864 -3184 -860 -3180
rect -852 -3184 -848 -3180
rect -840 -3184 -836 -3180
rect -831 -3184 -827 -3180
rect -822 -3184 -818 -3180
rect -754 -3184 -750 -3180
rect -745 -3184 -741 -3180
rect -736 -3184 -732 -3180
rect -728 -3184 -724 -3180
rect -719 -3184 -715 -3180
rect -710 -3184 -706 -3180
rect -702 -3184 -698 -3180
rect -694 -3184 -690 -3180
rect -676 -3184 -672 -3180
rect -666 -3184 -662 -3180
rect -658 -3184 -654 -3180
rect -641 -3184 -637 -3180
rect -632 -3184 -628 -3180
rect -624 -3184 -620 -3180
rect -615 -3184 -611 -3180
rect -597 -3184 -593 -3180
rect -588 -3184 -584 -3180
rect -580 -3184 -576 -3180
rect -564 -3184 -560 -3180
rect -556 -3184 -552 -3180
rect -544 -3184 -540 -3180
rect -532 -3184 -528 -3180
rect -523 -3184 -519 -3180
rect -514 -3184 -510 -3180
rect -446 -3184 -442 -3180
rect -437 -3184 -433 -3180
rect -428 -3184 -424 -3180
rect -420 -3184 -416 -3180
rect -411 -3184 -407 -3180
rect -402 -3184 -398 -3180
rect -394 -3184 -390 -3180
rect -386 -3184 -382 -3180
rect -368 -3184 -364 -3180
rect -358 -3184 -354 -3180
rect -350 -3184 -346 -3180
rect -333 -3184 -329 -3180
rect -324 -3184 -320 -3180
rect -316 -3184 -312 -3180
rect -307 -3184 -303 -3180
rect -289 -3184 -285 -3180
rect -280 -3184 -276 -3180
rect -272 -3184 -268 -3180
rect -256 -3184 -252 -3180
rect -248 -3184 -244 -3180
rect -236 -3184 -232 -3180
rect -224 -3184 -220 -3180
rect -215 -3184 -211 -3180
rect -206 -3184 -202 -3180
rect -138 -3184 -134 -3180
rect -129 -3184 -125 -3180
rect -120 -3184 -116 -3180
rect -112 -3184 -108 -3180
rect -103 -3184 -99 -3180
rect -94 -3184 -90 -3180
rect -86 -3184 -82 -3180
rect -78 -3184 -74 -3180
rect -60 -3184 -56 -3180
rect -50 -3184 -46 -3180
rect -42 -3184 -38 -3180
rect -25 -3184 -21 -3180
rect -16 -3184 -12 -3180
rect -8 -3184 -4 -3180
rect 1 -3184 5 -3180
rect 19 -3184 23 -3180
rect 28 -3184 32 -3180
rect 36 -3184 40 -3180
rect 52 -3184 56 -3180
rect 60 -3184 64 -3180
rect 72 -3184 76 -3180
rect 84 -3184 88 -3180
rect 93 -3184 97 -3180
rect 102 -3184 106 -3180
rect 170 -3184 174 -3180
rect 179 -3184 183 -3180
rect 188 -3184 192 -3180
rect 196 -3184 200 -3180
rect 205 -3184 209 -3180
rect 214 -3184 218 -3180
rect 222 -3184 226 -3180
rect 230 -3184 234 -3180
rect 248 -3184 252 -3180
rect 258 -3184 262 -3180
rect 266 -3184 270 -3180
rect 283 -3184 287 -3180
rect 292 -3184 296 -3180
rect 300 -3184 304 -3180
rect 309 -3184 313 -3180
rect 327 -3184 331 -3180
rect 336 -3184 340 -3180
rect 344 -3184 348 -3180
rect 360 -3184 364 -3180
rect 368 -3184 372 -3180
rect 380 -3184 384 -3180
rect 392 -3184 396 -3180
rect 401 -3184 405 -3180
rect 410 -3184 414 -3180
rect 478 -3184 482 -3180
rect 487 -3184 491 -3180
rect 496 -3184 500 -3180
rect 504 -3184 508 -3180
rect 513 -3184 517 -3180
rect 522 -3184 526 -3180
rect 530 -3184 534 -3180
rect 538 -3184 542 -3180
rect 556 -3184 560 -3180
rect 566 -3184 570 -3180
rect 574 -3184 578 -3180
rect 591 -3184 595 -3180
rect 600 -3184 604 -3180
rect 608 -3184 612 -3180
rect 617 -3184 621 -3180
rect 635 -3184 639 -3180
rect 644 -3184 648 -3180
rect 652 -3184 656 -3180
rect 668 -3184 672 -3180
rect 676 -3184 680 -3180
rect 688 -3184 692 -3180
rect 700 -3184 704 -3180
rect 709 -3184 713 -3180
rect 718 -3184 722 -3180
rect 786 -3184 790 -3180
rect 795 -3184 799 -3180
rect 804 -3184 808 -3180
rect 812 -3184 816 -3180
rect 821 -3184 825 -3180
rect 830 -3184 834 -3180
rect 838 -3184 842 -3180
rect 846 -3184 850 -3180
rect 864 -3184 868 -3180
rect 874 -3184 878 -3180
rect 882 -3184 886 -3180
rect 899 -3184 903 -3180
rect 908 -3184 912 -3180
rect 916 -3184 920 -3180
rect 925 -3184 929 -3180
rect 943 -3184 947 -3180
rect 952 -3184 956 -3180
rect 960 -3184 964 -3180
rect 976 -3184 980 -3180
rect 984 -3184 988 -3180
rect 996 -3184 1000 -3180
rect 1008 -3184 1012 -3180
rect 1017 -3184 1021 -3180
rect 1026 -3184 1030 -3180
<< pdcontact >>
rect -1307 -996 -1303 -988
rect -1299 -996 -1295 -988
rect -1290 -996 -1286 -988
rect -1281 -996 -1277 -988
rect -1063 -996 -1059 -988
rect -1055 -996 -1051 -988
rect -1046 -996 -1042 -988
rect -1037 -996 -1033 -988
rect -754 -996 -750 -988
rect -746 -996 -742 -988
rect -737 -996 -733 -988
rect -728 -996 -724 -988
rect -446 -996 -442 -988
rect -438 -996 -434 -988
rect -429 -996 -425 -988
rect -420 -996 -416 -988
rect -139 -996 -135 -988
rect -131 -996 -127 -988
rect -122 -996 -118 -988
rect -113 -996 -109 -988
rect 170 -996 174 -988
rect 178 -996 182 -988
rect 187 -996 191 -988
rect 196 -996 200 -988
rect 478 -996 482 -988
rect 486 -996 490 -988
rect 495 -996 499 -988
rect 504 -996 508 -988
rect 786 -996 790 -988
rect 794 -996 798 -988
rect 803 -996 807 -988
rect 812 -996 816 -988
rect -1309 -1146 -1305 -1138
rect -1301 -1146 -1297 -1138
rect -1292 -1146 -1288 -1138
rect -1283 -1146 -1279 -1138
rect -1062 -1146 -1058 -1138
rect -1054 -1146 -1050 -1138
rect -1045 -1146 -1041 -1138
rect -1036 -1146 -1032 -1138
rect -754 -1146 -750 -1138
rect -746 -1146 -742 -1138
rect -737 -1146 -733 -1138
rect -728 -1146 -724 -1138
rect -446 -1146 -442 -1138
rect -438 -1146 -434 -1138
rect -429 -1146 -425 -1138
rect -420 -1146 -416 -1138
rect -138 -1146 -134 -1138
rect -130 -1146 -126 -1138
rect -121 -1146 -117 -1138
rect -112 -1146 -108 -1138
rect 170 -1146 174 -1138
rect 178 -1146 182 -1138
rect 187 -1146 191 -1138
rect 196 -1146 200 -1138
rect 478 -1146 482 -1138
rect 486 -1146 490 -1138
rect 495 -1146 499 -1138
rect 504 -1146 508 -1138
rect 786 -1146 790 -1138
rect 794 -1146 798 -1138
rect 803 -1146 807 -1138
rect 812 -1146 816 -1138
rect -1230 -1310 -1226 -1302
rect -1221 -1310 -1217 -1302
rect -1212 -1310 -1208 -1302
rect -1204 -1310 -1200 -1302
rect -1186 -1310 -1182 -1302
rect -1164 -1310 -1160 -1302
rect -1152 -1310 -1148 -1302
rect -1143 -1310 -1139 -1302
rect -1134 -1310 -1130 -1302
rect -1062 -1310 -1058 -1302
rect -1053 -1310 -1049 -1302
rect -1044 -1310 -1040 -1302
rect -1036 -1310 -1032 -1302
rect -1027 -1310 -1023 -1302
rect -1018 -1310 -1014 -1302
rect -1010 -1310 -1006 -1302
rect -992 -1310 -988 -1302
rect -970 -1310 -966 -1302
rect -958 -1310 -954 -1302
rect -949 -1310 -945 -1302
rect -940 -1310 -936 -1302
rect -932 -1310 -928 -1302
rect -914 -1310 -910 -1302
rect -892 -1310 -888 -1302
rect -880 -1310 -876 -1302
rect -868 -1310 -864 -1302
rect -856 -1310 -852 -1302
rect -848 -1310 -844 -1302
rect -831 -1310 -827 -1302
rect -822 -1310 -818 -1302
rect -754 -1310 -750 -1302
rect -745 -1310 -741 -1302
rect -736 -1310 -732 -1302
rect -728 -1310 -724 -1302
rect -719 -1310 -715 -1302
rect -710 -1310 -706 -1302
rect -702 -1310 -698 -1302
rect -684 -1310 -680 -1302
rect -662 -1310 -658 -1302
rect -650 -1310 -646 -1302
rect -641 -1310 -637 -1302
rect -632 -1310 -628 -1302
rect -624 -1310 -620 -1302
rect -606 -1310 -602 -1302
rect -584 -1310 -580 -1302
rect -572 -1310 -568 -1302
rect -560 -1310 -556 -1302
rect -548 -1310 -544 -1302
rect -540 -1310 -536 -1302
rect -523 -1310 -519 -1302
rect -514 -1310 -510 -1302
rect -446 -1310 -442 -1302
rect -437 -1310 -433 -1302
rect -428 -1310 -424 -1302
rect -420 -1310 -416 -1302
rect -411 -1310 -407 -1302
rect -402 -1310 -398 -1302
rect -394 -1310 -390 -1302
rect -376 -1310 -372 -1302
rect -354 -1310 -350 -1302
rect -342 -1310 -338 -1302
rect -333 -1310 -329 -1302
rect -324 -1310 -320 -1302
rect -316 -1310 -312 -1302
rect -298 -1310 -294 -1302
rect -276 -1310 -272 -1302
rect -264 -1310 -260 -1302
rect -252 -1310 -248 -1302
rect -240 -1310 -236 -1302
rect -232 -1310 -228 -1302
rect -215 -1310 -211 -1302
rect -206 -1310 -202 -1302
rect -138 -1310 -134 -1302
rect -129 -1310 -125 -1302
rect -120 -1310 -116 -1302
rect -112 -1310 -108 -1302
rect -103 -1310 -99 -1302
rect -94 -1310 -90 -1302
rect -86 -1310 -82 -1302
rect -68 -1310 -64 -1302
rect -46 -1310 -42 -1302
rect -34 -1310 -30 -1302
rect -25 -1310 -21 -1302
rect -16 -1310 -12 -1302
rect -8 -1310 -4 -1302
rect 10 -1310 14 -1302
rect 32 -1310 36 -1302
rect 44 -1310 48 -1302
rect 56 -1310 60 -1302
rect 68 -1310 72 -1302
rect 76 -1310 80 -1302
rect 93 -1310 97 -1302
rect 102 -1310 106 -1302
rect 170 -1310 174 -1302
rect 179 -1310 183 -1302
rect 188 -1310 192 -1302
rect 196 -1310 200 -1302
rect 205 -1310 209 -1302
rect 214 -1310 218 -1302
rect 222 -1310 226 -1302
rect 240 -1310 244 -1302
rect 262 -1310 266 -1302
rect 274 -1310 278 -1302
rect 283 -1310 287 -1302
rect 292 -1310 296 -1302
rect 300 -1310 304 -1302
rect 318 -1310 322 -1302
rect 340 -1310 344 -1302
rect 352 -1310 356 -1302
rect 364 -1310 368 -1302
rect 376 -1310 380 -1302
rect 384 -1310 388 -1302
rect 401 -1310 405 -1302
rect 410 -1310 414 -1302
rect 478 -1310 482 -1302
rect 487 -1310 491 -1302
rect 496 -1310 500 -1302
rect 504 -1310 508 -1302
rect 513 -1310 517 -1302
rect 522 -1310 526 -1302
rect 530 -1310 534 -1302
rect 548 -1310 552 -1302
rect 570 -1310 574 -1302
rect 582 -1310 586 -1302
rect 591 -1310 595 -1302
rect 600 -1310 604 -1302
rect 608 -1310 612 -1302
rect 626 -1310 630 -1302
rect 648 -1310 652 -1302
rect 660 -1310 664 -1302
rect 672 -1310 676 -1302
rect 684 -1310 688 -1302
rect 692 -1310 696 -1302
rect 709 -1310 713 -1302
rect 718 -1310 722 -1302
rect 784 -1310 788 -1302
rect 793 -1310 797 -1302
rect 802 -1310 806 -1302
rect 810 -1310 814 -1302
rect 828 -1310 832 -1302
rect 850 -1310 854 -1302
rect 862 -1310 866 -1302
rect 871 -1310 875 -1302
rect 880 -1310 884 -1302
rect -1309 -1467 -1305 -1459
rect -1301 -1467 -1297 -1459
rect -1292 -1467 -1288 -1459
rect -1283 -1467 -1279 -1459
rect -1062 -1467 -1058 -1459
rect -1054 -1467 -1050 -1459
rect -1045 -1467 -1041 -1459
rect -1036 -1467 -1032 -1459
rect -754 -1467 -750 -1459
rect -746 -1467 -742 -1459
rect -737 -1467 -733 -1459
rect -728 -1467 -724 -1459
rect -446 -1467 -442 -1459
rect -438 -1467 -434 -1459
rect -429 -1467 -425 -1459
rect -420 -1467 -416 -1459
rect -138 -1467 -134 -1459
rect -130 -1467 -126 -1459
rect -121 -1467 -117 -1459
rect -112 -1467 -108 -1459
rect 170 -1467 174 -1459
rect 178 -1467 182 -1459
rect 187 -1467 191 -1459
rect 196 -1467 200 -1459
rect 478 -1467 482 -1459
rect 486 -1467 490 -1459
rect 495 -1467 499 -1459
rect 504 -1467 508 -1459
rect 786 -1467 790 -1459
rect 794 -1467 798 -1459
rect 803 -1467 807 -1459
rect 812 -1467 816 -1459
rect -1234 -1626 -1230 -1618
rect -1225 -1626 -1221 -1618
rect -1216 -1626 -1212 -1618
rect -1208 -1626 -1204 -1618
rect -1190 -1626 -1186 -1618
rect -1168 -1626 -1164 -1618
rect -1156 -1626 -1152 -1618
rect -1147 -1626 -1143 -1618
rect -1138 -1626 -1134 -1618
rect -1062 -1626 -1058 -1618
rect -1053 -1626 -1049 -1618
rect -1044 -1626 -1040 -1618
rect -1036 -1626 -1032 -1618
rect -1027 -1626 -1023 -1618
rect -1018 -1626 -1014 -1618
rect -1010 -1626 -1006 -1618
rect -992 -1626 -988 -1618
rect -970 -1626 -966 -1618
rect -958 -1626 -954 -1618
rect -949 -1626 -945 -1618
rect -940 -1626 -936 -1618
rect -932 -1626 -928 -1618
rect -914 -1626 -910 -1618
rect -892 -1626 -888 -1618
rect -880 -1626 -876 -1618
rect -868 -1626 -864 -1618
rect -856 -1626 -852 -1618
rect -848 -1626 -844 -1618
rect -831 -1626 -827 -1618
rect -822 -1626 -818 -1618
rect -754 -1626 -750 -1618
rect -745 -1626 -741 -1618
rect -736 -1626 -732 -1618
rect -728 -1626 -724 -1618
rect -719 -1626 -715 -1618
rect -710 -1626 -706 -1618
rect -702 -1626 -698 -1618
rect -684 -1626 -680 -1618
rect -662 -1626 -658 -1618
rect -650 -1626 -646 -1618
rect -641 -1626 -637 -1618
rect -632 -1626 -628 -1618
rect -624 -1626 -620 -1618
rect -606 -1626 -602 -1618
rect -584 -1626 -580 -1618
rect -572 -1626 -568 -1618
rect -560 -1626 -556 -1618
rect -548 -1626 -544 -1618
rect -540 -1626 -536 -1618
rect -523 -1626 -519 -1618
rect -514 -1626 -510 -1618
rect -446 -1626 -442 -1618
rect -437 -1626 -433 -1618
rect -428 -1626 -424 -1618
rect -420 -1626 -416 -1618
rect -411 -1626 -407 -1618
rect -402 -1626 -398 -1618
rect -394 -1626 -390 -1618
rect -376 -1626 -372 -1618
rect -354 -1626 -350 -1618
rect -342 -1626 -338 -1618
rect -333 -1626 -329 -1618
rect -324 -1626 -320 -1618
rect -316 -1626 -312 -1618
rect -298 -1626 -294 -1618
rect -276 -1626 -272 -1618
rect -264 -1626 -260 -1618
rect -252 -1626 -248 -1618
rect -240 -1626 -236 -1618
rect -232 -1626 -228 -1618
rect -215 -1626 -211 -1618
rect -206 -1626 -202 -1618
rect -138 -1626 -134 -1618
rect -129 -1626 -125 -1618
rect -120 -1626 -116 -1618
rect -112 -1626 -108 -1618
rect -103 -1626 -99 -1618
rect -94 -1626 -90 -1618
rect -86 -1626 -82 -1618
rect -68 -1626 -64 -1618
rect -46 -1626 -42 -1618
rect -34 -1626 -30 -1618
rect -25 -1626 -21 -1618
rect -16 -1626 -12 -1618
rect -8 -1626 -4 -1618
rect 10 -1626 14 -1618
rect 32 -1626 36 -1618
rect 44 -1626 48 -1618
rect 56 -1626 60 -1618
rect 68 -1626 72 -1618
rect 76 -1626 80 -1618
rect 93 -1626 97 -1618
rect 102 -1626 106 -1618
rect 170 -1626 174 -1618
rect 179 -1626 183 -1618
rect 188 -1626 192 -1618
rect 196 -1626 200 -1618
rect 205 -1626 209 -1618
rect 214 -1626 218 -1618
rect 222 -1626 226 -1618
rect 240 -1626 244 -1618
rect 262 -1626 266 -1618
rect 274 -1626 278 -1618
rect 283 -1626 287 -1618
rect 292 -1626 296 -1618
rect 300 -1626 304 -1618
rect 318 -1626 322 -1618
rect 340 -1626 344 -1618
rect 352 -1626 356 -1618
rect 364 -1626 368 -1618
rect 376 -1626 380 -1618
rect 384 -1626 388 -1618
rect 401 -1626 405 -1618
rect 410 -1626 414 -1618
rect 478 -1626 482 -1618
rect 487 -1626 491 -1618
rect 496 -1626 500 -1618
rect 504 -1626 508 -1618
rect 513 -1626 517 -1618
rect 522 -1626 526 -1618
rect 530 -1626 534 -1618
rect 548 -1626 552 -1618
rect 570 -1626 574 -1618
rect 582 -1626 586 -1618
rect 591 -1626 595 -1618
rect 600 -1626 604 -1618
rect 608 -1626 612 -1618
rect 626 -1626 630 -1618
rect 648 -1626 652 -1618
rect 660 -1626 664 -1618
rect 672 -1626 676 -1618
rect 684 -1626 688 -1618
rect 692 -1626 696 -1618
rect 709 -1626 713 -1618
rect 718 -1626 722 -1618
rect 786 -1626 790 -1618
rect 795 -1626 799 -1618
rect 804 -1626 808 -1618
rect 812 -1626 816 -1618
rect 821 -1626 825 -1618
rect 830 -1626 834 -1618
rect 838 -1626 842 -1618
rect 856 -1626 860 -1618
rect 878 -1626 882 -1618
rect 890 -1626 894 -1618
rect 899 -1626 903 -1618
rect 908 -1626 912 -1618
rect 916 -1626 920 -1618
rect 934 -1626 938 -1618
rect 956 -1626 960 -1618
rect 968 -1626 972 -1618
rect 980 -1626 984 -1618
rect 992 -1626 996 -1618
rect 1000 -1626 1004 -1618
rect 1017 -1626 1021 -1618
rect 1026 -1626 1030 -1618
rect -1309 -1758 -1305 -1750
rect -1301 -1758 -1297 -1750
rect -1292 -1758 -1288 -1750
rect -1283 -1758 -1279 -1750
rect -1062 -1758 -1058 -1750
rect -1054 -1758 -1050 -1750
rect -1045 -1758 -1041 -1750
rect -1036 -1758 -1032 -1750
rect -754 -1758 -750 -1750
rect -746 -1758 -742 -1750
rect -737 -1758 -733 -1750
rect -728 -1758 -724 -1750
rect -446 -1758 -442 -1750
rect -438 -1758 -434 -1750
rect -429 -1758 -425 -1750
rect -420 -1758 -416 -1750
rect -138 -1758 -134 -1750
rect -130 -1758 -126 -1750
rect -121 -1758 -117 -1750
rect -112 -1758 -108 -1750
rect 170 -1758 174 -1750
rect 178 -1758 182 -1750
rect 187 -1758 191 -1750
rect 196 -1758 200 -1750
rect 478 -1758 482 -1750
rect 486 -1758 490 -1750
rect 495 -1758 499 -1750
rect 504 -1758 508 -1750
rect 786 -1758 790 -1750
rect 794 -1758 798 -1750
rect 803 -1758 807 -1750
rect 812 -1758 816 -1750
rect -1234 -1917 -1230 -1909
rect -1225 -1917 -1221 -1909
rect -1216 -1917 -1212 -1909
rect -1208 -1917 -1204 -1909
rect -1190 -1917 -1186 -1909
rect -1168 -1917 -1164 -1909
rect -1156 -1917 -1152 -1909
rect -1147 -1917 -1143 -1909
rect -1138 -1917 -1134 -1909
rect -1062 -1917 -1058 -1909
rect -1053 -1917 -1049 -1909
rect -1044 -1917 -1040 -1909
rect -1036 -1917 -1032 -1909
rect -1027 -1917 -1023 -1909
rect -1018 -1917 -1014 -1909
rect -1010 -1917 -1006 -1909
rect -992 -1917 -988 -1909
rect -970 -1917 -966 -1909
rect -958 -1917 -954 -1909
rect -949 -1917 -945 -1909
rect -940 -1917 -936 -1909
rect -932 -1917 -928 -1909
rect -914 -1917 -910 -1909
rect -892 -1917 -888 -1909
rect -880 -1917 -876 -1909
rect -868 -1917 -864 -1909
rect -856 -1917 -852 -1909
rect -848 -1917 -844 -1909
rect -831 -1917 -827 -1909
rect -822 -1917 -818 -1909
rect -754 -1917 -750 -1909
rect -745 -1917 -741 -1909
rect -736 -1917 -732 -1909
rect -728 -1917 -724 -1909
rect -719 -1917 -715 -1909
rect -710 -1917 -706 -1909
rect -702 -1917 -698 -1909
rect -684 -1917 -680 -1909
rect -662 -1917 -658 -1909
rect -650 -1917 -646 -1909
rect -641 -1917 -637 -1909
rect -632 -1917 -628 -1909
rect -624 -1917 -620 -1909
rect -606 -1917 -602 -1909
rect -584 -1917 -580 -1909
rect -572 -1917 -568 -1909
rect -560 -1917 -556 -1909
rect -548 -1917 -544 -1909
rect -540 -1917 -536 -1909
rect -523 -1917 -519 -1909
rect -514 -1917 -510 -1909
rect -446 -1917 -442 -1909
rect -437 -1917 -433 -1909
rect -428 -1917 -424 -1909
rect -420 -1917 -416 -1909
rect -411 -1917 -407 -1909
rect -402 -1917 -398 -1909
rect -394 -1917 -390 -1909
rect -376 -1917 -372 -1909
rect -354 -1917 -350 -1909
rect -342 -1917 -338 -1909
rect -333 -1917 -329 -1909
rect -324 -1917 -320 -1909
rect -316 -1917 -312 -1909
rect -298 -1917 -294 -1909
rect -276 -1917 -272 -1909
rect -264 -1917 -260 -1909
rect -252 -1917 -248 -1909
rect -240 -1917 -236 -1909
rect -232 -1917 -228 -1909
rect -215 -1917 -211 -1909
rect -206 -1917 -202 -1909
rect -138 -1917 -134 -1909
rect -129 -1917 -125 -1909
rect -120 -1917 -116 -1909
rect -112 -1917 -108 -1909
rect -103 -1917 -99 -1909
rect -94 -1917 -90 -1909
rect -86 -1917 -82 -1909
rect -68 -1917 -64 -1909
rect -46 -1917 -42 -1909
rect -34 -1917 -30 -1909
rect -25 -1917 -21 -1909
rect -16 -1917 -12 -1909
rect -8 -1917 -4 -1909
rect 10 -1917 14 -1909
rect 32 -1917 36 -1909
rect 44 -1917 48 -1909
rect 56 -1917 60 -1909
rect 68 -1917 72 -1909
rect 76 -1917 80 -1909
rect 93 -1917 97 -1909
rect 102 -1917 106 -1909
rect 170 -1917 174 -1909
rect 179 -1917 183 -1909
rect 188 -1917 192 -1909
rect 196 -1917 200 -1909
rect 205 -1917 209 -1909
rect 214 -1917 218 -1909
rect 222 -1917 226 -1909
rect 240 -1917 244 -1909
rect 262 -1917 266 -1909
rect 274 -1917 278 -1909
rect 283 -1917 287 -1909
rect 292 -1917 296 -1909
rect 300 -1917 304 -1909
rect 318 -1917 322 -1909
rect 340 -1917 344 -1909
rect 352 -1917 356 -1909
rect 364 -1917 368 -1909
rect 376 -1917 380 -1909
rect 384 -1917 388 -1909
rect 401 -1917 405 -1909
rect 410 -1917 414 -1909
rect 478 -1917 482 -1909
rect 487 -1917 491 -1909
rect 496 -1917 500 -1909
rect 504 -1917 508 -1909
rect 513 -1917 517 -1909
rect 522 -1917 526 -1909
rect 530 -1917 534 -1909
rect 548 -1917 552 -1909
rect 570 -1917 574 -1909
rect 582 -1917 586 -1909
rect 591 -1917 595 -1909
rect 600 -1917 604 -1909
rect 608 -1917 612 -1909
rect 626 -1917 630 -1909
rect 648 -1917 652 -1909
rect 660 -1917 664 -1909
rect 672 -1917 676 -1909
rect 684 -1917 688 -1909
rect 692 -1917 696 -1909
rect 709 -1917 713 -1909
rect 718 -1917 722 -1909
rect 786 -1917 790 -1909
rect 795 -1917 799 -1909
rect 804 -1917 808 -1909
rect 812 -1917 816 -1909
rect 821 -1917 825 -1909
rect 830 -1917 834 -1909
rect 838 -1917 842 -1909
rect 856 -1917 860 -1909
rect 878 -1917 882 -1909
rect 890 -1917 894 -1909
rect 899 -1917 903 -1909
rect 908 -1917 912 -1909
rect 916 -1917 920 -1909
rect 934 -1917 938 -1909
rect 956 -1917 960 -1909
rect 968 -1917 972 -1909
rect 980 -1917 984 -1909
rect 992 -1917 996 -1909
rect 1000 -1917 1004 -1909
rect 1017 -1917 1021 -1909
rect 1026 -1917 1030 -1909
rect -1309 -2080 -1305 -2072
rect -1301 -2080 -1297 -2072
rect -1292 -2080 -1288 -2072
rect -1283 -2080 -1279 -2072
rect -1062 -2080 -1058 -2072
rect -1054 -2080 -1050 -2072
rect -1045 -2080 -1041 -2072
rect -1036 -2080 -1032 -2072
rect -754 -2080 -750 -2072
rect -746 -2080 -742 -2072
rect -737 -2080 -733 -2072
rect -728 -2080 -724 -2072
rect -446 -2080 -442 -2072
rect -438 -2080 -434 -2072
rect -429 -2080 -425 -2072
rect -420 -2080 -416 -2072
rect -138 -2080 -134 -2072
rect -130 -2080 -126 -2072
rect -121 -2080 -117 -2072
rect -112 -2080 -108 -2072
rect 170 -2080 174 -2072
rect 178 -2080 182 -2072
rect 187 -2080 191 -2072
rect 196 -2080 200 -2072
rect 478 -2080 482 -2072
rect 486 -2080 490 -2072
rect 495 -2080 499 -2072
rect 504 -2080 508 -2072
rect 786 -2080 790 -2072
rect 794 -2080 798 -2072
rect 803 -2080 807 -2072
rect 812 -2080 816 -2072
rect -1234 -2239 -1230 -2231
rect -1225 -2239 -1221 -2231
rect -1216 -2239 -1212 -2231
rect -1208 -2239 -1204 -2231
rect -1190 -2239 -1186 -2231
rect -1168 -2239 -1164 -2231
rect -1156 -2239 -1152 -2231
rect -1147 -2239 -1143 -2231
rect -1138 -2239 -1134 -2231
rect -1062 -2239 -1058 -2231
rect -1053 -2239 -1049 -2231
rect -1044 -2239 -1040 -2231
rect -1036 -2239 -1032 -2231
rect -1027 -2239 -1023 -2231
rect -1018 -2239 -1014 -2231
rect -1010 -2239 -1006 -2231
rect -992 -2239 -988 -2231
rect -970 -2239 -966 -2231
rect -958 -2239 -954 -2231
rect -949 -2239 -945 -2231
rect -940 -2239 -936 -2231
rect -932 -2239 -928 -2231
rect -914 -2239 -910 -2231
rect -892 -2239 -888 -2231
rect -880 -2239 -876 -2231
rect -868 -2239 -864 -2231
rect -856 -2239 -852 -2231
rect -848 -2239 -844 -2231
rect -831 -2239 -827 -2231
rect -822 -2239 -818 -2231
rect -754 -2239 -750 -2231
rect -745 -2239 -741 -2231
rect -736 -2239 -732 -2231
rect -728 -2239 -724 -2231
rect -719 -2239 -715 -2231
rect -710 -2239 -706 -2231
rect -702 -2239 -698 -2231
rect -684 -2239 -680 -2231
rect -662 -2239 -658 -2231
rect -650 -2239 -646 -2231
rect -641 -2239 -637 -2231
rect -632 -2239 -628 -2231
rect -624 -2239 -620 -2231
rect -606 -2239 -602 -2231
rect -584 -2239 -580 -2231
rect -572 -2239 -568 -2231
rect -560 -2239 -556 -2231
rect -548 -2239 -544 -2231
rect -540 -2239 -536 -2231
rect -523 -2239 -519 -2231
rect -514 -2239 -510 -2231
rect -446 -2239 -442 -2231
rect -437 -2239 -433 -2231
rect -428 -2239 -424 -2231
rect -420 -2239 -416 -2231
rect -411 -2239 -407 -2231
rect -402 -2239 -398 -2231
rect -394 -2239 -390 -2231
rect -376 -2239 -372 -2231
rect -354 -2239 -350 -2231
rect -342 -2239 -338 -2231
rect -333 -2239 -329 -2231
rect -324 -2239 -320 -2231
rect -316 -2239 -312 -2231
rect -298 -2239 -294 -2231
rect -276 -2239 -272 -2231
rect -264 -2239 -260 -2231
rect -252 -2239 -248 -2231
rect -240 -2239 -236 -2231
rect -232 -2239 -228 -2231
rect -215 -2239 -211 -2231
rect -206 -2239 -202 -2231
rect -138 -2239 -134 -2231
rect -129 -2239 -125 -2231
rect -120 -2239 -116 -2231
rect -112 -2239 -108 -2231
rect -103 -2239 -99 -2231
rect -94 -2239 -90 -2231
rect -86 -2239 -82 -2231
rect -68 -2239 -64 -2231
rect -46 -2239 -42 -2231
rect -34 -2239 -30 -2231
rect -25 -2239 -21 -2231
rect -16 -2239 -12 -2231
rect -8 -2239 -4 -2231
rect 10 -2239 14 -2231
rect 32 -2239 36 -2231
rect 44 -2239 48 -2231
rect 56 -2239 60 -2231
rect 68 -2239 72 -2231
rect 76 -2239 80 -2231
rect 93 -2239 97 -2231
rect 102 -2239 106 -2231
rect 170 -2239 174 -2231
rect 179 -2239 183 -2231
rect 188 -2239 192 -2231
rect 196 -2239 200 -2231
rect 205 -2239 209 -2231
rect 214 -2239 218 -2231
rect 222 -2239 226 -2231
rect 240 -2239 244 -2231
rect 262 -2239 266 -2231
rect 274 -2239 278 -2231
rect 283 -2239 287 -2231
rect 292 -2239 296 -2231
rect 300 -2239 304 -2231
rect 318 -2239 322 -2231
rect 340 -2239 344 -2231
rect 352 -2239 356 -2231
rect 364 -2239 368 -2231
rect 376 -2239 380 -2231
rect 384 -2239 388 -2231
rect 401 -2239 405 -2231
rect 410 -2239 414 -2231
rect 478 -2239 482 -2231
rect 487 -2239 491 -2231
rect 496 -2239 500 -2231
rect 504 -2239 508 -2231
rect 513 -2239 517 -2231
rect 522 -2239 526 -2231
rect 530 -2239 534 -2231
rect 548 -2239 552 -2231
rect 570 -2239 574 -2231
rect 582 -2239 586 -2231
rect 591 -2239 595 -2231
rect 600 -2239 604 -2231
rect 608 -2239 612 -2231
rect 626 -2239 630 -2231
rect 648 -2239 652 -2231
rect 660 -2239 664 -2231
rect 672 -2239 676 -2231
rect 684 -2239 688 -2231
rect 692 -2239 696 -2231
rect 709 -2239 713 -2231
rect 718 -2239 722 -2231
rect 786 -2239 790 -2231
rect 795 -2239 799 -2231
rect 804 -2239 808 -2231
rect 812 -2239 816 -2231
rect 821 -2239 825 -2231
rect 830 -2239 834 -2231
rect 838 -2239 842 -2231
rect 856 -2239 860 -2231
rect 878 -2239 882 -2231
rect 890 -2239 894 -2231
rect 899 -2239 903 -2231
rect 908 -2239 912 -2231
rect 916 -2239 920 -2231
rect 934 -2239 938 -2231
rect 956 -2239 960 -2231
rect 968 -2239 972 -2231
rect 980 -2239 984 -2231
rect 992 -2239 996 -2231
rect 1000 -2239 1004 -2231
rect 1017 -2239 1021 -2231
rect 1026 -2239 1030 -2231
rect -1309 -2371 -1305 -2363
rect -1301 -2371 -1297 -2363
rect -1292 -2371 -1288 -2363
rect -1283 -2371 -1279 -2363
rect -1062 -2371 -1058 -2363
rect -1054 -2371 -1050 -2363
rect -1045 -2371 -1041 -2363
rect -1036 -2371 -1032 -2363
rect -754 -2371 -750 -2363
rect -746 -2371 -742 -2363
rect -737 -2371 -733 -2363
rect -728 -2371 -724 -2363
rect -446 -2371 -442 -2363
rect -438 -2371 -434 -2363
rect -429 -2371 -425 -2363
rect -420 -2371 -416 -2363
rect -138 -2371 -134 -2363
rect -130 -2371 -126 -2363
rect -121 -2371 -117 -2363
rect -112 -2371 -108 -2363
rect 170 -2371 174 -2363
rect 178 -2371 182 -2363
rect 187 -2371 191 -2363
rect 196 -2371 200 -2363
rect 478 -2371 482 -2363
rect 486 -2371 490 -2363
rect 495 -2371 499 -2363
rect 504 -2371 508 -2363
rect 786 -2371 790 -2363
rect 794 -2371 798 -2363
rect 803 -2371 807 -2363
rect 812 -2371 816 -2363
rect -1234 -2530 -1230 -2522
rect -1225 -2530 -1221 -2522
rect -1216 -2530 -1212 -2522
rect -1208 -2530 -1204 -2522
rect -1190 -2530 -1186 -2522
rect -1168 -2530 -1164 -2522
rect -1156 -2530 -1152 -2522
rect -1147 -2530 -1143 -2522
rect -1138 -2530 -1134 -2522
rect -1062 -2530 -1058 -2522
rect -1053 -2530 -1049 -2522
rect -1044 -2530 -1040 -2522
rect -1036 -2530 -1032 -2522
rect -1027 -2530 -1023 -2522
rect -1018 -2530 -1014 -2522
rect -1010 -2530 -1006 -2522
rect -992 -2530 -988 -2522
rect -970 -2530 -966 -2522
rect -958 -2530 -954 -2522
rect -949 -2530 -945 -2522
rect -940 -2530 -936 -2522
rect -932 -2530 -928 -2522
rect -914 -2530 -910 -2522
rect -892 -2530 -888 -2522
rect -880 -2530 -876 -2522
rect -868 -2530 -864 -2522
rect -856 -2530 -852 -2522
rect -848 -2530 -844 -2522
rect -831 -2530 -827 -2522
rect -822 -2530 -818 -2522
rect -754 -2530 -750 -2522
rect -745 -2530 -741 -2522
rect -736 -2530 -732 -2522
rect -728 -2530 -724 -2522
rect -719 -2530 -715 -2522
rect -710 -2530 -706 -2522
rect -702 -2530 -698 -2522
rect -684 -2530 -680 -2522
rect -662 -2530 -658 -2522
rect -650 -2530 -646 -2522
rect -641 -2530 -637 -2522
rect -632 -2530 -628 -2522
rect -624 -2530 -620 -2522
rect -606 -2530 -602 -2522
rect -584 -2530 -580 -2522
rect -572 -2530 -568 -2522
rect -560 -2530 -556 -2522
rect -548 -2530 -544 -2522
rect -540 -2530 -536 -2522
rect -523 -2530 -519 -2522
rect -514 -2530 -510 -2522
rect -446 -2530 -442 -2522
rect -437 -2530 -433 -2522
rect -428 -2530 -424 -2522
rect -420 -2530 -416 -2522
rect -411 -2530 -407 -2522
rect -402 -2530 -398 -2522
rect -394 -2530 -390 -2522
rect -376 -2530 -372 -2522
rect -354 -2530 -350 -2522
rect -342 -2530 -338 -2522
rect -333 -2530 -329 -2522
rect -324 -2530 -320 -2522
rect -316 -2530 -312 -2522
rect -298 -2530 -294 -2522
rect -276 -2530 -272 -2522
rect -264 -2530 -260 -2522
rect -252 -2530 -248 -2522
rect -240 -2530 -236 -2522
rect -232 -2530 -228 -2522
rect -215 -2530 -211 -2522
rect -206 -2530 -202 -2522
rect -138 -2530 -134 -2522
rect -129 -2530 -125 -2522
rect -120 -2530 -116 -2522
rect -112 -2530 -108 -2522
rect -103 -2530 -99 -2522
rect -94 -2530 -90 -2522
rect -86 -2530 -82 -2522
rect -68 -2530 -64 -2522
rect -46 -2530 -42 -2522
rect -34 -2530 -30 -2522
rect -25 -2530 -21 -2522
rect -16 -2530 -12 -2522
rect -8 -2530 -4 -2522
rect 10 -2530 14 -2522
rect 32 -2530 36 -2522
rect 44 -2530 48 -2522
rect 56 -2530 60 -2522
rect 68 -2530 72 -2522
rect 76 -2530 80 -2522
rect 93 -2530 97 -2522
rect 102 -2530 106 -2522
rect 170 -2530 174 -2522
rect 179 -2530 183 -2522
rect 188 -2530 192 -2522
rect 196 -2530 200 -2522
rect 205 -2530 209 -2522
rect 214 -2530 218 -2522
rect 222 -2530 226 -2522
rect 240 -2530 244 -2522
rect 262 -2530 266 -2522
rect 274 -2530 278 -2522
rect 283 -2530 287 -2522
rect 292 -2530 296 -2522
rect 300 -2530 304 -2522
rect 318 -2530 322 -2522
rect 340 -2530 344 -2522
rect 352 -2530 356 -2522
rect 364 -2530 368 -2522
rect 376 -2530 380 -2522
rect 384 -2530 388 -2522
rect 401 -2530 405 -2522
rect 410 -2530 414 -2522
rect 478 -2530 482 -2522
rect 487 -2530 491 -2522
rect 496 -2530 500 -2522
rect 504 -2530 508 -2522
rect 513 -2530 517 -2522
rect 522 -2530 526 -2522
rect 530 -2530 534 -2522
rect 548 -2530 552 -2522
rect 570 -2530 574 -2522
rect 582 -2530 586 -2522
rect 591 -2530 595 -2522
rect 600 -2530 604 -2522
rect 608 -2530 612 -2522
rect 626 -2530 630 -2522
rect 648 -2530 652 -2522
rect 660 -2530 664 -2522
rect 672 -2530 676 -2522
rect 684 -2530 688 -2522
rect 692 -2530 696 -2522
rect 709 -2530 713 -2522
rect 718 -2530 722 -2522
rect 786 -2530 790 -2522
rect 795 -2530 799 -2522
rect 804 -2530 808 -2522
rect 812 -2530 816 -2522
rect 821 -2530 825 -2522
rect 830 -2530 834 -2522
rect 838 -2530 842 -2522
rect 856 -2530 860 -2522
rect 878 -2530 882 -2522
rect 890 -2530 894 -2522
rect 899 -2530 903 -2522
rect 908 -2530 912 -2522
rect 916 -2530 920 -2522
rect 934 -2530 938 -2522
rect 956 -2530 960 -2522
rect 968 -2530 972 -2522
rect 980 -2530 984 -2522
rect 992 -2530 996 -2522
rect 1000 -2530 1004 -2522
rect 1017 -2530 1021 -2522
rect 1026 -2530 1030 -2522
rect -1309 -2662 -1305 -2654
rect -1301 -2662 -1297 -2654
rect -1292 -2662 -1288 -2654
rect -1283 -2662 -1279 -2654
rect -1062 -2662 -1058 -2654
rect -1054 -2662 -1050 -2654
rect -1045 -2662 -1041 -2654
rect -1036 -2662 -1032 -2654
rect -754 -2662 -750 -2654
rect -746 -2662 -742 -2654
rect -737 -2662 -733 -2654
rect -728 -2662 -724 -2654
rect -446 -2662 -442 -2654
rect -438 -2662 -434 -2654
rect -429 -2662 -425 -2654
rect -420 -2662 -416 -2654
rect -138 -2662 -134 -2654
rect -130 -2662 -126 -2654
rect -121 -2662 -117 -2654
rect -112 -2662 -108 -2654
rect 170 -2662 174 -2654
rect 178 -2662 182 -2654
rect 187 -2662 191 -2654
rect 196 -2662 200 -2654
rect 478 -2662 482 -2654
rect 486 -2662 490 -2654
rect 495 -2662 499 -2654
rect 504 -2662 508 -2654
rect 786 -2662 790 -2654
rect 794 -2662 798 -2654
rect 803 -2662 807 -2654
rect 812 -2662 816 -2654
rect -1234 -2821 -1230 -2813
rect -1225 -2821 -1221 -2813
rect -1216 -2821 -1212 -2813
rect -1208 -2821 -1204 -2813
rect -1190 -2821 -1186 -2813
rect -1168 -2821 -1164 -2813
rect -1156 -2821 -1152 -2813
rect -1147 -2821 -1143 -2813
rect -1138 -2821 -1134 -2813
rect -1062 -2821 -1058 -2813
rect -1053 -2821 -1049 -2813
rect -1044 -2821 -1040 -2813
rect -1036 -2821 -1032 -2813
rect -1027 -2821 -1023 -2813
rect -1018 -2821 -1014 -2813
rect -1010 -2821 -1006 -2813
rect -992 -2821 -988 -2813
rect -970 -2821 -966 -2813
rect -958 -2821 -954 -2813
rect -949 -2821 -945 -2813
rect -940 -2821 -936 -2813
rect -932 -2821 -928 -2813
rect -914 -2821 -910 -2813
rect -892 -2821 -888 -2813
rect -880 -2821 -876 -2813
rect -868 -2821 -864 -2813
rect -856 -2821 -852 -2813
rect -848 -2821 -844 -2813
rect -831 -2821 -827 -2813
rect -822 -2821 -818 -2813
rect -754 -2821 -750 -2813
rect -745 -2821 -741 -2813
rect -736 -2821 -732 -2813
rect -728 -2821 -724 -2813
rect -719 -2821 -715 -2813
rect -710 -2821 -706 -2813
rect -702 -2821 -698 -2813
rect -684 -2821 -680 -2813
rect -662 -2821 -658 -2813
rect -650 -2821 -646 -2813
rect -641 -2821 -637 -2813
rect -632 -2821 -628 -2813
rect -624 -2821 -620 -2813
rect -606 -2821 -602 -2813
rect -584 -2821 -580 -2813
rect -572 -2821 -568 -2813
rect -560 -2821 -556 -2813
rect -548 -2821 -544 -2813
rect -540 -2821 -536 -2813
rect -523 -2821 -519 -2813
rect -514 -2821 -510 -2813
rect -446 -2821 -442 -2813
rect -437 -2821 -433 -2813
rect -428 -2821 -424 -2813
rect -420 -2821 -416 -2813
rect -411 -2821 -407 -2813
rect -402 -2821 -398 -2813
rect -394 -2821 -390 -2813
rect -376 -2821 -372 -2813
rect -354 -2821 -350 -2813
rect -342 -2821 -338 -2813
rect -333 -2821 -329 -2813
rect -324 -2821 -320 -2813
rect -316 -2821 -312 -2813
rect -298 -2821 -294 -2813
rect -276 -2821 -272 -2813
rect -264 -2821 -260 -2813
rect -252 -2821 -248 -2813
rect -240 -2821 -236 -2813
rect -232 -2821 -228 -2813
rect -215 -2821 -211 -2813
rect -206 -2821 -202 -2813
rect -138 -2821 -134 -2813
rect -129 -2821 -125 -2813
rect -120 -2821 -116 -2813
rect -112 -2821 -108 -2813
rect -103 -2821 -99 -2813
rect -94 -2821 -90 -2813
rect -86 -2821 -82 -2813
rect -68 -2821 -64 -2813
rect -46 -2821 -42 -2813
rect -34 -2821 -30 -2813
rect -25 -2821 -21 -2813
rect -16 -2821 -12 -2813
rect -8 -2821 -4 -2813
rect 10 -2821 14 -2813
rect 32 -2821 36 -2813
rect 44 -2821 48 -2813
rect 56 -2821 60 -2813
rect 68 -2821 72 -2813
rect 76 -2821 80 -2813
rect 93 -2821 97 -2813
rect 102 -2821 106 -2813
rect 170 -2821 174 -2813
rect 179 -2821 183 -2813
rect 188 -2821 192 -2813
rect 196 -2821 200 -2813
rect 205 -2821 209 -2813
rect 214 -2821 218 -2813
rect 222 -2821 226 -2813
rect 240 -2821 244 -2813
rect 262 -2821 266 -2813
rect 274 -2821 278 -2813
rect 283 -2821 287 -2813
rect 292 -2821 296 -2813
rect 300 -2821 304 -2813
rect 318 -2821 322 -2813
rect 340 -2821 344 -2813
rect 352 -2821 356 -2813
rect 364 -2821 368 -2813
rect 376 -2821 380 -2813
rect 384 -2821 388 -2813
rect 401 -2821 405 -2813
rect 410 -2821 414 -2813
rect 478 -2821 482 -2813
rect 487 -2821 491 -2813
rect 496 -2821 500 -2813
rect 504 -2821 508 -2813
rect 513 -2821 517 -2813
rect 522 -2821 526 -2813
rect 530 -2821 534 -2813
rect 548 -2821 552 -2813
rect 570 -2821 574 -2813
rect 582 -2821 586 -2813
rect 591 -2821 595 -2813
rect 600 -2821 604 -2813
rect 608 -2821 612 -2813
rect 626 -2821 630 -2813
rect 648 -2821 652 -2813
rect 660 -2821 664 -2813
rect 672 -2821 676 -2813
rect 684 -2821 688 -2813
rect 692 -2821 696 -2813
rect 709 -2821 713 -2813
rect 718 -2821 722 -2813
rect 786 -2821 790 -2813
rect 795 -2821 799 -2813
rect 804 -2821 808 -2813
rect 812 -2821 816 -2813
rect 821 -2821 825 -2813
rect 830 -2821 834 -2813
rect 838 -2821 842 -2813
rect 856 -2821 860 -2813
rect 878 -2821 882 -2813
rect 890 -2821 894 -2813
rect 899 -2821 903 -2813
rect 908 -2821 912 -2813
rect 916 -2821 920 -2813
rect 934 -2821 938 -2813
rect 956 -2821 960 -2813
rect 968 -2821 972 -2813
rect 980 -2821 984 -2813
rect 992 -2821 996 -2813
rect 1000 -2821 1004 -2813
rect 1017 -2821 1021 -2813
rect 1026 -2821 1030 -2813
rect -1309 -2953 -1305 -2945
rect -1301 -2953 -1297 -2945
rect -1292 -2953 -1288 -2945
rect -1283 -2953 -1279 -2945
rect -1062 -2953 -1058 -2945
rect -1054 -2953 -1050 -2945
rect -1045 -2953 -1041 -2945
rect -1036 -2953 -1032 -2945
rect -754 -2953 -750 -2945
rect -746 -2953 -742 -2945
rect -737 -2953 -733 -2945
rect -728 -2953 -724 -2945
rect -446 -2953 -442 -2945
rect -438 -2953 -434 -2945
rect -429 -2953 -425 -2945
rect -420 -2953 -416 -2945
rect -138 -2953 -134 -2945
rect -130 -2953 -126 -2945
rect -121 -2953 -117 -2945
rect -112 -2953 -108 -2945
rect 170 -2953 174 -2945
rect 178 -2953 182 -2945
rect 187 -2953 191 -2945
rect 196 -2953 200 -2945
rect 478 -2953 482 -2945
rect 486 -2953 490 -2945
rect 495 -2953 499 -2945
rect 504 -2953 508 -2945
rect 786 -2953 790 -2945
rect 794 -2953 798 -2945
rect 803 -2953 807 -2945
rect 812 -2953 816 -2945
rect -1234 -3112 -1230 -3104
rect -1225 -3112 -1221 -3104
rect -1216 -3112 -1212 -3104
rect -1208 -3112 -1204 -3104
rect -1190 -3112 -1186 -3104
rect -1168 -3112 -1164 -3104
rect -1156 -3112 -1152 -3104
rect -1147 -3112 -1143 -3104
rect -1138 -3112 -1134 -3104
rect -1062 -3112 -1058 -3104
rect -1053 -3112 -1049 -3104
rect -1044 -3112 -1040 -3104
rect -1036 -3112 -1032 -3104
rect -1027 -3112 -1023 -3104
rect -1018 -3112 -1014 -3104
rect -1010 -3112 -1006 -3104
rect -992 -3112 -988 -3104
rect -970 -3112 -966 -3104
rect -958 -3112 -954 -3104
rect -949 -3112 -945 -3104
rect -940 -3112 -936 -3104
rect -932 -3112 -928 -3104
rect -914 -3112 -910 -3104
rect -892 -3112 -888 -3104
rect -880 -3112 -876 -3104
rect -868 -3112 -864 -3104
rect -856 -3112 -852 -3104
rect -848 -3112 -844 -3104
rect -831 -3112 -827 -3104
rect -822 -3112 -818 -3104
rect -754 -3112 -750 -3104
rect -745 -3112 -741 -3104
rect -736 -3112 -732 -3104
rect -728 -3112 -724 -3104
rect -719 -3112 -715 -3104
rect -710 -3112 -706 -3104
rect -702 -3112 -698 -3104
rect -684 -3112 -680 -3104
rect -662 -3112 -658 -3104
rect -650 -3112 -646 -3104
rect -641 -3112 -637 -3104
rect -632 -3112 -628 -3104
rect -624 -3112 -620 -3104
rect -606 -3112 -602 -3104
rect -584 -3112 -580 -3104
rect -572 -3112 -568 -3104
rect -560 -3112 -556 -3104
rect -548 -3112 -544 -3104
rect -540 -3112 -536 -3104
rect -523 -3112 -519 -3104
rect -514 -3112 -510 -3104
rect -446 -3112 -442 -3104
rect -437 -3112 -433 -3104
rect -428 -3112 -424 -3104
rect -420 -3112 -416 -3104
rect -411 -3112 -407 -3104
rect -402 -3112 -398 -3104
rect -394 -3112 -390 -3104
rect -376 -3112 -372 -3104
rect -354 -3112 -350 -3104
rect -342 -3112 -338 -3104
rect -333 -3112 -329 -3104
rect -324 -3112 -320 -3104
rect -316 -3112 -312 -3104
rect -298 -3112 -294 -3104
rect -276 -3112 -272 -3104
rect -264 -3112 -260 -3104
rect -252 -3112 -248 -3104
rect -240 -3112 -236 -3104
rect -232 -3112 -228 -3104
rect -215 -3112 -211 -3104
rect -206 -3112 -202 -3104
rect -138 -3112 -134 -3104
rect -129 -3112 -125 -3104
rect -120 -3112 -116 -3104
rect -112 -3112 -108 -3104
rect -103 -3112 -99 -3104
rect -94 -3112 -90 -3104
rect -86 -3112 -82 -3104
rect -68 -3112 -64 -3104
rect -46 -3112 -42 -3104
rect -34 -3112 -30 -3104
rect -25 -3112 -21 -3104
rect -16 -3112 -12 -3104
rect -8 -3112 -4 -3104
rect 10 -3112 14 -3104
rect 32 -3112 36 -3104
rect 44 -3112 48 -3104
rect 56 -3112 60 -3104
rect 68 -3112 72 -3104
rect 76 -3112 80 -3104
rect 93 -3112 97 -3104
rect 102 -3112 106 -3104
rect 170 -3112 174 -3104
rect 179 -3112 183 -3104
rect 188 -3112 192 -3104
rect 196 -3112 200 -3104
rect 205 -3112 209 -3104
rect 214 -3112 218 -3104
rect 222 -3112 226 -3104
rect 240 -3112 244 -3104
rect 262 -3112 266 -3104
rect 274 -3112 278 -3104
rect 283 -3112 287 -3104
rect 292 -3112 296 -3104
rect 300 -3112 304 -3104
rect 318 -3112 322 -3104
rect 340 -3112 344 -3104
rect 352 -3112 356 -3104
rect 364 -3112 368 -3104
rect 376 -3112 380 -3104
rect 384 -3112 388 -3104
rect 401 -3112 405 -3104
rect 410 -3112 414 -3104
rect 478 -3112 482 -3104
rect 487 -3112 491 -3104
rect 496 -3112 500 -3104
rect 504 -3112 508 -3104
rect 513 -3112 517 -3104
rect 522 -3112 526 -3104
rect 530 -3112 534 -3104
rect 548 -3112 552 -3104
rect 570 -3112 574 -3104
rect 582 -3112 586 -3104
rect 591 -3112 595 -3104
rect 600 -3112 604 -3104
rect 608 -3112 612 -3104
rect 626 -3112 630 -3104
rect 648 -3112 652 -3104
rect 660 -3112 664 -3104
rect 672 -3112 676 -3104
rect 684 -3112 688 -3104
rect 692 -3112 696 -3104
rect 709 -3112 713 -3104
rect 718 -3112 722 -3104
rect 786 -3112 790 -3104
rect 795 -3112 799 -3104
rect 804 -3112 808 -3104
rect 812 -3112 816 -3104
rect 821 -3112 825 -3104
rect 830 -3112 834 -3104
rect 838 -3112 842 -3104
rect 856 -3112 860 -3104
rect 878 -3112 882 -3104
rect 890 -3112 894 -3104
rect 899 -3112 903 -3104
rect 908 -3112 912 -3104
rect 916 -3112 920 -3104
rect 934 -3112 938 -3104
rect 956 -3112 960 -3104
rect 968 -3112 972 -3104
rect 980 -3112 984 -3104
rect 992 -3112 996 -3104
rect 1000 -3112 1004 -3104
rect 1017 -3112 1021 -3104
rect 1026 -3112 1030 -3104
<< m2contact >>
rect -1307 -984 -1303 -980
rect -1290 -984 -1286 -980
rect -1063 -984 -1059 -980
rect -1046 -984 -1042 -980
rect -1091 -1032 -1087 -1028
rect -1251 -1040 -1247 -1036
rect -1290 -1076 -1286 -1072
rect -1309 -1134 -1305 -1130
rect -1292 -1134 -1288 -1130
rect -1292 -1226 -1288 -1222
rect -1103 -1187 -1099 -1183
rect -1221 -1298 -1217 -1294
rect -1204 -1298 -1200 -1294
rect -1164 -1298 -1160 -1294
rect -1143 -1298 -1139 -1294
rect -1251 -1354 -1247 -1350
rect -1230 -1347 -1226 -1343
rect -1283 -1361 -1279 -1357
rect -1186 -1368 -1182 -1364
rect -1134 -1346 -1130 -1342
rect -1204 -1375 -1200 -1371
rect -1168 -1375 -1164 -1371
rect -1091 -1338 -1087 -1334
rect -754 -984 -750 -980
rect -737 -984 -733 -980
rect -1037 -1040 -1033 -1036
rect -782 -1040 -778 -1036
rect -1046 -1076 -1042 -1072
rect -1062 -1134 -1058 -1130
rect -1045 -1134 -1041 -1130
rect -1103 -1353 -1099 -1349
rect -1221 -1390 -1217 -1386
rect -1177 -1390 -1173 -1386
rect -1143 -1390 -1139 -1386
rect -1257 -1397 -1253 -1393
rect -1309 -1455 -1305 -1451
rect -1292 -1455 -1288 -1451
rect -1292 -1547 -1288 -1543
rect -1113 -1404 -1109 -1400
rect -1225 -1614 -1221 -1610
rect -1208 -1614 -1204 -1610
rect -1168 -1614 -1164 -1610
rect -1147 -1614 -1143 -1610
rect -1257 -1670 -1253 -1666
rect -1234 -1663 -1230 -1659
rect -1283 -1677 -1279 -1673
rect -1190 -1684 -1186 -1680
rect -1036 -1187 -1032 -1183
rect -795 -1187 -791 -1183
rect -1045 -1226 -1041 -1222
rect -1053 -1298 -1049 -1294
rect -1027 -1298 -1023 -1294
rect -1010 -1298 -1006 -1294
rect -970 -1298 -966 -1294
rect -949 -1298 -945 -1294
rect -932 -1298 -928 -1294
rect -892 -1298 -888 -1294
rect -868 -1298 -864 -1294
rect -831 -1298 -827 -1294
rect -1062 -1331 -1058 -1327
rect -1044 -1324 -1040 -1320
rect -1018 -1346 -1014 -1342
rect -1036 -1353 -1032 -1349
rect -992 -1338 -988 -1334
rect -940 -1331 -936 -1327
rect -1010 -1375 -1006 -1371
rect -974 -1375 -970 -1371
rect -914 -1346 -910 -1342
rect -932 -1375 -928 -1371
rect -896 -1375 -892 -1371
rect -822 -1338 -818 -1334
rect -815 -1346 -811 -1342
rect -1053 -1390 -1049 -1386
rect -1027 -1390 -1023 -1386
rect -984 -1390 -980 -1386
rect -949 -1390 -945 -1386
rect -905 -1390 -901 -1386
rect -888 -1390 -884 -1386
rect -852 -1390 -848 -1386
rect -831 -1390 -827 -1386
rect -782 -1338 -778 -1334
rect -446 -984 -442 -980
rect -429 -984 -425 -980
rect -728 -1032 -724 -1028
rect -471 -1032 -467 -1028
rect -737 -1076 -733 -1072
rect -754 -1134 -750 -1130
rect -737 -1134 -733 -1130
rect -795 -1353 -791 -1349
rect -815 -1397 -811 -1393
rect -782 -1411 -778 -1407
rect -1062 -1455 -1058 -1451
rect -1045 -1455 -1041 -1451
rect -1113 -1654 -1109 -1650
rect -1095 -1508 -1091 -1504
rect -1138 -1662 -1134 -1658
rect -1208 -1691 -1204 -1687
rect -1172 -1691 -1168 -1687
rect -1095 -1669 -1091 -1665
rect -1225 -1706 -1221 -1702
rect -1181 -1706 -1177 -1702
rect -1147 -1706 -1143 -1702
rect -1257 -1713 -1253 -1709
rect -1309 -1746 -1305 -1742
rect -1292 -1746 -1288 -1742
rect -1292 -1838 -1288 -1834
rect -1090 -1720 -1086 -1716
rect -1106 -1799 -1102 -1795
rect -1225 -1905 -1221 -1901
rect -1208 -1905 -1204 -1901
rect -1168 -1905 -1164 -1901
rect -1147 -1905 -1143 -1901
rect -1257 -1961 -1253 -1957
rect -1234 -1954 -1230 -1950
rect -1283 -1968 -1279 -1964
rect -1190 -1975 -1186 -1971
rect -1106 -1945 -1102 -1941
rect -1138 -1953 -1134 -1949
rect -1208 -1982 -1204 -1978
rect -1172 -1982 -1168 -1978
rect -1090 -1960 -1086 -1956
rect -1036 -1508 -1032 -1504
rect -795 -1508 -791 -1504
rect -1045 -1547 -1041 -1543
rect -1053 -1614 -1049 -1610
rect -1027 -1614 -1023 -1610
rect -1010 -1614 -1006 -1610
rect -970 -1614 -966 -1610
rect -949 -1614 -945 -1610
rect -932 -1614 -928 -1610
rect -892 -1614 -888 -1610
rect -868 -1614 -864 -1610
rect -831 -1614 -827 -1610
rect -1062 -1647 -1058 -1643
rect -1044 -1640 -1040 -1636
rect -1018 -1662 -1014 -1658
rect -1036 -1669 -1032 -1665
rect -992 -1654 -988 -1650
rect -940 -1647 -936 -1643
rect -1010 -1691 -1006 -1687
rect -974 -1691 -970 -1687
rect -914 -1662 -910 -1658
rect -932 -1691 -928 -1687
rect -896 -1691 -892 -1687
rect -822 -1654 -818 -1650
rect -814 -1662 -810 -1658
rect -1053 -1706 -1049 -1702
rect -1027 -1706 -1023 -1702
rect -984 -1706 -980 -1702
rect -949 -1706 -945 -1702
rect -905 -1706 -901 -1702
rect -888 -1706 -884 -1702
rect -852 -1706 -848 -1702
rect -831 -1706 -827 -1702
rect -782 -1654 -778 -1650
rect -728 -1187 -724 -1183
rect -494 -1187 -490 -1183
rect -737 -1226 -733 -1222
rect -745 -1298 -741 -1294
rect -719 -1298 -715 -1294
rect -702 -1298 -698 -1294
rect -662 -1298 -658 -1294
rect -641 -1298 -637 -1294
rect -624 -1298 -620 -1294
rect -584 -1298 -580 -1294
rect -560 -1298 -556 -1294
rect -523 -1298 -519 -1294
rect -754 -1331 -750 -1327
rect -736 -1324 -732 -1320
rect -710 -1346 -706 -1342
rect -728 -1353 -724 -1349
rect -684 -1338 -680 -1334
rect -632 -1331 -628 -1327
rect -702 -1375 -698 -1371
rect -666 -1375 -662 -1371
rect -606 -1346 -602 -1342
rect -624 -1375 -620 -1371
rect -588 -1375 -584 -1371
rect -514 -1338 -510 -1334
rect -505 -1346 -501 -1342
rect -745 -1390 -741 -1386
rect -719 -1390 -715 -1386
rect -676 -1390 -672 -1386
rect -641 -1390 -637 -1386
rect -597 -1390 -593 -1386
rect -580 -1390 -576 -1386
rect -544 -1390 -540 -1386
rect -523 -1390 -519 -1386
rect -471 -1338 -467 -1334
rect -139 -984 -135 -980
rect -122 -984 -118 -980
rect -420 -1040 -416 -1036
rect -170 -1040 -166 -1036
rect -429 -1076 -425 -1072
rect -446 -1134 -442 -1130
rect -429 -1134 -425 -1130
rect -494 -1353 -490 -1349
rect -505 -1404 -501 -1400
rect -471 -1404 -467 -1400
rect -754 -1455 -750 -1451
rect -737 -1455 -733 -1451
rect -795 -1669 -791 -1665
rect -814 -1713 -810 -1709
rect -780 -1713 -776 -1709
rect -1062 -1746 -1058 -1742
rect -1045 -1746 -1041 -1742
rect -1225 -1997 -1221 -1993
rect -1181 -1997 -1177 -1993
rect -1147 -1997 -1143 -1993
rect -1257 -2004 -1253 -2000
rect -1309 -2068 -1305 -2064
rect -1292 -2068 -1288 -2064
rect -1292 -2160 -1288 -2156
rect -1090 -2011 -1086 -2007
rect -1106 -2121 -1102 -2117
rect -1225 -2227 -1221 -2223
rect -1208 -2227 -1204 -2223
rect -1168 -2227 -1164 -2223
rect -1147 -2227 -1143 -2223
rect -1257 -2283 -1253 -2279
rect -1234 -2276 -1230 -2272
rect -1283 -2290 -1279 -2286
rect -1190 -2297 -1186 -2293
rect -1106 -2267 -1102 -2263
rect -1138 -2275 -1134 -2271
rect -1208 -2304 -1204 -2300
rect -1172 -2304 -1168 -2300
rect -1090 -2282 -1086 -2278
rect -1036 -1799 -1032 -1795
rect -793 -1799 -789 -1795
rect -1045 -1838 -1041 -1834
rect -1053 -1905 -1049 -1901
rect -1027 -1905 -1023 -1901
rect -1010 -1905 -1006 -1901
rect -970 -1905 -966 -1901
rect -949 -1905 -945 -1901
rect -932 -1905 -928 -1901
rect -892 -1905 -888 -1901
rect -868 -1905 -864 -1901
rect -831 -1905 -827 -1901
rect -1062 -1938 -1058 -1934
rect -1044 -1931 -1040 -1927
rect -1018 -1953 -1014 -1949
rect -1036 -1960 -1032 -1956
rect -992 -1945 -988 -1941
rect -940 -1938 -936 -1934
rect -1010 -1982 -1006 -1978
rect -974 -1982 -970 -1978
rect -914 -1953 -910 -1949
rect -932 -1982 -928 -1978
rect -896 -1982 -892 -1978
rect -822 -1945 -818 -1941
rect -815 -1953 -811 -1949
rect -1053 -1997 -1049 -1993
rect -1027 -1997 -1023 -1993
rect -984 -1997 -980 -1993
rect -949 -1997 -945 -1993
rect -905 -1997 -901 -1993
rect -888 -1997 -884 -1993
rect -852 -1997 -848 -1993
rect -831 -1997 -827 -1993
rect -780 -1945 -776 -1941
rect -728 -1508 -724 -1504
rect -489 -1508 -485 -1504
rect -737 -1547 -733 -1543
rect -745 -1614 -741 -1610
rect -719 -1614 -715 -1610
rect -702 -1614 -698 -1610
rect -662 -1614 -658 -1610
rect -641 -1614 -637 -1610
rect -624 -1614 -620 -1610
rect -584 -1614 -580 -1610
rect -560 -1614 -556 -1610
rect -523 -1614 -519 -1610
rect -754 -1647 -750 -1643
rect -736 -1640 -732 -1636
rect -710 -1662 -706 -1658
rect -728 -1669 -724 -1665
rect -684 -1654 -680 -1650
rect -632 -1647 -628 -1643
rect -702 -1691 -698 -1687
rect -666 -1691 -662 -1687
rect -606 -1662 -602 -1658
rect -624 -1691 -620 -1687
rect -588 -1691 -584 -1687
rect -514 -1651 -510 -1647
rect -505 -1662 -501 -1658
rect -745 -1706 -741 -1702
rect -719 -1706 -715 -1702
rect -676 -1706 -672 -1702
rect -641 -1706 -637 -1702
rect -597 -1706 -593 -1702
rect -580 -1706 -576 -1702
rect -544 -1706 -540 -1702
rect -523 -1706 -519 -1702
rect -471 -1654 -467 -1650
rect -420 -1187 -416 -1183
rect -186 -1187 -182 -1183
rect -429 -1226 -425 -1222
rect -437 -1298 -433 -1294
rect -411 -1298 -407 -1294
rect -394 -1298 -390 -1294
rect -354 -1298 -350 -1294
rect -333 -1298 -329 -1294
rect -316 -1298 -312 -1294
rect -276 -1298 -272 -1294
rect -252 -1298 -248 -1294
rect -215 -1298 -211 -1294
rect -446 -1331 -442 -1327
rect -428 -1324 -424 -1320
rect -402 -1346 -398 -1342
rect -420 -1353 -416 -1349
rect -376 -1338 -372 -1334
rect -324 -1331 -320 -1327
rect -394 -1375 -390 -1371
rect -358 -1375 -354 -1371
rect -298 -1346 -294 -1342
rect -316 -1375 -312 -1371
rect -280 -1375 -276 -1371
rect -206 -1338 -202 -1334
rect -198 -1346 -194 -1342
rect -437 -1390 -433 -1386
rect -411 -1390 -407 -1386
rect -368 -1390 -364 -1386
rect -333 -1390 -329 -1386
rect -289 -1390 -285 -1386
rect -272 -1390 -268 -1386
rect -236 -1390 -232 -1386
rect -215 -1390 -211 -1386
rect -170 -1338 -166 -1334
rect 170 -984 174 -980
rect 187 -984 191 -980
rect -113 -1032 -109 -1028
rect 145 -1032 149 -1028
rect -122 -1076 -118 -1072
rect -138 -1134 -134 -1130
rect -121 -1134 -117 -1130
rect -186 -1353 -182 -1349
rect -198 -1411 -194 -1407
rect -170 -1411 -166 -1407
rect -446 -1455 -442 -1451
rect -429 -1455 -425 -1451
rect -489 -1669 -485 -1665
rect -505 -1720 -501 -1716
rect -476 -1720 -472 -1716
rect -754 -1746 -750 -1742
rect -737 -1746 -733 -1742
rect -793 -1960 -789 -1956
rect -815 -2004 -811 -2000
rect -780 -2004 -776 -2000
rect -1062 -2068 -1058 -2064
rect -1045 -2068 -1041 -2064
rect -1225 -2319 -1221 -2315
rect -1181 -2319 -1177 -2315
rect -1147 -2319 -1143 -2315
rect -1257 -2326 -1253 -2322
rect -1309 -2359 -1305 -2355
rect -1292 -2359 -1288 -2355
rect -1292 -2451 -1288 -2447
rect -1090 -2333 -1086 -2329
rect -1106 -2412 -1102 -2408
rect -1225 -2518 -1221 -2514
rect -1208 -2518 -1204 -2514
rect -1168 -2518 -1164 -2514
rect -1147 -2518 -1143 -2514
rect -1257 -2574 -1253 -2570
rect -1234 -2567 -1230 -2563
rect -1283 -2581 -1279 -2577
rect -1190 -2588 -1186 -2584
rect -1106 -2558 -1102 -2554
rect -1138 -2566 -1134 -2562
rect -1208 -2595 -1204 -2591
rect -1172 -2595 -1168 -2591
rect -1090 -2573 -1086 -2569
rect -1036 -2121 -1032 -2117
rect -793 -2121 -789 -2117
rect -1045 -2160 -1041 -2156
rect -1053 -2227 -1049 -2223
rect -1027 -2227 -1023 -2223
rect -1010 -2227 -1006 -2223
rect -970 -2227 -966 -2223
rect -949 -2227 -945 -2223
rect -932 -2227 -928 -2223
rect -892 -2227 -888 -2223
rect -868 -2227 -864 -2223
rect -831 -2227 -827 -2223
rect -1062 -2260 -1058 -2256
rect -1044 -2253 -1040 -2249
rect -1018 -2275 -1014 -2271
rect -1036 -2282 -1032 -2278
rect -992 -2267 -988 -2263
rect -940 -2260 -936 -2256
rect -1010 -2304 -1006 -2300
rect -974 -2304 -970 -2300
rect -914 -2275 -910 -2271
rect -932 -2304 -928 -2300
rect -896 -2304 -892 -2300
rect -822 -2267 -818 -2263
rect -814 -2275 -810 -2271
rect -1053 -2319 -1049 -2315
rect -1027 -2319 -1023 -2315
rect -984 -2319 -980 -2315
rect -949 -2319 -945 -2315
rect -905 -2319 -901 -2315
rect -888 -2319 -884 -2315
rect -852 -2319 -848 -2315
rect -831 -2319 -827 -2315
rect -780 -2267 -776 -2263
rect -728 -1799 -724 -1795
rect -490 -1799 -486 -1795
rect -737 -1838 -733 -1834
rect -745 -1905 -741 -1901
rect -719 -1905 -715 -1901
rect -702 -1905 -698 -1901
rect -662 -1905 -658 -1901
rect -641 -1905 -637 -1901
rect -624 -1905 -620 -1901
rect -584 -1905 -580 -1901
rect -560 -1905 -556 -1901
rect -523 -1905 -519 -1901
rect -754 -1938 -750 -1934
rect -736 -1931 -732 -1927
rect -710 -1953 -706 -1949
rect -728 -1960 -724 -1956
rect -684 -1945 -680 -1941
rect -632 -1938 -628 -1934
rect -702 -1982 -698 -1978
rect -666 -1982 -662 -1978
rect -606 -1953 -602 -1949
rect -624 -1982 -620 -1978
rect -588 -1982 -584 -1978
rect -514 -1944 -510 -1940
rect -506 -1953 -502 -1949
rect -745 -1997 -741 -1993
rect -719 -1997 -715 -1993
rect -676 -1997 -672 -1993
rect -641 -1997 -637 -1993
rect -597 -1997 -593 -1993
rect -580 -1997 -576 -1993
rect -544 -1997 -540 -1993
rect -523 -1997 -519 -1993
rect -476 -1945 -472 -1941
rect -420 -1508 -416 -1504
rect -184 -1508 -180 -1504
rect -429 -1547 -425 -1543
rect -437 -1614 -433 -1610
rect -411 -1614 -407 -1610
rect -394 -1614 -390 -1610
rect -354 -1614 -350 -1610
rect -333 -1614 -329 -1610
rect -316 -1614 -312 -1610
rect -276 -1614 -272 -1610
rect -252 -1614 -248 -1610
rect -215 -1614 -211 -1610
rect -446 -1647 -442 -1643
rect -428 -1640 -424 -1636
rect -402 -1662 -398 -1658
rect -420 -1669 -416 -1665
rect -376 -1654 -372 -1650
rect -324 -1647 -320 -1643
rect -394 -1691 -390 -1687
rect -358 -1691 -354 -1687
rect -298 -1662 -294 -1658
rect -316 -1691 -312 -1687
rect -280 -1691 -276 -1687
rect -206 -1654 -202 -1650
rect -198 -1662 -194 -1658
rect -437 -1706 -433 -1702
rect -411 -1706 -407 -1702
rect -368 -1706 -364 -1702
rect -333 -1706 -329 -1702
rect -289 -1706 -285 -1702
rect -272 -1706 -268 -1702
rect -236 -1706 -232 -1702
rect -215 -1706 -211 -1702
rect -170 -1654 -166 -1650
rect -112 -1187 -108 -1183
rect 122 -1187 126 -1183
rect -121 -1226 -117 -1222
rect -129 -1298 -125 -1294
rect -103 -1298 -99 -1294
rect -86 -1298 -82 -1294
rect -46 -1298 -42 -1294
rect -25 -1298 -21 -1294
rect -8 -1298 -4 -1294
rect 32 -1298 36 -1294
rect 56 -1298 60 -1294
rect 93 -1298 97 -1294
rect -138 -1331 -134 -1327
rect -120 -1324 -116 -1320
rect -94 -1346 -90 -1342
rect -112 -1353 -108 -1349
rect -68 -1338 -64 -1334
rect -16 -1331 -12 -1327
rect -86 -1375 -82 -1371
rect -50 -1375 -46 -1371
rect 10 -1346 14 -1342
rect -8 -1375 -4 -1371
rect 28 -1375 32 -1371
rect 102 -1338 106 -1334
rect 109 -1346 113 -1342
rect -129 -1390 -125 -1386
rect -103 -1390 -99 -1386
rect -60 -1390 -56 -1386
rect -25 -1390 -21 -1386
rect 19 -1390 23 -1386
rect 36 -1390 40 -1386
rect 72 -1390 76 -1386
rect 93 -1390 97 -1386
rect 145 -1338 149 -1334
rect 478 -984 482 -980
rect 495 -984 499 -980
rect 196 -1040 200 -1036
rect 446 -1040 450 -1036
rect 187 -1076 191 -1072
rect 170 -1134 174 -1130
rect 187 -1134 191 -1130
rect 122 -1353 126 -1349
rect 109 -1404 113 -1400
rect 145 -1404 149 -1400
rect -138 -1455 -134 -1451
rect -121 -1455 -117 -1451
rect -184 -1669 -180 -1665
rect -198 -1713 -194 -1709
rect -166 -1713 -162 -1709
rect -446 -1746 -442 -1742
rect -429 -1746 -425 -1742
rect -490 -1960 -486 -1956
rect -506 -2011 -502 -2007
rect -476 -2011 -472 -2007
rect -754 -2068 -750 -2064
rect -737 -2068 -733 -2064
rect -793 -2282 -789 -2278
rect -814 -2326 -810 -2322
rect -780 -2326 -776 -2322
rect -1062 -2359 -1058 -2355
rect -1045 -2359 -1041 -2355
rect -1225 -2610 -1221 -2606
rect -1181 -2610 -1177 -2606
rect -1147 -2610 -1143 -2606
rect -1257 -2617 -1253 -2613
rect -1309 -2650 -1305 -2646
rect -1292 -2650 -1288 -2646
rect -1292 -2742 -1288 -2738
rect -1090 -2624 -1086 -2620
rect -1106 -2703 -1102 -2699
rect -1225 -2809 -1221 -2805
rect -1208 -2809 -1204 -2805
rect -1168 -2809 -1164 -2805
rect -1147 -2809 -1143 -2805
rect -1257 -2865 -1253 -2861
rect -1234 -2858 -1230 -2854
rect -1283 -2872 -1279 -2868
rect -1190 -2879 -1186 -2875
rect -1106 -2849 -1102 -2845
rect -1138 -2857 -1134 -2853
rect -1208 -2886 -1204 -2882
rect -1172 -2886 -1168 -2882
rect -1090 -2864 -1086 -2860
rect -1036 -2412 -1032 -2408
rect -793 -2412 -789 -2408
rect -1045 -2451 -1041 -2447
rect -1053 -2518 -1049 -2514
rect -1027 -2518 -1023 -2514
rect -1010 -2518 -1006 -2514
rect -970 -2518 -966 -2514
rect -949 -2518 -945 -2514
rect -932 -2518 -928 -2514
rect -892 -2518 -888 -2514
rect -868 -2518 -864 -2514
rect -831 -2518 -827 -2514
rect -1062 -2551 -1058 -2547
rect -1044 -2544 -1040 -2540
rect -1018 -2566 -1014 -2562
rect -1036 -2573 -1032 -2569
rect -992 -2558 -988 -2554
rect -940 -2551 -936 -2547
rect -1010 -2595 -1006 -2591
rect -974 -2595 -970 -2591
rect -914 -2566 -910 -2562
rect -932 -2595 -928 -2591
rect -896 -2595 -892 -2591
rect -822 -2558 -818 -2554
rect -814 -2566 -810 -2562
rect -1053 -2610 -1049 -2606
rect -1027 -2610 -1023 -2606
rect -984 -2610 -980 -2606
rect -949 -2610 -945 -2606
rect -905 -2610 -901 -2606
rect -888 -2610 -884 -2606
rect -852 -2610 -848 -2606
rect -831 -2610 -827 -2606
rect -780 -2558 -776 -2554
rect -728 -2121 -724 -2117
rect -490 -2121 -486 -2117
rect -737 -2160 -733 -2156
rect -745 -2227 -741 -2223
rect -719 -2227 -715 -2223
rect -702 -2227 -698 -2223
rect -662 -2227 -658 -2223
rect -641 -2227 -637 -2223
rect -624 -2227 -620 -2223
rect -584 -2227 -580 -2223
rect -560 -2227 -556 -2223
rect -523 -2227 -519 -2223
rect -754 -2260 -750 -2256
rect -736 -2253 -732 -2249
rect -710 -2275 -706 -2271
rect -728 -2282 -724 -2278
rect -684 -2267 -680 -2263
rect -632 -2260 -628 -2256
rect -702 -2304 -698 -2300
rect -666 -2304 -662 -2300
rect -606 -2275 -602 -2271
rect -624 -2304 -620 -2300
rect -588 -2304 -584 -2300
rect -514 -2266 -510 -2262
rect -505 -2275 -501 -2271
rect -745 -2319 -741 -2315
rect -719 -2319 -715 -2315
rect -676 -2319 -672 -2315
rect -641 -2319 -637 -2315
rect -597 -2319 -593 -2315
rect -580 -2319 -576 -2315
rect -544 -2319 -540 -2315
rect -523 -2319 -519 -2315
rect -476 -2267 -472 -2263
rect -420 -1799 -416 -1795
rect -180 -1799 -176 -1795
rect -429 -1838 -425 -1834
rect -437 -1905 -433 -1901
rect -411 -1905 -407 -1901
rect -394 -1905 -390 -1901
rect -354 -1905 -350 -1901
rect -333 -1905 -329 -1901
rect -316 -1905 -312 -1901
rect -276 -1905 -272 -1901
rect -252 -1905 -248 -1901
rect -215 -1905 -211 -1901
rect -446 -1938 -442 -1934
rect -428 -1931 -424 -1927
rect -402 -1953 -398 -1949
rect -420 -1960 -416 -1956
rect -376 -1945 -372 -1941
rect -324 -1938 -320 -1934
rect -394 -1982 -390 -1978
rect -358 -1982 -354 -1978
rect -298 -1953 -294 -1949
rect -316 -1982 -312 -1978
rect -280 -1982 -276 -1978
rect -206 -1945 -202 -1941
rect -199 -1953 -195 -1949
rect -437 -1997 -433 -1993
rect -411 -1997 -407 -1993
rect -368 -1997 -364 -1993
rect -333 -1997 -329 -1993
rect -289 -1997 -285 -1993
rect -272 -1997 -268 -1993
rect -236 -1997 -232 -1993
rect -215 -1997 -211 -1993
rect -166 -1945 -162 -1941
rect -112 -1508 -108 -1504
rect 126 -1508 130 -1504
rect -121 -1547 -117 -1543
rect -129 -1614 -125 -1610
rect -103 -1614 -99 -1610
rect -86 -1614 -82 -1610
rect -46 -1614 -42 -1610
rect -25 -1614 -21 -1610
rect -8 -1614 -4 -1610
rect 32 -1614 36 -1610
rect 56 -1614 60 -1610
rect 93 -1614 97 -1610
rect -138 -1647 -134 -1643
rect -120 -1640 -116 -1636
rect -94 -1662 -90 -1658
rect -112 -1669 -108 -1665
rect -68 -1654 -64 -1650
rect -16 -1647 -12 -1643
rect -86 -1691 -82 -1687
rect -50 -1691 -46 -1687
rect 10 -1662 14 -1658
rect -8 -1691 -4 -1687
rect 28 -1691 32 -1687
rect 102 -1654 106 -1650
rect 111 -1662 115 -1658
rect -129 -1706 -125 -1702
rect -103 -1706 -99 -1702
rect -60 -1706 -56 -1702
rect -25 -1706 -21 -1702
rect 19 -1706 23 -1702
rect 36 -1706 40 -1702
rect 72 -1706 76 -1702
rect 93 -1706 97 -1702
rect 145 -1654 149 -1650
rect 196 -1187 200 -1183
rect 430 -1187 434 -1183
rect 187 -1226 191 -1222
rect 179 -1298 183 -1294
rect 205 -1298 209 -1294
rect 222 -1298 226 -1294
rect 262 -1298 266 -1294
rect 283 -1298 287 -1294
rect 300 -1298 304 -1294
rect 340 -1298 344 -1294
rect 364 -1298 368 -1294
rect 401 -1298 405 -1294
rect 170 -1331 174 -1327
rect 188 -1324 192 -1320
rect 214 -1346 218 -1342
rect 196 -1353 200 -1349
rect 240 -1338 244 -1334
rect 292 -1331 296 -1327
rect 222 -1375 226 -1371
rect 258 -1375 262 -1371
rect 318 -1346 322 -1342
rect 300 -1375 304 -1371
rect 336 -1375 340 -1371
rect 410 -1338 414 -1334
rect 417 -1346 421 -1342
rect 179 -1390 183 -1386
rect 205 -1390 209 -1386
rect 248 -1390 252 -1386
rect 283 -1390 287 -1386
rect 327 -1390 331 -1386
rect 344 -1390 348 -1386
rect 380 -1390 384 -1386
rect 401 -1390 405 -1386
rect 446 -1338 450 -1334
rect 504 -1032 508 -1028
rect 786 -984 790 -980
rect 803 -984 807 -980
rect 495 -1076 499 -1072
rect 478 -1134 482 -1130
rect 495 -1134 499 -1130
rect 430 -1353 434 -1349
rect 417 -1411 421 -1407
rect 448 -1411 452 -1407
rect 170 -1455 174 -1451
rect 187 -1455 191 -1451
rect 126 -1669 130 -1665
rect 111 -1720 115 -1716
rect 140 -1720 144 -1716
rect -138 -1746 -134 -1742
rect -121 -1746 -117 -1742
rect -180 -1960 -176 -1956
rect -199 -2004 -195 -2000
rect -166 -2004 -162 -2000
rect -446 -2068 -442 -2064
rect -429 -2068 -425 -2064
rect -490 -2282 -486 -2278
rect -505 -2333 -501 -2329
rect -476 -2333 -472 -2329
rect -754 -2359 -750 -2355
rect -737 -2359 -733 -2355
rect -793 -2573 -789 -2569
rect -814 -2617 -810 -2613
rect -780 -2617 -776 -2613
rect -1062 -2650 -1058 -2646
rect -1045 -2650 -1041 -2646
rect -1225 -2901 -1221 -2897
rect -1181 -2901 -1177 -2897
rect -1147 -2901 -1143 -2897
rect -1257 -2908 -1253 -2904
rect -1309 -2941 -1305 -2937
rect -1292 -2941 -1288 -2937
rect -1292 -3033 -1288 -3029
rect -1090 -2915 -1086 -2911
rect -1106 -2994 -1102 -2990
rect -1225 -3100 -1221 -3096
rect -1208 -3100 -1204 -3096
rect -1168 -3100 -1164 -3096
rect -1147 -3100 -1143 -3096
rect -1257 -3156 -1253 -3152
rect -1234 -3149 -1230 -3145
rect -1283 -3163 -1279 -3159
rect -1190 -3170 -1186 -3166
rect -1106 -3140 -1102 -3136
rect -1138 -3148 -1134 -3144
rect -1208 -3177 -1204 -3173
rect -1172 -3177 -1168 -3173
rect -1036 -2703 -1032 -2699
rect -793 -2703 -789 -2699
rect -1045 -2742 -1041 -2738
rect -1053 -2809 -1049 -2805
rect -1027 -2809 -1023 -2805
rect -1010 -2809 -1006 -2805
rect -970 -2809 -966 -2805
rect -949 -2809 -945 -2805
rect -932 -2809 -928 -2805
rect -892 -2809 -888 -2805
rect -868 -2809 -864 -2805
rect -831 -2809 -827 -2805
rect -1062 -2842 -1058 -2838
rect -1044 -2835 -1040 -2831
rect -1018 -2857 -1014 -2853
rect -1036 -2864 -1032 -2860
rect -992 -2849 -988 -2845
rect -940 -2842 -936 -2838
rect -1010 -2886 -1006 -2882
rect -974 -2886 -970 -2882
rect -914 -2857 -910 -2853
rect -932 -2886 -928 -2882
rect -896 -2886 -892 -2882
rect -822 -2849 -818 -2845
rect -814 -2857 -810 -2853
rect -1053 -2901 -1049 -2897
rect -1027 -2901 -1023 -2897
rect -984 -2901 -980 -2897
rect -949 -2901 -945 -2897
rect -905 -2901 -901 -2897
rect -888 -2901 -884 -2897
rect -852 -2901 -848 -2897
rect -831 -2901 -827 -2897
rect -780 -2849 -776 -2845
rect -728 -2412 -724 -2408
rect -490 -2412 -486 -2408
rect -737 -2451 -733 -2447
rect -745 -2518 -741 -2514
rect -719 -2518 -715 -2514
rect -702 -2518 -698 -2514
rect -662 -2518 -658 -2514
rect -641 -2518 -637 -2514
rect -624 -2518 -620 -2514
rect -584 -2518 -580 -2514
rect -560 -2518 -556 -2514
rect -523 -2518 -519 -2514
rect -754 -2551 -750 -2547
rect -736 -2544 -732 -2540
rect -710 -2566 -706 -2562
rect -728 -2573 -724 -2569
rect -684 -2558 -680 -2554
rect -632 -2551 -628 -2547
rect -702 -2595 -698 -2591
rect -666 -2595 -662 -2591
rect -606 -2566 -602 -2562
rect -624 -2595 -620 -2591
rect -588 -2595 -584 -2591
rect -514 -2557 -510 -2553
rect -505 -2566 -501 -2562
rect -745 -2610 -741 -2606
rect -719 -2610 -715 -2606
rect -676 -2610 -672 -2606
rect -641 -2610 -637 -2606
rect -597 -2610 -593 -2606
rect -580 -2610 -576 -2606
rect -544 -2610 -540 -2606
rect -523 -2610 -519 -2606
rect -476 -2558 -472 -2554
rect -420 -2121 -416 -2117
rect -180 -2121 -176 -2117
rect -429 -2160 -425 -2156
rect -437 -2227 -433 -2223
rect -411 -2227 -407 -2223
rect -394 -2227 -390 -2223
rect -354 -2227 -350 -2223
rect -333 -2227 -329 -2223
rect -316 -2227 -312 -2223
rect -276 -2227 -272 -2223
rect -252 -2227 -248 -2223
rect -215 -2227 -211 -2223
rect -446 -2260 -442 -2256
rect -428 -2253 -424 -2249
rect -402 -2275 -398 -2271
rect -420 -2282 -416 -2278
rect -376 -2267 -372 -2263
rect -324 -2260 -320 -2256
rect -394 -2304 -390 -2300
rect -358 -2304 -354 -2300
rect -298 -2275 -294 -2271
rect -316 -2304 -312 -2300
rect -280 -2304 -276 -2300
rect -206 -2267 -202 -2263
rect -198 -2275 -194 -2271
rect -437 -2319 -433 -2315
rect -411 -2319 -407 -2315
rect -368 -2319 -364 -2315
rect -333 -2319 -329 -2315
rect -289 -2319 -285 -2315
rect -272 -2319 -268 -2315
rect -236 -2319 -232 -2315
rect -215 -2319 -211 -2315
rect -166 -2267 -162 -2263
rect -112 -1799 -108 -1795
rect 126 -1799 130 -1795
rect -121 -1838 -117 -1834
rect -129 -1905 -125 -1901
rect -103 -1905 -99 -1901
rect -86 -1905 -82 -1901
rect -46 -1905 -42 -1901
rect -25 -1905 -21 -1901
rect -8 -1905 -4 -1901
rect 32 -1905 36 -1901
rect 56 -1905 60 -1901
rect 93 -1905 97 -1901
rect -138 -1938 -134 -1934
rect -120 -1931 -116 -1927
rect -94 -1953 -90 -1949
rect -112 -1960 -108 -1956
rect -68 -1945 -64 -1941
rect -16 -1938 -12 -1934
rect -86 -1982 -82 -1978
rect -50 -1982 -46 -1978
rect 10 -1953 14 -1949
rect -8 -1982 -4 -1978
rect 28 -1982 32 -1978
rect 102 -1945 106 -1941
rect 112 -1953 116 -1949
rect -129 -1997 -125 -1993
rect -103 -1997 -99 -1993
rect -60 -1997 -56 -1993
rect -25 -1997 -21 -1993
rect 19 -1997 23 -1993
rect 36 -1997 40 -1993
rect 72 -1997 76 -1993
rect 93 -1997 97 -1993
rect 140 -1945 144 -1941
rect 196 -1508 200 -1504
rect 434 -1508 438 -1504
rect 187 -1547 191 -1543
rect 179 -1614 183 -1610
rect 205 -1614 209 -1610
rect 222 -1614 226 -1610
rect 262 -1614 266 -1610
rect 283 -1614 287 -1610
rect 300 -1614 304 -1610
rect 340 -1614 344 -1610
rect 364 -1614 368 -1610
rect 401 -1614 405 -1610
rect 170 -1647 174 -1643
rect 188 -1640 192 -1636
rect 214 -1662 218 -1658
rect 196 -1669 200 -1665
rect 240 -1654 244 -1650
rect 292 -1647 296 -1643
rect 222 -1691 226 -1687
rect 258 -1691 262 -1687
rect 318 -1662 322 -1658
rect 300 -1691 304 -1687
rect 336 -1691 340 -1687
rect 410 -1654 414 -1650
rect 418 -1662 422 -1658
rect 179 -1706 183 -1702
rect 205 -1706 209 -1702
rect 248 -1706 252 -1702
rect 283 -1706 287 -1702
rect 327 -1706 331 -1702
rect 344 -1706 348 -1702
rect 380 -1706 384 -1702
rect 401 -1706 405 -1702
rect 448 -1654 452 -1650
rect 812 -1040 816 -1036
rect 803 -1076 807 -1072
rect 786 -1134 790 -1130
rect 803 -1134 807 -1130
rect 504 -1187 508 -1183
rect 738 -1187 742 -1183
rect 495 -1226 499 -1222
rect 487 -1298 491 -1294
rect 513 -1298 517 -1294
rect 530 -1298 534 -1294
rect 570 -1298 574 -1294
rect 591 -1298 595 -1294
rect 608 -1298 612 -1294
rect 648 -1298 652 -1294
rect 672 -1298 676 -1294
rect 709 -1298 713 -1294
rect 478 -1331 482 -1327
rect 496 -1324 500 -1320
rect 522 -1346 526 -1342
rect 504 -1353 508 -1349
rect 548 -1338 552 -1334
rect 600 -1331 604 -1327
rect 530 -1375 534 -1371
rect 566 -1375 570 -1371
rect 626 -1346 630 -1342
rect 608 -1375 612 -1371
rect 644 -1375 648 -1371
rect 718 -1354 722 -1350
rect 725 -1346 729 -1342
rect 487 -1390 491 -1386
rect 513 -1390 517 -1386
rect 556 -1390 560 -1386
rect 591 -1390 595 -1386
rect 635 -1390 639 -1386
rect 652 -1390 656 -1386
rect 688 -1390 692 -1386
rect 709 -1390 713 -1386
rect 738 -1361 742 -1357
rect 725 -1404 729 -1400
rect 759 -1404 763 -1400
rect 478 -1455 482 -1451
rect 495 -1455 499 -1451
rect 434 -1669 438 -1665
rect 418 -1713 422 -1709
rect 449 -1713 453 -1709
rect 170 -1746 174 -1742
rect 187 -1746 191 -1742
rect 126 -1960 130 -1956
rect 112 -2011 116 -2007
rect 140 -2011 144 -2007
rect -138 -2068 -134 -2064
rect -121 -2068 -117 -2064
rect -180 -2282 -176 -2278
rect -198 -2326 -194 -2322
rect -166 -2326 -162 -2322
rect -446 -2359 -442 -2355
rect -429 -2359 -425 -2355
rect -490 -2573 -486 -2569
rect -505 -2624 -501 -2620
rect -476 -2624 -472 -2620
rect -754 -2650 -750 -2646
rect -737 -2650 -733 -2646
rect -793 -2864 -789 -2860
rect -814 -2908 -810 -2904
rect -780 -2908 -776 -2904
rect -1062 -2941 -1058 -2937
rect -1045 -2941 -1041 -2937
rect -1036 -2994 -1032 -2990
rect -793 -2994 -789 -2990
rect -1045 -3033 -1041 -3029
rect -1090 -3155 -1086 -3151
rect -1225 -3192 -1221 -3188
rect -1181 -3192 -1177 -3188
rect -1147 -3192 -1143 -3188
rect -1053 -3100 -1049 -3096
rect -1027 -3100 -1023 -3096
rect -1010 -3100 -1006 -3096
rect -970 -3100 -966 -3096
rect -949 -3100 -945 -3096
rect -932 -3100 -928 -3096
rect -892 -3100 -888 -3096
rect -868 -3100 -864 -3096
rect -831 -3100 -827 -3096
rect -1062 -3133 -1058 -3129
rect -1044 -3126 -1040 -3122
rect -1018 -3148 -1014 -3144
rect -1036 -3155 -1032 -3151
rect -992 -3140 -988 -3136
rect -940 -3133 -936 -3129
rect -1010 -3177 -1006 -3173
rect -974 -3177 -970 -3173
rect -914 -3148 -910 -3144
rect -932 -3177 -928 -3173
rect -896 -3177 -892 -3173
rect -822 -3140 -818 -3136
rect -728 -2703 -724 -2699
rect -490 -2703 -486 -2699
rect -737 -2742 -733 -2738
rect -745 -2809 -741 -2805
rect -719 -2809 -715 -2805
rect -702 -2809 -698 -2805
rect -662 -2809 -658 -2805
rect -641 -2809 -637 -2805
rect -624 -2809 -620 -2805
rect -584 -2809 -580 -2805
rect -560 -2809 -556 -2805
rect -523 -2809 -519 -2805
rect -754 -2842 -750 -2838
rect -736 -2835 -732 -2831
rect -710 -2857 -706 -2853
rect -728 -2864 -724 -2860
rect -684 -2849 -680 -2845
rect -632 -2842 -628 -2838
rect -702 -2886 -698 -2882
rect -666 -2886 -662 -2882
rect -606 -2857 -602 -2853
rect -624 -2886 -620 -2882
rect -588 -2886 -584 -2882
rect -514 -2848 -510 -2844
rect -505 -2857 -501 -2853
rect -745 -2901 -741 -2897
rect -719 -2901 -715 -2897
rect -676 -2901 -672 -2897
rect -641 -2901 -637 -2897
rect -597 -2901 -593 -2897
rect -580 -2901 -576 -2897
rect -544 -2901 -540 -2897
rect -523 -2901 -519 -2897
rect -476 -2849 -472 -2845
rect -420 -2412 -416 -2408
rect -180 -2412 -176 -2408
rect -429 -2451 -425 -2447
rect -437 -2518 -433 -2514
rect -411 -2518 -407 -2514
rect -394 -2518 -390 -2514
rect -354 -2518 -350 -2514
rect -333 -2518 -329 -2514
rect -316 -2518 -312 -2514
rect -276 -2518 -272 -2514
rect -252 -2518 -248 -2514
rect -215 -2518 -211 -2514
rect -446 -2551 -442 -2547
rect -428 -2544 -424 -2540
rect -402 -2566 -398 -2562
rect -420 -2573 -416 -2569
rect -376 -2558 -372 -2554
rect -324 -2551 -320 -2547
rect -394 -2595 -390 -2591
rect -358 -2595 -354 -2591
rect -298 -2566 -294 -2562
rect -316 -2595 -312 -2591
rect -280 -2595 -276 -2591
rect -206 -2558 -202 -2554
rect -198 -2566 -194 -2562
rect -437 -2610 -433 -2606
rect -411 -2610 -407 -2606
rect -368 -2610 -364 -2606
rect -333 -2610 -329 -2606
rect -289 -2610 -285 -2606
rect -272 -2610 -268 -2606
rect -236 -2610 -232 -2606
rect -215 -2610 -211 -2606
rect -166 -2558 -162 -2554
rect -112 -2121 -108 -2117
rect 126 -2121 130 -2117
rect -121 -2160 -117 -2156
rect -129 -2227 -125 -2223
rect -103 -2227 -99 -2223
rect -86 -2227 -82 -2223
rect -46 -2227 -42 -2223
rect -25 -2227 -21 -2223
rect -8 -2227 -4 -2223
rect 32 -2227 36 -2223
rect 56 -2227 60 -2223
rect 93 -2227 97 -2223
rect -138 -2260 -134 -2256
rect -120 -2253 -116 -2249
rect -94 -2275 -90 -2271
rect -112 -2282 -108 -2278
rect -68 -2267 -64 -2263
rect -16 -2260 -12 -2256
rect -86 -2304 -82 -2300
rect -50 -2304 -46 -2300
rect 10 -2275 14 -2271
rect -8 -2304 -4 -2300
rect 28 -2304 32 -2300
rect 102 -2267 106 -2263
rect 111 -2275 115 -2271
rect -129 -2319 -125 -2315
rect -103 -2319 -99 -2315
rect -60 -2319 -56 -2315
rect -25 -2319 -21 -2315
rect 19 -2319 23 -2315
rect 36 -2319 40 -2315
rect 72 -2319 76 -2315
rect 93 -2319 97 -2315
rect 140 -2267 144 -2263
rect 196 -1799 200 -1795
rect 435 -1799 439 -1795
rect 187 -1838 191 -1834
rect 179 -1905 183 -1901
rect 205 -1905 209 -1901
rect 222 -1905 226 -1901
rect 262 -1905 266 -1901
rect 283 -1905 287 -1901
rect 300 -1905 304 -1901
rect 340 -1905 344 -1901
rect 364 -1905 368 -1901
rect 401 -1905 405 -1901
rect 170 -1938 174 -1934
rect 188 -1931 192 -1927
rect 214 -1953 218 -1949
rect 196 -1960 200 -1956
rect 240 -1945 244 -1941
rect 292 -1938 296 -1934
rect 222 -1982 226 -1978
rect 258 -1982 262 -1978
rect 318 -1953 322 -1949
rect 300 -1982 304 -1978
rect 336 -1982 340 -1978
rect 410 -1945 414 -1941
rect 417 -1953 421 -1949
rect 179 -1997 183 -1993
rect 205 -1997 209 -1993
rect 248 -1997 252 -1993
rect 283 -1997 287 -1993
rect 327 -1997 331 -1993
rect 344 -1997 348 -1993
rect 380 -1997 384 -1993
rect 401 -1997 405 -1993
rect 449 -1945 453 -1941
rect 504 -1508 508 -1504
rect 742 -1508 746 -1504
rect 495 -1547 499 -1543
rect 487 -1614 491 -1610
rect 513 -1614 517 -1610
rect 530 -1614 534 -1610
rect 570 -1614 574 -1610
rect 591 -1614 595 -1610
rect 608 -1614 612 -1610
rect 648 -1614 652 -1610
rect 672 -1614 676 -1610
rect 709 -1614 713 -1610
rect 478 -1647 482 -1643
rect 496 -1640 500 -1636
rect 522 -1662 526 -1658
rect 504 -1669 508 -1665
rect 548 -1654 552 -1650
rect 600 -1647 604 -1643
rect 530 -1691 534 -1687
rect 566 -1691 570 -1687
rect 626 -1662 630 -1658
rect 608 -1691 612 -1687
rect 644 -1691 648 -1687
rect 718 -1652 722 -1648
rect 742 -1654 746 -1650
rect 718 -1670 722 -1666
rect 726 -1662 730 -1658
rect 487 -1706 491 -1702
rect 513 -1706 517 -1702
rect 556 -1706 560 -1702
rect 591 -1706 595 -1702
rect 635 -1706 639 -1702
rect 652 -1706 656 -1702
rect 688 -1706 692 -1702
rect 709 -1706 713 -1702
rect 759 -1669 763 -1665
rect 812 -1187 816 -1183
rect 803 -1226 807 -1222
rect 793 -1298 797 -1294
rect 810 -1298 814 -1294
rect 850 -1298 854 -1294
rect 871 -1298 875 -1294
rect 784 -1347 788 -1343
rect 828 -1368 832 -1364
rect 880 -1346 884 -1342
rect 810 -1375 814 -1371
rect 846 -1375 850 -1371
rect 897 -1368 901 -1364
rect 793 -1390 797 -1386
rect 837 -1390 841 -1386
rect 871 -1390 875 -1386
rect 904 -1404 908 -1400
rect 897 -1411 901 -1407
rect 786 -1455 790 -1451
rect 803 -1455 807 -1451
rect 726 -1720 730 -1716
rect 759 -1720 763 -1716
rect 478 -1746 482 -1742
rect 495 -1746 499 -1742
rect 435 -1960 439 -1956
rect 417 -2004 421 -2000
rect 448 -2004 452 -2000
rect 170 -2068 174 -2064
rect 187 -2068 191 -2064
rect 126 -2282 130 -2278
rect 111 -2333 115 -2329
rect 140 -2333 144 -2329
rect -138 -2359 -134 -2355
rect -121 -2359 -117 -2355
rect -180 -2573 -176 -2569
rect -198 -2617 -194 -2613
rect -166 -2617 -162 -2613
rect -446 -2650 -442 -2646
rect -429 -2650 -425 -2646
rect -490 -2864 -486 -2860
rect -505 -2915 -501 -2911
rect -476 -2915 -472 -2911
rect -754 -2941 -750 -2937
rect -737 -2941 -733 -2937
rect -728 -2994 -724 -2990
rect -490 -2994 -486 -2990
rect -737 -3033 -733 -3029
rect -745 -3100 -741 -3096
rect -719 -3100 -715 -3096
rect -702 -3100 -698 -3096
rect -662 -3100 -658 -3096
rect -641 -3100 -637 -3096
rect -624 -3100 -620 -3096
rect -584 -3100 -580 -3096
rect -560 -3100 -556 -3096
rect -523 -3100 -519 -3096
rect -780 -3140 -776 -3136
rect -754 -3133 -750 -3129
rect -793 -3155 -789 -3151
rect -736 -3126 -732 -3122
rect -710 -3148 -706 -3144
rect -728 -3155 -724 -3151
rect -684 -3140 -680 -3136
rect -632 -3133 -628 -3129
rect -702 -3177 -698 -3173
rect -666 -3177 -662 -3173
rect -606 -3148 -602 -3144
rect -624 -3177 -620 -3173
rect -588 -3177 -584 -3173
rect -514 -3139 -510 -3135
rect -420 -2703 -416 -2699
rect -180 -2703 -176 -2699
rect -429 -2742 -425 -2738
rect -437 -2809 -433 -2805
rect -411 -2809 -407 -2805
rect -394 -2809 -390 -2805
rect -354 -2809 -350 -2805
rect -333 -2809 -329 -2805
rect -316 -2809 -312 -2805
rect -276 -2809 -272 -2805
rect -252 -2809 -248 -2805
rect -215 -2809 -211 -2805
rect -446 -2842 -442 -2838
rect -428 -2835 -424 -2831
rect -402 -2857 -398 -2853
rect -420 -2864 -416 -2860
rect -376 -2849 -372 -2845
rect -324 -2842 -320 -2838
rect -394 -2886 -390 -2882
rect -358 -2886 -354 -2882
rect -298 -2857 -294 -2853
rect -316 -2886 -312 -2882
rect -280 -2886 -276 -2882
rect -206 -2849 -202 -2845
rect -198 -2857 -194 -2853
rect -437 -2901 -433 -2897
rect -411 -2901 -407 -2897
rect -368 -2901 -364 -2897
rect -333 -2901 -329 -2897
rect -289 -2901 -285 -2897
rect -272 -2901 -268 -2897
rect -236 -2901 -232 -2897
rect -215 -2901 -211 -2897
rect -166 -2849 -162 -2845
rect -112 -2412 -108 -2408
rect 126 -2412 130 -2408
rect -121 -2451 -117 -2447
rect -129 -2518 -125 -2514
rect -103 -2518 -99 -2514
rect -86 -2518 -82 -2514
rect -46 -2518 -42 -2514
rect -25 -2518 -21 -2514
rect -8 -2518 -4 -2514
rect 32 -2518 36 -2514
rect 56 -2518 60 -2514
rect 93 -2518 97 -2514
rect -138 -2551 -134 -2547
rect -120 -2544 -116 -2540
rect -94 -2566 -90 -2562
rect -112 -2573 -108 -2569
rect -68 -2558 -64 -2554
rect -16 -2551 -12 -2547
rect -86 -2595 -82 -2591
rect -50 -2595 -46 -2591
rect 10 -2566 14 -2562
rect -8 -2595 -4 -2591
rect 28 -2595 32 -2591
rect 102 -2558 106 -2554
rect 111 -2566 115 -2562
rect -129 -2610 -125 -2606
rect -103 -2610 -99 -2606
rect -60 -2610 -56 -2606
rect -25 -2610 -21 -2606
rect 19 -2610 23 -2606
rect 36 -2610 40 -2606
rect 72 -2610 76 -2606
rect 93 -2610 97 -2606
rect 140 -2558 144 -2554
rect 196 -2121 200 -2117
rect 434 -2121 438 -2117
rect 187 -2160 191 -2156
rect 504 -1799 508 -1795
rect 742 -1799 746 -1795
rect 495 -1838 499 -1834
rect 487 -1905 491 -1901
rect 513 -1905 517 -1901
rect 530 -1905 534 -1901
rect 570 -1905 574 -1901
rect 591 -1905 595 -1901
rect 608 -1905 612 -1901
rect 648 -1905 652 -1901
rect 672 -1905 676 -1901
rect 709 -1905 713 -1901
rect 478 -1938 482 -1934
rect 496 -1931 500 -1927
rect 522 -1953 526 -1949
rect 504 -1960 508 -1956
rect 548 -1945 552 -1941
rect 600 -1938 604 -1934
rect 530 -1982 534 -1978
rect 566 -1982 570 -1978
rect 626 -1953 630 -1949
rect 608 -1982 612 -1978
rect 644 -1982 648 -1978
rect 718 -1943 722 -1939
rect 742 -1945 746 -1941
rect 718 -1961 722 -1957
rect 728 -1953 732 -1949
rect 487 -1997 491 -1993
rect 513 -1997 517 -1993
rect 556 -1997 560 -1993
rect 591 -1997 595 -1993
rect 635 -1997 639 -1993
rect 652 -1997 656 -1993
rect 688 -1997 692 -1993
rect 709 -1997 713 -1993
rect 759 -1960 763 -1956
rect 812 -1508 816 -1504
rect 803 -1547 807 -1543
rect 795 -1614 799 -1610
rect 821 -1614 825 -1610
rect 838 -1614 842 -1610
rect 878 -1614 882 -1610
rect 899 -1614 903 -1610
rect 916 -1614 920 -1610
rect 956 -1614 960 -1610
rect 980 -1614 984 -1610
rect 1017 -1614 1021 -1610
rect 786 -1647 790 -1643
rect 804 -1640 808 -1636
rect 830 -1662 834 -1658
rect 812 -1669 816 -1665
rect 856 -1654 860 -1650
rect 908 -1647 912 -1643
rect 838 -1691 842 -1687
rect 874 -1691 878 -1687
rect 934 -1662 938 -1658
rect 916 -1691 920 -1687
rect 952 -1691 956 -1687
rect 795 -1706 799 -1702
rect 821 -1706 825 -1702
rect 864 -1706 868 -1702
rect 899 -1706 903 -1702
rect 943 -1706 947 -1702
rect 960 -1706 964 -1702
rect 996 -1706 1000 -1702
rect 1017 -1706 1021 -1702
rect 1041 -1662 1045 -1658
rect 1041 -1713 1045 -1709
rect 1026 -1720 1030 -1716
rect 786 -1746 790 -1742
rect 803 -1746 807 -1742
rect 728 -2011 732 -2007
rect 759 -2011 763 -2007
rect 478 -2068 482 -2064
rect 495 -2068 499 -2064
rect 179 -2227 183 -2223
rect 205 -2227 209 -2223
rect 222 -2227 226 -2223
rect 262 -2227 266 -2223
rect 283 -2227 287 -2223
rect 300 -2227 304 -2223
rect 340 -2227 344 -2223
rect 364 -2227 368 -2223
rect 401 -2227 405 -2223
rect 170 -2260 174 -2256
rect 188 -2253 192 -2249
rect 214 -2275 218 -2271
rect 196 -2282 200 -2278
rect 240 -2267 244 -2263
rect 292 -2260 296 -2256
rect 222 -2304 226 -2300
rect 258 -2304 262 -2300
rect 318 -2275 322 -2271
rect 300 -2304 304 -2300
rect 336 -2304 340 -2300
rect 410 -2267 414 -2263
rect 418 -2275 422 -2271
rect 179 -2319 183 -2315
rect 205 -2319 209 -2315
rect 248 -2319 252 -2315
rect 283 -2319 287 -2315
rect 327 -2319 331 -2315
rect 344 -2319 348 -2315
rect 380 -2319 384 -2315
rect 401 -2319 405 -2315
rect 449 -2267 453 -2263
rect 435 -2282 439 -2278
rect 418 -2326 422 -2322
rect 449 -2326 453 -2322
rect 170 -2359 174 -2355
rect 187 -2359 191 -2355
rect 126 -2573 130 -2569
rect 111 -2624 115 -2620
rect 140 -2624 144 -2620
rect -138 -2650 -134 -2646
rect -121 -2650 -117 -2646
rect -180 -2864 -176 -2860
rect -198 -2908 -194 -2904
rect -169 -2908 -165 -2904
rect -446 -2941 -442 -2937
rect -429 -2941 -425 -2937
rect -420 -2994 -416 -2990
rect -180 -2994 -176 -2990
rect -429 -3033 -425 -3029
rect -476 -3140 -472 -3136
rect -490 -3155 -486 -3151
rect -1053 -3192 -1049 -3188
rect -1027 -3192 -1023 -3188
rect -984 -3192 -980 -3188
rect -949 -3192 -945 -3188
rect -905 -3192 -901 -3188
rect -888 -3192 -884 -3188
rect -852 -3192 -848 -3188
rect -831 -3192 -827 -3188
rect -745 -3192 -741 -3188
rect -719 -3192 -715 -3188
rect -676 -3192 -672 -3188
rect -641 -3192 -637 -3188
rect -597 -3192 -593 -3188
rect -580 -3192 -576 -3188
rect -544 -3192 -540 -3188
rect -523 -3192 -519 -3188
rect -437 -3100 -433 -3096
rect -411 -3100 -407 -3096
rect -394 -3100 -390 -3096
rect -354 -3100 -350 -3096
rect -333 -3100 -329 -3096
rect -316 -3100 -312 -3096
rect -276 -3100 -272 -3096
rect -252 -3100 -248 -3096
rect -215 -3100 -211 -3096
rect -446 -3133 -442 -3129
rect -428 -3126 -424 -3122
rect -402 -3148 -398 -3144
rect -420 -3155 -416 -3151
rect -376 -3140 -372 -3136
rect -324 -3133 -320 -3129
rect -394 -3177 -390 -3173
rect -358 -3177 -354 -3173
rect -298 -3148 -294 -3144
rect -316 -3177 -312 -3173
rect -280 -3177 -276 -3173
rect -206 -3140 -202 -3136
rect -112 -2703 -108 -2699
rect 126 -2703 130 -2699
rect -121 -2742 -117 -2738
rect -129 -2809 -125 -2805
rect -103 -2809 -99 -2805
rect -86 -2809 -82 -2805
rect -46 -2809 -42 -2805
rect -25 -2809 -21 -2805
rect -8 -2809 -4 -2805
rect 32 -2809 36 -2805
rect 56 -2809 60 -2805
rect 93 -2809 97 -2805
rect -138 -2842 -134 -2838
rect -120 -2835 -116 -2831
rect -94 -2857 -90 -2853
rect -112 -2864 -108 -2860
rect -68 -2849 -64 -2845
rect -16 -2842 -12 -2838
rect -86 -2886 -82 -2882
rect -50 -2886 -46 -2882
rect 10 -2857 14 -2853
rect -8 -2886 -4 -2882
rect 28 -2886 32 -2882
rect 102 -2849 106 -2845
rect 111 -2857 115 -2853
rect -129 -2901 -125 -2897
rect -103 -2901 -99 -2897
rect -60 -2901 -56 -2897
rect -25 -2901 -21 -2897
rect 19 -2901 23 -2897
rect 36 -2901 40 -2897
rect 72 -2901 76 -2897
rect 93 -2901 97 -2897
rect 140 -2849 144 -2845
rect 196 -2412 200 -2408
rect 435 -2412 439 -2408
rect 187 -2451 191 -2447
rect 179 -2518 183 -2514
rect 205 -2518 209 -2514
rect 222 -2518 226 -2514
rect 262 -2518 266 -2514
rect 283 -2518 287 -2514
rect 300 -2518 304 -2514
rect 340 -2518 344 -2514
rect 364 -2518 368 -2514
rect 401 -2518 405 -2514
rect 170 -2551 174 -2547
rect 188 -2544 192 -2540
rect 214 -2566 218 -2562
rect 196 -2573 200 -2569
rect 240 -2558 244 -2554
rect 292 -2551 296 -2547
rect 222 -2595 226 -2591
rect 258 -2595 262 -2591
rect 318 -2566 322 -2562
rect 300 -2595 304 -2591
rect 336 -2595 340 -2591
rect 410 -2558 414 -2554
rect 418 -2566 422 -2562
rect 179 -2610 183 -2606
rect 205 -2610 209 -2606
rect 248 -2610 252 -2606
rect 283 -2610 287 -2606
rect 327 -2610 331 -2606
rect 344 -2610 348 -2606
rect 380 -2610 384 -2606
rect 401 -2610 405 -2606
rect 449 -2558 453 -2554
rect 504 -2121 508 -2117
rect 742 -2121 746 -2117
rect 495 -2160 499 -2156
rect 487 -2227 491 -2223
rect 513 -2227 517 -2223
rect 530 -2227 534 -2223
rect 570 -2227 574 -2223
rect 591 -2227 595 -2223
rect 608 -2227 612 -2223
rect 648 -2227 652 -2223
rect 672 -2227 676 -2223
rect 709 -2227 713 -2223
rect 478 -2260 482 -2256
rect 496 -2253 500 -2249
rect 522 -2275 526 -2271
rect 504 -2282 508 -2278
rect 548 -2267 552 -2263
rect 600 -2260 604 -2256
rect 530 -2304 534 -2300
rect 566 -2304 570 -2300
rect 626 -2275 630 -2271
rect 608 -2304 612 -2300
rect 644 -2304 648 -2300
rect 718 -2265 722 -2261
rect 742 -2267 746 -2263
rect 726 -2275 730 -2271
rect 487 -2319 491 -2315
rect 513 -2319 517 -2315
rect 556 -2319 560 -2315
rect 591 -2319 595 -2315
rect 635 -2319 639 -2315
rect 652 -2319 656 -2315
rect 688 -2319 692 -2315
rect 709 -2319 713 -2315
rect 759 -2282 763 -2278
rect 812 -1799 816 -1795
rect 803 -1838 807 -1834
rect 795 -1905 799 -1901
rect 821 -1905 825 -1901
rect 838 -1905 842 -1901
rect 878 -1905 882 -1901
rect 899 -1905 903 -1901
rect 916 -1905 920 -1901
rect 956 -1905 960 -1901
rect 980 -1905 984 -1901
rect 1017 -1905 1021 -1901
rect 786 -1938 790 -1934
rect 804 -1931 808 -1927
rect 830 -1953 834 -1949
rect 812 -1960 816 -1956
rect 856 -1945 860 -1941
rect 908 -1938 912 -1934
rect 838 -1982 842 -1978
rect 874 -1982 878 -1978
rect 934 -1953 938 -1949
rect 916 -1982 920 -1978
rect 952 -1982 956 -1978
rect 795 -1997 799 -1993
rect 821 -1997 825 -1993
rect 864 -1997 868 -1993
rect 899 -1997 903 -1993
rect 943 -1997 947 -1993
rect 960 -1997 964 -1993
rect 996 -1997 1000 -1993
rect 1017 -1997 1021 -1993
rect 1042 -1953 1046 -1949
rect 1042 -2004 1046 -2000
rect 1026 -2011 1030 -2007
rect 786 -2068 790 -2064
rect 803 -2068 807 -2064
rect 726 -2333 730 -2329
rect 759 -2333 763 -2329
rect 478 -2359 482 -2355
rect 495 -2359 499 -2355
rect 435 -2573 439 -2569
rect 418 -2617 422 -2613
rect 449 -2617 453 -2613
rect 170 -2650 174 -2646
rect 187 -2650 191 -2646
rect 126 -2864 130 -2860
rect 111 -2915 115 -2911
rect 139 -2915 143 -2911
rect -138 -2941 -134 -2937
rect -121 -2941 -117 -2937
rect -112 -2994 -108 -2990
rect 126 -2994 130 -2990
rect -121 -3033 -117 -3029
rect -169 -3140 -165 -3136
rect -180 -3155 -176 -3151
rect -437 -3192 -433 -3188
rect -411 -3192 -407 -3188
rect -368 -3192 -364 -3188
rect -333 -3192 -329 -3188
rect -289 -3192 -285 -3188
rect -272 -3192 -268 -3188
rect -236 -3192 -232 -3188
rect -215 -3192 -211 -3188
rect -129 -3100 -125 -3096
rect -103 -3100 -99 -3096
rect -86 -3100 -82 -3096
rect -46 -3100 -42 -3096
rect -25 -3100 -21 -3096
rect -8 -3100 -4 -3096
rect 32 -3100 36 -3096
rect 56 -3100 60 -3096
rect 93 -3100 97 -3096
rect -138 -3133 -134 -3129
rect -120 -3126 -116 -3122
rect -94 -3148 -90 -3144
rect -112 -3155 -108 -3151
rect -68 -3140 -64 -3136
rect -16 -3133 -12 -3129
rect -86 -3177 -82 -3173
rect -50 -3177 -46 -3173
rect 10 -3148 14 -3144
rect -8 -3177 -4 -3173
rect 28 -3177 32 -3173
rect 102 -3140 106 -3136
rect 196 -2703 200 -2699
rect 435 -2703 439 -2699
rect 187 -2742 191 -2738
rect 179 -2809 183 -2805
rect 205 -2809 209 -2805
rect 222 -2809 226 -2805
rect 262 -2809 266 -2805
rect 283 -2809 287 -2805
rect 300 -2809 304 -2805
rect 340 -2809 344 -2805
rect 364 -2809 368 -2805
rect 401 -2809 405 -2805
rect 170 -2842 174 -2838
rect 188 -2835 192 -2831
rect 214 -2857 218 -2853
rect 196 -2864 200 -2860
rect 240 -2849 244 -2845
rect 292 -2842 296 -2838
rect 222 -2886 226 -2882
rect 258 -2886 262 -2882
rect 318 -2857 322 -2853
rect 300 -2886 304 -2882
rect 336 -2886 340 -2882
rect 410 -2849 414 -2845
rect 418 -2857 422 -2853
rect 179 -2901 183 -2897
rect 205 -2901 209 -2897
rect 248 -2901 252 -2897
rect 283 -2901 287 -2897
rect 327 -2901 331 -2897
rect 344 -2901 348 -2897
rect 380 -2901 384 -2897
rect 401 -2901 405 -2897
rect 449 -2849 453 -2845
rect 504 -2412 508 -2408
rect 742 -2412 746 -2408
rect 495 -2451 499 -2447
rect 487 -2518 491 -2514
rect 513 -2518 517 -2514
rect 530 -2518 534 -2514
rect 570 -2518 574 -2514
rect 591 -2518 595 -2514
rect 608 -2518 612 -2514
rect 648 -2518 652 -2514
rect 672 -2518 676 -2514
rect 709 -2518 713 -2514
rect 478 -2551 482 -2547
rect 496 -2544 500 -2540
rect 522 -2566 526 -2562
rect 504 -2573 508 -2569
rect 548 -2558 552 -2554
rect 600 -2551 604 -2547
rect 530 -2595 534 -2591
rect 566 -2595 570 -2591
rect 626 -2566 630 -2562
rect 608 -2595 612 -2591
rect 644 -2595 648 -2591
rect 718 -2556 722 -2552
rect 742 -2558 746 -2554
rect 726 -2566 730 -2562
rect 487 -2610 491 -2606
rect 513 -2610 517 -2606
rect 556 -2610 560 -2606
rect 591 -2610 595 -2606
rect 635 -2610 639 -2606
rect 652 -2610 656 -2606
rect 688 -2610 692 -2606
rect 709 -2610 713 -2606
rect 759 -2573 763 -2569
rect 812 -2121 816 -2117
rect 803 -2160 807 -2156
rect 795 -2227 799 -2223
rect 821 -2227 825 -2223
rect 838 -2227 842 -2223
rect 878 -2227 882 -2223
rect 899 -2227 903 -2223
rect 916 -2227 920 -2223
rect 956 -2227 960 -2223
rect 980 -2227 984 -2223
rect 1017 -2227 1021 -2223
rect 786 -2260 790 -2256
rect 804 -2253 808 -2249
rect 830 -2275 834 -2271
rect 812 -2282 816 -2278
rect 856 -2267 860 -2263
rect 908 -2260 912 -2256
rect 838 -2304 842 -2300
rect 874 -2304 878 -2300
rect 934 -2275 938 -2271
rect 916 -2304 920 -2300
rect 952 -2304 956 -2300
rect 795 -2319 799 -2315
rect 821 -2319 825 -2315
rect 864 -2319 868 -2315
rect 899 -2319 903 -2315
rect 943 -2319 947 -2315
rect 960 -2319 964 -2315
rect 996 -2319 1000 -2315
rect 1017 -2319 1021 -2315
rect 1039 -2275 1043 -2271
rect 1039 -2326 1043 -2322
rect 1026 -2333 1030 -2329
rect 786 -2359 790 -2355
rect 803 -2359 807 -2355
rect 726 -2624 730 -2620
rect 759 -2624 763 -2620
rect 478 -2650 482 -2646
rect 495 -2650 499 -2646
rect 435 -2864 439 -2860
rect 418 -2908 422 -2904
rect 447 -2908 451 -2904
rect 170 -2941 174 -2937
rect 187 -2941 191 -2937
rect 196 -2994 200 -2990
rect 435 -2994 439 -2990
rect 187 -3033 191 -3029
rect 179 -3100 183 -3096
rect 205 -3100 209 -3096
rect 222 -3100 226 -3096
rect 262 -3100 266 -3096
rect 283 -3100 287 -3096
rect 300 -3100 304 -3096
rect 340 -3100 344 -3096
rect 364 -3100 368 -3096
rect 401 -3100 405 -3096
rect 139 -3140 143 -3136
rect 170 -3133 174 -3129
rect 126 -3155 130 -3151
rect 188 -3126 192 -3122
rect 214 -3148 218 -3144
rect 196 -3155 200 -3151
rect 240 -3140 244 -3136
rect 292 -3133 296 -3129
rect 222 -3177 226 -3173
rect 258 -3177 262 -3173
rect 318 -3148 322 -3144
rect 300 -3177 304 -3173
rect 336 -3177 340 -3173
rect 410 -3140 414 -3136
rect 504 -2703 508 -2699
rect 742 -2703 746 -2699
rect 495 -2742 499 -2738
rect 487 -2809 491 -2805
rect 513 -2809 517 -2805
rect 530 -2809 534 -2805
rect 570 -2809 574 -2805
rect 591 -2809 595 -2805
rect 608 -2809 612 -2805
rect 648 -2809 652 -2805
rect 672 -2809 676 -2805
rect 709 -2809 713 -2805
rect 478 -2842 482 -2838
rect 496 -2835 500 -2831
rect 522 -2857 526 -2853
rect 504 -2864 508 -2860
rect 548 -2849 552 -2845
rect 600 -2842 604 -2838
rect 530 -2886 534 -2882
rect 566 -2886 570 -2882
rect 626 -2857 630 -2853
rect 608 -2886 612 -2882
rect 644 -2886 648 -2882
rect 718 -2847 722 -2843
rect 742 -2849 746 -2845
rect 726 -2857 730 -2853
rect 487 -2901 491 -2897
rect 513 -2901 517 -2897
rect 556 -2901 560 -2897
rect 591 -2901 595 -2897
rect 635 -2901 639 -2897
rect 652 -2901 656 -2897
rect 688 -2901 692 -2897
rect 709 -2901 713 -2897
rect 759 -2864 763 -2860
rect 812 -2412 816 -2408
rect 803 -2451 807 -2447
rect 795 -2518 799 -2514
rect 821 -2518 825 -2514
rect 838 -2518 842 -2514
rect 878 -2518 882 -2514
rect 899 -2518 903 -2514
rect 916 -2518 920 -2514
rect 956 -2518 960 -2514
rect 980 -2518 984 -2514
rect 1017 -2518 1021 -2514
rect 786 -2551 790 -2547
rect 804 -2544 808 -2540
rect 830 -2566 834 -2562
rect 812 -2573 816 -2569
rect 856 -2558 860 -2554
rect 908 -2551 912 -2547
rect 838 -2595 842 -2591
rect 874 -2595 878 -2591
rect 934 -2566 938 -2562
rect 916 -2595 920 -2591
rect 952 -2595 956 -2591
rect 795 -2610 799 -2606
rect 821 -2610 825 -2606
rect 864 -2610 868 -2606
rect 899 -2610 903 -2606
rect 943 -2610 947 -2606
rect 960 -2610 964 -2606
rect 996 -2610 1000 -2606
rect 1017 -2610 1021 -2606
rect 1039 -2566 1043 -2562
rect 1039 -2617 1043 -2613
rect 1026 -2624 1030 -2620
rect 786 -2650 790 -2646
rect 803 -2650 807 -2646
rect 726 -2915 730 -2911
rect 752 -2915 756 -2911
rect 478 -2941 482 -2937
rect 495 -2941 499 -2937
rect 504 -2994 508 -2990
rect 742 -2994 746 -2990
rect 495 -3033 499 -3029
rect 487 -3100 491 -3096
rect 513 -3100 517 -3096
rect 530 -3100 534 -3096
rect 570 -3100 574 -3096
rect 591 -3100 595 -3096
rect 608 -3100 612 -3096
rect 648 -3100 652 -3096
rect 672 -3100 676 -3096
rect 709 -3100 713 -3096
rect 447 -3140 451 -3136
rect 478 -3133 482 -3129
rect 435 -3155 439 -3151
rect 496 -3126 500 -3122
rect 522 -3148 526 -3144
rect 504 -3155 508 -3151
rect 548 -3140 552 -3136
rect 600 -3133 604 -3129
rect 530 -3177 534 -3173
rect 566 -3177 570 -3173
rect 626 -3148 630 -3144
rect 608 -3177 612 -3173
rect 644 -3177 648 -3173
rect 718 -3138 722 -3134
rect 742 -3140 746 -3136
rect 812 -2703 816 -2699
rect 803 -2742 807 -2738
rect 795 -2809 799 -2805
rect 821 -2809 825 -2805
rect 838 -2809 842 -2805
rect 878 -2809 882 -2805
rect 899 -2809 903 -2805
rect 916 -2809 920 -2805
rect 956 -2809 960 -2805
rect 980 -2809 984 -2805
rect 1017 -2809 1021 -2805
rect 786 -2842 790 -2838
rect 804 -2835 808 -2831
rect 830 -2857 834 -2853
rect 812 -2864 816 -2860
rect 856 -2849 860 -2845
rect 908 -2842 912 -2838
rect 838 -2886 842 -2882
rect 874 -2886 878 -2882
rect 934 -2857 938 -2853
rect 916 -2886 920 -2882
rect 952 -2886 956 -2882
rect 795 -2901 799 -2897
rect 821 -2901 825 -2897
rect 864 -2901 868 -2897
rect 899 -2901 903 -2897
rect 943 -2901 947 -2897
rect 960 -2901 964 -2897
rect 996 -2901 1000 -2897
rect 1017 -2901 1021 -2897
rect 1039 -2857 1043 -2853
rect 1039 -2908 1043 -2904
rect 1026 -2915 1030 -2911
rect 786 -2941 790 -2937
rect 803 -2941 807 -2937
rect 812 -2994 816 -2990
rect 803 -3033 807 -3029
rect 795 -3100 799 -3096
rect 821 -3100 825 -3096
rect 838 -3100 842 -3096
rect 878 -3100 882 -3096
rect 899 -3100 903 -3096
rect 916 -3100 920 -3096
rect 956 -3100 960 -3096
rect 980 -3100 984 -3096
rect 1017 -3100 1021 -3096
rect 752 -3155 756 -3151
rect 786 -3133 790 -3129
rect 804 -3126 808 -3122
rect 830 -3148 834 -3144
rect 812 -3155 816 -3151
rect 856 -3140 860 -3136
rect 908 -3133 912 -3129
rect 838 -3177 842 -3173
rect 874 -3177 878 -3173
rect 934 -3148 938 -3144
rect 916 -3177 920 -3173
rect 952 -3177 956 -3173
rect -129 -3192 -125 -3188
rect -103 -3192 -99 -3188
rect -60 -3192 -56 -3188
rect -25 -3192 -21 -3188
rect 19 -3192 23 -3188
rect 36 -3192 40 -3188
rect 72 -3192 76 -3188
rect 93 -3192 97 -3188
rect 179 -3192 183 -3188
rect 205 -3192 209 -3188
rect 248 -3192 252 -3188
rect 283 -3192 287 -3188
rect 327 -3192 331 -3188
rect 344 -3192 348 -3188
rect 380 -3192 384 -3188
rect 401 -3192 405 -3188
rect 487 -3192 491 -3188
rect 513 -3192 517 -3188
rect 556 -3192 560 -3188
rect 591 -3192 595 -3188
rect 635 -3192 639 -3188
rect 652 -3192 656 -3188
rect 688 -3192 692 -3188
rect 709 -3192 713 -3188
rect 795 -3192 799 -3188
rect 821 -3192 825 -3188
rect 864 -3192 868 -3188
rect 899 -3192 903 -3188
rect 943 -3192 947 -3188
rect 960 -3192 964 -3188
rect 996 -3192 1000 -3188
rect 1017 -3192 1021 -3188
<< pad >>
rect -1295 -1024 -1291 -1020
rect -1051 -1024 -1047 -1020
rect -742 -1024 -738 -1020
rect -434 -1024 -430 -1020
rect -127 -1024 -123 -1020
rect 182 -1024 186 -1020
rect 490 -1024 494 -1020
rect 798 -1024 802 -1020
rect -1297 -1174 -1293 -1170
rect -1050 -1174 -1046 -1170
rect -742 -1174 -738 -1170
rect -434 -1174 -430 -1170
rect -126 -1174 -122 -1170
rect 182 -1174 186 -1170
rect 490 -1174 494 -1170
rect 798 -1174 802 -1170
rect -1051 -1317 -1047 -1313
rect -985 -1317 -981 -1313
rect -951 -1317 -947 -1313
rect -907 -1317 -903 -1313
rect -873 -1317 -869 -1313
rect -743 -1317 -739 -1313
rect -677 -1317 -673 -1313
rect -643 -1317 -639 -1313
rect -599 -1317 -595 -1313
rect -565 -1317 -561 -1313
rect -435 -1317 -431 -1313
rect -369 -1317 -365 -1313
rect -335 -1317 -331 -1313
rect -291 -1317 -287 -1313
rect -257 -1317 -253 -1313
rect -127 -1317 -123 -1313
rect -61 -1317 -57 -1313
rect -27 -1317 -23 -1313
rect 17 -1317 21 -1313
rect 51 -1317 55 -1313
rect 181 -1317 185 -1313
rect 247 -1317 251 -1313
rect 281 -1317 285 -1313
rect 325 -1317 329 -1313
rect 359 -1317 363 -1313
rect 489 -1317 493 -1313
rect 555 -1317 559 -1313
rect 589 -1317 593 -1313
rect 633 -1317 637 -1313
rect 667 -1317 671 -1313
rect -1009 -1324 -1005 -1320
rect -701 -1324 -697 -1320
rect -393 -1324 -389 -1320
rect -85 -1324 -81 -1320
rect 223 -1324 227 -1320
rect 531 -1324 535 -1320
rect -975 -1331 -971 -1327
rect -833 -1331 -829 -1327
rect -667 -1331 -663 -1327
rect -525 -1331 -521 -1327
rect -359 -1331 -355 -1327
rect -217 -1331 -213 -1327
rect -51 -1331 -47 -1327
rect 91 -1331 95 -1327
rect 257 -1331 261 -1327
rect 399 -1331 403 -1327
rect 565 -1331 569 -1327
rect 707 -1331 711 -1327
rect -1055 -1338 -1051 -1334
rect -1025 -1338 -1021 -1334
rect -907 -1338 -903 -1334
rect -747 -1338 -743 -1334
rect -717 -1338 -713 -1334
rect -599 -1338 -595 -1334
rect -439 -1338 -435 -1334
rect -409 -1338 -405 -1334
rect -291 -1338 -287 -1334
rect -131 -1338 -127 -1334
rect -101 -1338 -97 -1334
rect 17 -1338 21 -1334
rect 177 -1338 181 -1334
rect 207 -1338 211 -1334
rect 325 -1338 329 -1334
rect 485 -1338 489 -1334
rect 515 -1338 519 -1334
rect 633 -1338 637 -1334
rect -1169 -1347 -1165 -1343
rect -1029 -1346 -1025 -1342
rect -931 -1346 -927 -1342
rect -721 -1346 -717 -1342
rect -623 -1346 -619 -1342
rect -413 -1346 -409 -1342
rect -315 -1346 -311 -1342
rect -105 -1346 -101 -1342
rect -7 -1346 -3 -1342
rect 203 -1346 207 -1342
rect 301 -1346 305 -1342
rect 511 -1346 515 -1342
rect 609 -1346 613 -1342
rect 845 -1347 849 -1343
rect -1219 -1354 -1215 -1350
rect -1179 -1354 -1175 -1350
rect -1159 -1354 -1155 -1350
rect -1051 -1353 -1047 -1349
rect -903 -1353 -899 -1349
rect -743 -1353 -739 -1349
rect -595 -1353 -591 -1349
rect -435 -1353 -431 -1349
rect -287 -1353 -283 -1349
rect -127 -1353 -123 -1349
rect 21 -1353 25 -1349
rect 181 -1353 185 -1349
rect 329 -1353 333 -1349
rect 489 -1353 493 -1349
rect 637 -1353 641 -1349
rect 795 -1354 799 -1350
rect 835 -1354 839 -1350
rect 855 -1354 859 -1350
rect -1223 -1361 -1219 -1357
rect -1193 -1361 -1189 -1357
rect -1145 -1361 -1141 -1357
rect -1029 -1360 -1025 -1356
rect -921 -1360 -917 -1356
rect -887 -1360 -883 -1356
rect -721 -1360 -717 -1356
rect -613 -1360 -609 -1356
rect -579 -1360 -575 -1356
rect -413 -1360 -409 -1356
rect -305 -1360 -301 -1356
rect -271 -1360 -267 -1356
rect -105 -1360 -101 -1356
rect 3 -1360 7 -1356
rect 37 -1360 41 -1356
rect 203 -1360 207 -1356
rect 311 -1360 315 -1356
rect 345 -1360 349 -1356
rect 511 -1360 515 -1356
rect 619 -1360 623 -1356
rect 653 -1360 657 -1356
rect 791 -1361 795 -1357
rect 821 -1361 825 -1357
rect 869 -1361 873 -1357
rect -1055 -1367 -1051 -1363
rect -999 -1367 -995 -1363
rect -965 -1367 -961 -1363
rect -747 -1367 -743 -1363
rect -691 -1367 -687 -1363
rect -657 -1367 -653 -1363
rect -439 -1367 -435 -1363
rect -383 -1367 -379 -1363
rect -349 -1367 -345 -1363
rect -131 -1367 -127 -1363
rect -75 -1367 -71 -1363
rect -41 -1367 -37 -1363
rect 177 -1367 181 -1363
rect 233 -1367 237 -1363
rect 267 -1367 271 -1363
rect 485 -1367 489 -1363
rect 541 -1367 545 -1363
rect 575 -1367 579 -1363
rect -1297 -1495 -1293 -1491
rect -1050 -1495 -1046 -1491
rect -742 -1495 -738 -1491
rect -434 -1495 -430 -1491
rect -126 -1495 -122 -1491
rect 182 -1495 186 -1491
rect 490 -1495 494 -1491
rect 798 -1495 802 -1491
rect -1051 -1633 -1047 -1629
rect -985 -1633 -981 -1629
rect -951 -1633 -947 -1629
rect -907 -1633 -903 -1629
rect -873 -1633 -869 -1629
rect -743 -1633 -739 -1629
rect -677 -1633 -673 -1629
rect -643 -1633 -639 -1629
rect -599 -1633 -595 -1629
rect -565 -1633 -561 -1629
rect -435 -1633 -431 -1629
rect -369 -1633 -365 -1629
rect -335 -1633 -331 -1629
rect -291 -1633 -287 -1629
rect -257 -1633 -253 -1629
rect -127 -1633 -123 -1629
rect -61 -1633 -57 -1629
rect -27 -1633 -23 -1629
rect 17 -1633 21 -1629
rect 51 -1633 55 -1629
rect 181 -1633 185 -1629
rect 247 -1633 251 -1629
rect 281 -1633 285 -1629
rect 325 -1633 329 -1629
rect 359 -1633 363 -1629
rect 489 -1633 493 -1629
rect 555 -1633 559 -1629
rect 589 -1633 593 -1629
rect 633 -1633 637 -1629
rect 667 -1633 671 -1629
rect 797 -1633 801 -1629
rect 863 -1633 867 -1629
rect 897 -1633 901 -1629
rect 941 -1633 945 -1629
rect 975 -1633 979 -1629
rect -1009 -1640 -1005 -1636
rect -701 -1640 -697 -1636
rect -393 -1640 -389 -1636
rect -85 -1640 -81 -1636
rect 223 -1640 227 -1636
rect 531 -1640 535 -1636
rect 839 -1640 843 -1636
rect -975 -1647 -971 -1643
rect -833 -1647 -829 -1643
rect -667 -1647 -663 -1643
rect -525 -1647 -521 -1643
rect -359 -1647 -355 -1643
rect -217 -1647 -213 -1643
rect -51 -1647 -47 -1643
rect 91 -1647 95 -1643
rect 257 -1647 261 -1643
rect 399 -1647 403 -1643
rect 565 -1647 569 -1643
rect 707 -1647 711 -1643
rect 873 -1647 877 -1643
rect 1015 -1647 1019 -1643
rect -1055 -1654 -1051 -1650
rect -1025 -1654 -1021 -1650
rect -907 -1654 -903 -1650
rect -747 -1654 -743 -1650
rect -717 -1654 -713 -1650
rect -599 -1654 -595 -1650
rect -439 -1654 -435 -1650
rect -409 -1654 -405 -1650
rect -291 -1654 -287 -1650
rect -131 -1654 -127 -1650
rect -101 -1654 -97 -1650
rect 17 -1654 21 -1650
rect 177 -1654 181 -1650
rect 207 -1654 211 -1650
rect 325 -1654 329 -1650
rect 485 -1654 489 -1650
rect 515 -1654 519 -1650
rect 633 -1654 637 -1650
rect 793 -1654 797 -1650
rect 823 -1654 827 -1650
rect 941 -1654 945 -1650
rect -1173 -1663 -1169 -1659
rect -1029 -1662 -1025 -1658
rect -931 -1662 -927 -1658
rect -721 -1662 -717 -1658
rect -623 -1662 -619 -1658
rect -413 -1662 -409 -1658
rect -315 -1662 -311 -1658
rect -105 -1662 -101 -1658
rect -7 -1662 -3 -1658
rect 203 -1662 207 -1658
rect 301 -1662 305 -1658
rect 511 -1662 515 -1658
rect 609 -1662 613 -1658
rect 819 -1662 823 -1658
rect 917 -1662 921 -1658
rect -1223 -1670 -1219 -1666
rect -1183 -1670 -1179 -1666
rect -1163 -1670 -1159 -1666
rect -1051 -1669 -1047 -1665
rect -903 -1669 -899 -1665
rect -743 -1669 -739 -1665
rect -595 -1669 -591 -1665
rect -435 -1669 -431 -1665
rect -287 -1669 -283 -1665
rect -127 -1669 -123 -1665
rect 21 -1669 25 -1665
rect 181 -1669 185 -1665
rect 329 -1669 333 -1665
rect 489 -1669 493 -1665
rect 637 -1669 641 -1665
rect 797 -1669 801 -1665
rect 945 -1669 949 -1665
rect -1227 -1677 -1223 -1673
rect -1197 -1677 -1193 -1673
rect -1149 -1677 -1145 -1673
rect -1029 -1676 -1025 -1672
rect -921 -1676 -917 -1672
rect -887 -1676 -883 -1672
rect -721 -1676 -717 -1672
rect -613 -1676 -609 -1672
rect -579 -1676 -575 -1672
rect -413 -1676 -409 -1672
rect -305 -1676 -301 -1672
rect -271 -1676 -267 -1672
rect -105 -1676 -101 -1672
rect 3 -1676 7 -1672
rect 37 -1676 41 -1672
rect 203 -1676 207 -1672
rect 311 -1676 315 -1672
rect 345 -1676 349 -1672
rect 511 -1676 515 -1672
rect 619 -1676 623 -1672
rect 653 -1676 657 -1672
rect 819 -1676 823 -1672
rect 927 -1676 931 -1672
rect 961 -1676 965 -1672
rect -1055 -1683 -1051 -1679
rect -999 -1683 -995 -1679
rect -965 -1683 -961 -1679
rect -747 -1683 -743 -1679
rect -691 -1683 -687 -1679
rect -657 -1683 -653 -1679
rect -439 -1683 -435 -1679
rect -383 -1683 -379 -1679
rect -349 -1683 -345 -1679
rect -131 -1683 -127 -1679
rect -75 -1683 -71 -1679
rect -41 -1683 -37 -1679
rect 177 -1683 181 -1679
rect 233 -1683 237 -1679
rect 267 -1683 271 -1679
rect 485 -1683 489 -1679
rect 541 -1683 545 -1679
rect 575 -1683 579 -1679
rect 793 -1683 797 -1679
rect 849 -1683 853 -1679
rect 883 -1683 887 -1679
rect -1297 -1786 -1293 -1782
rect -1050 -1786 -1046 -1782
rect -742 -1786 -738 -1782
rect -434 -1786 -430 -1782
rect -126 -1786 -122 -1782
rect 182 -1786 186 -1782
rect 490 -1786 494 -1782
rect 798 -1786 802 -1782
rect -1051 -1924 -1047 -1920
rect -985 -1924 -981 -1920
rect -951 -1924 -947 -1920
rect -907 -1924 -903 -1920
rect -873 -1924 -869 -1920
rect -743 -1924 -739 -1920
rect -677 -1924 -673 -1920
rect -643 -1924 -639 -1920
rect -599 -1924 -595 -1920
rect -565 -1924 -561 -1920
rect -435 -1924 -431 -1920
rect -369 -1924 -365 -1920
rect -335 -1924 -331 -1920
rect -291 -1924 -287 -1920
rect -257 -1924 -253 -1920
rect -127 -1924 -123 -1920
rect -61 -1924 -57 -1920
rect -27 -1924 -23 -1920
rect 17 -1924 21 -1920
rect 51 -1924 55 -1920
rect 181 -1924 185 -1920
rect 247 -1924 251 -1920
rect 281 -1924 285 -1920
rect 325 -1924 329 -1920
rect 359 -1924 363 -1920
rect 489 -1924 493 -1920
rect 555 -1924 559 -1920
rect 589 -1924 593 -1920
rect 633 -1924 637 -1920
rect 667 -1924 671 -1920
rect 797 -1924 801 -1920
rect 863 -1924 867 -1920
rect 897 -1924 901 -1920
rect 941 -1924 945 -1920
rect 975 -1924 979 -1920
rect -1009 -1931 -1005 -1927
rect -701 -1931 -697 -1927
rect -393 -1931 -389 -1927
rect -85 -1931 -81 -1927
rect 223 -1931 227 -1927
rect 531 -1931 535 -1927
rect 839 -1931 843 -1927
rect -975 -1938 -971 -1934
rect -833 -1938 -829 -1934
rect -667 -1938 -663 -1934
rect -525 -1938 -521 -1934
rect -359 -1938 -355 -1934
rect -217 -1938 -213 -1934
rect -51 -1938 -47 -1934
rect 91 -1938 95 -1934
rect 257 -1938 261 -1934
rect 399 -1938 403 -1934
rect 565 -1938 569 -1934
rect 707 -1938 711 -1934
rect 873 -1938 877 -1934
rect 1015 -1938 1019 -1934
rect -1055 -1945 -1051 -1941
rect -1025 -1945 -1021 -1941
rect -907 -1945 -903 -1941
rect -747 -1945 -743 -1941
rect -717 -1945 -713 -1941
rect -599 -1945 -595 -1941
rect -439 -1945 -435 -1941
rect -409 -1945 -405 -1941
rect -291 -1945 -287 -1941
rect -131 -1945 -127 -1941
rect -101 -1945 -97 -1941
rect 17 -1945 21 -1941
rect 177 -1945 181 -1941
rect 207 -1945 211 -1941
rect 325 -1945 329 -1941
rect 485 -1945 489 -1941
rect 515 -1945 519 -1941
rect 633 -1945 637 -1941
rect 793 -1945 797 -1941
rect 823 -1945 827 -1941
rect 941 -1945 945 -1941
rect -1173 -1954 -1169 -1950
rect -1029 -1953 -1025 -1949
rect -931 -1953 -927 -1949
rect -721 -1953 -717 -1949
rect -623 -1953 -619 -1949
rect -413 -1953 -409 -1949
rect -315 -1953 -311 -1949
rect -105 -1953 -101 -1949
rect -7 -1953 -3 -1949
rect 203 -1953 207 -1949
rect 301 -1953 305 -1949
rect 511 -1953 515 -1949
rect 609 -1953 613 -1949
rect 819 -1953 823 -1949
rect 917 -1953 921 -1949
rect -1223 -1961 -1219 -1957
rect -1183 -1961 -1179 -1957
rect -1163 -1961 -1159 -1957
rect -1051 -1960 -1047 -1956
rect -903 -1960 -899 -1956
rect -743 -1960 -739 -1956
rect -595 -1960 -591 -1956
rect -435 -1960 -431 -1956
rect -287 -1960 -283 -1956
rect -127 -1960 -123 -1956
rect 21 -1960 25 -1956
rect 181 -1960 185 -1956
rect 329 -1960 333 -1956
rect 489 -1960 493 -1956
rect 637 -1960 641 -1956
rect 797 -1960 801 -1956
rect 945 -1960 949 -1956
rect -1227 -1968 -1223 -1964
rect -1197 -1968 -1193 -1964
rect -1149 -1968 -1145 -1964
rect -1029 -1967 -1025 -1963
rect -921 -1967 -917 -1963
rect -887 -1967 -883 -1963
rect -721 -1967 -717 -1963
rect -613 -1967 -609 -1963
rect -579 -1967 -575 -1963
rect -413 -1967 -409 -1963
rect -305 -1967 -301 -1963
rect -271 -1967 -267 -1963
rect -105 -1967 -101 -1963
rect 3 -1967 7 -1963
rect 37 -1967 41 -1963
rect 203 -1967 207 -1963
rect 311 -1967 315 -1963
rect 345 -1967 349 -1963
rect 511 -1967 515 -1963
rect 619 -1967 623 -1963
rect 653 -1967 657 -1963
rect 819 -1967 823 -1963
rect 927 -1967 931 -1963
rect 961 -1967 965 -1963
rect -1055 -1974 -1051 -1970
rect -999 -1974 -995 -1970
rect -965 -1974 -961 -1970
rect -747 -1974 -743 -1970
rect -691 -1974 -687 -1970
rect -657 -1974 -653 -1970
rect -439 -1974 -435 -1970
rect -383 -1974 -379 -1970
rect -349 -1974 -345 -1970
rect -131 -1974 -127 -1970
rect -75 -1974 -71 -1970
rect -41 -1974 -37 -1970
rect 177 -1974 181 -1970
rect 233 -1974 237 -1970
rect 267 -1974 271 -1970
rect 485 -1974 489 -1970
rect 541 -1974 545 -1970
rect 575 -1974 579 -1970
rect 793 -1974 797 -1970
rect 849 -1974 853 -1970
rect 883 -1974 887 -1970
rect -1297 -2108 -1293 -2104
rect -1050 -2108 -1046 -2104
rect -742 -2108 -738 -2104
rect -434 -2108 -430 -2104
rect -126 -2108 -122 -2104
rect 182 -2108 186 -2104
rect 490 -2108 494 -2104
rect 798 -2108 802 -2104
rect -1051 -2246 -1047 -2242
rect -985 -2246 -981 -2242
rect -951 -2246 -947 -2242
rect -907 -2246 -903 -2242
rect -873 -2246 -869 -2242
rect -743 -2246 -739 -2242
rect -677 -2246 -673 -2242
rect -643 -2246 -639 -2242
rect -599 -2246 -595 -2242
rect -565 -2246 -561 -2242
rect -435 -2246 -431 -2242
rect -369 -2246 -365 -2242
rect -335 -2246 -331 -2242
rect -291 -2246 -287 -2242
rect -257 -2246 -253 -2242
rect -127 -2246 -123 -2242
rect -61 -2246 -57 -2242
rect -27 -2246 -23 -2242
rect 17 -2246 21 -2242
rect 51 -2246 55 -2242
rect 181 -2246 185 -2242
rect 247 -2246 251 -2242
rect 281 -2246 285 -2242
rect 325 -2246 329 -2242
rect 359 -2246 363 -2242
rect 489 -2246 493 -2242
rect 555 -2246 559 -2242
rect 589 -2246 593 -2242
rect 633 -2246 637 -2242
rect 667 -2246 671 -2242
rect 797 -2246 801 -2242
rect 863 -2246 867 -2242
rect 897 -2246 901 -2242
rect 941 -2246 945 -2242
rect 975 -2246 979 -2242
rect -1009 -2253 -1005 -2249
rect -701 -2253 -697 -2249
rect -393 -2253 -389 -2249
rect -85 -2253 -81 -2249
rect 223 -2253 227 -2249
rect 531 -2253 535 -2249
rect 839 -2253 843 -2249
rect -975 -2260 -971 -2256
rect -833 -2260 -829 -2256
rect -667 -2260 -663 -2256
rect -525 -2260 -521 -2256
rect -359 -2260 -355 -2256
rect -217 -2260 -213 -2256
rect -51 -2260 -47 -2256
rect 91 -2260 95 -2256
rect 257 -2260 261 -2256
rect 399 -2260 403 -2256
rect 565 -2260 569 -2256
rect 707 -2260 711 -2256
rect 873 -2260 877 -2256
rect 1015 -2260 1019 -2256
rect -1055 -2267 -1051 -2263
rect -1025 -2267 -1021 -2263
rect -907 -2267 -903 -2263
rect -747 -2267 -743 -2263
rect -717 -2267 -713 -2263
rect -599 -2267 -595 -2263
rect -439 -2267 -435 -2263
rect -409 -2267 -405 -2263
rect -291 -2267 -287 -2263
rect -131 -2267 -127 -2263
rect -101 -2267 -97 -2263
rect 17 -2267 21 -2263
rect 177 -2267 181 -2263
rect 207 -2267 211 -2263
rect 325 -2267 329 -2263
rect 485 -2267 489 -2263
rect 515 -2267 519 -2263
rect 633 -2267 637 -2263
rect 793 -2267 797 -2263
rect 823 -2267 827 -2263
rect 941 -2267 945 -2263
rect -1173 -2276 -1169 -2272
rect -1029 -2275 -1025 -2271
rect -931 -2275 -927 -2271
rect -721 -2275 -717 -2271
rect -623 -2275 -619 -2271
rect -413 -2275 -409 -2271
rect -315 -2275 -311 -2271
rect -105 -2275 -101 -2271
rect -7 -2275 -3 -2271
rect 203 -2275 207 -2271
rect 301 -2275 305 -2271
rect 511 -2275 515 -2271
rect 609 -2275 613 -2271
rect 819 -2275 823 -2271
rect 917 -2275 921 -2271
rect -1223 -2283 -1219 -2279
rect -1183 -2283 -1179 -2279
rect -1163 -2283 -1159 -2279
rect -1051 -2282 -1047 -2278
rect -903 -2282 -899 -2278
rect -743 -2282 -739 -2278
rect -595 -2282 -591 -2278
rect -435 -2282 -431 -2278
rect -287 -2282 -283 -2278
rect -127 -2282 -123 -2278
rect 21 -2282 25 -2278
rect 181 -2282 185 -2278
rect 329 -2282 333 -2278
rect 489 -2282 493 -2278
rect 637 -2282 641 -2278
rect 797 -2282 801 -2278
rect 945 -2282 949 -2278
rect -1227 -2290 -1223 -2286
rect -1197 -2290 -1193 -2286
rect -1149 -2290 -1145 -2286
rect -1029 -2289 -1025 -2285
rect -921 -2289 -917 -2285
rect -887 -2289 -883 -2285
rect -721 -2289 -717 -2285
rect -613 -2289 -609 -2285
rect -579 -2289 -575 -2285
rect -413 -2289 -409 -2285
rect -305 -2289 -301 -2285
rect -271 -2289 -267 -2285
rect -105 -2289 -101 -2285
rect 3 -2289 7 -2285
rect 37 -2289 41 -2285
rect 203 -2289 207 -2285
rect 311 -2289 315 -2285
rect 345 -2289 349 -2285
rect 511 -2289 515 -2285
rect 619 -2289 623 -2285
rect 653 -2289 657 -2285
rect 819 -2289 823 -2285
rect 927 -2289 931 -2285
rect 961 -2289 965 -2285
rect -1055 -2296 -1051 -2292
rect -999 -2296 -995 -2292
rect -965 -2296 -961 -2292
rect -747 -2296 -743 -2292
rect -691 -2296 -687 -2292
rect -657 -2296 -653 -2292
rect -439 -2296 -435 -2292
rect -383 -2296 -379 -2292
rect -349 -2296 -345 -2292
rect -131 -2296 -127 -2292
rect -75 -2296 -71 -2292
rect -41 -2296 -37 -2292
rect 177 -2296 181 -2292
rect 233 -2296 237 -2292
rect 267 -2296 271 -2292
rect 485 -2296 489 -2292
rect 541 -2296 545 -2292
rect 575 -2296 579 -2292
rect 793 -2296 797 -2292
rect 849 -2296 853 -2292
rect 883 -2296 887 -2292
rect -1297 -2399 -1293 -2395
rect -1050 -2399 -1046 -2395
rect -742 -2399 -738 -2395
rect -434 -2399 -430 -2395
rect -126 -2399 -122 -2395
rect 182 -2399 186 -2395
rect 490 -2399 494 -2395
rect 798 -2399 802 -2395
rect -1051 -2537 -1047 -2533
rect -985 -2537 -981 -2533
rect -951 -2537 -947 -2533
rect -907 -2537 -903 -2533
rect -873 -2537 -869 -2533
rect -743 -2537 -739 -2533
rect -677 -2537 -673 -2533
rect -643 -2537 -639 -2533
rect -599 -2537 -595 -2533
rect -565 -2537 -561 -2533
rect -435 -2537 -431 -2533
rect -369 -2537 -365 -2533
rect -335 -2537 -331 -2533
rect -291 -2537 -287 -2533
rect -257 -2537 -253 -2533
rect -127 -2537 -123 -2533
rect -61 -2537 -57 -2533
rect -27 -2537 -23 -2533
rect 17 -2537 21 -2533
rect 51 -2537 55 -2533
rect 181 -2537 185 -2533
rect 247 -2537 251 -2533
rect 281 -2537 285 -2533
rect 325 -2537 329 -2533
rect 359 -2537 363 -2533
rect 489 -2537 493 -2533
rect 555 -2537 559 -2533
rect 589 -2537 593 -2533
rect 633 -2537 637 -2533
rect 667 -2537 671 -2533
rect 797 -2537 801 -2533
rect 863 -2537 867 -2533
rect 897 -2537 901 -2533
rect 941 -2537 945 -2533
rect 975 -2537 979 -2533
rect -1009 -2544 -1005 -2540
rect -701 -2544 -697 -2540
rect -393 -2544 -389 -2540
rect -85 -2544 -81 -2540
rect 223 -2544 227 -2540
rect 531 -2544 535 -2540
rect 839 -2544 843 -2540
rect -975 -2551 -971 -2547
rect -833 -2551 -829 -2547
rect -667 -2551 -663 -2547
rect -525 -2551 -521 -2547
rect -359 -2551 -355 -2547
rect -217 -2551 -213 -2547
rect -51 -2551 -47 -2547
rect 91 -2551 95 -2547
rect 257 -2551 261 -2547
rect 399 -2551 403 -2547
rect 565 -2551 569 -2547
rect 707 -2551 711 -2547
rect 873 -2551 877 -2547
rect 1015 -2551 1019 -2547
rect -1055 -2558 -1051 -2554
rect -1025 -2558 -1021 -2554
rect -907 -2558 -903 -2554
rect -747 -2558 -743 -2554
rect -717 -2558 -713 -2554
rect -599 -2558 -595 -2554
rect -439 -2558 -435 -2554
rect -409 -2558 -405 -2554
rect -291 -2558 -287 -2554
rect -131 -2558 -127 -2554
rect -101 -2558 -97 -2554
rect 17 -2558 21 -2554
rect 177 -2558 181 -2554
rect 207 -2558 211 -2554
rect 325 -2558 329 -2554
rect 485 -2558 489 -2554
rect 515 -2558 519 -2554
rect 633 -2558 637 -2554
rect 793 -2558 797 -2554
rect 823 -2558 827 -2554
rect 941 -2558 945 -2554
rect -1173 -2567 -1169 -2563
rect -1029 -2566 -1025 -2562
rect -931 -2566 -927 -2562
rect -721 -2566 -717 -2562
rect -623 -2566 -619 -2562
rect -413 -2566 -409 -2562
rect -315 -2566 -311 -2562
rect -105 -2566 -101 -2562
rect -7 -2566 -3 -2562
rect 203 -2566 207 -2562
rect 301 -2566 305 -2562
rect 511 -2566 515 -2562
rect 609 -2566 613 -2562
rect 819 -2566 823 -2562
rect 917 -2566 921 -2562
rect -1223 -2574 -1219 -2570
rect -1183 -2574 -1179 -2570
rect -1163 -2574 -1159 -2570
rect -1051 -2573 -1047 -2569
rect -903 -2573 -899 -2569
rect -743 -2573 -739 -2569
rect -595 -2573 -591 -2569
rect -435 -2573 -431 -2569
rect -287 -2573 -283 -2569
rect -127 -2573 -123 -2569
rect 21 -2573 25 -2569
rect 181 -2573 185 -2569
rect 329 -2573 333 -2569
rect 489 -2573 493 -2569
rect 637 -2573 641 -2569
rect 797 -2573 801 -2569
rect 945 -2573 949 -2569
rect -1227 -2581 -1223 -2577
rect -1197 -2581 -1193 -2577
rect -1149 -2581 -1145 -2577
rect -1029 -2580 -1025 -2576
rect -921 -2580 -917 -2576
rect -887 -2580 -883 -2576
rect -721 -2580 -717 -2576
rect -613 -2580 -609 -2576
rect -579 -2580 -575 -2576
rect -413 -2580 -409 -2576
rect -305 -2580 -301 -2576
rect -271 -2580 -267 -2576
rect -105 -2580 -101 -2576
rect 3 -2580 7 -2576
rect 37 -2580 41 -2576
rect 203 -2580 207 -2576
rect 311 -2580 315 -2576
rect 345 -2580 349 -2576
rect 511 -2580 515 -2576
rect 619 -2580 623 -2576
rect 653 -2580 657 -2576
rect 819 -2580 823 -2576
rect 927 -2580 931 -2576
rect 961 -2580 965 -2576
rect -1055 -2587 -1051 -2583
rect -999 -2587 -995 -2583
rect -965 -2587 -961 -2583
rect -747 -2587 -743 -2583
rect -691 -2587 -687 -2583
rect -657 -2587 -653 -2583
rect -439 -2587 -435 -2583
rect -383 -2587 -379 -2583
rect -349 -2587 -345 -2583
rect -131 -2587 -127 -2583
rect -75 -2587 -71 -2583
rect -41 -2587 -37 -2583
rect 177 -2587 181 -2583
rect 233 -2587 237 -2583
rect 267 -2587 271 -2583
rect 485 -2587 489 -2583
rect 541 -2587 545 -2583
rect 575 -2587 579 -2583
rect 793 -2587 797 -2583
rect 849 -2587 853 -2583
rect 883 -2587 887 -2583
rect -1297 -2690 -1293 -2686
rect -1050 -2690 -1046 -2686
rect -742 -2690 -738 -2686
rect -434 -2690 -430 -2686
rect -126 -2690 -122 -2686
rect 182 -2690 186 -2686
rect 490 -2690 494 -2686
rect 798 -2690 802 -2686
rect -1051 -2828 -1047 -2824
rect -985 -2828 -981 -2824
rect -951 -2828 -947 -2824
rect -907 -2828 -903 -2824
rect -873 -2828 -869 -2824
rect -743 -2828 -739 -2824
rect -677 -2828 -673 -2824
rect -643 -2828 -639 -2824
rect -599 -2828 -595 -2824
rect -565 -2828 -561 -2824
rect -435 -2828 -431 -2824
rect -369 -2828 -365 -2824
rect -335 -2828 -331 -2824
rect -291 -2828 -287 -2824
rect -257 -2828 -253 -2824
rect -127 -2828 -123 -2824
rect -61 -2828 -57 -2824
rect -27 -2828 -23 -2824
rect 17 -2828 21 -2824
rect 51 -2828 55 -2824
rect 181 -2828 185 -2824
rect 247 -2828 251 -2824
rect 281 -2828 285 -2824
rect 325 -2828 329 -2824
rect 359 -2828 363 -2824
rect 489 -2828 493 -2824
rect 555 -2828 559 -2824
rect 589 -2828 593 -2824
rect 633 -2828 637 -2824
rect 667 -2828 671 -2824
rect 797 -2828 801 -2824
rect 863 -2828 867 -2824
rect 897 -2828 901 -2824
rect 941 -2828 945 -2824
rect 975 -2828 979 -2824
rect -1009 -2835 -1005 -2831
rect -701 -2835 -697 -2831
rect -393 -2835 -389 -2831
rect -85 -2835 -81 -2831
rect 223 -2835 227 -2831
rect 531 -2835 535 -2831
rect 839 -2835 843 -2831
rect -975 -2842 -971 -2838
rect -833 -2842 -829 -2838
rect -667 -2842 -663 -2838
rect -525 -2842 -521 -2838
rect -359 -2842 -355 -2838
rect -217 -2842 -213 -2838
rect -51 -2842 -47 -2838
rect 91 -2842 95 -2838
rect 257 -2842 261 -2838
rect 399 -2842 403 -2838
rect 565 -2842 569 -2838
rect 707 -2842 711 -2838
rect 873 -2842 877 -2838
rect 1015 -2842 1019 -2838
rect -1055 -2849 -1051 -2845
rect -1025 -2849 -1021 -2845
rect -907 -2849 -903 -2845
rect -747 -2849 -743 -2845
rect -717 -2849 -713 -2845
rect -599 -2849 -595 -2845
rect -439 -2849 -435 -2845
rect -409 -2849 -405 -2845
rect -291 -2849 -287 -2845
rect -131 -2849 -127 -2845
rect -101 -2849 -97 -2845
rect 17 -2849 21 -2845
rect 177 -2849 181 -2845
rect 207 -2849 211 -2845
rect 325 -2849 329 -2845
rect 485 -2849 489 -2845
rect 515 -2849 519 -2845
rect 633 -2849 637 -2845
rect 793 -2849 797 -2845
rect 823 -2849 827 -2845
rect 941 -2849 945 -2845
rect -1173 -2858 -1169 -2854
rect -1029 -2857 -1025 -2853
rect -931 -2857 -927 -2853
rect -721 -2857 -717 -2853
rect -623 -2857 -619 -2853
rect -413 -2857 -409 -2853
rect -315 -2857 -311 -2853
rect -105 -2857 -101 -2853
rect -7 -2857 -3 -2853
rect 203 -2857 207 -2853
rect 301 -2857 305 -2853
rect 511 -2857 515 -2853
rect 609 -2857 613 -2853
rect 819 -2857 823 -2853
rect 917 -2857 921 -2853
rect -1223 -2865 -1219 -2861
rect -1183 -2865 -1179 -2861
rect -1163 -2865 -1159 -2861
rect -1051 -2864 -1047 -2860
rect -903 -2864 -899 -2860
rect -743 -2864 -739 -2860
rect -595 -2864 -591 -2860
rect -435 -2864 -431 -2860
rect -287 -2864 -283 -2860
rect -127 -2864 -123 -2860
rect 21 -2864 25 -2860
rect 181 -2864 185 -2860
rect 329 -2864 333 -2860
rect 489 -2864 493 -2860
rect 637 -2864 641 -2860
rect 797 -2864 801 -2860
rect 945 -2864 949 -2860
rect -1227 -2872 -1223 -2868
rect -1197 -2872 -1193 -2868
rect -1149 -2872 -1145 -2868
rect -1029 -2871 -1025 -2867
rect -921 -2871 -917 -2867
rect -887 -2871 -883 -2867
rect -721 -2871 -717 -2867
rect -613 -2871 -609 -2867
rect -579 -2871 -575 -2867
rect -413 -2871 -409 -2867
rect -305 -2871 -301 -2867
rect -271 -2871 -267 -2867
rect -105 -2871 -101 -2867
rect 3 -2871 7 -2867
rect 37 -2871 41 -2867
rect 203 -2871 207 -2867
rect 311 -2871 315 -2867
rect 345 -2871 349 -2867
rect 511 -2871 515 -2867
rect 619 -2871 623 -2867
rect 653 -2871 657 -2867
rect 819 -2871 823 -2867
rect 927 -2871 931 -2867
rect 961 -2871 965 -2867
rect -1055 -2878 -1051 -2874
rect -999 -2878 -995 -2874
rect -965 -2878 -961 -2874
rect -747 -2878 -743 -2874
rect -691 -2878 -687 -2874
rect -657 -2878 -653 -2874
rect -439 -2878 -435 -2874
rect -383 -2878 -379 -2874
rect -349 -2878 -345 -2874
rect -131 -2878 -127 -2874
rect -75 -2878 -71 -2874
rect -41 -2878 -37 -2874
rect 177 -2878 181 -2874
rect 233 -2878 237 -2874
rect 267 -2878 271 -2874
rect 485 -2878 489 -2874
rect 541 -2878 545 -2874
rect 575 -2878 579 -2874
rect 793 -2878 797 -2874
rect 849 -2878 853 -2874
rect 883 -2878 887 -2874
rect -1297 -2981 -1293 -2977
rect -1050 -2981 -1046 -2977
rect -742 -2981 -738 -2977
rect -434 -2981 -430 -2977
rect -126 -2981 -122 -2977
rect 182 -2981 186 -2977
rect 490 -2981 494 -2977
rect 798 -2981 802 -2977
rect -1051 -3119 -1047 -3115
rect -985 -3119 -981 -3115
rect -951 -3119 -947 -3115
rect -907 -3119 -903 -3115
rect -873 -3119 -869 -3115
rect -743 -3119 -739 -3115
rect -677 -3119 -673 -3115
rect -643 -3119 -639 -3115
rect -599 -3119 -595 -3115
rect -565 -3119 -561 -3115
rect -435 -3119 -431 -3115
rect -369 -3119 -365 -3115
rect -335 -3119 -331 -3115
rect -291 -3119 -287 -3115
rect -257 -3119 -253 -3115
rect -127 -3119 -123 -3115
rect -61 -3119 -57 -3115
rect -27 -3119 -23 -3115
rect 17 -3119 21 -3115
rect 51 -3119 55 -3115
rect 181 -3119 185 -3115
rect 247 -3119 251 -3115
rect 281 -3119 285 -3115
rect 325 -3119 329 -3115
rect 359 -3119 363 -3115
rect 489 -3119 493 -3115
rect 555 -3119 559 -3115
rect 589 -3119 593 -3115
rect 633 -3119 637 -3115
rect 667 -3119 671 -3115
rect 797 -3119 801 -3115
rect 863 -3119 867 -3115
rect 897 -3119 901 -3115
rect 941 -3119 945 -3115
rect 975 -3119 979 -3115
rect -1009 -3126 -1005 -3122
rect -701 -3126 -697 -3122
rect -393 -3126 -389 -3122
rect -85 -3126 -81 -3122
rect 223 -3126 227 -3122
rect 531 -3126 535 -3122
rect 839 -3126 843 -3122
rect -975 -3133 -971 -3129
rect -833 -3133 -829 -3129
rect -667 -3133 -663 -3129
rect -525 -3133 -521 -3129
rect -359 -3133 -355 -3129
rect -217 -3133 -213 -3129
rect -51 -3133 -47 -3129
rect 91 -3133 95 -3129
rect 257 -3133 261 -3129
rect 399 -3133 403 -3129
rect 565 -3133 569 -3129
rect 707 -3133 711 -3129
rect 873 -3133 877 -3129
rect 1015 -3133 1019 -3129
rect -1055 -3140 -1051 -3136
rect -1025 -3140 -1021 -3136
rect -907 -3140 -903 -3136
rect -747 -3140 -743 -3136
rect -717 -3140 -713 -3136
rect -599 -3140 -595 -3136
rect -439 -3140 -435 -3136
rect -409 -3140 -405 -3136
rect -291 -3140 -287 -3136
rect -131 -3140 -127 -3136
rect -101 -3140 -97 -3136
rect 17 -3140 21 -3136
rect 177 -3140 181 -3136
rect 207 -3140 211 -3136
rect 325 -3140 329 -3136
rect 485 -3140 489 -3136
rect 515 -3140 519 -3136
rect 633 -3140 637 -3136
rect 793 -3140 797 -3136
rect 823 -3140 827 -3136
rect 941 -3140 945 -3136
rect -1173 -3149 -1169 -3145
rect -1029 -3148 -1025 -3144
rect -931 -3148 -927 -3144
rect -721 -3148 -717 -3144
rect -623 -3148 -619 -3144
rect -413 -3148 -409 -3144
rect -315 -3148 -311 -3144
rect -105 -3148 -101 -3144
rect -7 -3148 -3 -3144
rect 203 -3148 207 -3144
rect 301 -3148 305 -3144
rect 511 -3148 515 -3144
rect 609 -3148 613 -3144
rect 819 -3148 823 -3144
rect 917 -3148 921 -3144
rect -1223 -3156 -1219 -3152
rect -1183 -3156 -1179 -3152
rect -1163 -3156 -1159 -3152
rect -1051 -3155 -1047 -3151
rect -903 -3155 -899 -3151
rect -743 -3155 -739 -3151
rect -595 -3155 -591 -3151
rect -435 -3155 -431 -3151
rect -287 -3155 -283 -3151
rect -127 -3155 -123 -3151
rect 21 -3155 25 -3151
rect 181 -3155 185 -3151
rect 329 -3155 333 -3151
rect 489 -3155 493 -3151
rect 637 -3155 641 -3151
rect 797 -3155 801 -3151
rect 945 -3155 949 -3151
rect -1227 -3163 -1223 -3159
rect -1197 -3163 -1193 -3159
rect -1149 -3163 -1145 -3159
rect -1029 -3162 -1025 -3158
rect -921 -3162 -917 -3158
rect -887 -3162 -883 -3158
rect -721 -3162 -717 -3158
rect -613 -3162 -609 -3158
rect -579 -3162 -575 -3158
rect -413 -3162 -409 -3158
rect -305 -3162 -301 -3158
rect -271 -3162 -267 -3158
rect -105 -3162 -101 -3158
rect 3 -3162 7 -3158
rect 37 -3162 41 -3158
rect 203 -3162 207 -3158
rect 311 -3162 315 -3158
rect 345 -3162 349 -3158
rect 511 -3162 515 -3158
rect 619 -3162 623 -3158
rect 653 -3162 657 -3158
rect 819 -3162 823 -3158
rect 927 -3162 931 -3158
rect 961 -3162 965 -3158
rect -1055 -3169 -1051 -3165
rect -999 -3169 -995 -3165
rect -965 -3169 -961 -3165
rect -747 -3169 -743 -3165
rect -691 -3169 -687 -3165
rect -657 -3169 -653 -3165
rect -439 -3169 -435 -3165
rect -383 -3169 -379 -3165
rect -349 -3169 -345 -3165
rect -131 -3169 -127 -3165
rect -75 -3169 -71 -3165
rect -41 -3169 -37 -3165
rect 177 -3169 181 -3165
rect 233 -3169 237 -3165
rect 267 -3169 271 -3165
rect 485 -3169 489 -3165
rect 541 -3169 545 -3165
rect 575 -3169 579 -3165
rect 793 -3169 797 -3165
rect 849 -3169 853 -3165
rect 883 -3169 887 -3165
<< labels >>
rlabel metal1 -1319 -948 -1315 -948 5 X0
rlabel metal1 -1076 -948 -1072 -948 5 X1
rlabel metal1 -768 -949 -764 -949 5 X2
rlabel metal1 -460 -948 -456 -948 5 X3
rlabel metal1 -152 -948 -148 -948 5 X4
rlabel metal1 156 -948 160 -948 5 X5
rlabel metal1 464 -948 468 -948 5 X6
rlabel metal1 772 -948 776 -948 5 X7
rlabel metal2 -1411 -1024 -1411 -1020 1 Y0
rlabel metal2 -1411 -1174 -1411 -1170 1 Y1
rlabel metal2 -1119 -1368 -1119 -1364 1 Z1
rlabel metal2 -1122 -1684 -1122 -1680 1 Z2
rlabel metal2 -1441 -2225 -1441 -2225 1 VDD!
rlabel metal2 1193 -2317 1193 -2317 1 GND!
rlabel metal2 -1411 -1495 -1411 -1491 1 Y2
rlabel metal2 -1411 -1786 -1411 -1782 1 Y3
rlabel metal2 -1411 -2108 -1411 -2104 1 Y4
rlabel metal2 -1411 -2399 -1411 -2395 1 Y5
rlabel metal2 -1411 -2690 -1411 -2686 1 Y6
rlabel metal2 -1411 -2981 -1411 -2977 1 Y7
rlabel metal2 -1122 -1975 -1122 -1971 1 Z3
rlabel metal2 -1122 -2297 -1122 -2293 1 Z4
rlabel metal2 -1122 -2588 -1122 -2584 1 Z5
rlabel metal2 -1122 -2879 -1122 -2875 1 Z6
rlabel metal2 -1122 -3170 -1122 -3166 1 Z7
rlabel metal2 -814 -3148 -814 -3144 1 Z8
rlabel metal2 -505 -3148 -505 -3144 1 Z9
rlabel metal2 -198 -3148 -198 -3144 1 Z10
rlabel metal2 111 -3148 111 -3144 1 Z11
rlabel metal2 418 -3148 418 -3144 1 Z12
rlabel metal2 726 -3148 726 -3144 1 Z13
rlabel metal2 1034 -3148 1034 -3144 1 Z14
rlabel metal1 1034 -3141 1034 -3137 1 Z15
rlabel metal1 -1277 -1033 -1277 -1029 1 Z0
<< end >>
