magic
tech scmos
timestamp 1615652171
<< ntransistor >>
rect -102 -30 -100 -26
rect -86 -30 -84 -26
rect -70 -30 -68 -26
rect -62 -30 -60 -26
rect -54 -30 -52 -26
rect -46 -30 -44 -26
rect -28 -30 -26 -26
rect -20 -30 -18 -26
rect -1 -30 1 -26
rect 15 -30 17 -26
rect 31 -30 33 -26
rect 47 -30 49 -26
rect 55 -30 57 -26
rect 63 -30 65 -26
rect 71 -30 73 -26
rect 87 -30 89 -26
rect 95 -30 97 -26
rect 114 -30 116 -26
rect 130 -30 132 -26
rect 138 -30 140 -26
rect 157 -30 159 -26
<< ptransistor >>
rect -102 26 -100 35
rect -86 26 -84 35
rect -70 26 -68 35
rect -62 26 -60 35
rect -54 26 -52 35
rect -46 26 -44 35
rect -28 26 -26 35
rect -20 26 -18 35
rect -1 26 1 35
rect 15 26 17 35
rect 31 26 33 35
rect 47 26 49 35
rect 55 26 57 35
rect 63 26 65 35
rect 71 26 73 35
rect 87 26 89 35
rect 95 26 97 35
rect 114 26 116 35
rect 130 26 132 35
rect 138 26 140 35
rect 157 26 159 35
<< ndiffusion >>
rect -103 -30 -102 -26
rect -100 -30 -99 -26
rect -87 -30 -86 -26
rect -84 -30 -83 -26
rect -71 -30 -70 -26
rect -68 -30 -62 -26
rect -60 -30 -59 -26
rect -55 -30 -54 -26
rect -52 -30 -46 -26
rect -44 -30 -43 -26
rect -29 -30 -28 -26
rect -26 -30 -20 -26
rect -18 -30 -17 -26
rect -2 -30 -1 -26
rect 1 -30 2 -26
rect 14 -30 15 -26
rect 17 -30 18 -26
rect 30 -30 31 -26
rect 33 -30 34 -26
rect 46 -30 47 -26
rect 49 -30 55 -26
rect 57 -30 58 -26
rect 62 -30 63 -26
rect 65 -30 71 -26
rect 73 -30 74 -26
rect 86 -30 87 -26
rect 89 -30 95 -26
rect 97 -30 98 -26
rect 113 -30 114 -26
rect 116 -30 117 -26
rect 129 -30 130 -26
rect 132 -30 133 -26
rect 137 -30 138 -26
rect 140 -30 146 -26
rect 150 -30 157 -26
rect 159 -30 160 -26
<< pdiffusion >>
rect -103 26 -102 35
rect -100 26 -99 35
rect -87 26 -86 35
rect -84 26 -83 35
rect -71 26 -70 35
rect -68 26 -67 35
rect -63 26 -62 35
rect -60 26 -54 35
rect -52 26 -51 35
rect -47 26 -46 35
rect -44 26 -43 35
rect -29 26 -28 35
rect -26 26 -25 35
rect -21 26 -20 35
rect -18 26 -11 35
rect -7 26 -1 35
rect 1 26 2 35
rect 14 26 15 35
rect 17 26 18 35
rect 30 26 31 35
rect 33 26 34 35
rect 46 26 47 35
rect 49 26 50 35
rect 54 26 55 35
rect 57 26 63 35
rect 65 26 66 35
rect 70 26 71 35
rect 73 26 74 35
rect 86 26 87 35
rect 89 26 90 35
rect 94 26 95 35
rect 97 26 104 35
rect 108 26 114 35
rect 116 26 117 35
rect 129 26 130 35
rect 132 26 138 35
rect 140 26 141 35
rect 156 26 157 35
rect 159 26 160 35
<< ndcontact >>
rect -107 -30 -103 -26
rect -99 -30 -95 -26
rect -91 -30 -87 -26
rect -83 -30 -79 -26
rect -59 -30 -55 -26
rect -33 -30 -29 -26
rect -17 -30 -13 -26
rect -6 -30 -2 -26
rect 2 -30 6 -26
rect 10 -30 14 -26
rect 18 -30 22 -26
rect 26 -30 30 -26
rect 34 -30 38 -26
rect 58 -30 62 -26
rect 82 -30 86 -26
rect 98 -30 102 -26
rect 109 -30 113 -26
rect 117 -30 121 -26
rect 125 -30 129 -26
rect 133 -30 137 -26
rect 146 -30 150 -26
rect 160 -30 164 -26
<< pdcontact >>
rect -107 26 -103 35
rect -99 26 -95 35
rect -91 26 -87 35
rect -83 26 -79 35
rect -75 26 -71 35
rect -67 26 -63 35
rect -43 26 -39 35
rect -33 26 -29 35
rect -25 26 -21 35
rect -11 26 -7 35
rect 2 26 6 35
rect 10 26 14 35
rect 18 26 22 35
rect 26 26 30 35
rect 34 26 38 35
rect 42 26 46 35
rect 50 26 54 35
rect 74 26 78 35
rect 82 26 86 35
rect 90 26 94 35
rect 104 26 108 35
rect 117 26 121 35
rect 125 26 129 35
rect 141 26 145 35
rect 152 26 156 35
rect 160 26 164 35
<< psubstratepcontact >>
rect -107 -38 -103 -34
rect -91 -38 -87 -34
rect -59 -38 -55 -34
rect -33 -38 -29 -34
rect -6 -38 -2 -34
rect 10 -38 14 -34
rect 26 -38 30 -34
rect 58 -38 62 -34
rect 82 -38 86 -34
rect 109 -38 113 -34
rect 125 -38 129 -34
rect 146 -38 150 -34
<< nsubstratencontact >>
rect -107 39 -103 43
rect -91 39 -87 43
rect -67 39 -63 43
rect -33 39 -29 43
rect -11 39 -7 43
rect 10 39 14 43
rect 26 39 30 43
rect 50 39 54 43
rect 82 39 86 43
rect 104 39 108 43
rect 125 39 129 43
rect 152 39 156 43
<< polysilicon >>
rect -102 35 -100 37
rect -86 35 -84 37
rect -70 35 -68 37
rect -62 35 -60 37
rect -54 35 -52 37
rect -46 35 -44 37
rect -28 35 -26 37
rect -20 35 -18 37
rect -1 35 1 37
rect 15 35 17 37
rect 31 35 33 37
rect 47 35 49 37
rect 55 35 57 37
rect 63 35 65 37
rect 71 35 73 37
rect 87 35 89 37
rect 95 35 97 37
rect 114 35 116 37
rect 130 35 132 37
rect 138 35 140 37
rect 157 35 159 37
rect -102 -26 -100 26
rect -86 -26 -84 26
rect -70 -5 -68 26
rect -62 16 -60 26
rect -70 -26 -68 -9
rect -62 -26 -60 12
rect -54 2 -52 26
rect -46 9 -44 26
rect -54 -26 -52 -2
rect -46 -26 -44 5
rect -28 -26 -26 26
rect -20 2 -18 26
rect -1 9 1 26
rect -2 5 1 9
rect -20 -26 -18 -2
rect -1 -26 1 5
rect 15 -26 17 26
rect 31 -26 33 26
rect 47 -5 49 26
rect 55 16 57 26
rect 47 -26 49 -9
rect 55 -26 57 12
rect 63 2 65 26
rect 71 9 73 26
rect 63 -26 65 -2
rect 71 -26 73 5
rect 87 -26 89 26
rect 95 2 97 26
rect 114 9 116 26
rect 130 9 132 26
rect 113 5 116 9
rect 95 -26 97 -2
rect 114 -26 116 5
rect 130 -26 132 5
rect 138 2 140 26
rect 157 9 159 26
rect 156 5 159 9
rect 138 -26 140 -2
rect 157 -26 159 5
rect -102 -32 -100 -30
rect -86 -32 -84 -30
rect -70 -32 -68 -30
rect -62 -32 -60 -30
rect -54 -32 -52 -30
rect -46 -32 -44 -30
rect -28 -32 -26 -30
rect -20 -32 -18 -30
rect -1 -32 1 -30
rect 15 -32 17 -30
rect 31 -32 33 -30
rect 47 -32 49 -30
rect 55 -32 57 -30
rect 63 -32 65 -30
rect 71 -32 73 -30
rect 87 -32 89 -30
rect 95 -32 97 -30
rect 114 -32 116 -30
rect 130 -32 132 -30
rect 138 -32 140 -30
rect 157 -32 159 -30
<< polycontact >>
rect -72 -9 -68 -5
rect -32 5 -28 9
rect -6 5 -2 9
rect -22 -2 -18 2
rect 45 -9 49 -5
rect 83 5 87 9
rect 109 5 113 9
rect 128 5 132 9
rect 93 -2 97 2
rect 152 5 156 9
rect 136 -2 140 2
<< metal1 >>
rect -111 39 -107 43
rect -103 39 -91 43
rect -87 39 -67 43
rect -63 39 -33 43
rect -29 39 -11 43
rect -7 39 10 43
rect 14 39 26 43
rect 30 39 50 43
rect 54 39 82 43
rect 86 39 104 43
rect 108 39 125 43
rect 129 39 152 43
rect 156 39 168 43
rect -107 35 -103 39
rect -91 35 -87 39
rect -67 35 -63 39
rect -33 35 -29 39
rect -11 35 -7 39
rect 10 35 14 39
rect 26 35 30 39
rect 50 35 54 39
rect 82 35 86 39
rect 104 35 108 39
rect 125 35 129 39
rect 152 35 156 39
rect -99 16 -95 26
rect -99 -26 -95 12
rect -83 -5 -79 26
rect -75 23 -71 26
rect -43 23 -39 26
rect -75 19 -39 23
rect -25 9 -21 26
rect -44 5 -32 9
rect -25 5 -6 9
rect -52 -2 -22 2
rect -83 -9 -72 -5
rect -55 -9 -32 -5
rect -83 -26 -79 -9
rect -13 -30 -9 5
rect 2 -12 6 26
rect 18 16 22 26
rect 11 -5 15 5
rect 2 -26 6 -16
rect 18 -26 22 12
rect 34 -5 38 26
rect 42 23 46 26
rect 74 23 78 26
rect 42 19 78 23
rect 90 9 94 26
rect 117 9 121 26
rect 145 9 149 35
rect 160 9 164 26
rect 73 5 83 9
rect 90 5 109 9
rect 117 5 128 9
rect 145 5 152 9
rect 160 5 168 9
rect 65 -2 93 2
rect 34 -9 45 -5
rect 70 -9 90 -5
rect 34 -26 38 -9
rect 102 -30 106 5
rect 117 -26 121 5
rect 136 -5 140 -2
rect 129 -9 140 -5
rect 145 -19 149 5
rect 133 -23 149 -19
rect 133 -26 137 -23
rect 160 -26 164 5
rect -107 -34 -103 -30
rect -91 -34 -87 -30
rect -59 -34 -55 -30
rect -33 -34 -29 -30
rect -6 -34 -2 -30
rect 10 -34 14 -30
rect 26 -34 30 -30
rect 58 -34 62 -30
rect 82 -34 86 -30
rect 109 -34 113 -30
rect 125 -34 129 -30
rect 146 -34 150 -30
rect -111 -38 -107 -34
rect -103 -38 -91 -34
rect -87 -38 -59 -34
rect -55 -38 -33 -34
rect -29 -38 -6 -34
rect -2 -38 10 -34
rect 14 -38 26 -34
rect 30 -38 58 -34
rect 62 -38 82 -34
rect 86 -38 109 -34
rect 113 -38 125 -34
rect 129 -38 146 -34
rect 150 -38 168 -34
<< m2contact >>
rect -99 12 -95 16
rect -59 -9 -55 -5
rect -32 -9 -28 -5
rect 18 12 22 16
rect 11 -9 15 -5
rect 2 -16 6 -12
rect 66 -9 70 -5
rect 90 -9 94 -5
rect 125 -9 129 -5
<< pm12contact >>
rect -106 5 -102 9
rect -90 -2 -86 2
rect -64 12 -60 16
rect -48 5 -44 9
rect -56 -2 -52 2
rect 11 5 15 9
rect 27 -2 31 2
rect 53 12 57 16
rect 69 5 73 9
rect 61 -2 65 2
<< pdm12contact >>
rect -51 26 -47 35
rect 66 26 70 35
<< ndm12contact >>
rect -75 -30 -71 -26
rect -43 -30 -39 -26
rect 42 -30 46 -26
rect 74 -30 78 -26
<< metal2 >>
rect -51 23 -47 26
rect 66 23 70 26
rect -51 19 -35 23
rect 66 19 82 23
rect -95 12 -64 16
rect -110 5 -106 9
rect -102 5 -48 9
rect -39 2 -35 19
rect 22 12 53 16
rect 15 5 69 9
rect 78 2 82 19
rect -110 -2 -90 2
rect -86 -2 -56 2
rect -39 -2 27 2
rect 31 -2 61 2
rect 78 -2 168 2
rect -110 -9 -59 -5
rect -39 -19 -35 -2
rect -28 -9 11 -5
rect 18 -9 66 -5
rect 18 -12 22 -9
rect 6 -16 22 -12
rect 78 -19 82 -2
rect 94 -9 125 -5
rect -75 -23 -35 -19
rect -75 -26 -71 -23
rect -39 -30 -35 -23
rect 42 -23 82 -19
rect 42 -26 46 -23
rect 78 -30 82 -23
<< labels >>
rlabel metal2 -110 -2 -110 2 3 B
rlabel metal2 -110 5 -110 9 3 A
rlabel metal2 -110 -9 -110 -5 3 CIN
rlabel metal2 168 -2 168 2 1 SUM
rlabel metal1 168 5 168 9 1 COUT
rlabel metal1 40 41 41 41 5 VDD!
rlabel metal1 40 -36 41 -36 1 GND!
<< end >>
