magic
tech scmos
timestamp 1618504402
<< polysilicon >>
rect -1302 -788 -1300 -786
rect -1294 -788 -1292 -786
rect -1284 -788 -1282 -786
rect -931 -788 -929 -786
rect -923 -788 -921 -786
rect -913 -788 -911 -786
rect -572 -788 -570 -786
rect -564 -788 -562 -786
rect -554 -788 -552 -786
rect -214 -788 -212 -786
rect -206 -788 -204 -786
rect -196 -788 -194 -786
rect 143 -788 145 -786
rect 151 -788 153 -786
rect 161 -788 163 -786
rect 500 -788 502 -786
rect 508 -788 510 -786
rect 518 -788 520 -786
rect 858 -788 860 -786
rect 866 -788 868 -786
rect 876 -788 878 -786
rect 1216 -788 1218 -786
rect 1224 -788 1226 -786
rect 1234 -788 1236 -786
rect -1302 -864 -1300 -796
rect -1294 -820 -1292 -796
rect -1294 -864 -1292 -824
rect -1284 -864 -1282 -796
rect -931 -864 -929 -796
rect -923 -820 -921 -796
rect -923 -864 -921 -824
rect -913 -864 -911 -796
rect -572 -864 -570 -796
rect -564 -820 -562 -796
rect -564 -864 -562 -824
rect -554 -864 -552 -796
rect -214 -864 -212 -796
rect -206 -820 -204 -796
rect -206 -864 -204 -824
rect -196 -864 -194 -796
rect 143 -864 145 -796
rect 151 -820 153 -796
rect 151 -864 153 -824
rect 161 -864 163 -796
rect 500 -864 502 -796
rect 508 -820 510 -796
rect 508 -864 510 -824
rect 518 -864 520 -796
rect 858 -864 860 -796
rect 866 -820 868 -796
rect 866 -864 868 -824
rect 876 -864 878 -796
rect 1216 -864 1218 -796
rect 1224 -820 1226 -796
rect 1224 -864 1226 -824
rect 1234 -864 1236 -796
rect -1302 -870 -1300 -868
rect -1294 -870 -1292 -868
rect -1284 -870 -1282 -868
rect -931 -870 -929 -868
rect -923 -870 -921 -868
rect -913 -870 -911 -868
rect -572 -870 -570 -868
rect -564 -870 -562 -868
rect -554 -870 -552 -868
rect -214 -870 -212 -868
rect -206 -870 -204 -868
rect -196 -870 -194 -868
rect 143 -870 145 -868
rect 151 -870 153 -868
rect 161 -870 163 -868
rect 500 -870 502 -868
rect 508 -870 510 -868
rect 518 -870 520 -868
rect 858 -870 860 -868
rect 866 -870 868 -868
rect 876 -870 878 -868
rect 1216 -870 1218 -868
rect 1224 -870 1226 -868
rect 1234 -870 1236 -868
rect -1225 -1022 -1223 -1020
rect -1215 -1022 -1213 -1020
rect -1199 -1022 -1197 -1020
rect -1191 -1022 -1189 -1020
rect -1175 -1022 -1173 -1020
rect -1167 -1022 -1165 -1020
rect -1157 -1022 -1155 -1020
rect -1149 -1022 -1147 -1020
rect -1133 -1022 -1131 -1020
rect -1125 -1022 -1123 -1020
rect -1115 -1022 -1113 -1020
rect -1107 -1022 -1105 -1020
rect -1091 -1022 -1089 -1020
rect -1083 -1022 -1081 -1020
rect -1073 -1022 -1071 -1020
rect -1065 -1022 -1063 -1020
rect -1049 -1022 -1047 -1020
rect -1041 -1022 -1039 -1020
rect -930 -1022 -928 -1020
rect -920 -1022 -918 -1020
rect -904 -1022 -902 -1020
rect -896 -1022 -894 -1020
rect -880 -1022 -878 -1020
rect -872 -1022 -870 -1020
rect -862 -1022 -860 -1020
rect -854 -1022 -852 -1020
rect -838 -1022 -836 -1020
rect -830 -1022 -828 -1020
rect -820 -1022 -818 -1020
rect -812 -1022 -810 -1020
rect -796 -1022 -794 -1020
rect -788 -1022 -786 -1020
rect -778 -1022 -776 -1020
rect -770 -1022 -768 -1020
rect -754 -1022 -752 -1020
rect -746 -1022 -744 -1020
rect -572 -1022 -570 -1020
rect -562 -1022 -560 -1020
rect -546 -1022 -544 -1020
rect -538 -1022 -536 -1020
rect -522 -1022 -520 -1020
rect -514 -1022 -512 -1020
rect -504 -1022 -502 -1020
rect -496 -1022 -494 -1020
rect -480 -1022 -478 -1020
rect -472 -1022 -470 -1020
rect -462 -1022 -460 -1020
rect -454 -1022 -452 -1020
rect -438 -1022 -436 -1020
rect -430 -1022 -428 -1020
rect -420 -1022 -418 -1020
rect -412 -1022 -410 -1020
rect -396 -1022 -394 -1020
rect -388 -1022 -386 -1020
rect -214 -1022 -212 -1020
rect -204 -1022 -202 -1020
rect -188 -1022 -186 -1020
rect -180 -1022 -178 -1020
rect -164 -1022 -162 -1020
rect -156 -1022 -154 -1020
rect -146 -1022 -144 -1020
rect -138 -1022 -136 -1020
rect -122 -1022 -120 -1020
rect -114 -1022 -112 -1020
rect -104 -1022 -102 -1020
rect -96 -1022 -94 -1020
rect -80 -1022 -78 -1020
rect -72 -1022 -70 -1020
rect -62 -1022 -60 -1020
rect -54 -1022 -52 -1020
rect -38 -1022 -36 -1020
rect -30 -1022 -28 -1020
rect 144 -1022 146 -1020
rect 154 -1022 156 -1020
rect 170 -1022 172 -1020
rect 178 -1022 180 -1020
rect 194 -1022 196 -1020
rect 202 -1022 204 -1020
rect 212 -1022 214 -1020
rect 220 -1022 222 -1020
rect 236 -1022 238 -1020
rect 244 -1022 246 -1020
rect 254 -1022 256 -1020
rect 262 -1022 264 -1020
rect 278 -1022 280 -1020
rect 286 -1022 288 -1020
rect 296 -1022 298 -1020
rect 304 -1022 306 -1020
rect 320 -1022 322 -1020
rect 328 -1022 330 -1020
rect 500 -1022 502 -1020
rect 510 -1022 512 -1020
rect 526 -1022 528 -1020
rect 534 -1022 536 -1020
rect 550 -1022 552 -1020
rect 558 -1022 560 -1020
rect 568 -1022 570 -1020
rect 576 -1022 578 -1020
rect 592 -1022 594 -1020
rect 600 -1022 602 -1020
rect 610 -1022 612 -1020
rect 618 -1022 620 -1020
rect 634 -1022 636 -1020
rect 642 -1022 644 -1020
rect 652 -1022 654 -1020
rect 660 -1022 662 -1020
rect 676 -1022 678 -1020
rect 684 -1022 686 -1020
rect 858 -1022 860 -1020
rect 868 -1022 870 -1020
rect 884 -1022 886 -1020
rect 892 -1022 894 -1020
rect 908 -1022 910 -1020
rect 916 -1022 918 -1020
rect 926 -1022 928 -1020
rect 934 -1022 936 -1020
rect 950 -1022 952 -1020
rect 958 -1022 960 -1020
rect 968 -1022 970 -1020
rect 976 -1022 978 -1020
rect 992 -1022 994 -1020
rect 1000 -1022 1002 -1020
rect 1010 -1022 1012 -1020
rect 1018 -1022 1020 -1020
rect 1034 -1022 1036 -1020
rect 1042 -1022 1044 -1020
rect -1225 -1098 -1223 -1030
rect -1215 -1098 -1213 -1030
rect -1199 -1098 -1197 -1030
rect -1191 -1098 -1189 -1030
rect -1175 -1098 -1173 -1030
rect -1167 -1098 -1165 -1030
rect -1157 -1098 -1155 -1030
rect -1149 -1098 -1147 -1030
rect -1133 -1098 -1131 -1030
rect -1125 -1063 -1123 -1030
rect -1115 -1063 -1113 -1030
rect -1125 -1065 -1113 -1063
rect -1125 -1098 -1123 -1065
rect -1115 -1098 -1113 -1065
rect -1107 -1098 -1105 -1030
rect -1091 -1098 -1089 -1030
rect -1083 -1098 -1081 -1030
rect -1073 -1098 -1071 -1030
rect -1065 -1098 -1063 -1030
rect -1049 -1098 -1047 -1030
rect -1041 -1098 -1039 -1030
rect -930 -1098 -928 -1030
rect -920 -1098 -918 -1030
rect -904 -1098 -902 -1030
rect -896 -1098 -894 -1030
rect -880 -1098 -878 -1030
rect -872 -1098 -870 -1030
rect -862 -1098 -860 -1030
rect -854 -1098 -852 -1030
rect -838 -1098 -836 -1030
rect -830 -1063 -828 -1030
rect -820 -1063 -818 -1030
rect -830 -1065 -818 -1063
rect -830 -1098 -828 -1065
rect -820 -1098 -818 -1065
rect -812 -1098 -810 -1030
rect -796 -1098 -794 -1030
rect -788 -1098 -786 -1030
rect -778 -1098 -776 -1030
rect -770 -1098 -768 -1030
rect -754 -1098 -752 -1030
rect -746 -1098 -744 -1030
rect -572 -1098 -570 -1030
rect -562 -1098 -560 -1030
rect -546 -1098 -544 -1030
rect -538 -1098 -536 -1030
rect -522 -1098 -520 -1030
rect -514 -1098 -512 -1030
rect -504 -1098 -502 -1030
rect -496 -1098 -494 -1030
rect -480 -1098 -478 -1030
rect -472 -1063 -470 -1030
rect -462 -1063 -460 -1030
rect -472 -1065 -460 -1063
rect -472 -1098 -470 -1065
rect -462 -1098 -460 -1065
rect -454 -1098 -452 -1030
rect -438 -1098 -436 -1030
rect -430 -1098 -428 -1030
rect -420 -1098 -418 -1030
rect -412 -1098 -410 -1030
rect -396 -1098 -394 -1030
rect -388 -1098 -386 -1030
rect -214 -1098 -212 -1030
rect -204 -1098 -202 -1030
rect -188 -1098 -186 -1030
rect -180 -1098 -178 -1030
rect -164 -1098 -162 -1030
rect -156 -1098 -154 -1030
rect -146 -1098 -144 -1030
rect -138 -1098 -136 -1030
rect -122 -1098 -120 -1030
rect -114 -1063 -112 -1030
rect -104 -1063 -102 -1030
rect -114 -1065 -102 -1063
rect -114 -1098 -112 -1065
rect -104 -1098 -102 -1065
rect -96 -1098 -94 -1030
rect -80 -1098 -78 -1030
rect -72 -1098 -70 -1030
rect -62 -1098 -60 -1030
rect -54 -1098 -52 -1030
rect -38 -1098 -36 -1030
rect -30 -1098 -28 -1030
rect 144 -1098 146 -1030
rect 154 -1098 156 -1030
rect 170 -1098 172 -1030
rect 178 -1098 180 -1030
rect 194 -1098 196 -1030
rect 202 -1098 204 -1030
rect 212 -1098 214 -1030
rect 220 -1098 222 -1030
rect 236 -1098 238 -1030
rect 244 -1063 246 -1030
rect 254 -1063 256 -1030
rect 244 -1065 256 -1063
rect 244 -1098 246 -1065
rect 254 -1098 256 -1065
rect 262 -1098 264 -1030
rect 278 -1098 280 -1030
rect 286 -1098 288 -1030
rect 296 -1098 298 -1030
rect 304 -1098 306 -1030
rect 320 -1098 322 -1030
rect 328 -1098 330 -1030
rect 500 -1098 502 -1030
rect 510 -1098 512 -1030
rect 526 -1098 528 -1030
rect 534 -1098 536 -1030
rect 550 -1098 552 -1030
rect 558 -1098 560 -1030
rect 568 -1098 570 -1030
rect 576 -1098 578 -1030
rect 592 -1098 594 -1030
rect 600 -1063 602 -1030
rect 610 -1063 612 -1030
rect 600 -1065 612 -1063
rect 600 -1098 602 -1065
rect 610 -1098 612 -1065
rect 618 -1098 620 -1030
rect 634 -1098 636 -1030
rect 642 -1098 644 -1030
rect 652 -1098 654 -1030
rect 660 -1098 662 -1030
rect 676 -1098 678 -1030
rect 684 -1098 686 -1030
rect 858 -1098 860 -1030
rect 868 -1098 870 -1030
rect 884 -1098 886 -1030
rect 892 -1098 894 -1030
rect 908 -1098 910 -1030
rect 916 -1098 918 -1030
rect 926 -1098 928 -1030
rect 934 -1098 936 -1030
rect 950 -1098 952 -1030
rect 958 -1063 960 -1030
rect 968 -1063 970 -1030
rect 958 -1065 970 -1063
rect 958 -1098 960 -1065
rect 968 -1098 970 -1065
rect 976 -1098 978 -1030
rect 992 -1098 994 -1030
rect 1000 -1098 1002 -1030
rect 1010 -1098 1012 -1030
rect 1018 -1098 1020 -1030
rect 1034 -1098 1036 -1030
rect 1042 -1098 1044 -1030
rect -1225 -1104 -1223 -1102
rect -1215 -1104 -1213 -1102
rect -1199 -1104 -1197 -1102
rect -1191 -1104 -1189 -1102
rect -1175 -1104 -1173 -1102
rect -1167 -1104 -1165 -1102
rect -1157 -1104 -1155 -1102
rect -1149 -1104 -1147 -1102
rect -1133 -1104 -1131 -1102
rect -1125 -1104 -1123 -1102
rect -1115 -1104 -1113 -1102
rect -1107 -1104 -1105 -1102
rect -1091 -1104 -1089 -1102
rect -1083 -1104 -1081 -1102
rect -1073 -1104 -1071 -1102
rect -1065 -1104 -1063 -1102
rect -1049 -1104 -1047 -1102
rect -1041 -1104 -1039 -1102
rect -930 -1104 -928 -1102
rect -920 -1104 -918 -1102
rect -904 -1104 -902 -1102
rect -896 -1104 -894 -1102
rect -880 -1104 -878 -1102
rect -872 -1104 -870 -1102
rect -862 -1104 -860 -1102
rect -854 -1104 -852 -1102
rect -838 -1104 -836 -1102
rect -830 -1104 -828 -1102
rect -820 -1104 -818 -1102
rect -812 -1104 -810 -1102
rect -796 -1104 -794 -1102
rect -788 -1104 -786 -1102
rect -778 -1104 -776 -1102
rect -770 -1104 -768 -1102
rect -754 -1104 -752 -1102
rect -746 -1104 -744 -1102
rect -572 -1104 -570 -1102
rect -562 -1104 -560 -1102
rect -546 -1104 -544 -1102
rect -538 -1104 -536 -1102
rect -522 -1104 -520 -1102
rect -514 -1104 -512 -1102
rect -504 -1104 -502 -1102
rect -496 -1104 -494 -1102
rect -480 -1104 -478 -1102
rect -472 -1104 -470 -1102
rect -462 -1104 -460 -1102
rect -454 -1104 -452 -1102
rect -438 -1104 -436 -1102
rect -430 -1104 -428 -1102
rect -420 -1104 -418 -1102
rect -412 -1104 -410 -1102
rect -396 -1104 -394 -1102
rect -388 -1104 -386 -1102
rect -214 -1104 -212 -1102
rect -204 -1104 -202 -1102
rect -188 -1104 -186 -1102
rect -180 -1104 -178 -1102
rect -164 -1104 -162 -1102
rect -156 -1104 -154 -1102
rect -146 -1104 -144 -1102
rect -138 -1104 -136 -1102
rect -122 -1104 -120 -1102
rect -114 -1104 -112 -1102
rect -104 -1104 -102 -1102
rect -96 -1104 -94 -1102
rect -80 -1104 -78 -1102
rect -72 -1104 -70 -1102
rect -62 -1104 -60 -1102
rect -54 -1104 -52 -1102
rect -38 -1104 -36 -1102
rect -30 -1104 -28 -1102
rect 144 -1104 146 -1102
rect 154 -1104 156 -1102
rect 170 -1104 172 -1102
rect 178 -1104 180 -1102
rect 194 -1104 196 -1102
rect 202 -1104 204 -1102
rect 212 -1104 214 -1102
rect 220 -1104 222 -1102
rect 236 -1104 238 -1102
rect 244 -1104 246 -1102
rect 254 -1104 256 -1102
rect 262 -1104 264 -1102
rect 278 -1104 280 -1102
rect 286 -1104 288 -1102
rect 296 -1104 298 -1102
rect 304 -1104 306 -1102
rect 320 -1104 322 -1102
rect 328 -1104 330 -1102
rect 500 -1104 502 -1102
rect 510 -1104 512 -1102
rect 526 -1104 528 -1102
rect 534 -1104 536 -1102
rect 550 -1104 552 -1102
rect 558 -1104 560 -1102
rect 568 -1104 570 -1102
rect 576 -1104 578 -1102
rect 592 -1104 594 -1102
rect 600 -1104 602 -1102
rect 610 -1104 612 -1102
rect 618 -1104 620 -1102
rect 634 -1104 636 -1102
rect 642 -1104 644 -1102
rect 652 -1104 654 -1102
rect 660 -1104 662 -1102
rect 676 -1104 678 -1102
rect 684 -1104 686 -1102
rect 858 -1104 860 -1102
rect 868 -1104 870 -1102
rect 884 -1104 886 -1102
rect 892 -1104 894 -1102
rect 908 -1104 910 -1102
rect 916 -1104 918 -1102
rect 926 -1104 928 -1102
rect 934 -1104 936 -1102
rect 950 -1104 952 -1102
rect 958 -1104 960 -1102
rect 968 -1104 970 -1102
rect 976 -1104 978 -1102
rect 992 -1104 994 -1102
rect 1000 -1104 1002 -1102
rect 1010 -1104 1012 -1102
rect 1018 -1104 1020 -1102
rect 1034 -1104 1036 -1102
rect 1042 -1104 1044 -1102
rect -1304 -1138 -1302 -1136
rect -1296 -1138 -1294 -1136
rect -1286 -1138 -1284 -1136
rect -930 -1138 -928 -1136
rect -922 -1138 -920 -1136
rect -912 -1138 -910 -1136
rect -572 -1138 -570 -1136
rect -564 -1138 -562 -1136
rect -554 -1138 -552 -1136
rect -214 -1138 -212 -1136
rect -206 -1138 -204 -1136
rect -196 -1138 -194 -1136
rect 144 -1138 146 -1136
rect 152 -1138 154 -1136
rect 162 -1138 164 -1136
rect 500 -1138 502 -1136
rect 508 -1138 510 -1136
rect 518 -1138 520 -1136
rect 858 -1138 860 -1136
rect 866 -1138 868 -1136
rect 876 -1138 878 -1136
rect 1216 -1138 1218 -1136
rect 1224 -1138 1226 -1136
rect 1234 -1138 1236 -1136
rect -1304 -1214 -1302 -1146
rect -1296 -1170 -1294 -1146
rect -1296 -1214 -1294 -1174
rect -1286 -1214 -1284 -1146
rect -930 -1214 -928 -1146
rect -922 -1170 -920 -1146
rect -922 -1214 -920 -1174
rect -912 -1214 -910 -1146
rect -572 -1214 -570 -1146
rect -564 -1170 -562 -1146
rect -564 -1214 -562 -1174
rect -554 -1214 -552 -1146
rect -214 -1214 -212 -1146
rect -206 -1170 -204 -1146
rect -206 -1214 -204 -1174
rect -196 -1214 -194 -1146
rect 144 -1214 146 -1146
rect 152 -1170 154 -1146
rect 152 -1214 154 -1174
rect 162 -1214 164 -1146
rect 500 -1214 502 -1146
rect 508 -1170 510 -1146
rect 508 -1214 510 -1174
rect 518 -1214 520 -1146
rect 858 -1214 860 -1146
rect 866 -1170 868 -1146
rect 866 -1214 868 -1174
rect 876 -1214 878 -1146
rect 1216 -1214 1218 -1146
rect 1224 -1170 1226 -1146
rect 1224 -1214 1226 -1174
rect 1234 -1214 1236 -1146
rect -1304 -1220 -1302 -1218
rect -1296 -1220 -1294 -1218
rect -1286 -1220 -1284 -1218
rect -930 -1220 -928 -1218
rect -922 -1220 -920 -1218
rect -912 -1220 -910 -1218
rect -572 -1220 -570 -1218
rect -564 -1220 -562 -1218
rect -554 -1220 -552 -1218
rect -214 -1220 -212 -1218
rect -206 -1220 -204 -1218
rect -196 -1220 -194 -1218
rect 144 -1220 146 -1218
rect 152 -1220 154 -1218
rect 162 -1220 164 -1218
rect 500 -1220 502 -1218
rect 508 -1220 510 -1218
rect 518 -1220 520 -1218
rect 858 -1220 860 -1218
rect 866 -1220 868 -1218
rect 876 -1220 878 -1218
rect 1216 -1220 1218 -1218
rect 1224 -1220 1226 -1218
rect 1234 -1220 1236 -1218
rect -1225 -1302 -1223 -1300
rect -1215 -1302 -1213 -1300
rect -1199 -1302 -1197 -1300
rect -1189 -1302 -1187 -1300
rect -1181 -1302 -1179 -1300
rect -1171 -1302 -1169 -1300
rect -1155 -1302 -1153 -1300
rect -1147 -1302 -1145 -1300
rect -1137 -1302 -1135 -1300
rect -930 -1302 -928 -1300
rect -920 -1302 -918 -1300
rect -904 -1302 -902 -1300
rect -894 -1302 -892 -1300
rect -878 -1302 -876 -1300
rect -868 -1302 -866 -1300
rect -860 -1302 -858 -1300
rect -850 -1302 -848 -1300
rect -834 -1302 -832 -1300
rect -826 -1302 -824 -1300
rect -816 -1302 -814 -1300
rect -800 -1302 -798 -1300
rect -790 -1302 -788 -1300
rect -782 -1302 -780 -1300
rect -772 -1302 -770 -1300
rect -756 -1302 -754 -1300
rect -748 -1302 -746 -1300
rect -732 -1302 -730 -1300
rect -716 -1302 -714 -1300
rect -708 -1302 -706 -1300
rect -698 -1302 -696 -1300
rect -572 -1302 -570 -1300
rect -562 -1302 -560 -1300
rect -546 -1302 -544 -1300
rect -536 -1302 -534 -1300
rect -520 -1302 -518 -1300
rect -510 -1302 -508 -1300
rect -502 -1302 -500 -1300
rect -492 -1302 -490 -1300
rect -476 -1302 -474 -1300
rect -468 -1302 -466 -1300
rect -458 -1302 -456 -1300
rect -442 -1302 -440 -1300
rect -432 -1302 -430 -1300
rect -424 -1302 -422 -1300
rect -414 -1302 -412 -1300
rect -398 -1302 -396 -1300
rect -390 -1302 -388 -1300
rect -374 -1302 -372 -1300
rect -358 -1302 -356 -1300
rect -350 -1302 -348 -1300
rect -340 -1302 -338 -1300
rect -214 -1302 -212 -1300
rect -204 -1302 -202 -1300
rect -188 -1302 -186 -1300
rect -178 -1302 -176 -1300
rect -162 -1302 -160 -1300
rect -152 -1302 -150 -1300
rect -144 -1302 -142 -1300
rect -134 -1302 -132 -1300
rect -118 -1302 -116 -1300
rect -110 -1302 -108 -1300
rect -100 -1302 -98 -1300
rect -84 -1302 -82 -1300
rect -74 -1302 -72 -1300
rect -66 -1302 -64 -1300
rect -56 -1302 -54 -1300
rect -40 -1302 -38 -1300
rect -32 -1302 -30 -1300
rect -16 -1302 -14 -1300
rect 0 -1302 2 -1300
rect 8 -1302 10 -1300
rect 18 -1302 20 -1300
rect 144 -1302 146 -1300
rect 154 -1302 156 -1300
rect 170 -1302 172 -1300
rect 180 -1302 182 -1300
rect 196 -1302 198 -1300
rect 206 -1302 208 -1300
rect 214 -1302 216 -1300
rect 224 -1302 226 -1300
rect 240 -1302 242 -1300
rect 248 -1302 250 -1300
rect 258 -1302 260 -1300
rect 274 -1302 276 -1300
rect 284 -1302 286 -1300
rect 292 -1302 294 -1300
rect 302 -1302 304 -1300
rect 318 -1302 320 -1300
rect 326 -1302 328 -1300
rect 342 -1302 344 -1300
rect 358 -1302 360 -1300
rect 366 -1302 368 -1300
rect 376 -1302 378 -1300
rect 500 -1302 502 -1300
rect 510 -1302 512 -1300
rect 526 -1302 528 -1300
rect 536 -1302 538 -1300
rect 552 -1302 554 -1300
rect 562 -1302 564 -1300
rect 570 -1302 572 -1300
rect 580 -1302 582 -1300
rect 596 -1302 598 -1300
rect 604 -1302 606 -1300
rect 614 -1302 616 -1300
rect 630 -1302 632 -1300
rect 640 -1302 642 -1300
rect 648 -1302 650 -1300
rect 658 -1302 660 -1300
rect 674 -1302 676 -1300
rect 682 -1302 684 -1300
rect 698 -1302 700 -1300
rect 714 -1302 716 -1300
rect 722 -1302 724 -1300
rect 732 -1302 734 -1300
rect 858 -1302 860 -1300
rect 868 -1302 870 -1300
rect 884 -1302 886 -1300
rect 894 -1302 896 -1300
rect 910 -1302 912 -1300
rect 920 -1302 922 -1300
rect 928 -1302 930 -1300
rect 938 -1302 940 -1300
rect 954 -1302 956 -1300
rect 962 -1302 964 -1300
rect 972 -1302 974 -1300
rect 988 -1302 990 -1300
rect 998 -1302 1000 -1300
rect 1006 -1302 1008 -1300
rect 1016 -1302 1018 -1300
rect 1032 -1302 1034 -1300
rect 1040 -1302 1042 -1300
rect 1056 -1302 1058 -1300
rect 1072 -1302 1074 -1300
rect 1080 -1302 1082 -1300
rect 1090 -1302 1092 -1300
rect 1216 -1302 1218 -1300
rect 1226 -1302 1228 -1300
rect 1242 -1302 1244 -1300
rect 1252 -1302 1254 -1300
rect 1260 -1302 1262 -1300
rect 1270 -1302 1272 -1300
rect 1286 -1302 1288 -1300
rect 1294 -1302 1296 -1300
rect 1304 -1302 1306 -1300
rect -1225 -1378 -1223 -1310
rect -1215 -1378 -1213 -1310
rect -1199 -1378 -1197 -1310
rect -1189 -1378 -1187 -1310
rect -1181 -1378 -1179 -1310
rect -1171 -1378 -1169 -1310
rect -1155 -1378 -1153 -1310
rect -1147 -1378 -1145 -1310
rect -1137 -1378 -1135 -1310
rect -930 -1378 -928 -1310
rect -920 -1378 -918 -1310
rect -904 -1378 -902 -1310
rect -894 -1378 -892 -1310
rect -878 -1378 -876 -1310
rect -868 -1378 -866 -1310
rect -860 -1378 -858 -1310
rect -850 -1378 -848 -1310
rect -834 -1378 -832 -1310
rect -826 -1378 -824 -1310
rect -816 -1378 -814 -1310
rect -800 -1378 -798 -1310
rect -790 -1378 -788 -1310
rect -782 -1378 -780 -1310
rect -772 -1378 -770 -1310
rect -756 -1378 -754 -1310
rect -748 -1378 -746 -1310
rect -732 -1378 -730 -1310
rect -716 -1378 -714 -1310
rect -708 -1378 -706 -1310
rect -698 -1378 -696 -1310
rect -572 -1378 -570 -1310
rect -562 -1378 -560 -1310
rect -546 -1378 -544 -1310
rect -536 -1378 -534 -1310
rect -520 -1378 -518 -1310
rect -510 -1378 -508 -1310
rect -502 -1378 -500 -1310
rect -492 -1378 -490 -1310
rect -476 -1378 -474 -1310
rect -468 -1378 -466 -1310
rect -458 -1378 -456 -1310
rect -442 -1378 -440 -1310
rect -432 -1378 -430 -1310
rect -424 -1378 -422 -1310
rect -414 -1378 -412 -1310
rect -398 -1378 -396 -1310
rect -390 -1378 -388 -1310
rect -374 -1378 -372 -1310
rect -358 -1378 -356 -1310
rect -350 -1378 -348 -1310
rect -340 -1378 -338 -1310
rect -214 -1378 -212 -1310
rect -204 -1378 -202 -1310
rect -188 -1378 -186 -1310
rect -178 -1378 -176 -1310
rect -162 -1378 -160 -1310
rect -152 -1378 -150 -1310
rect -144 -1378 -142 -1310
rect -134 -1378 -132 -1310
rect -118 -1378 -116 -1310
rect -110 -1378 -108 -1310
rect -100 -1378 -98 -1310
rect -84 -1378 -82 -1310
rect -74 -1378 -72 -1310
rect -66 -1378 -64 -1310
rect -56 -1378 -54 -1310
rect -40 -1378 -38 -1310
rect -32 -1378 -30 -1310
rect -16 -1378 -14 -1310
rect 0 -1378 2 -1310
rect 8 -1378 10 -1310
rect 18 -1378 20 -1310
rect 144 -1378 146 -1310
rect 154 -1378 156 -1310
rect 170 -1378 172 -1310
rect 180 -1378 182 -1310
rect 196 -1378 198 -1310
rect 206 -1378 208 -1310
rect 214 -1378 216 -1310
rect 224 -1378 226 -1310
rect 240 -1378 242 -1310
rect 248 -1378 250 -1310
rect 258 -1378 260 -1310
rect 274 -1378 276 -1310
rect 284 -1378 286 -1310
rect 292 -1378 294 -1310
rect 302 -1378 304 -1310
rect 318 -1378 320 -1310
rect 326 -1378 328 -1310
rect 342 -1378 344 -1310
rect 358 -1378 360 -1310
rect 366 -1378 368 -1310
rect 376 -1378 378 -1310
rect 500 -1378 502 -1310
rect 510 -1378 512 -1310
rect 526 -1378 528 -1310
rect 536 -1378 538 -1310
rect 552 -1378 554 -1310
rect 562 -1378 564 -1310
rect 570 -1378 572 -1310
rect 580 -1378 582 -1310
rect 596 -1378 598 -1310
rect 604 -1378 606 -1310
rect 614 -1378 616 -1310
rect 630 -1378 632 -1310
rect 640 -1378 642 -1310
rect 648 -1378 650 -1310
rect 658 -1378 660 -1310
rect 674 -1378 676 -1310
rect 682 -1378 684 -1310
rect 698 -1378 700 -1310
rect 714 -1378 716 -1310
rect 722 -1378 724 -1310
rect 732 -1378 734 -1310
rect 858 -1378 860 -1310
rect 868 -1378 870 -1310
rect 884 -1378 886 -1310
rect 894 -1378 896 -1310
rect 910 -1378 912 -1310
rect 920 -1378 922 -1310
rect 928 -1378 930 -1310
rect 938 -1378 940 -1310
rect 954 -1378 956 -1310
rect 962 -1378 964 -1310
rect 972 -1378 974 -1310
rect 988 -1378 990 -1310
rect 998 -1378 1000 -1310
rect 1006 -1378 1008 -1310
rect 1016 -1378 1018 -1310
rect 1032 -1378 1034 -1310
rect 1040 -1378 1042 -1310
rect 1056 -1378 1058 -1310
rect 1072 -1378 1074 -1310
rect 1080 -1378 1082 -1310
rect 1090 -1378 1092 -1310
rect 1216 -1378 1218 -1310
rect 1226 -1378 1228 -1310
rect 1242 -1378 1244 -1310
rect 1252 -1378 1254 -1310
rect 1260 -1378 1262 -1310
rect 1270 -1378 1272 -1310
rect 1286 -1378 1288 -1310
rect 1294 -1378 1296 -1310
rect 1304 -1378 1306 -1310
rect -1225 -1384 -1223 -1382
rect -1215 -1384 -1213 -1382
rect -1199 -1384 -1197 -1382
rect -1189 -1384 -1187 -1382
rect -1181 -1384 -1179 -1382
rect -1171 -1384 -1169 -1382
rect -1155 -1384 -1153 -1382
rect -1147 -1384 -1145 -1382
rect -1137 -1384 -1135 -1382
rect -930 -1384 -928 -1382
rect -920 -1384 -918 -1382
rect -904 -1384 -902 -1382
rect -894 -1384 -892 -1382
rect -878 -1384 -876 -1382
rect -868 -1384 -866 -1382
rect -860 -1384 -858 -1382
rect -850 -1384 -848 -1382
rect -834 -1384 -832 -1382
rect -826 -1384 -824 -1382
rect -816 -1384 -814 -1382
rect -800 -1384 -798 -1382
rect -790 -1384 -788 -1382
rect -782 -1384 -780 -1382
rect -772 -1384 -770 -1382
rect -756 -1384 -754 -1382
rect -748 -1384 -746 -1382
rect -732 -1384 -730 -1382
rect -716 -1384 -714 -1382
rect -708 -1384 -706 -1382
rect -698 -1384 -696 -1382
rect -572 -1384 -570 -1382
rect -562 -1384 -560 -1382
rect -546 -1384 -544 -1382
rect -536 -1384 -534 -1382
rect -520 -1384 -518 -1382
rect -510 -1384 -508 -1382
rect -502 -1384 -500 -1382
rect -492 -1384 -490 -1382
rect -476 -1384 -474 -1382
rect -468 -1384 -466 -1382
rect -458 -1384 -456 -1382
rect -442 -1384 -440 -1382
rect -432 -1384 -430 -1382
rect -424 -1384 -422 -1382
rect -414 -1384 -412 -1382
rect -398 -1384 -396 -1382
rect -390 -1384 -388 -1382
rect -374 -1384 -372 -1382
rect -358 -1384 -356 -1382
rect -350 -1384 -348 -1382
rect -340 -1384 -338 -1382
rect -214 -1384 -212 -1382
rect -204 -1384 -202 -1382
rect -188 -1384 -186 -1382
rect -178 -1384 -176 -1382
rect -162 -1384 -160 -1382
rect -152 -1384 -150 -1382
rect -144 -1384 -142 -1382
rect -134 -1384 -132 -1382
rect -118 -1384 -116 -1382
rect -110 -1384 -108 -1382
rect -100 -1384 -98 -1382
rect -84 -1384 -82 -1382
rect -74 -1384 -72 -1382
rect -66 -1384 -64 -1382
rect -56 -1384 -54 -1382
rect -40 -1384 -38 -1382
rect -32 -1384 -30 -1382
rect -16 -1384 -14 -1382
rect 0 -1384 2 -1382
rect 8 -1384 10 -1382
rect 18 -1384 20 -1382
rect 144 -1384 146 -1382
rect 154 -1384 156 -1382
rect 170 -1384 172 -1382
rect 180 -1384 182 -1382
rect 196 -1384 198 -1382
rect 206 -1384 208 -1382
rect 214 -1384 216 -1382
rect 224 -1384 226 -1382
rect 240 -1384 242 -1382
rect 248 -1384 250 -1382
rect 258 -1384 260 -1382
rect 274 -1384 276 -1382
rect 284 -1384 286 -1382
rect 292 -1384 294 -1382
rect 302 -1384 304 -1382
rect 318 -1384 320 -1382
rect 326 -1384 328 -1382
rect 342 -1384 344 -1382
rect 358 -1384 360 -1382
rect 366 -1384 368 -1382
rect 376 -1384 378 -1382
rect 500 -1384 502 -1382
rect 510 -1384 512 -1382
rect 526 -1384 528 -1382
rect 536 -1384 538 -1382
rect 552 -1384 554 -1382
rect 562 -1384 564 -1382
rect 570 -1384 572 -1382
rect 580 -1384 582 -1382
rect 596 -1384 598 -1382
rect 604 -1384 606 -1382
rect 614 -1384 616 -1382
rect 630 -1384 632 -1382
rect 640 -1384 642 -1382
rect 648 -1384 650 -1382
rect 658 -1384 660 -1382
rect 674 -1384 676 -1382
rect 682 -1384 684 -1382
rect 698 -1384 700 -1382
rect 714 -1384 716 -1382
rect 722 -1384 724 -1382
rect 732 -1384 734 -1382
rect 858 -1384 860 -1382
rect 868 -1384 870 -1382
rect 884 -1384 886 -1382
rect 894 -1384 896 -1382
rect 910 -1384 912 -1382
rect 920 -1384 922 -1382
rect 928 -1384 930 -1382
rect 938 -1384 940 -1382
rect 954 -1384 956 -1382
rect 962 -1384 964 -1382
rect 972 -1384 974 -1382
rect 988 -1384 990 -1382
rect 998 -1384 1000 -1382
rect 1006 -1384 1008 -1382
rect 1016 -1384 1018 -1382
rect 1032 -1384 1034 -1382
rect 1040 -1384 1042 -1382
rect 1056 -1384 1058 -1382
rect 1072 -1384 1074 -1382
rect 1080 -1384 1082 -1382
rect 1090 -1384 1092 -1382
rect 1216 -1384 1218 -1382
rect 1226 -1384 1228 -1382
rect 1242 -1384 1244 -1382
rect 1252 -1384 1254 -1382
rect 1260 -1384 1262 -1382
rect 1270 -1384 1272 -1382
rect 1286 -1384 1288 -1382
rect 1294 -1384 1296 -1382
rect 1304 -1384 1306 -1382
rect -1225 -1425 -1223 -1423
rect -1215 -1425 -1213 -1423
rect -1199 -1425 -1197 -1423
rect -1191 -1425 -1189 -1423
rect -1175 -1425 -1173 -1423
rect -1167 -1425 -1165 -1423
rect -1157 -1425 -1155 -1423
rect -1149 -1425 -1147 -1423
rect -1133 -1425 -1131 -1423
rect -1125 -1425 -1123 -1423
rect -1115 -1425 -1113 -1423
rect -1107 -1425 -1105 -1423
rect -1091 -1425 -1089 -1423
rect -1083 -1425 -1081 -1423
rect -1073 -1425 -1071 -1423
rect -1065 -1425 -1063 -1423
rect -1049 -1425 -1047 -1423
rect -1041 -1425 -1039 -1423
rect -930 -1425 -928 -1423
rect -920 -1425 -918 -1423
rect -904 -1425 -902 -1423
rect -896 -1425 -894 -1423
rect -880 -1425 -878 -1423
rect -872 -1425 -870 -1423
rect -862 -1425 -860 -1423
rect -854 -1425 -852 -1423
rect -838 -1425 -836 -1423
rect -830 -1425 -828 -1423
rect -820 -1425 -818 -1423
rect -812 -1425 -810 -1423
rect -796 -1425 -794 -1423
rect -788 -1425 -786 -1423
rect -778 -1425 -776 -1423
rect -770 -1425 -768 -1423
rect -754 -1425 -752 -1423
rect -746 -1425 -744 -1423
rect -572 -1425 -570 -1423
rect -562 -1425 -560 -1423
rect -546 -1425 -544 -1423
rect -538 -1425 -536 -1423
rect -522 -1425 -520 -1423
rect -514 -1425 -512 -1423
rect -504 -1425 -502 -1423
rect -496 -1425 -494 -1423
rect -480 -1425 -478 -1423
rect -472 -1425 -470 -1423
rect -462 -1425 -460 -1423
rect -454 -1425 -452 -1423
rect -438 -1425 -436 -1423
rect -430 -1425 -428 -1423
rect -420 -1425 -418 -1423
rect -412 -1425 -410 -1423
rect -396 -1425 -394 -1423
rect -388 -1425 -386 -1423
rect -214 -1425 -212 -1423
rect -204 -1425 -202 -1423
rect -188 -1425 -186 -1423
rect -180 -1425 -178 -1423
rect -164 -1425 -162 -1423
rect -156 -1425 -154 -1423
rect -146 -1425 -144 -1423
rect -138 -1425 -136 -1423
rect -122 -1425 -120 -1423
rect -114 -1425 -112 -1423
rect -104 -1425 -102 -1423
rect -96 -1425 -94 -1423
rect -80 -1425 -78 -1423
rect -72 -1425 -70 -1423
rect -62 -1425 -60 -1423
rect -54 -1425 -52 -1423
rect -38 -1425 -36 -1423
rect -30 -1425 -28 -1423
rect 144 -1425 146 -1423
rect 154 -1425 156 -1423
rect 170 -1425 172 -1423
rect 178 -1425 180 -1423
rect 194 -1425 196 -1423
rect 202 -1425 204 -1423
rect 212 -1425 214 -1423
rect 220 -1425 222 -1423
rect 236 -1425 238 -1423
rect 244 -1425 246 -1423
rect 254 -1425 256 -1423
rect 262 -1425 264 -1423
rect 278 -1425 280 -1423
rect 286 -1425 288 -1423
rect 296 -1425 298 -1423
rect 304 -1425 306 -1423
rect 320 -1425 322 -1423
rect 328 -1425 330 -1423
rect 500 -1425 502 -1423
rect 510 -1425 512 -1423
rect 526 -1425 528 -1423
rect 534 -1425 536 -1423
rect 550 -1425 552 -1423
rect 558 -1425 560 -1423
rect 568 -1425 570 -1423
rect 576 -1425 578 -1423
rect 592 -1425 594 -1423
rect 600 -1425 602 -1423
rect 610 -1425 612 -1423
rect 618 -1425 620 -1423
rect 634 -1425 636 -1423
rect 642 -1425 644 -1423
rect 652 -1425 654 -1423
rect 660 -1425 662 -1423
rect 676 -1425 678 -1423
rect 684 -1425 686 -1423
rect 858 -1425 860 -1423
rect 868 -1425 870 -1423
rect 884 -1425 886 -1423
rect 892 -1425 894 -1423
rect 908 -1425 910 -1423
rect 916 -1425 918 -1423
rect 926 -1425 928 -1423
rect 934 -1425 936 -1423
rect 950 -1425 952 -1423
rect 958 -1425 960 -1423
rect 968 -1425 970 -1423
rect 976 -1425 978 -1423
rect 992 -1425 994 -1423
rect 1000 -1425 1002 -1423
rect 1010 -1425 1012 -1423
rect 1018 -1425 1020 -1423
rect 1034 -1425 1036 -1423
rect 1042 -1425 1044 -1423
rect -1225 -1501 -1223 -1433
rect -1215 -1501 -1213 -1433
rect -1199 -1501 -1197 -1433
rect -1191 -1501 -1189 -1433
rect -1175 -1501 -1173 -1433
rect -1167 -1501 -1165 -1433
rect -1157 -1501 -1155 -1433
rect -1149 -1501 -1147 -1433
rect -1133 -1501 -1131 -1433
rect -1125 -1466 -1123 -1433
rect -1115 -1466 -1113 -1433
rect -1125 -1468 -1113 -1466
rect -1125 -1501 -1123 -1468
rect -1115 -1501 -1113 -1468
rect -1107 -1501 -1105 -1433
rect -1091 -1501 -1089 -1433
rect -1083 -1501 -1081 -1433
rect -1073 -1501 -1071 -1433
rect -1065 -1501 -1063 -1433
rect -1049 -1501 -1047 -1433
rect -1041 -1501 -1039 -1433
rect -930 -1501 -928 -1433
rect -920 -1501 -918 -1433
rect -904 -1501 -902 -1433
rect -896 -1501 -894 -1433
rect -880 -1501 -878 -1433
rect -872 -1501 -870 -1433
rect -862 -1501 -860 -1433
rect -854 -1501 -852 -1433
rect -838 -1501 -836 -1433
rect -830 -1466 -828 -1433
rect -820 -1466 -818 -1433
rect -830 -1468 -818 -1466
rect -830 -1501 -828 -1468
rect -820 -1501 -818 -1468
rect -812 -1501 -810 -1433
rect -796 -1501 -794 -1433
rect -788 -1501 -786 -1433
rect -778 -1501 -776 -1433
rect -770 -1501 -768 -1433
rect -754 -1501 -752 -1433
rect -746 -1501 -744 -1433
rect -572 -1501 -570 -1433
rect -562 -1501 -560 -1433
rect -546 -1501 -544 -1433
rect -538 -1501 -536 -1433
rect -522 -1501 -520 -1433
rect -514 -1501 -512 -1433
rect -504 -1501 -502 -1433
rect -496 -1501 -494 -1433
rect -480 -1501 -478 -1433
rect -472 -1466 -470 -1433
rect -462 -1466 -460 -1433
rect -472 -1468 -460 -1466
rect -472 -1501 -470 -1468
rect -462 -1501 -460 -1468
rect -454 -1501 -452 -1433
rect -438 -1501 -436 -1433
rect -430 -1501 -428 -1433
rect -420 -1501 -418 -1433
rect -412 -1501 -410 -1433
rect -396 -1501 -394 -1433
rect -388 -1501 -386 -1433
rect -214 -1501 -212 -1433
rect -204 -1501 -202 -1433
rect -188 -1501 -186 -1433
rect -180 -1501 -178 -1433
rect -164 -1501 -162 -1433
rect -156 -1501 -154 -1433
rect -146 -1501 -144 -1433
rect -138 -1501 -136 -1433
rect -122 -1501 -120 -1433
rect -114 -1466 -112 -1433
rect -104 -1466 -102 -1433
rect -114 -1468 -102 -1466
rect -114 -1501 -112 -1468
rect -104 -1501 -102 -1468
rect -96 -1501 -94 -1433
rect -80 -1501 -78 -1433
rect -72 -1501 -70 -1433
rect -62 -1501 -60 -1433
rect -54 -1501 -52 -1433
rect -38 -1501 -36 -1433
rect -30 -1501 -28 -1433
rect 144 -1501 146 -1433
rect 154 -1501 156 -1433
rect 170 -1501 172 -1433
rect 178 -1501 180 -1433
rect 194 -1501 196 -1433
rect 202 -1501 204 -1433
rect 212 -1501 214 -1433
rect 220 -1501 222 -1433
rect 236 -1501 238 -1433
rect 244 -1466 246 -1433
rect 254 -1466 256 -1433
rect 244 -1468 256 -1466
rect 244 -1501 246 -1468
rect 254 -1501 256 -1468
rect 262 -1501 264 -1433
rect 278 -1501 280 -1433
rect 286 -1501 288 -1433
rect 296 -1501 298 -1433
rect 304 -1501 306 -1433
rect 320 -1501 322 -1433
rect 328 -1501 330 -1433
rect 500 -1501 502 -1433
rect 510 -1501 512 -1433
rect 526 -1501 528 -1433
rect 534 -1501 536 -1433
rect 550 -1501 552 -1433
rect 558 -1501 560 -1433
rect 568 -1501 570 -1433
rect 576 -1501 578 -1433
rect 592 -1501 594 -1433
rect 600 -1466 602 -1433
rect 610 -1466 612 -1433
rect 600 -1468 612 -1466
rect 600 -1501 602 -1468
rect 610 -1501 612 -1468
rect 618 -1501 620 -1433
rect 634 -1501 636 -1433
rect 642 -1501 644 -1433
rect 652 -1501 654 -1433
rect 660 -1501 662 -1433
rect 676 -1501 678 -1433
rect 684 -1501 686 -1433
rect 858 -1501 860 -1433
rect 868 -1501 870 -1433
rect 884 -1501 886 -1433
rect 892 -1501 894 -1433
rect 908 -1501 910 -1433
rect 916 -1501 918 -1433
rect 926 -1501 928 -1433
rect 934 -1501 936 -1433
rect 950 -1501 952 -1433
rect 958 -1466 960 -1433
rect 968 -1466 970 -1433
rect 958 -1468 970 -1466
rect 958 -1501 960 -1468
rect 968 -1501 970 -1468
rect 976 -1501 978 -1433
rect 992 -1501 994 -1433
rect 1000 -1501 1002 -1433
rect 1010 -1501 1012 -1433
rect 1018 -1501 1020 -1433
rect 1034 -1501 1036 -1433
rect 1042 -1501 1044 -1433
rect -1225 -1507 -1223 -1505
rect -1215 -1507 -1213 -1505
rect -1199 -1507 -1197 -1505
rect -1191 -1507 -1189 -1505
rect -1175 -1507 -1173 -1505
rect -1167 -1507 -1165 -1505
rect -1157 -1507 -1155 -1505
rect -1149 -1507 -1147 -1505
rect -1133 -1507 -1131 -1505
rect -1125 -1507 -1123 -1505
rect -1115 -1507 -1113 -1505
rect -1107 -1507 -1105 -1505
rect -1091 -1507 -1089 -1505
rect -1083 -1507 -1081 -1505
rect -1073 -1507 -1071 -1505
rect -1065 -1507 -1063 -1505
rect -1049 -1507 -1047 -1505
rect -1041 -1507 -1039 -1505
rect -930 -1507 -928 -1505
rect -920 -1507 -918 -1505
rect -904 -1507 -902 -1505
rect -896 -1507 -894 -1505
rect -880 -1507 -878 -1505
rect -872 -1507 -870 -1505
rect -862 -1507 -860 -1505
rect -854 -1507 -852 -1505
rect -838 -1507 -836 -1505
rect -830 -1507 -828 -1505
rect -820 -1507 -818 -1505
rect -812 -1507 -810 -1505
rect -796 -1507 -794 -1505
rect -788 -1507 -786 -1505
rect -778 -1507 -776 -1505
rect -770 -1507 -768 -1505
rect -754 -1507 -752 -1505
rect -746 -1507 -744 -1505
rect -572 -1507 -570 -1505
rect -562 -1507 -560 -1505
rect -546 -1507 -544 -1505
rect -538 -1507 -536 -1505
rect -522 -1507 -520 -1505
rect -514 -1507 -512 -1505
rect -504 -1507 -502 -1505
rect -496 -1507 -494 -1505
rect -480 -1507 -478 -1505
rect -472 -1507 -470 -1505
rect -462 -1507 -460 -1505
rect -454 -1507 -452 -1505
rect -438 -1507 -436 -1505
rect -430 -1507 -428 -1505
rect -420 -1507 -418 -1505
rect -412 -1507 -410 -1505
rect -396 -1507 -394 -1505
rect -388 -1507 -386 -1505
rect -214 -1507 -212 -1505
rect -204 -1507 -202 -1505
rect -188 -1507 -186 -1505
rect -180 -1507 -178 -1505
rect -164 -1507 -162 -1505
rect -156 -1507 -154 -1505
rect -146 -1507 -144 -1505
rect -138 -1507 -136 -1505
rect -122 -1507 -120 -1505
rect -114 -1507 -112 -1505
rect -104 -1507 -102 -1505
rect -96 -1507 -94 -1505
rect -80 -1507 -78 -1505
rect -72 -1507 -70 -1505
rect -62 -1507 -60 -1505
rect -54 -1507 -52 -1505
rect -38 -1507 -36 -1505
rect -30 -1507 -28 -1505
rect 144 -1507 146 -1505
rect 154 -1507 156 -1505
rect 170 -1507 172 -1505
rect 178 -1507 180 -1505
rect 194 -1507 196 -1505
rect 202 -1507 204 -1505
rect 212 -1507 214 -1505
rect 220 -1507 222 -1505
rect 236 -1507 238 -1505
rect 244 -1507 246 -1505
rect 254 -1507 256 -1505
rect 262 -1507 264 -1505
rect 278 -1507 280 -1505
rect 286 -1507 288 -1505
rect 296 -1507 298 -1505
rect 304 -1507 306 -1505
rect 320 -1507 322 -1505
rect 328 -1507 330 -1505
rect 500 -1507 502 -1505
rect 510 -1507 512 -1505
rect 526 -1507 528 -1505
rect 534 -1507 536 -1505
rect 550 -1507 552 -1505
rect 558 -1507 560 -1505
rect 568 -1507 570 -1505
rect 576 -1507 578 -1505
rect 592 -1507 594 -1505
rect 600 -1507 602 -1505
rect 610 -1507 612 -1505
rect 618 -1507 620 -1505
rect 634 -1507 636 -1505
rect 642 -1507 644 -1505
rect 652 -1507 654 -1505
rect 660 -1507 662 -1505
rect 676 -1507 678 -1505
rect 684 -1507 686 -1505
rect 858 -1507 860 -1505
rect 868 -1507 870 -1505
rect 884 -1507 886 -1505
rect 892 -1507 894 -1505
rect 908 -1507 910 -1505
rect 916 -1507 918 -1505
rect 926 -1507 928 -1505
rect 934 -1507 936 -1505
rect 950 -1507 952 -1505
rect 958 -1507 960 -1505
rect 968 -1507 970 -1505
rect 976 -1507 978 -1505
rect 992 -1507 994 -1505
rect 1000 -1507 1002 -1505
rect 1010 -1507 1012 -1505
rect 1018 -1507 1020 -1505
rect 1034 -1507 1036 -1505
rect 1042 -1507 1044 -1505
rect -1225 -1596 -1223 -1594
rect -1215 -1596 -1213 -1594
rect -1199 -1596 -1197 -1594
rect -1191 -1596 -1189 -1594
rect -1175 -1596 -1173 -1594
rect -1167 -1596 -1165 -1594
rect -1157 -1596 -1155 -1594
rect -1149 -1596 -1147 -1594
rect -1133 -1596 -1131 -1594
rect -1125 -1596 -1123 -1594
rect -1115 -1596 -1113 -1594
rect -1107 -1596 -1105 -1594
rect -1091 -1596 -1089 -1594
rect -1083 -1596 -1081 -1594
rect -1073 -1596 -1071 -1594
rect -1065 -1596 -1063 -1594
rect -1049 -1596 -1047 -1594
rect -1041 -1596 -1039 -1594
rect -930 -1596 -928 -1594
rect -920 -1596 -918 -1594
rect -904 -1596 -902 -1594
rect -896 -1596 -894 -1594
rect -880 -1596 -878 -1594
rect -872 -1596 -870 -1594
rect -862 -1596 -860 -1594
rect -854 -1596 -852 -1594
rect -838 -1596 -836 -1594
rect -830 -1596 -828 -1594
rect -820 -1596 -818 -1594
rect -812 -1596 -810 -1594
rect -796 -1596 -794 -1594
rect -788 -1596 -786 -1594
rect -778 -1596 -776 -1594
rect -770 -1596 -768 -1594
rect -754 -1596 -752 -1594
rect -746 -1596 -744 -1594
rect -572 -1596 -570 -1594
rect -562 -1596 -560 -1594
rect -546 -1596 -544 -1594
rect -538 -1596 -536 -1594
rect -522 -1596 -520 -1594
rect -514 -1596 -512 -1594
rect -504 -1596 -502 -1594
rect -496 -1596 -494 -1594
rect -480 -1596 -478 -1594
rect -472 -1596 -470 -1594
rect -462 -1596 -460 -1594
rect -454 -1596 -452 -1594
rect -438 -1596 -436 -1594
rect -430 -1596 -428 -1594
rect -420 -1596 -418 -1594
rect -412 -1596 -410 -1594
rect -396 -1596 -394 -1594
rect -388 -1596 -386 -1594
rect -214 -1596 -212 -1594
rect -204 -1596 -202 -1594
rect -188 -1596 -186 -1594
rect -180 -1596 -178 -1594
rect -164 -1596 -162 -1594
rect -156 -1596 -154 -1594
rect -146 -1596 -144 -1594
rect -138 -1596 -136 -1594
rect -122 -1596 -120 -1594
rect -114 -1596 -112 -1594
rect -104 -1596 -102 -1594
rect -96 -1596 -94 -1594
rect -80 -1596 -78 -1594
rect -72 -1596 -70 -1594
rect -62 -1596 -60 -1594
rect -54 -1596 -52 -1594
rect -38 -1596 -36 -1594
rect -30 -1596 -28 -1594
rect 144 -1596 146 -1594
rect 154 -1596 156 -1594
rect 170 -1596 172 -1594
rect 178 -1596 180 -1594
rect 194 -1596 196 -1594
rect 202 -1596 204 -1594
rect 212 -1596 214 -1594
rect 220 -1596 222 -1594
rect 236 -1596 238 -1594
rect 244 -1596 246 -1594
rect 254 -1596 256 -1594
rect 262 -1596 264 -1594
rect 278 -1596 280 -1594
rect 286 -1596 288 -1594
rect 296 -1596 298 -1594
rect 304 -1596 306 -1594
rect 320 -1596 322 -1594
rect 328 -1596 330 -1594
rect 500 -1596 502 -1594
rect 510 -1596 512 -1594
rect 526 -1596 528 -1594
rect 534 -1596 536 -1594
rect 550 -1596 552 -1594
rect 558 -1596 560 -1594
rect 568 -1596 570 -1594
rect 576 -1596 578 -1594
rect 592 -1596 594 -1594
rect 600 -1596 602 -1594
rect 610 -1596 612 -1594
rect 618 -1596 620 -1594
rect 634 -1596 636 -1594
rect 642 -1596 644 -1594
rect 652 -1596 654 -1594
rect 660 -1596 662 -1594
rect 676 -1596 678 -1594
rect 684 -1596 686 -1594
rect 858 -1596 860 -1594
rect 868 -1596 870 -1594
rect 884 -1596 886 -1594
rect 892 -1596 894 -1594
rect 908 -1596 910 -1594
rect 916 -1596 918 -1594
rect 926 -1596 928 -1594
rect 934 -1596 936 -1594
rect 950 -1596 952 -1594
rect 958 -1596 960 -1594
rect 968 -1596 970 -1594
rect 976 -1596 978 -1594
rect 992 -1596 994 -1594
rect 1000 -1596 1002 -1594
rect 1010 -1596 1012 -1594
rect 1018 -1596 1020 -1594
rect 1034 -1596 1036 -1594
rect 1042 -1596 1044 -1594
rect 1216 -1596 1218 -1594
rect 1226 -1596 1228 -1594
rect 1242 -1596 1244 -1594
rect 1250 -1596 1252 -1594
rect 1266 -1596 1268 -1594
rect 1274 -1596 1276 -1594
rect 1284 -1596 1286 -1594
rect 1292 -1596 1294 -1594
rect 1308 -1596 1310 -1594
rect 1316 -1596 1318 -1594
rect 1326 -1596 1328 -1594
rect 1334 -1596 1336 -1594
rect 1350 -1596 1352 -1594
rect 1358 -1596 1360 -1594
rect 1368 -1596 1370 -1594
rect 1376 -1596 1378 -1594
rect 1392 -1596 1394 -1594
rect 1400 -1596 1402 -1594
rect -1225 -1672 -1223 -1604
rect -1215 -1672 -1213 -1604
rect -1199 -1672 -1197 -1604
rect -1191 -1672 -1189 -1604
rect -1175 -1672 -1173 -1604
rect -1167 -1672 -1165 -1604
rect -1157 -1672 -1155 -1604
rect -1149 -1672 -1147 -1604
rect -1133 -1672 -1131 -1604
rect -1125 -1637 -1123 -1604
rect -1115 -1637 -1113 -1604
rect -1125 -1639 -1113 -1637
rect -1125 -1672 -1123 -1639
rect -1115 -1672 -1113 -1639
rect -1107 -1672 -1105 -1604
rect -1091 -1672 -1089 -1604
rect -1083 -1672 -1081 -1604
rect -1073 -1672 -1071 -1604
rect -1065 -1672 -1063 -1604
rect -1049 -1672 -1047 -1604
rect -1041 -1672 -1039 -1604
rect -930 -1672 -928 -1604
rect -920 -1672 -918 -1604
rect -904 -1672 -902 -1604
rect -896 -1672 -894 -1604
rect -880 -1672 -878 -1604
rect -872 -1672 -870 -1604
rect -862 -1672 -860 -1604
rect -854 -1672 -852 -1604
rect -838 -1672 -836 -1604
rect -830 -1637 -828 -1604
rect -820 -1637 -818 -1604
rect -830 -1639 -818 -1637
rect -830 -1672 -828 -1639
rect -820 -1672 -818 -1639
rect -812 -1672 -810 -1604
rect -796 -1672 -794 -1604
rect -788 -1672 -786 -1604
rect -778 -1672 -776 -1604
rect -770 -1672 -768 -1604
rect -754 -1672 -752 -1604
rect -746 -1672 -744 -1604
rect -572 -1672 -570 -1604
rect -562 -1672 -560 -1604
rect -546 -1672 -544 -1604
rect -538 -1672 -536 -1604
rect -522 -1672 -520 -1604
rect -514 -1672 -512 -1604
rect -504 -1672 -502 -1604
rect -496 -1672 -494 -1604
rect -480 -1672 -478 -1604
rect -472 -1637 -470 -1604
rect -462 -1637 -460 -1604
rect -472 -1639 -460 -1637
rect -472 -1672 -470 -1639
rect -462 -1672 -460 -1639
rect -454 -1672 -452 -1604
rect -438 -1672 -436 -1604
rect -430 -1672 -428 -1604
rect -420 -1672 -418 -1604
rect -412 -1672 -410 -1604
rect -396 -1672 -394 -1604
rect -388 -1672 -386 -1604
rect -214 -1672 -212 -1604
rect -204 -1672 -202 -1604
rect -188 -1672 -186 -1604
rect -180 -1672 -178 -1604
rect -164 -1672 -162 -1604
rect -156 -1672 -154 -1604
rect -146 -1672 -144 -1604
rect -138 -1672 -136 -1604
rect -122 -1672 -120 -1604
rect -114 -1637 -112 -1604
rect -104 -1637 -102 -1604
rect -114 -1639 -102 -1637
rect -114 -1672 -112 -1639
rect -104 -1672 -102 -1639
rect -96 -1672 -94 -1604
rect -80 -1672 -78 -1604
rect -72 -1672 -70 -1604
rect -62 -1672 -60 -1604
rect -54 -1672 -52 -1604
rect -38 -1672 -36 -1604
rect -30 -1672 -28 -1604
rect 144 -1672 146 -1604
rect 154 -1672 156 -1604
rect 170 -1672 172 -1604
rect 178 -1672 180 -1604
rect 194 -1672 196 -1604
rect 202 -1672 204 -1604
rect 212 -1672 214 -1604
rect 220 -1672 222 -1604
rect 236 -1672 238 -1604
rect 244 -1637 246 -1604
rect 254 -1637 256 -1604
rect 244 -1639 256 -1637
rect 244 -1672 246 -1639
rect 254 -1672 256 -1639
rect 262 -1672 264 -1604
rect 278 -1672 280 -1604
rect 286 -1672 288 -1604
rect 296 -1672 298 -1604
rect 304 -1672 306 -1604
rect 320 -1672 322 -1604
rect 328 -1672 330 -1604
rect 500 -1672 502 -1604
rect 510 -1672 512 -1604
rect 526 -1672 528 -1604
rect 534 -1672 536 -1604
rect 550 -1672 552 -1604
rect 558 -1672 560 -1604
rect 568 -1672 570 -1604
rect 576 -1672 578 -1604
rect 592 -1672 594 -1604
rect 600 -1637 602 -1604
rect 610 -1637 612 -1604
rect 600 -1639 612 -1637
rect 600 -1672 602 -1639
rect 610 -1672 612 -1639
rect 618 -1672 620 -1604
rect 634 -1672 636 -1604
rect 642 -1672 644 -1604
rect 652 -1672 654 -1604
rect 660 -1672 662 -1604
rect 676 -1672 678 -1604
rect 684 -1672 686 -1604
rect 858 -1672 860 -1604
rect 868 -1672 870 -1604
rect 884 -1672 886 -1604
rect 892 -1672 894 -1604
rect 908 -1672 910 -1604
rect 916 -1672 918 -1604
rect 926 -1672 928 -1604
rect 934 -1672 936 -1604
rect 950 -1672 952 -1604
rect 958 -1637 960 -1604
rect 968 -1637 970 -1604
rect 958 -1639 970 -1637
rect 958 -1672 960 -1639
rect 968 -1672 970 -1639
rect 976 -1672 978 -1604
rect 992 -1672 994 -1604
rect 1000 -1672 1002 -1604
rect 1010 -1672 1012 -1604
rect 1018 -1672 1020 -1604
rect 1034 -1672 1036 -1604
rect 1042 -1672 1044 -1604
rect 1216 -1672 1218 -1604
rect 1226 -1672 1228 -1604
rect 1242 -1672 1244 -1604
rect 1250 -1672 1252 -1604
rect 1266 -1672 1268 -1604
rect 1274 -1672 1276 -1604
rect 1284 -1672 1286 -1604
rect 1292 -1672 1294 -1604
rect 1308 -1672 1310 -1604
rect 1316 -1637 1318 -1604
rect 1326 -1637 1328 -1604
rect 1316 -1639 1328 -1637
rect 1316 -1672 1318 -1639
rect 1326 -1672 1328 -1639
rect 1334 -1672 1336 -1604
rect 1350 -1672 1352 -1604
rect 1358 -1672 1360 -1604
rect 1368 -1672 1370 -1604
rect 1376 -1672 1378 -1604
rect 1392 -1672 1394 -1604
rect 1400 -1672 1402 -1604
rect -1225 -1678 -1223 -1676
rect -1215 -1678 -1213 -1676
rect -1199 -1678 -1197 -1676
rect -1191 -1678 -1189 -1676
rect -1175 -1678 -1173 -1676
rect -1167 -1678 -1165 -1676
rect -1157 -1678 -1155 -1676
rect -1149 -1678 -1147 -1676
rect -1133 -1678 -1131 -1676
rect -1125 -1678 -1123 -1676
rect -1115 -1678 -1113 -1676
rect -1107 -1678 -1105 -1676
rect -1091 -1678 -1089 -1676
rect -1083 -1678 -1081 -1676
rect -1073 -1678 -1071 -1676
rect -1065 -1678 -1063 -1676
rect -1049 -1678 -1047 -1676
rect -1041 -1678 -1039 -1676
rect -930 -1678 -928 -1676
rect -920 -1678 -918 -1676
rect -904 -1678 -902 -1676
rect -896 -1678 -894 -1676
rect -880 -1678 -878 -1676
rect -872 -1678 -870 -1676
rect -862 -1678 -860 -1676
rect -854 -1678 -852 -1676
rect -838 -1678 -836 -1676
rect -830 -1678 -828 -1676
rect -820 -1678 -818 -1676
rect -812 -1678 -810 -1676
rect -796 -1678 -794 -1676
rect -788 -1678 -786 -1676
rect -778 -1678 -776 -1676
rect -770 -1678 -768 -1676
rect -754 -1678 -752 -1676
rect -746 -1678 -744 -1676
rect -572 -1678 -570 -1676
rect -562 -1678 -560 -1676
rect -546 -1678 -544 -1676
rect -538 -1678 -536 -1676
rect -522 -1678 -520 -1676
rect -514 -1678 -512 -1676
rect -504 -1678 -502 -1676
rect -496 -1678 -494 -1676
rect -480 -1678 -478 -1676
rect -472 -1678 -470 -1676
rect -462 -1678 -460 -1676
rect -454 -1678 -452 -1676
rect -438 -1678 -436 -1676
rect -430 -1678 -428 -1676
rect -420 -1678 -418 -1676
rect -412 -1678 -410 -1676
rect -396 -1678 -394 -1676
rect -388 -1678 -386 -1676
rect -214 -1678 -212 -1676
rect -204 -1678 -202 -1676
rect -188 -1678 -186 -1676
rect -180 -1678 -178 -1676
rect -164 -1678 -162 -1676
rect -156 -1678 -154 -1676
rect -146 -1678 -144 -1676
rect -138 -1678 -136 -1676
rect -122 -1678 -120 -1676
rect -114 -1678 -112 -1676
rect -104 -1678 -102 -1676
rect -96 -1678 -94 -1676
rect -80 -1678 -78 -1676
rect -72 -1678 -70 -1676
rect -62 -1678 -60 -1676
rect -54 -1678 -52 -1676
rect -38 -1678 -36 -1676
rect -30 -1678 -28 -1676
rect 144 -1678 146 -1676
rect 154 -1678 156 -1676
rect 170 -1678 172 -1676
rect 178 -1678 180 -1676
rect 194 -1678 196 -1676
rect 202 -1678 204 -1676
rect 212 -1678 214 -1676
rect 220 -1678 222 -1676
rect 236 -1678 238 -1676
rect 244 -1678 246 -1676
rect 254 -1678 256 -1676
rect 262 -1678 264 -1676
rect 278 -1678 280 -1676
rect 286 -1678 288 -1676
rect 296 -1678 298 -1676
rect 304 -1678 306 -1676
rect 320 -1678 322 -1676
rect 328 -1678 330 -1676
rect 500 -1678 502 -1676
rect 510 -1678 512 -1676
rect 526 -1678 528 -1676
rect 534 -1678 536 -1676
rect 550 -1678 552 -1676
rect 558 -1678 560 -1676
rect 568 -1678 570 -1676
rect 576 -1678 578 -1676
rect 592 -1678 594 -1676
rect 600 -1678 602 -1676
rect 610 -1678 612 -1676
rect 618 -1678 620 -1676
rect 634 -1678 636 -1676
rect 642 -1678 644 -1676
rect 652 -1678 654 -1676
rect 660 -1678 662 -1676
rect 676 -1678 678 -1676
rect 684 -1678 686 -1676
rect 858 -1678 860 -1676
rect 868 -1678 870 -1676
rect 884 -1678 886 -1676
rect 892 -1678 894 -1676
rect 908 -1678 910 -1676
rect 916 -1678 918 -1676
rect 926 -1678 928 -1676
rect 934 -1678 936 -1676
rect 950 -1678 952 -1676
rect 958 -1678 960 -1676
rect 968 -1678 970 -1676
rect 976 -1678 978 -1676
rect 992 -1678 994 -1676
rect 1000 -1678 1002 -1676
rect 1010 -1678 1012 -1676
rect 1018 -1678 1020 -1676
rect 1034 -1678 1036 -1676
rect 1042 -1678 1044 -1676
rect 1216 -1678 1218 -1676
rect 1226 -1678 1228 -1676
rect 1242 -1678 1244 -1676
rect 1250 -1678 1252 -1676
rect 1266 -1678 1268 -1676
rect 1274 -1678 1276 -1676
rect 1284 -1678 1286 -1676
rect 1292 -1678 1294 -1676
rect 1308 -1678 1310 -1676
rect 1316 -1678 1318 -1676
rect 1326 -1678 1328 -1676
rect 1334 -1678 1336 -1676
rect 1350 -1678 1352 -1676
rect 1358 -1678 1360 -1676
rect 1368 -1678 1370 -1676
rect 1376 -1678 1378 -1676
rect 1392 -1678 1394 -1676
rect 1400 -1678 1402 -1676
rect -1554 -1767 -1552 -1765
rect -1544 -1767 -1542 -1765
rect -1528 -1767 -1526 -1765
rect -1520 -1767 -1518 -1765
rect -1504 -1767 -1502 -1765
rect -1496 -1767 -1494 -1765
rect -1486 -1767 -1484 -1765
rect -1478 -1767 -1476 -1765
rect -1462 -1767 -1460 -1765
rect -1454 -1767 -1452 -1765
rect -1444 -1767 -1442 -1765
rect -1436 -1767 -1434 -1765
rect -1420 -1767 -1418 -1765
rect -1412 -1767 -1410 -1765
rect -1402 -1767 -1400 -1765
rect -1394 -1767 -1392 -1765
rect -1378 -1767 -1376 -1765
rect -1370 -1767 -1368 -1765
rect -1225 -1767 -1223 -1765
rect -1215 -1767 -1213 -1765
rect -1199 -1767 -1197 -1765
rect -1191 -1767 -1189 -1765
rect -1175 -1767 -1173 -1765
rect -1167 -1767 -1165 -1765
rect -1157 -1767 -1155 -1765
rect -1149 -1767 -1147 -1765
rect -1133 -1767 -1131 -1765
rect -1125 -1767 -1123 -1765
rect -1115 -1767 -1113 -1765
rect -1107 -1767 -1105 -1765
rect -1091 -1767 -1089 -1765
rect -1083 -1767 -1081 -1765
rect -1073 -1767 -1071 -1765
rect -1065 -1767 -1063 -1765
rect -1049 -1767 -1047 -1765
rect -1041 -1767 -1039 -1765
rect -930 -1767 -928 -1765
rect -920 -1767 -918 -1765
rect -904 -1767 -902 -1765
rect -896 -1767 -894 -1765
rect -880 -1767 -878 -1765
rect -872 -1767 -870 -1765
rect -862 -1767 -860 -1765
rect -854 -1767 -852 -1765
rect -838 -1767 -836 -1765
rect -830 -1767 -828 -1765
rect -820 -1767 -818 -1765
rect -812 -1767 -810 -1765
rect -796 -1767 -794 -1765
rect -788 -1767 -786 -1765
rect -778 -1767 -776 -1765
rect -770 -1767 -768 -1765
rect -754 -1767 -752 -1765
rect -746 -1767 -744 -1765
rect -572 -1767 -570 -1765
rect -562 -1767 -560 -1765
rect -546 -1767 -544 -1765
rect -538 -1767 -536 -1765
rect -522 -1767 -520 -1765
rect -514 -1767 -512 -1765
rect -504 -1767 -502 -1765
rect -496 -1767 -494 -1765
rect -480 -1767 -478 -1765
rect -472 -1767 -470 -1765
rect -462 -1767 -460 -1765
rect -454 -1767 -452 -1765
rect -438 -1767 -436 -1765
rect -430 -1767 -428 -1765
rect -420 -1767 -418 -1765
rect -412 -1767 -410 -1765
rect -396 -1767 -394 -1765
rect -388 -1767 -386 -1765
rect -214 -1767 -212 -1765
rect -204 -1767 -202 -1765
rect -188 -1767 -186 -1765
rect -180 -1767 -178 -1765
rect -164 -1767 -162 -1765
rect -156 -1767 -154 -1765
rect -146 -1767 -144 -1765
rect -138 -1767 -136 -1765
rect -122 -1767 -120 -1765
rect -114 -1767 -112 -1765
rect -104 -1767 -102 -1765
rect -96 -1767 -94 -1765
rect -80 -1767 -78 -1765
rect -72 -1767 -70 -1765
rect -62 -1767 -60 -1765
rect -54 -1767 -52 -1765
rect -38 -1767 -36 -1765
rect -30 -1767 -28 -1765
rect 144 -1767 146 -1765
rect 154 -1767 156 -1765
rect 170 -1767 172 -1765
rect 178 -1767 180 -1765
rect 194 -1767 196 -1765
rect 202 -1767 204 -1765
rect 212 -1767 214 -1765
rect 220 -1767 222 -1765
rect 236 -1767 238 -1765
rect 244 -1767 246 -1765
rect 254 -1767 256 -1765
rect 262 -1767 264 -1765
rect 278 -1767 280 -1765
rect 286 -1767 288 -1765
rect 296 -1767 298 -1765
rect 304 -1767 306 -1765
rect 320 -1767 322 -1765
rect 328 -1767 330 -1765
rect 500 -1767 502 -1765
rect 510 -1767 512 -1765
rect 526 -1767 528 -1765
rect 534 -1767 536 -1765
rect 550 -1767 552 -1765
rect 558 -1767 560 -1765
rect 568 -1767 570 -1765
rect 576 -1767 578 -1765
rect 592 -1767 594 -1765
rect 600 -1767 602 -1765
rect 610 -1767 612 -1765
rect 618 -1767 620 -1765
rect 634 -1767 636 -1765
rect 642 -1767 644 -1765
rect 652 -1767 654 -1765
rect 660 -1767 662 -1765
rect 676 -1767 678 -1765
rect 684 -1767 686 -1765
rect 858 -1767 860 -1765
rect 868 -1767 870 -1765
rect 884 -1767 886 -1765
rect 892 -1767 894 -1765
rect 908 -1767 910 -1765
rect 916 -1767 918 -1765
rect 926 -1767 928 -1765
rect 934 -1767 936 -1765
rect 950 -1767 952 -1765
rect 958 -1767 960 -1765
rect 968 -1767 970 -1765
rect 976 -1767 978 -1765
rect 992 -1767 994 -1765
rect 1000 -1767 1002 -1765
rect 1010 -1767 1012 -1765
rect 1018 -1767 1020 -1765
rect 1034 -1767 1036 -1765
rect 1042 -1767 1044 -1765
rect 1216 -1767 1218 -1765
rect 1226 -1767 1228 -1765
rect 1242 -1767 1244 -1765
rect 1250 -1767 1252 -1765
rect 1266 -1767 1268 -1765
rect 1274 -1767 1276 -1765
rect 1284 -1767 1286 -1765
rect 1292 -1767 1294 -1765
rect 1308 -1767 1310 -1765
rect 1316 -1767 1318 -1765
rect 1326 -1767 1328 -1765
rect 1334 -1767 1336 -1765
rect 1350 -1767 1352 -1765
rect 1358 -1767 1360 -1765
rect 1368 -1767 1370 -1765
rect 1376 -1767 1378 -1765
rect 1392 -1767 1394 -1765
rect 1400 -1767 1402 -1765
rect -1554 -1843 -1552 -1775
rect -1544 -1843 -1542 -1775
rect -1528 -1843 -1526 -1775
rect -1520 -1843 -1518 -1775
rect -1504 -1843 -1502 -1775
rect -1496 -1843 -1494 -1775
rect -1486 -1843 -1484 -1775
rect -1478 -1843 -1476 -1775
rect -1462 -1843 -1460 -1775
rect -1454 -1808 -1452 -1775
rect -1444 -1808 -1442 -1775
rect -1454 -1810 -1442 -1808
rect -1454 -1843 -1452 -1810
rect -1444 -1843 -1442 -1810
rect -1436 -1843 -1434 -1775
rect -1420 -1843 -1418 -1775
rect -1412 -1843 -1410 -1775
rect -1402 -1843 -1400 -1775
rect -1394 -1843 -1392 -1775
rect -1378 -1843 -1376 -1775
rect -1370 -1843 -1368 -1775
rect -1225 -1843 -1223 -1775
rect -1215 -1843 -1213 -1775
rect -1199 -1843 -1197 -1775
rect -1191 -1843 -1189 -1775
rect -1175 -1843 -1173 -1775
rect -1167 -1843 -1165 -1775
rect -1157 -1843 -1155 -1775
rect -1149 -1843 -1147 -1775
rect -1133 -1843 -1131 -1775
rect -1125 -1808 -1123 -1775
rect -1115 -1808 -1113 -1775
rect -1125 -1810 -1113 -1808
rect -1125 -1843 -1123 -1810
rect -1115 -1843 -1113 -1810
rect -1107 -1843 -1105 -1775
rect -1091 -1843 -1089 -1775
rect -1083 -1843 -1081 -1775
rect -1073 -1843 -1071 -1775
rect -1065 -1843 -1063 -1775
rect -1049 -1843 -1047 -1775
rect -1041 -1843 -1039 -1775
rect -930 -1843 -928 -1775
rect -920 -1843 -918 -1775
rect -904 -1843 -902 -1775
rect -896 -1843 -894 -1775
rect -880 -1843 -878 -1775
rect -872 -1843 -870 -1775
rect -862 -1843 -860 -1775
rect -854 -1843 -852 -1775
rect -838 -1843 -836 -1775
rect -830 -1808 -828 -1775
rect -820 -1808 -818 -1775
rect -830 -1810 -818 -1808
rect -830 -1843 -828 -1810
rect -820 -1843 -818 -1810
rect -812 -1843 -810 -1775
rect -796 -1843 -794 -1775
rect -788 -1843 -786 -1775
rect -778 -1843 -776 -1775
rect -770 -1843 -768 -1775
rect -754 -1843 -752 -1775
rect -746 -1843 -744 -1775
rect -572 -1843 -570 -1775
rect -562 -1843 -560 -1775
rect -546 -1843 -544 -1775
rect -538 -1843 -536 -1775
rect -522 -1843 -520 -1775
rect -514 -1843 -512 -1775
rect -504 -1843 -502 -1775
rect -496 -1843 -494 -1775
rect -480 -1843 -478 -1775
rect -472 -1808 -470 -1775
rect -462 -1808 -460 -1775
rect -472 -1810 -460 -1808
rect -472 -1843 -470 -1810
rect -462 -1843 -460 -1810
rect -454 -1843 -452 -1775
rect -438 -1843 -436 -1775
rect -430 -1843 -428 -1775
rect -420 -1843 -418 -1775
rect -412 -1843 -410 -1775
rect -396 -1843 -394 -1775
rect -388 -1843 -386 -1775
rect -214 -1843 -212 -1775
rect -204 -1843 -202 -1775
rect -188 -1843 -186 -1775
rect -180 -1843 -178 -1775
rect -164 -1843 -162 -1775
rect -156 -1843 -154 -1775
rect -146 -1843 -144 -1775
rect -138 -1843 -136 -1775
rect -122 -1843 -120 -1775
rect -114 -1808 -112 -1775
rect -104 -1808 -102 -1775
rect -114 -1810 -102 -1808
rect -114 -1843 -112 -1810
rect -104 -1843 -102 -1810
rect -96 -1843 -94 -1775
rect -80 -1843 -78 -1775
rect -72 -1843 -70 -1775
rect -62 -1843 -60 -1775
rect -54 -1843 -52 -1775
rect -38 -1843 -36 -1775
rect -30 -1843 -28 -1775
rect 144 -1843 146 -1775
rect 154 -1843 156 -1775
rect 170 -1843 172 -1775
rect 178 -1843 180 -1775
rect 194 -1843 196 -1775
rect 202 -1843 204 -1775
rect 212 -1843 214 -1775
rect 220 -1843 222 -1775
rect 236 -1843 238 -1775
rect 244 -1808 246 -1775
rect 254 -1808 256 -1775
rect 244 -1810 256 -1808
rect 244 -1843 246 -1810
rect 254 -1843 256 -1810
rect 262 -1843 264 -1775
rect 278 -1843 280 -1775
rect 286 -1843 288 -1775
rect 296 -1843 298 -1775
rect 304 -1843 306 -1775
rect 320 -1843 322 -1775
rect 328 -1843 330 -1775
rect 500 -1843 502 -1775
rect 510 -1843 512 -1775
rect 526 -1843 528 -1775
rect 534 -1843 536 -1775
rect 550 -1843 552 -1775
rect 558 -1843 560 -1775
rect 568 -1843 570 -1775
rect 576 -1843 578 -1775
rect 592 -1843 594 -1775
rect 600 -1808 602 -1775
rect 610 -1808 612 -1775
rect 600 -1810 612 -1808
rect 600 -1843 602 -1810
rect 610 -1843 612 -1810
rect 618 -1843 620 -1775
rect 634 -1843 636 -1775
rect 642 -1843 644 -1775
rect 652 -1843 654 -1775
rect 660 -1843 662 -1775
rect 676 -1843 678 -1775
rect 684 -1843 686 -1775
rect 858 -1843 860 -1775
rect 868 -1843 870 -1775
rect 884 -1843 886 -1775
rect 892 -1843 894 -1775
rect 908 -1843 910 -1775
rect 916 -1843 918 -1775
rect 926 -1843 928 -1775
rect 934 -1843 936 -1775
rect 950 -1843 952 -1775
rect 958 -1808 960 -1775
rect 968 -1808 970 -1775
rect 958 -1810 970 -1808
rect 958 -1843 960 -1810
rect 968 -1843 970 -1810
rect 976 -1843 978 -1775
rect 992 -1843 994 -1775
rect 1000 -1843 1002 -1775
rect 1010 -1843 1012 -1775
rect 1018 -1843 1020 -1775
rect 1034 -1843 1036 -1775
rect 1042 -1843 1044 -1775
rect 1216 -1843 1218 -1775
rect 1226 -1843 1228 -1775
rect 1242 -1843 1244 -1775
rect 1250 -1843 1252 -1775
rect 1266 -1843 1268 -1775
rect 1274 -1843 1276 -1775
rect 1284 -1843 1286 -1775
rect 1292 -1843 1294 -1775
rect 1308 -1843 1310 -1775
rect 1316 -1808 1318 -1775
rect 1326 -1808 1328 -1775
rect 1316 -1810 1328 -1808
rect 1316 -1843 1318 -1810
rect 1326 -1843 1328 -1810
rect 1334 -1843 1336 -1775
rect 1350 -1843 1352 -1775
rect 1358 -1843 1360 -1775
rect 1368 -1843 1370 -1775
rect 1376 -1843 1378 -1775
rect 1392 -1843 1394 -1775
rect 1400 -1843 1402 -1775
rect -1554 -1849 -1552 -1847
rect -1544 -1849 -1542 -1847
rect -1528 -1849 -1526 -1847
rect -1520 -1849 -1518 -1847
rect -1504 -1849 -1502 -1847
rect -1496 -1849 -1494 -1847
rect -1486 -1849 -1484 -1847
rect -1478 -1849 -1476 -1847
rect -1462 -1849 -1460 -1847
rect -1454 -1849 -1452 -1847
rect -1444 -1849 -1442 -1847
rect -1436 -1849 -1434 -1847
rect -1420 -1849 -1418 -1847
rect -1412 -1849 -1410 -1847
rect -1402 -1849 -1400 -1847
rect -1394 -1849 -1392 -1847
rect -1378 -1849 -1376 -1847
rect -1370 -1849 -1368 -1847
rect -1225 -1849 -1223 -1847
rect -1215 -1849 -1213 -1847
rect -1199 -1849 -1197 -1847
rect -1191 -1849 -1189 -1847
rect -1175 -1849 -1173 -1847
rect -1167 -1849 -1165 -1847
rect -1157 -1849 -1155 -1847
rect -1149 -1849 -1147 -1847
rect -1133 -1849 -1131 -1847
rect -1125 -1849 -1123 -1847
rect -1115 -1849 -1113 -1847
rect -1107 -1849 -1105 -1847
rect -1091 -1849 -1089 -1847
rect -1083 -1849 -1081 -1847
rect -1073 -1849 -1071 -1847
rect -1065 -1849 -1063 -1847
rect -1049 -1849 -1047 -1847
rect -1041 -1849 -1039 -1847
rect -930 -1849 -928 -1847
rect -920 -1849 -918 -1847
rect -904 -1849 -902 -1847
rect -896 -1849 -894 -1847
rect -880 -1849 -878 -1847
rect -872 -1849 -870 -1847
rect -862 -1849 -860 -1847
rect -854 -1849 -852 -1847
rect -838 -1849 -836 -1847
rect -830 -1849 -828 -1847
rect -820 -1849 -818 -1847
rect -812 -1849 -810 -1847
rect -796 -1849 -794 -1847
rect -788 -1849 -786 -1847
rect -778 -1849 -776 -1847
rect -770 -1849 -768 -1847
rect -754 -1849 -752 -1847
rect -746 -1849 -744 -1847
rect -572 -1849 -570 -1847
rect -562 -1849 -560 -1847
rect -546 -1849 -544 -1847
rect -538 -1849 -536 -1847
rect -522 -1849 -520 -1847
rect -514 -1849 -512 -1847
rect -504 -1849 -502 -1847
rect -496 -1849 -494 -1847
rect -480 -1849 -478 -1847
rect -472 -1849 -470 -1847
rect -462 -1849 -460 -1847
rect -454 -1849 -452 -1847
rect -438 -1849 -436 -1847
rect -430 -1849 -428 -1847
rect -420 -1849 -418 -1847
rect -412 -1849 -410 -1847
rect -396 -1849 -394 -1847
rect -388 -1849 -386 -1847
rect -214 -1849 -212 -1847
rect -204 -1849 -202 -1847
rect -188 -1849 -186 -1847
rect -180 -1849 -178 -1847
rect -164 -1849 -162 -1847
rect -156 -1849 -154 -1847
rect -146 -1849 -144 -1847
rect -138 -1849 -136 -1847
rect -122 -1849 -120 -1847
rect -114 -1849 -112 -1847
rect -104 -1849 -102 -1847
rect -96 -1849 -94 -1847
rect -80 -1849 -78 -1847
rect -72 -1849 -70 -1847
rect -62 -1849 -60 -1847
rect -54 -1849 -52 -1847
rect -38 -1849 -36 -1847
rect -30 -1849 -28 -1847
rect 144 -1849 146 -1847
rect 154 -1849 156 -1847
rect 170 -1849 172 -1847
rect 178 -1849 180 -1847
rect 194 -1849 196 -1847
rect 202 -1849 204 -1847
rect 212 -1849 214 -1847
rect 220 -1849 222 -1847
rect 236 -1849 238 -1847
rect 244 -1849 246 -1847
rect 254 -1849 256 -1847
rect 262 -1849 264 -1847
rect 278 -1849 280 -1847
rect 286 -1849 288 -1847
rect 296 -1849 298 -1847
rect 304 -1849 306 -1847
rect 320 -1849 322 -1847
rect 328 -1849 330 -1847
rect 500 -1849 502 -1847
rect 510 -1849 512 -1847
rect 526 -1849 528 -1847
rect 534 -1849 536 -1847
rect 550 -1849 552 -1847
rect 558 -1849 560 -1847
rect 568 -1849 570 -1847
rect 576 -1849 578 -1847
rect 592 -1849 594 -1847
rect 600 -1849 602 -1847
rect 610 -1849 612 -1847
rect 618 -1849 620 -1847
rect 634 -1849 636 -1847
rect 642 -1849 644 -1847
rect 652 -1849 654 -1847
rect 660 -1849 662 -1847
rect 676 -1849 678 -1847
rect 684 -1849 686 -1847
rect 858 -1849 860 -1847
rect 868 -1849 870 -1847
rect 884 -1849 886 -1847
rect 892 -1849 894 -1847
rect 908 -1849 910 -1847
rect 916 -1849 918 -1847
rect 926 -1849 928 -1847
rect 934 -1849 936 -1847
rect 950 -1849 952 -1847
rect 958 -1849 960 -1847
rect 968 -1849 970 -1847
rect 976 -1849 978 -1847
rect 992 -1849 994 -1847
rect 1000 -1849 1002 -1847
rect 1010 -1849 1012 -1847
rect 1018 -1849 1020 -1847
rect 1034 -1849 1036 -1847
rect 1042 -1849 1044 -1847
rect 1216 -1849 1218 -1847
rect 1226 -1849 1228 -1847
rect 1242 -1849 1244 -1847
rect 1250 -1849 1252 -1847
rect 1266 -1849 1268 -1847
rect 1274 -1849 1276 -1847
rect 1284 -1849 1286 -1847
rect 1292 -1849 1294 -1847
rect 1308 -1849 1310 -1847
rect 1316 -1849 1318 -1847
rect 1326 -1849 1328 -1847
rect 1334 -1849 1336 -1847
rect 1350 -1849 1352 -1847
rect 1358 -1849 1360 -1847
rect 1368 -1849 1370 -1847
rect 1376 -1849 1378 -1847
rect 1392 -1849 1394 -1847
rect 1400 -1849 1402 -1847
rect -1304 -1874 -1302 -1872
rect -1296 -1874 -1294 -1872
rect -1286 -1874 -1284 -1872
rect -930 -1874 -928 -1872
rect -922 -1874 -920 -1872
rect -912 -1874 -910 -1872
rect -572 -1874 -570 -1872
rect -564 -1874 -562 -1872
rect -554 -1874 -552 -1872
rect -214 -1874 -212 -1872
rect -206 -1874 -204 -1872
rect -196 -1874 -194 -1872
rect 144 -1874 146 -1872
rect 152 -1874 154 -1872
rect 162 -1874 164 -1872
rect 500 -1874 502 -1872
rect 508 -1874 510 -1872
rect 518 -1874 520 -1872
rect 858 -1874 860 -1872
rect 866 -1874 868 -1872
rect 876 -1874 878 -1872
rect 1216 -1874 1218 -1872
rect 1224 -1874 1226 -1872
rect 1234 -1874 1236 -1872
rect -1304 -1950 -1302 -1882
rect -1296 -1906 -1294 -1882
rect -1296 -1950 -1294 -1910
rect -1286 -1950 -1284 -1882
rect -930 -1950 -928 -1882
rect -922 -1906 -920 -1882
rect -922 -1950 -920 -1910
rect -912 -1950 -910 -1882
rect -572 -1950 -570 -1882
rect -564 -1906 -562 -1882
rect -564 -1950 -562 -1910
rect -554 -1950 -552 -1882
rect -214 -1950 -212 -1882
rect -206 -1906 -204 -1882
rect -206 -1950 -204 -1910
rect -196 -1950 -194 -1882
rect 144 -1950 146 -1882
rect 152 -1906 154 -1882
rect 152 -1950 154 -1910
rect 162 -1950 164 -1882
rect 500 -1950 502 -1882
rect 508 -1906 510 -1882
rect 508 -1950 510 -1910
rect 518 -1950 520 -1882
rect 858 -1950 860 -1882
rect 866 -1906 868 -1882
rect 866 -1950 868 -1910
rect 876 -1950 878 -1882
rect 1216 -1950 1218 -1882
rect 1224 -1906 1226 -1882
rect 1224 -1950 1226 -1910
rect 1234 -1950 1236 -1882
rect -1304 -1956 -1302 -1954
rect -1296 -1956 -1294 -1954
rect -1286 -1956 -1284 -1954
rect -930 -1956 -928 -1954
rect -922 -1956 -920 -1954
rect -912 -1956 -910 -1954
rect -572 -1956 -570 -1954
rect -564 -1956 -562 -1954
rect -554 -1956 -552 -1954
rect -214 -1956 -212 -1954
rect -206 -1956 -204 -1954
rect -196 -1956 -194 -1954
rect 144 -1956 146 -1954
rect 152 -1956 154 -1954
rect 162 -1956 164 -1954
rect 500 -1956 502 -1954
rect 508 -1956 510 -1954
rect 518 -1956 520 -1954
rect 858 -1956 860 -1954
rect 866 -1956 868 -1954
rect 876 -1956 878 -1954
rect 1216 -1956 1218 -1954
rect 1224 -1956 1226 -1954
rect 1234 -1956 1236 -1954
rect -1229 -2033 -1227 -2031
rect -1219 -2033 -1217 -2031
rect -1203 -2033 -1201 -2031
rect -1193 -2033 -1191 -2031
rect -1185 -2033 -1183 -2031
rect -1175 -2033 -1173 -2031
rect -1159 -2033 -1157 -2031
rect -1151 -2033 -1149 -2031
rect -1141 -2033 -1139 -2031
rect -930 -2033 -928 -2031
rect -920 -2033 -918 -2031
rect -904 -2033 -902 -2031
rect -894 -2033 -892 -2031
rect -878 -2033 -876 -2031
rect -868 -2033 -866 -2031
rect -860 -2033 -858 -2031
rect -850 -2033 -848 -2031
rect -834 -2033 -832 -2031
rect -826 -2033 -824 -2031
rect -816 -2033 -814 -2031
rect -800 -2033 -798 -2031
rect -790 -2033 -788 -2031
rect -782 -2033 -780 -2031
rect -772 -2033 -770 -2031
rect -756 -2033 -754 -2031
rect -748 -2033 -746 -2031
rect -732 -2033 -730 -2031
rect -716 -2033 -714 -2031
rect -708 -2033 -706 -2031
rect -698 -2033 -696 -2031
rect -572 -2033 -570 -2031
rect -562 -2033 -560 -2031
rect -546 -2033 -544 -2031
rect -536 -2033 -534 -2031
rect -520 -2033 -518 -2031
rect -510 -2033 -508 -2031
rect -502 -2033 -500 -2031
rect -492 -2033 -490 -2031
rect -476 -2033 -474 -2031
rect -468 -2033 -466 -2031
rect -458 -2033 -456 -2031
rect -442 -2033 -440 -2031
rect -432 -2033 -430 -2031
rect -424 -2033 -422 -2031
rect -414 -2033 -412 -2031
rect -398 -2033 -396 -2031
rect -390 -2033 -388 -2031
rect -374 -2033 -372 -2031
rect -358 -2033 -356 -2031
rect -350 -2033 -348 -2031
rect -340 -2033 -338 -2031
rect -214 -2033 -212 -2031
rect -204 -2033 -202 -2031
rect -188 -2033 -186 -2031
rect -178 -2033 -176 -2031
rect -162 -2033 -160 -2031
rect -152 -2033 -150 -2031
rect -144 -2033 -142 -2031
rect -134 -2033 -132 -2031
rect -118 -2033 -116 -2031
rect -110 -2033 -108 -2031
rect -100 -2033 -98 -2031
rect -84 -2033 -82 -2031
rect -74 -2033 -72 -2031
rect -66 -2033 -64 -2031
rect -56 -2033 -54 -2031
rect -40 -2033 -38 -2031
rect -32 -2033 -30 -2031
rect -16 -2033 -14 -2031
rect 0 -2033 2 -2031
rect 8 -2033 10 -2031
rect 18 -2033 20 -2031
rect 144 -2033 146 -2031
rect 154 -2033 156 -2031
rect 170 -2033 172 -2031
rect 180 -2033 182 -2031
rect 196 -2033 198 -2031
rect 206 -2033 208 -2031
rect 214 -2033 216 -2031
rect 224 -2033 226 -2031
rect 240 -2033 242 -2031
rect 248 -2033 250 -2031
rect 258 -2033 260 -2031
rect 274 -2033 276 -2031
rect 284 -2033 286 -2031
rect 292 -2033 294 -2031
rect 302 -2033 304 -2031
rect 318 -2033 320 -2031
rect 326 -2033 328 -2031
rect 342 -2033 344 -2031
rect 358 -2033 360 -2031
rect 366 -2033 368 -2031
rect 376 -2033 378 -2031
rect 500 -2033 502 -2031
rect 510 -2033 512 -2031
rect 526 -2033 528 -2031
rect 536 -2033 538 -2031
rect 552 -2033 554 -2031
rect 562 -2033 564 -2031
rect 570 -2033 572 -2031
rect 580 -2033 582 -2031
rect 596 -2033 598 -2031
rect 604 -2033 606 -2031
rect 614 -2033 616 -2031
rect 630 -2033 632 -2031
rect 640 -2033 642 -2031
rect 648 -2033 650 -2031
rect 658 -2033 660 -2031
rect 674 -2033 676 -2031
rect 682 -2033 684 -2031
rect 698 -2033 700 -2031
rect 714 -2033 716 -2031
rect 722 -2033 724 -2031
rect 732 -2033 734 -2031
rect 858 -2033 860 -2031
rect 868 -2033 870 -2031
rect 884 -2033 886 -2031
rect 894 -2033 896 -2031
rect 910 -2033 912 -2031
rect 920 -2033 922 -2031
rect 928 -2033 930 -2031
rect 938 -2033 940 -2031
rect 954 -2033 956 -2031
rect 962 -2033 964 -2031
rect 972 -2033 974 -2031
rect 988 -2033 990 -2031
rect 998 -2033 1000 -2031
rect 1006 -2033 1008 -2031
rect 1016 -2033 1018 -2031
rect 1032 -2033 1034 -2031
rect 1040 -2033 1042 -2031
rect 1056 -2033 1058 -2031
rect 1072 -2033 1074 -2031
rect 1080 -2033 1082 -2031
rect 1090 -2033 1092 -2031
rect 1216 -2033 1218 -2031
rect 1226 -2033 1228 -2031
rect 1242 -2033 1244 -2031
rect 1252 -2033 1254 -2031
rect 1268 -2033 1270 -2031
rect 1278 -2033 1280 -2031
rect 1286 -2033 1288 -2031
rect 1296 -2033 1298 -2031
rect 1312 -2033 1314 -2031
rect 1320 -2033 1322 -2031
rect 1330 -2033 1332 -2031
rect 1346 -2033 1348 -2031
rect 1356 -2033 1358 -2031
rect 1364 -2033 1366 -2031
rect 1374 -2033 1376 -2031
rect 1390 -2033 1392 -2031
rect 1398 -2033 1400 -2031
rect 1414 -2033 1416 -2031
rect 1430 -2033 1432 -2031
rect 1438 -2033 1440 -2031
rect 1448 -2033 1450 -2031
rect -1229 -2109 -1227 -2041
rect -1219 -2109 -1217 -2041
rect -1203 -2109 -1201 -2041
rect -1193 -2109 -1191 -2041
rect -1185 -2109 -1183 -2041
rect -1175 -2109 -1173 -2041
rect -1159 -2109 -1157 -2041
rect -1151 -2109 -1149 -2041
rect -1141 -2109 -1139 -2041
rect -930 -2109 -928 -2041
rect -920 -2109 -918 -2041
rect -904 -2109 -902 -2041
rect -894 -2109 -892 -2041
rect -878 -2109 -876 -2041
rect -868 -2109 -866 -2041
rect -860 -2109 -858 -2041
rect -850 -2109 -848 -2041
rect -834 -2109 -832 -2041
rect -826 -2109 -824 -2041
rect -816 -2109 -814 -2041
rect -800 -2109 -798 -2041
rect -790 -2109 -788 -2041
rect -782 -2109 -780 -2041
rect -772 -2109 -770 -2041
rect -756 -2109 -754 -2041
rect -748 -2109 -746 -2041
rect -732 -2109 -730 -2041
rect -716 -2109 -714 -2041
rect -708 -2109 -706 -2041
rect -698 -2109 -696 -2041
rect -572 -2109 -570 -2041
rect -562 -2109 -560 -2041
rect -546 -2109 -544 -2041
rect -536 -2109 -534 -2041
rect -520 -2109 -518 -2041
rect -510 -2109 -508 -2041
rect -502 -2109 -500 -2041
rect -492 -2109 -490 -2041
rect -476 -2109 -474 -2041
rect -468 -2109 -466 -2041
rect -458 -2109 -456 -2041
rect -442 -2109 -440 -2041
rect -432 -2109 -430 -2041
rect -424 -2109 -422 -2041
rect -414 -2109 -412 -2041
rect -398 -2109 -396 -2041
rect -390 -2109 -388 -2041
rect -374 -2109 -372 -2041
rect -358 -2109 -356 -2041
rect -350 -2109 -348 -2041
rect -340 -2109 -338 -2041
rect -214 -2109 -212 -2041
rect -204 -2109 -202 -2041
rect -188 -2109 -186 -2041
rect -178 -2109 -176 -2041
rect -162 -2109 -160 -2041
rect -152 -2109 -150 -2041
rect -144 -2109 -142 -2041
rect -134 -2109 -132 -2041
rect -118 -2109 -116 -2041
rect -110 -2109 -108 -2041
rect -100 -2109 -98 -2041
rect -84 -2109 -82 -2041
rect -74 -2109 -72 -2041
rect -66 -2109 -64 -2041
rect -56 -2109 -54 -2041
rect -40 -2109 -38 -2041
rect -32 -2109 -30 -2041
rect -16 -2109 -14 -2041
rect 0 -2109 2 -2041
rect 8 -2109 10 -2041
rect 18 -2109 20 -2041
rect 144 -2109 146 -2041
rect 154 -2109 156 -2041
rect 170 -2109 172 -2041
rect 180 -2109 182 -2041
rect 196 -2109 198 -2041
rect 206 -2109 208 -2041
rect 214 -2109 216 -2041
rect 224 -2109 226 -2041
rect 240 -2109 242 -2041
rect 248 -2109 250 -2041
rect 258 -2109 260 -2041
rect 274 -2109 276 -2041
rect 284 -2109 286 -2041
rect 292 -2109 294 -2041
rect 302 -2109 304 -2041
rect 318 -2109 320 -2041
rect 326 -2109 328 -2041
rect 342 -2109 344 -2041
rect 358 -2109 360 -2041
rect 366 -2109 368 -2041
rect 376 -2109 378 -2041
rect 500 -2109 502 -2041
rect 510 -2109 512 -2041
rect 526 -2109 528 -2041
rect 536 -2109 538 -2041
rect 552 -2109 554 -2041
rect 562 -2109 564 -2041
rect 570 -2109 572 -2041
rect 580 -2109 582 -2041
rect 596 -2109 598 -2041
rect 604 -2109 606 -2041
rect 614 -2109 616 -2041
rect 630 -2109 632 -2041
rect 640 -2109 642 -2041
rect 648 -2109 650 -2041
rect 658 -2109 660 -2041
rect 674 -2109 676 -2041
rect 682 -2109 684 -2041
rect 698 -2109 700 -2041
rect 714 -2109 716 -2041
rect 722 -2109 724 -2041
rect 732 -2109 734 -2041
rect 858 -2109 860 -2041
rect 868 -2109 870 -2041
rect 884 -2109 886 -2041
rect 894 -2109 896 -2041
rect 910 -2109 912 -2041
rect 920 -2109 922 -2041
rect 928 -2109 930 -2041
rect 938 -2109 940 -2041
rect 954 -2109 956 -2041
rect 962 -2109 964 -2041
rect 972 -2109 974 -2041
rect 988 -2109 990 -2041
rect 998 -2109 1000 -2041
rect 1006 -2109 1008 -2041
rect 1016 -2109 1018 -2041
rect 1032 -2109 1034 -2041
rect 1040 -2109 1042 -2041
rect 1056 -2109 1058 -2041
rect 1072 -2109 1074 -2041
rect 1080 -2109 1082 -2041
rect 1090 -2109 1092 -2041
rect 1216 -2109 1218 -2041
rect 1226 -2109 1228 -2041
rect 1242 -2109 1244 -2041
rect 1252 -2109 1254 -2041
rect 1268 -2109 1270 -2041
rect 1278 -2109 1280 -2041
rect 1286 -2109 1288 -2041
rect 1296 -2109 1298 -2041
rect 1312 -2109 1314 -2041
rect 1320 -2109 1322 -2041
rect 1330 -2109 1332 -2041
rect 1346 -2109 1348 -2041
rect 1356 -2109 1358 -2041
rect 1364 -2109 1366 -2041
rect 1374 -2109 1376 -2041
rect 1390 -2109 1392 -2041
rect 1398 -2109 1400 -2041
rect 1414 -2109 1416 -2041
rect 1430 -2109 1432 -2041
rect 1438 -2109 1440 -2041
rect 1448 -2109 1450 -2041
rect -1229 -2115 -1227 -2113
rect -1219 -2115 -1217 -2113
rect -1203 -2115 -1201 -2113
rect -1193 -2115 -1191 -2113
rect -1185 -2115 -1183 -2113
rect -1175 -2115 -1173 -2113
rect -1159 -2115 -1157 -2113
rect -1151 -2115 -1149 -2113
rect -1141 -2115 -1139 -2113
rect -930 -2115 -928 -2113
rect -920 -2115 -918 -2113
rect -904 -2115 -902 -2113
rect -894 -2115 -892 -2113
rect -878 -2115 -876 -2113
rect -868 -2115 -866 -2113
rect -860 -2115 -858 -2113
rect -850 -2115 -848 -2113
rect -834 -2115 -832 -2113
rect -826 -2115 -824 -2113
rect -816 -2115 -814 -2113
rect -800 -2115 -798 -2113
rect -790 -2115 -788 -2113
rect -782 -2115 -780 -2113
rect -772 -2115 -770 -2113
rect -756 -2115 -754 -2113
rect -748 -2115 -746 -2113
rect -732 -2115 -730 -2113
rect -716 -2115 -714 -2113
rect -708 -2115 -706 -2113
rect -698 -2115 -696 -2113
rect -572 -2115 -570 -2113
rect -562 -2115 -560 -2113
rect -546 -2115 -544 -2113
rect -536 -2115 -534 -2113
rect -520 -2115 -518 -2113
rect -510 -2115 -508 -2113
rect -502 -2115 -500 -2113
rect -492 -2115 -490 -2113
rect -476 -2115 -474 -2113
rect -468 -2115 -466 -2113
rect -458 -2115 -456 -2113
rect -442 -2115 -440 -2113
rect -432 -2115 -430 -2113
rect -424 -2115 -422 -2113
rect -414 -2115 -412 -2113
rect -398 -2115 -396 -2113
rect -390 -2115 -388 -2113
rect -374 -2115 -372 -2113
rect -358 -2115 -356 -2113
rect -350 -2115 -348 -2113
rect -340 -2115 -338 -2113
rect -214 -2115 -212 -2113
rect -204 -2115 -202 -2113
rect -188 -2115 -186 -2113
rect -178 -2115 -176 -2113
rect -162 -2115 -160 -2113
rect -152 -2115 -150 -2113
rect -144 -2115 -142 -2113
rect -134 -2115 -132 -2113
rect -118 -2115 -116 -2113
rect -110 -2115 -108 -2113
rect -100 -2115 -98 -2113
rect -84 -2115 -82 -2113
rect -74 -2115 -72 -2113
rect -66 -2115 -64 -2113
rect -56 -2115 -54 -2113
rect -40 -2115 -38 -2113
rect -32 -2115 -30 -2113
rect -16 -2115 -14 -2113
rect 0 -2115 2 -2113
rect 8 -2115 10 -2113
rect 18 -2115 20 -2113
rect 144 -2115 146 -2113
rect 154 -2115 156 -2113
rect 170 -2115 172 -2113
rect 180 -2115 182 -2113
rect 196 -2115 198 -2113
rect 206 -2115 208 -2113
rect 214 -2115 216 -2113
rect 224 -2115 226 -2113
rect 240 -2115 242 -2113
rect 248 -2115 250 -2113
rect 258 -2115 260 -2113
rect 274 -2115 276 -2113
rect 284 -2115 286 -2113
rect 292 -2115 294 -2113
rect 302 -2115 304 -2113
rect 318 -2115 320 -2113
rect 326 -2115 328 -2113
rect 342 -2115 344 -2113
rect 358 -2115 360 -2113
rect 366 -2115 368 -2113
rect 376 -2115 378 -2113
rect 500 -2115 502 -2113
rect 510 -2115 512 -2113
rect 526 -2115 528 -2113
rect 536 -2115 538 -2113
rect 552 -2115 554 -2113
rect 562 -2115 564 -2113
rect 570 -2115 572 -2113
rect 580 -2115 582 -2113
rect 596 -2115 598 -2113
rect 604 -2115 606 -2113
rect 614 -2115 616 -2113
rect 630 -2115 632 -2113
rect 640 -2115 642 -2113
rect 648 -2115 650 -2113
rect 658 -2115 660 -2113
rect 674 -2115 676 -2113
rect 682 -2115 684 -2113
rect 698 -2115 700 -2113
rect 714 -2115 716 -2113
rect 722 -2115 724 -2113
rect 732 -2115 734 -2113
rect 858 -2115 860 -2113
rect 868 -2115 870 -2113
rect 884 -2115 886 -2113
rect 894 -2115 896 -2113
rect 910 -2115 912 -2113
rect 920 -2115 922 -2113
rect 928 -2115 930 -2113
rect 938 -2115 940 -2113
rect 954 -2115 956 -2113
rect 962 -2115 964 -2113
rect 972 -2115 974 -2113
rect 988 -2115 990 -2113
rect 998 -2115 1000 -2113
rect 1006 -2115 1008 -2113
rect 1016 -2115 1018 -2113
rect 1032 -2115 1034 -2113
rect 1040 -2115 1042 -2113
rect 1056 -2115 1058 -2113
rect 1072 -2115 1074 -2113
rect 1080 -2115 1082 -2113
rect 1090 -2115 1092 -2113
rect 1216 -2115 1218 -2113
rect 1226 -2115 1228 -2113
rect 1242 -2115 1244 -2113
rect 1252 -2115 1254 -2113
rect 1268 -2115 1270 -2113
rect 1278 -2115 1280 -2113
rect 1286 -2115 1288 -2113
rect 1296 -2115 1298 -2113
rect 1312 -2115 1314 -2113
rect 1320 -2115 1322 -2113
rect 1330 -2115 1332 -2113
rect 1346 -2115 1348 -2113
rect 1356 -2115 1358 -2113
rect 1364 -2115 1366 -2113
rect 1374 -2115 1376 -2113
rect 1390 -2115 1392 -2113
rect 1398 -2115 1400 -2113
rect 1414 -2115 1416 -2113
rect 1430 -2115 1432 -2113
rect 1438 -2115 1440 -2113
rect 1448 -2115 1450 -2113
rect -1229 -2177 -1227 -2175
rect -1219 -2177 -1217 -2175
rect -1203 -2177 -1201 -2175
rect -1195 -2177 -1193 -2175
rect -1179 -2177 -1177 -2175
rect -1171 -2177 -1169 -2175
rect -1161 -2177 -1159 -2175
rect -1153 -2177 -1151 -2175
rect -1137 -2177 -1135 -2175
rect -1129 -2177 -1127 -2175
rect -1119 -2177 -1117 -2175
rect -1111 -2177 -1109 -2175
rect -1095 -2177 -1093 -2175
rect -1087 -2177 -1085 -2175
rect -1077 -2177 -1075 -2175
rect -1069 -2177 -1067 -2175
rect -1053 -2177 -1051 -2175
rect -1045 -2177 -1043 -2175
rect -930 -2177 -928 -2175
rect -920 -2177 -918 -2175
rect -904 -2177 -902 -2175
rect -896 -2177 -894 -2175
rect -880 -2177 -878 -2175
rect -872 -2177 -870 -2175
rect -862 -2177 -860 -2175
rect -854 -2177 -852 -2175
rect -838 -2177 -836 -2175
rect -830 -2177 -828 -2175
rect -820 -2177 -818 -2175
rect -812 -2177 -810 -2175
rect -796 -2177 -794 -2175
rect -788 -2177 -786 -2175
rect -778 -2177 -776 -2175
rect -770 -2177 -768 -2175
rect -754 -2177 -752 -2175
rect -746 -2177 -744 -2175
rect -572 -2177 -570 -2175
rect -562 -2177 -560 -2175
rect -546 -2177 -544 -2175
rect -538 -2177 -536 -2175
rect -522 -2177 -520 -2175
rect -514 -2177 -512 -2175
rect -504 -2177 -502 -2175
rect -496 -2177 -494 -2175
rect -480 -2177 -478 -2175
rect -472 -2177 -470 -2175
rect -462 -2177 -460 -2175
rect -454 -2177 -452 -2175
rect -438 -2177 -436 -2175
rect -430 -2177 -428 -2175
rect -420 -2177 -418 -2175
rect -412 -2177 -410 -2175
rect -396 -2177 -394 -2175
rect -388 -2177 -386 -2175
rect -214 -2177 -212 -2175
rect -204 -2177 -202 -2175
rect -188 -2177 -186 -2175
rect -180 -2177 -178 -2175
rect -164 -2177 -162 -2175
rect -156 -2177 -154 -2175
rect -146 -2177 -144 -2175
rect -138 -2177 -136 -2175
rect -122 -2177 -120 -2175
rect -114 -2177 -112 -2175
rect -104 -2177 -102 -2175
rect -96 -2177 -94 -2175
rect -80 -2177 -78 -2175
rect -72 -2177 -70 -2175
rect -62 -2177 -60 -2175
rect -54 -2177 -52 -2175
rect -38 -2177 -36 -2175
rect -30 -2177 -28 -2175
rect 144 -2177 146 -2175
rect 154 -2177 156 -2175
rect 170 -2177 172 -2175
rect 178 -2177 180 -2175
rect 194 -2177 196 -2175
rect 202 -2177 204 -2175
rect 212 -2177 214 -2175
rect 220 -2177 222 -2175
rect 236 -2177 238 -2175
rect 244 -2177 246 -2175
rect 254 -2177 256 -2175
rect 262 -2177 264 -2175
rect 278 -2177 280 -2175
rect 286 -2177 288 -2175
rect 296 -2177 298 -2175
rect 304 -2177 306 -2175
rect 320 -2177 322 -2175
rect 328 -2177 330 -2175
rect 500 -2177 502 -2175
rect 510 -2177 512 -2175
rect 526 -2177 528 -2175
rect 534 -2177 536 -2175
rect 550 -2177 552 -2175
rect 558 -2177 560 -2175
rect 568 -2177 570 -2175
rect 576 -2177 578 -2175
rect 592 -2177 594 -2175
rect 600 -2177 602 -2175
rect 610 -2177 612 -2175
rect 618 -2177 620 -2175
rect 634 -2177 636 -2175
rect 642 -2177 644 -2175
rect 652 -2177 654 -2175
rect 660 -2177 662 -2175
rect 676 -2177 678 -2175
rect 684 -2177 686 -2175
rect -1229 -2253 -1227 -2185
rect -1219 -2253 -1217 -2185
rect -1203 -2253 -1201 -2185
rect -1195 -2253 -1193 -2185
rect -1179 -2253 -1177 -2185
rect -1171 -2253 -1169 -2185
rect -1161 -2253 -1159 -2185
rect -1153 -2253 -1151 -2185
rect -1137 -2253 -1135 -2185
rect -1129 -2218 -1127 -2185
rect -1119 -2218 -1117 -2185
rect -1129 -2220 -1117 -2218
rect -1129 -2253 -1127 -2220
rect -1119 -2253 -1117 -2220
rect -1111 -2253 -1109 -2185
rect -1095 -2253 -1093 -2185
rect -1087 -2253 -1085 -2185
rect -1077 -2253 -1075 -2185
rect -1069 -2253 -1067 -2185
rect -1053 -2253 -1051 -2185
rect -1045 -2253 -1043 -2185
rect -930 -2253 -928 -2185
rect -920 -2253 -918 -2185
rect -904 -2253 -902 -2185
rect -896 -2253 -894 -2185
rect -880 -2253 -878 -2185
rect -872 -2253 -870 -2185
rect -862 -2253 -860 -2185
rect -854 -2253 -852 -2185
rect -838 -2253 -836 -2185
rect -830 -2218 -828 -2185
rect -820 -2218 -818 -2185
rect -830 -2220 -818 -2218
rect -830 -2253 -828 -2220
rect -820 -2253 -818 -2220
rect -812 -2253 -810 -2185
rect -796 -2253 -794 -2185
rect -788 -2253 -786 -2185
rect -778 -2253 -776 -2185
rect -770 -2253 -768 -2185
rect -754 -2253 -752 -2185
rect -746 -2253 -744 -2185
rect -572 -2253 -570 -2185
rect -562 -2253 -560 -2185
rect -546 -2253 -544 -2185
rect -538 -2253 -536 -2185
rect -522 -2253 -520 -2185
rect -514 -2253 -512 -2185
rect -504 -2253 -502 -2185
rect -496 -2253 -494 -2185
rect -480 -2253 -478 -2185
rect -472 -2218 -470 -2185
rect -462 -2218 -460 -2185
rect -472 -2220 -460 -2218
rect -472 -2253 -470 -2220
rect -462 -2253 -460 -2220
rect -454 -2253 -452 -2185
rect -438 -2253 -436 -2185
rect -430 -2253 -428 -2185
rect -420 -2253 -418 -2185
rect -412 -2253 -410 -2185
rect -396 -2253 -394 -2185
rect -388 -2253 -386 -2185
rect -214 -2253 -212 -2185
rect -204 -2253 -202 -2185
rect -188 -2253 -186 -2185
rect -180 -2253 -178 -2185
rect -164 -2253 -162 -2185
rect -156 -2253 -154 -2185
rect -146 -2253 -144 -2185
rect -138 -2253 -136 -2185
rect -122 -2253 -120 -2185
rect -114 -2218 -112 -2185
rect -104 -2218 -102 -2185
rect -114 -2220 -102 -2218
rect -114 -2253 -112 -2220
rect -104 -2253 -102 -2220
rect -96 -2253 -94 -2185
rect -80 -2253 -78 -2185
rect -72 -2253 -70 -2185
rect -62 -2253 -60 -2185
rect -54 -2253 -52 -2185
rect -38 -2253 -36 -2185
rect -30 -2253 -28 -2185
rect 144 -2253 146 -2185
rect 154 -2253 156 -2185
rect 170 -2253 172 -2185
rect 178 -2253 180 -2185
rect 194 -2253 196 -2185
rect 202 -2253 204 -2185
rect 212 -2253 214 -2185
rect 220 -2253 222 -2185
rect 236 -2253 238 -2185
rect 244 -2218 246 -2185
rect 254 -2218 256 -2185
rect 244 -2220 256 -2218
rect 244 -2253 246 -2220
rect 254 -2253 256 -2220
rect 262 -2253 264 -2185
rect 278 -2253 280 -2185
rect 286 -2253 288 -2185
rect 296 -2253 298 -2185
rect 304 -2253 306 -2185
rect 320 -2253 322 -2185
rect 328 -2253 330 -2185
rect 500 -2253 502 -2185
rect 510 -2253 512 -2185
rect 526 -2253 528 -2185
rect 534 -2253 536 -2185
rect 550 -2253 552 -2185
rect 558 -2253 560 -2185
rect 568 -2253 570 -2185
rect 576 -2253 578 -2185
rect 592 -2253 594 -2185
rect 600 -2218 602 -2185
rect 610 -2218 612 -2185
rect 600 -2220 612 -2218
rect 600 -2253 602 -2220
rect 610 -2253 612 -2220
rect 618 -2253 620 -2185
rect 634 -2253 636 -2185
rect 642 -2253 644 -2185
rect 652 -2253 654 -2185
rect 660 -2253 662 -2185
rect 676 -2253 678 -2185
rect 684 -2253 686 -2185
rect -1229 -2259 -1227 -2257
rect -1219 -2259 -1217 -2257
rect -1203 -2259 -1201 -2257
rect -1195 -2259 -1193 -2257
rect -1179 -2259 -1177 -2257
rect -1171 -2259 -1169 -2257
rect -1161 -2259 -1159 -2257
rect -1153 -2259 -1151 -2257
rect -1137 -2259 -1135 -2257
rect -1129 -2259 -1127 -2257
rect -1119 -2259 -1117 -2257
rect -1111 -2259 -1109 -2257
rect -1095 -2259 -1093 -2257
rect -1087 -2259 -1085 -2257
rect -1077 -2259 -1075 -2257
rect -1069 -2259 -1067 -2257
rect -1053 -2259 -1051 -2257
rect -1045 -2259 -1043 -2257
rect -930 -2259 -928 -2257
rect -920 -2259 -918 -2257
rect -904 -2259 -902 -2257
rect -896 -2259 -894 -2257
rect -880 -2259 -878 -2257
rect -872 -2259 -870 -2257
rect -862 -2259 -860 -2257
rect -854 -2259 -852 -2257
rect -838 -2259 -836 -2257
rect -830 -2259 -828 -2257
rect -820 -2259 -818 -2257
rect -812 -2259 -810 -2257
rect -796 -2259 -794 -2257
rect -788 -2259 -786 -2257
rect -778 -2259 -776 -2257
rect -770 -2259 -768 -2257
rect -754 -2259 -752 -2257
rect -746 -2259 -744 -2257
rect -572 -2259 -570 -2257
rect -562 -2259 -560 -2257
rect -546 -2259 -544 -2257
rect -538 -2259 -536 -2257
rect -522 -2259 -520 -2257
rect -514 -2259 -512 -2257
rect -504 -2259 -502 -2257
rect -496 -2259 -494 -2257
rect -480 -2259 -478 -2257
rect -472 -2259 -470 -2257
rect -462 -2259 -460 -2257
rect -454 -2259 -452 -2257
rect -438 -2259 -436 -2257
rect -430 -2259 -428 -2257
rect -420 -2259 -418 -2257
rect -412 -2259 -410 -2257
rect -396 -2259 -394 -2257
rect -388 -2259 -386 -2257
rect -214 -2259 -212 -2257
rect -204 -2259 -202 -2257
rect -188 -2259 -186 -2257
rect -180 -2259 -178 -2257
rect -164 -2259 -162 -2257
rect -156 -2259 -154 -2257
rect -146 -2259 -144 -2257
rect -138 -2259 -136 -2257
rect -122 -2259 -120 -2257
rect -114 -2259 -112 -2257
rect -104 -2259 -102 -2257
rect -96 -2259 -94 -2257
rect -80 -2259 -78 -2257
rect -72 -2259 -70 -2257
rect -62 -2259 -60 -2257
rect -54 -2259 -52 -2257
rect -38 -2259 -36 -2257
rect -30 -2259 -28 -2257
rect 144 -2259 146 -2257
rect 154 -2259 156 -2257
rect 170 -2259 172 -2257
rect 178 -2259 180 -2257
rect 194 -2259 196 -2257
rect 202 -2259 204 -2257
rect 212 -2259 214 -2257
rect 220 -2259 222 -2257
rect 236 -2259 238 -2257
rect 244 -2259 246 -2257
rect 254 -2259 256 -2257
rect 262 -2259 264 -2257
rect 278 -2259 280 -2257
rect 286 -2259 288 -2257
rect 296 -2259 298 -2257
rect 304 -2259 306 -2257
rect 320 -2259 322 -2257
rect 328 -2259 330 -2257
rect 500 -2259 502 -2257
rect 510 -2259 512 -2257
rect 526 -2259 528 -2257
rect 534 -2259 536 -2257
rect 550 -2259 552 -2257
rect 558 -2259 560 -2257
rect 568 -2259 570 -2257
rect 576 -2259 578 -2257
rect 592 -2259 594 -2257
rect 600 -2259 602 -2257
rect 610 -2259 612 -2257
rect 618 -2259 620 -2257
rect 634 -2259 636 -2257
rect 642 -2259 644 -2257
rect 652 -2259 654 -2257
rect 660 -2259 662 -2257
rect 676 -2259 678 -2257
rect 684 -2259 686 -2257
rect -1554 -2348 -1552 -2346
rect -1544 -2348 -1542 -2346
rect -1528 -2348 -1526 -2346
rect -1520 -2348 -1518 -2346
rect -1504 -2348 -1502 -2346
rect -1496 -2348 -1494 -2346
rect -1486 -2348 -1484 -2346
rect -1478 -2348 -1476 -2346
rect -1462 -2348 -1460 -2346
rect -1454 -2348 -1452 -2346
rect -1444 -2348 -1442 -2346
rect -1436 -2348 -1434 -2346
rect -1420 -2348 -1418 -2346
rect -1412 -2348 -1410 -2346
rect -1402 -2348 -1400 -2346
rect -1394 -2348 -1392 -2346
rect -1378 -2348 -1376 -2346
rect -1370 -2348 -1368 -2346
rect -1229 -2348 -1227 -2346
rect -1219 -2348 -1217 -2346
rect -1203 -2348 -1201 -2346
rect -1195 -2348 -1193 -2346
rect -1179 -2348 -1177 -2346
rect -1171 -2348 -1169 -2346
rect -1161 -2348 -1159 -2346
rect -1153 -2348 -1151 -2346
rect -1137 -2348 -1135 -2346
rect -1129 -2348 -1127 -2346
rect -1119 -2348 -1117 -2346
rect -1111 -2348 -1109 -2346
rect -1095 -2348 -1093 -2346
rect -1087 -2348 -1085 -2346
rect -1077 -2348 -1075 -2346
rect -1069 -2348 -1067 -2346
rect -1053 -2348 -1051 -2346
rect -1045 -2348 -1043 -2346
rect -930 -2348 -928 -2346
rect -920 -2348 -918 -2346
rect -904 -2348 -902 -2346
rect -896 -2348 -894 -2346
rect -880 -2348 -878 -2346
rect -872 -2348 -870 -2346
rect -862 -2348 -860 -2346
rect -854 -2348 -852 -2346
rect -838 -2348 -836 -2346
rect -830 -2348 -828 -2346
rect -820 -2348 -818 -2346
rect -812 -2348 -810 -2346
rect -796 -2348 -794 -2346
rect -788 -2348 -786 -2346
rect -778 -2348 -776 -2346
rect -770 -2348 -768 -2346
rect -754 -2348 -752 -2346
rect -746 -2348 -744 -2346
rect -572 -2348 -570 -2346
rect -562 -2348 -560 -2346
rect -546 -2348 -544 -2346
rect -538 -2348 -536 -2346
rect -522 -2348 -520 -2346
rect -514 -2348 -512 -2346
rect -504 -2348 -502 -2346
rect -496 -2348 -494 -2346
rect -480 -2348 -478 -2346
rect -472 -2348 -470 -2346
rect -462 -2348 -460 -2346
rect -454 -2348 -452 -2346
rect -438 -2348 -436 -2346
rect -430 -2348 -428 -2346
rect -420 -2348 -418 -2346
rect -412 -2348 -410 -2346
rect -396 -2348 -394 -2346
rect -388 -2348 -386 -2346
rect -214 -2348 -212 -2346
rect -204 -2348 -202 -2346
rect -188 -2348 -186 -2346
rect -180 -2348 -178 -2346
rect -164 -2348 -162 -2346
rect -156 -2348 -154 -2346
rect -146 -2348 -144 -2346
rect -138 -2348 -136 -2346
rect -122 -2348 -120 -2346
rect -114 -2348 -112 -2346
rect -104 -2348 -102 -2346
rect -96 -2348 -94 -2346
rect -80 -2348 -78 -2346
rect -72 -2348 -70 -2346
rect -62 -2348 -60 -2346
rect -54 -2348 -52 -2346
rect -38 -2348 -36 -2346
rect -30 -2348 -28 -2346
rect 144 -2348 146 -2346
rect 154 -2348 156 -2346
rect 170 -2348 172 -2346
rect 178 -2348 180 -2346
rect 194 -2348 196 -2346
rect 202 -2348 204 -2346
rect 212 -2348 214 -2346
rect 220 -2348 222 -2346
rect 236 -2348 238 -2346
rect 244 -2348 246 -2346
rect 254 -2348 256 -2346
rect 262 -2348 264 -2346
rect 278 -2348 280 -2346
rect 286 -2348 288 -2346
rect 296 -2348 298 -2346
rect 304 -2348 306 -2346
rect 320 -2348 322 -2346
rect 328 -2348 330 -2346
rect 500 -2348 502 -2346
rect 510 -2348 512 -2346
rect 526 -2348 528 -2346
rect 534 -2348 536 -2346
rect 550 -2348 552 -2346
rect 558 -2348 560 -2346
rect 568 -2348 570 -2346
rect 576 -2348 578 -2346
rect 592 -2348 594 -2346
rect 600 -2348 602 -2346
rect 610 -2348 612 -2346
rect 618 -2348 620 -2346
rect 634 -2348 636 -2346
rect 642 -2348 644 -2346
rect 652 -2348 654 -2346
rect 660 -2348 662 -2346
rect 676 -2348 678 -2346
rect 684 -2348 686 -2346
rect 858 -2348 860 -2346
rect 868 -2348 870 -2346
rect 884 -2348 886 -2346
rect 892 -2348 894 -2346
rect 908 -2348 910 -2346
rect 916 -2348 918 -2346
rect 926 -2348 928 -2346
rect 934 -2348 936 -2346
rect 950 -2348 952 -2346
rect 958 -2348 960 -2346
rect 968 -2348 970 -2346
rect 976 -2348 978 -2346
rect 992 -2348 994 -2346
rect 1000 -2348 1002 -2346
rect 1010 -2348 1012 -2346
rect 1018 -2348 1020 -2346
rect 1034 -2348 1036 -2346
rect 1042 -2348 1044 -2346
rect 1216 -2348 1218 -2346
rect 1226 -2348 1228 -2346
rect 1242 -2348 1244 -2346
rect 1250 -2348 1252 -2346
rect 1266 -2348 1268 -2346
rect 1274 -2348 1276 -2346
rect 1284 -2348 1286 -2346
rect 1292 -2348 1294 -2346
rect 1308 -2348 1310 -2346
rect 1316 -2348 1318 -2346
rect 1326 -2348 1328 -2346
rect 1334 -2348 1336 -2346
rect 1350 -2348 1352 -2346
rect 1358 -2348 1360 -2346
rect 1368 -2348 1370 -2346
rect 1376 -2348 1378 -2346
rect 1392 -2348 1394 -2346
rect 1400 -2348 1402 -2346
rect -1554 -2424 -1552 -2356
rect -1544 -2424 -1542 -2356
rect -1528 -2424 -1526 -2356
rect -1520 -2424 -1518 -2356
rect -1504 -2424 -1502 -2356
rect -1496 -2424 -1494 -2356
rect -1486 -2424 -1484 -2356
rect -1478 -2424 -1476 -2356
rect -1462 -2424 -1460 -2356
rect -1454 -2389 -1452 -2356
rect -1444 -2389 -1442 -2356
rect -1454 -2391 -1442 -2389
rect -1454 -2424 -1452 -2391
rect -1444 -2424 -1442 -2391
rect -1436 -2424 -1434 -2356
rect -1420 -2424 -1418 -2356
rect -1412 -2424 -1410 -2356
rect -1402 -2424 -1400 -2356
rect -1394 -2424 -1392 -2356
rect -1378 -2424 -1376 -2356
rect -1370 -2424 -1368 -2356
rect -1229 -2424 -1227 -2356
rect -1219 -2424 -1217 -2356
rect -1203 -2424 -1201 -2356
rect -1195 -2424 -1193 -2356
rect -1179 -2424 -1177 -2356
rect -1171 -2424 -1169 -2356
rect -1161 -2424 -1159 -2356
rect -1153 -2424 -1151 -2356
rect -1137 -2424 -1135 -2356
rect -1129 -2389 -1127 -2356
rect -1119 -2389 -1117 -2356
rect -1129 -2391 -1117 -2389
rect -1129 -2424 -1127 -2391
rect -1119 -2424 -1117 -2391
rect -1111 -2424 -1109 -2356
rect -1095 -2424 -1093 -2356
rect -1087 -2424 -1085 -2356
rect -1077 -2424 -1075 -2356
rect -1069 -2424 -1067 -2356
rect -1053 -2424 -1051 -2356
rect -1045 -2424 -1043 -2356
rect -930 -2424 -928 -2356
rect -920 -2424 -918 -2356
rect -904 -2424 -902 -2356
rect -896 -2424 -894 -2356
rect -880 -2424 -878 -2356
rect -872 -2424 -870 -2356
rect -862 -2424 -860 -2356
rect -854 -2424 -852 -2356
rect -838 -2424 -836 -2356
rect -830 -2389 -828 -2356
rect -820 -2389 -818 -2356
rect -830 -2391 -818 -2389
rect -830 -2424 -828 -2391
rect -820 -2424 -818 -2391
rect -812 -2424 -810 -2356
rect -796 -2424 -794 -2356
rect -788 -2424 -786 -2356
rect -778 -2424 -776 -2356
rect -770 -2424 -768 -2356
rect -754 -2424 -752 -2356
rect -746 -2424 -744 -2356
rect -572 -2424 -570 -2356
rect -562 -2424 -560 -2356
rect -546 -2424 -544 -2356
rect -538 -2424 -536 -2356
rect -522 -2424 -520 -2356
rect -514 -2424 -512 -2356
rect -504 -2424 -502 -2356
rect -496 -2424 -494 -2356
rect -480 -2424 -478 -2356
rect -472 -2389 -470 -2356
rect -462 -2389 -460 -2356
rect -472 -2391 -460 -2389
rect -472 -2424 -470 -2391
rect -462 -2424 -460 -2391
rect -454 -2424 -452 -2356
rect -438 -2424 -436 -2356
rect -430 -2424 -428 -2356
rect -420 -2424 -418 -2356
rect -412 -2424 -410 -2356
rect -396 -2424 -394 -2356
rect -388 -2424 -386 -2356
rect -214 -2424 -212 -2356
rect -204 -2424 -202 -2356
rect -188 -2424 -186 -2356
rect -180 -2424 -178 -2356
rect -164 -2424 -162 -2356
rect -156 -2424 -154 -2356
rect -146 -2424 -144 -2356
rect -138 -2424 -136 -2356
rect -122 -2424 -120 -2356
rect -114 -2389 -112 -2356
rect -104 -2389 -102 -2356
rect -114 -2391 -102 -2389
rect -114 -2424 -112 -2391
rect -104 -2424 -102 -2391
rect -96 -2424 -94 -2356
rect -80 -2424 -78 -2356
rect -72 -2424 -70 -2356
rect -62 -2424 -60 -2356
rect -54 -2424 -52 -2356
rect -38 -2424 -36 -2356
rect -30 -2424 -28 -2356
rect 144 -2424 146 -2356
rect 154 -2424 156 -2356
rect 170 -2424 172 -2356
rect 178 -2424 180 -2356
rect 194 -2424 196 -2356
rect 202 -2424 204 -2356
rect 212 -2424 214 -2356
rect 220 -2424 222 -2356
rect 236 -2424 238 -2356
rect 244 -2389 246 -2356
rect 254 -2389 256 -2356
rect 244 -2391 256 -2389
rect 244 -2424 246 -2391
rect 254 -2424 256 -2391
rect 262 -2424 264 -2356
rect 278 -2424 280 -2356
rect 286 -2424 288 -2356
rect 296 -2424 298 -2356
rect 304 -2424 306 -2356
rect 320 -2424 322 -2356
rect 328 -2424 330 -2356
rect 500 -2424 502 -2356
rect 510 -2424 512 -2356
rect 526 -2424 528 -2356
rect 534 -2424 536 -2356
rect 550 -2424 552 -2356
rect 558 -2424 560 -2356
rect 568 -2424 570 -2356
rect 576 -2424 578 -2356
rect 592 -2424 594 -2356
rect 600 -2389 602 -2356
rect 610 -2389 612 -2356
rect 600 -2391 612 -2389
rect 600 -2424 602 -2391
rect 610 -2424 612 -2391
rect 618 -2424 620 -2356
rect 634 -2424 636 -2356
rect 642 -2424 644 -2356
rect 652 -2424 654 -2356
rect 660 -2424 662 -2356
rect 676 -2424 678 -2356
rect 684 -2424 686 -2356
rect 858 -2424 860 -2356
rect 868 -2424 870 -2356
rect 884 -2424 886 -2356
rect 892 -2424 894 -2356
rect 908 -2424 910 -2356
rect 916 -2424 918 -2356
rect 926 -2424 928 -2356
rect 934 -2424 936 -2356
rect 950 -2424 952 -2356
rect 958 -2389 960 -2356
rect 968 -2389 970 -2356
rect 958 -2391 970 -2389
rect 958 -2424 960 -2391
rect 968 -2424 970 -2391
rect 976 -2424 978 -2356
rect 992 -2424 994 -2356
rect 1000 -2424 1002 -2356
rect 1010 -2424 1012 -2356
rect 1018 -2424 1020 -2356
rect 1034 -2424 1036 -2356
rect 1042 -2424 1044 -2356
rect 1216 -2424 1218 -2356
rect 1226 -2424 1228 -2356
rect 1242 -2424 1244 -2356
rect 1250 -2424 1252 -2356
rect 1266 -2424 1268 -2356
rect 1274 -2424 1276 -2356
rect 1284 -2424 1286 -2356
rect 1292 -2424 1294 -2356
rect 1308 -2424 1310 -2356
rect 1316 -2389 1318 -2356
rect 1326 -2389 1328 -2356
rect 1316 -2391 1328 -2389
rect 1316 -2424 1318 -2391
rect 1326 -2424 1328 -2391
rect 1334 -2424 1336 -2356
rect 1350 -2424 1352 -2356
rect 1358 -2424 1360 -2356
rect 1368 -2424 1370 -2356
rect 1376 -2424 1378 -2356
rect 1392 -2424 1394 -2356
rect 1400 -2424 1402 -2356
rect -1554 -2430 -1552 -2428
rect -1544 -2430 -1542 -2428
rect -1528 -2430 -1526 -2428
rect -1520 -2430 -1518 -2428
rect -1504 -2430 -1502 -2428
rect -1496 -2430 -1494 -2428
rect -1486 -2430 -1484 -2428
rect -1478 -2430 -1476 -2428
rect -1462 -2430 -1460 -2428
rect -1454 -2430 -1452 -2428
rect -1444 -2430 -1442 -2428
rect -1436 -2430 -1434 -2428
rect -1420 -2430 -1418 -2428
rect -1412 -2430 -1410 -2428
rect -1402 -2430 -1400 -2428
rect -1394 -2430 -1392 -2428
rect -1378 -2430 -1376 -2428
rect -1370 -2430 -1368 -2428
rect -1229 -2430 -1227 -2428
rect -1219 -2430 -1217 -2428
rect -1203 -2430 -1201 -2428
rect -1195 -2430 -1193 -2428
rect -1179 -2430 -1177 -2428
rect -1171 -2430 -1169 -2428
rect -1161 -2430 -1159 -2428
rect -1153 -2430 -1151 -2428
rect -1137 -2430 -1135 -2428
rect -1129 -2430 -1127 -2428
rect -1119 -2430 -1117 -2428
rect -1111 -2430 -1109 -2428
rect -1095 -2430 -1093 -2428
rect -1087 -2430 -1085 -2428
rect -1077 -2430 -1075 -2428
rect -1069 -2430 -1067 -2428
rect -1053 -2430 -1051 -2428
rect -1045 -2430 -1043 -2428
rect -930 -2430 -928 -2428
rect -920 -2430 -918 -2428
rect -904 -2430 -902 -2428
rect -896 -2430 -894 -2428
rect -880 -2430 -878 -2428
rect -872 -2430 -870 -2428
rect -862 -2430 -860 -2428
rect -854 -2430 -852 -2428
rect -838 -2430 -836 -2428
rect -830 -2430 -828 -2428
rect -820 -2430 -818 -2428
rect -812 -2430 -810 -2428
rect -796 -2430 -794 -2428
rect -788 -2430 -786 -2428
rect -778 -2430 -776 -2428
rect -770 -2430 -768 -2428
rect -754 -2430 -752 -2428
rect -746 -2430 -744 -2428
rect -572 -2430 -570 -2428
rect -562 -2430 -560 -2428
rect -546 -2430 -544 -2428
rect -538 -2430 -536 -2428
rect -522 -2430 -520 -2428
rect -514 -2430 -512 -2428
rect -504 -2430 -502 -2428
rect -496 -2430 -494 -2428
rect -480 -2430 -478 -2428
rect -472 -2430 -470 -2428
rect -462 -2430 -460 -2428
rect -454 -2430 -452 -2428
rect -438 -2430 -436 -2428
rect -430 -2430 -428 -2428
rect -420 -2430 -418 -2428
rect -412 -2430 -410 -2428
rect -396 -2430 -394 -2428
rect -388 -2430 -386 -2428
rect -214 -2430 -212 -2428
rect -204 -2430 -202 -2428
rect -188 -2430 -186 -2428
rect -180 -2430 -178 -2428
rect -164 -2430 -162 -2428
rect -156 -2430 -154 -2428
rect -146 -2430 -144 -2428
rect -138 -2430 -136 -2428
rect -122 -2430 -120 -2428
rect -114 -2430 -112 -2428
rect -104 -2430 -102 -2428
rect -96 -2430 -94 -2428
rect -80 -2430 -78 -2428
rect -72 -2430 -70 -2428
rect -62 -2430 -60 -2428
rect -54 -2430 -52 -2428
rect -38 -2430 -36 -2428
rect -30 -2430 -28 -2428
rect 144 -2430 146 -2428
rect 154 -2430 156 -2428
rect 170 -2430 172 -2428
rect 178 -2430 180 -2428
rect 194 -2430 196 -2428
rect 202 -2430 204 -2428
rect 212 -2430 214 -2428
rect 220 -2430 222 -2428
rect 236 -2430 238 -2428
rect 244 -2430 246 -2428
rect 254 -2430 256 -2428
rect 262 -2430 264 -2428
rect 278 -2430 280 -2428
rect 286 -2430 288 -2428
rect 296 -2430 298 -2428
rect 304 -2430 306 -2428
rect 320 -2430 322 -2428
rect 328 -2430 330 -2428
rect 500 -2430 502 -2428
rect 510 -2430 512 -2428
rect 526 -2430 528 -2428
rect 534 -2430 536 -2428
rect 550 -2430 552 -2428
rect 558 -2430 560 -2428
rect 568 -2430 570 -2428
rect 576 -2430 578 -2428
rect 592 -2430 594 -2428
rect 600 -2430 602 -2428
rect 610 -2430 612 -2428
rect 618 -2430 620 -2428
rect 634 -2430 636 -2428
rect 642 -2430 644 -2428
rect 652 -2430 654 -2428
rect 660 -2430 662 -2428
rect 676 -2430 678 -2428
rect 684 -2430 686 -2428
rect 858 -2430 860 -2428
rect 868 -2430 870 -2428
rect 884 -2430 886 -2428
rect 892 -2430 894 -2428
rect 908 -2430 910 -2428
rect 916 -2430 918 -2428
rect 926 -2430 928 -2428
rect 934 -2430 936 -2428
rect 950 -2430 952 -2428
rect 958 -2430 960 -2428
rect 968 -2430 970 -2428
rect 976 -2430 978 -2428
rect 992 -2430 994 -2428
rect 1000 -2430 1002 -2428
rect 1010 -2430 1012 -2428
rect 1018 -2430 1020 -2428
rect 1034 -2430 1036 -2428
rect 1042 -2430 1044 -2428
rect 1216 -2430 1218 -2428
rect 1226 -2430 1228 -2428
rect 1242 -2430 1244 -2428
rect 1250 -2430 1252 -2428
rect 1266 -2430 1268 -2428
rect 1274 -2430 1276 -2428
rect 1284 -2430 1286 -2428
rect 1292 -2430 1294 -2428
rect 1308 -2430 1310 -2428
rect 1316 -2430 1318 -2428
rect 1326 -2430 1328 -2428
rect 1334 -2430 1336 -2428
rect 1350 -2430 1352 -2428
rect 1358 -2430 1360 -2428
rect 1368 -2430 1370 -2428
rect 1376 -2430 1378 -2428
rect 1392 -2430 1394 -2428
rect 1400 -2430 1402 -2428
rect -1554 -2519 -1552 -2517
rect -1544 -2519 -1542 -2517
rect -1528 -2519 -1526 -2517
rect -1520 -2519 -1518 -2517
rect -1504 -2519 -1502 -2517
rect -1496 -2519 -1494 -2517
rect -1486 -2519 -1484 -2517
rect -1478 -2519 -1476 -2517
rect -1462 -2519 -1460 -2517
rect -1454 -2519 -1452 -2517
rect -1444 -2519 -1442 -2517
rect -1436 -2519 -1434 -2517
rect -1420 -2519 -1418 -2517
rect -1412 -2519 -1410 -2517
rect -1402 -2519 -1400 -2517
rect -1394 -2519 -1392 -2517
rect -1378 -2519 -1376 -2517
rect -1370 -2519 -1368 -2517
rect -1229 -2519 -1227 -2517
rect -1219 -2519 -1217 -2517
rect -1203 -2519 -1201 -2517
rect -1195 -2519 -1193 -2517
rect -1179 -2519 -1177 -2517
rect -1171 -2519 -1169 -2517
rect -1161 -2519 -1159 -2517
rect -1153 -2519 -1151 -2517
rect -1137 -2519 -1135 -2517
rect -1129 -2519 -1127 -2517
rect -1119 -2519 -1117 -2517
rect -1111 -2519 -1109 -2517
rect -1095 -2519 -1093 -2517
rect -1087 -2519 -1085 -2517
rect -1077 -2519 -1075 -2517
rect -1069 -2519 -1067 -2517
rect -1053 -2519 -1051 -2517
rect -1045 -2519 -1043 -2517
rect -930 -2519 -928 -2517
rect -920 -2519 -918 -2517
rect -904 -2519 -902 -2517
rect -896 -2519 -894 -2517
rect -880 -2519 -878 -2517
rect -872 -2519 -870 -2517
rect -862 -2519 -860 -2517
rect -854 -2519 -852 -2517
rect -838 -2519 -836 -2517
rect -830 -2519 -828 -2517
rect -820 -2519 -818 -2517
rect -812 -2519 -810 -2517
rect -796 -2519 -794 -2517
rect -788 -2519 -786 -2517
rect -778 -2519 -776 -2517
rect -770 -2519 -768 -2517
rect -754 -2519 -752 -2517
rect -746 -2519 -744 -2517
rect -572 -2519 -570 -2517
rect -562 -2519 -560 -2517
rect -546 -2519 -544 -2517
rect -538 -2519 -536 -2517
rect -522 -2519 -520 -2517
rect -514 -2519 -512 -2517
rect -504 -2519 -502 -2517
rect -496 -2519 -494 -2517
rect -480 -2519 -478 -2517
rect -472 -2519 -470 -2517
rect -462 -2519 -460 -2517
rect -454 -2519 -452 -2517
rect -438 -2519 -436 -2517
rect -430 -2519 -428 -2517
rect -420 -2519 -418 -2517
rect -412 -2519 -410 -2517
rect -396 -2519 -394 -2517
rect -388 -2519 -386 -2517
rect -215 -2519 -213 -2517
rect -205 -2519 -203 -2517
rect -189 -2519 -187 -2517
rect -181 -2519 -179 -2517
rect -165 -2519 -163 -2517
rect -157 -2519 -155 -2517
rect -147 -2519 -145 -2517
rect -139 -2519 -137 -2517
rect -123 -2519 -121 -2517
rect -115 -2519 -113 -2517
rect -105 -2519 -103 -2517
rect -97 -2519 -95 -2517
rect -81 -2519 -79 -2517
rect -73 -2519 -71 -2517
rect -63 -2519 -61 -2517
rect -55 -2519 -53 -2517
rect -39 -2519 -37 -2517
rect -31 -2519 -29 -2517
rect 144 -2519 146 -2517
rect 154 -2519 156 -2517
rect 170 -2519 172 -2517
rect 178 -2519 180 -2517
rect 194 -2519 196 -2517
rect 202 -2519 204 -2517
rect 212 -2519 214 -2517
rect 220 -2519 222 -2517
rect 236 -2519 238 -2517
rect 244 -2519 246 -2517
rect 254 -2519 256 -2517
rect 262 -2519 264 -2517
rect 278 -2519 280 -2517
rect 286 -2519 288 -2517
rect 296 -2519 298 -2517
rect 304 -2519 306 -2517
rect 320 -2519 322 -2517
rect 328 -2519 330 -2517
rect 500 -2519 502 -2517
rect 510 -2519 512 -2517
rect 526 -2519 528 -2517
rect 534 -2519 536 -2517
rect 550 -2519 552 -2517
rect 558 -2519 560 -2517
rect 568 -2519 570 -2517
rect 576 -2519 578 -2517
rect 592 -2519 594 -2517
rect 600 -2519 602 -2517
rect 610 -2519 612 -2517
rect 618 -2519 620 -2517
rect 634 -2519 636 -2517
rect 642 -2519 644 -2517
rect 652 -2519 654 -2517
rect 660 -2519 662 -2517
rect 676 -2519 678 -2517
rect 684 -2519 686 -2517
rect 858 -2519 860 -2517
rect 868 -2519 870 -2517
rect 884 -2519 886 -2517
rect 892 -2519 894 -2517
rect 908 -2519 910 -2517
rect 916 -2519 918 -2517
rect 926 -2519 928 -2517
rect 934 -2519 936 -2517
rect 950 -2519 952 -2517
rect 958 -2519 960 -2517
rect 968 -2519 970 -2517
rect 976 -2519 978 -2517
rect 992 -2519 994 -2517
rect 1000 -2519 1002 -2517
rect 1010 -2519 1012 -2517
rect 1018 -2519 1020 -2517
rect 1034 -2519 1036 -2517
rect 1042 -2519 1044 -2517
rect 1216 -2519 1218 -2517
rect 1226 -2519 1228 -2517
rect 1242 -2519 1244 -2517
rect 1250 -2519 1252 -2517
rect 1266 -2519 1268 -2517
rect 1274 -2519 1276 -2517
rect 1284 -2519 1286 -2517
rect 1292 -2519 1294 -2517
rect 1308 -2519 1310 -2517
rect 1316 -2519 1318 -2517
rect 1326 -2519 1328 -2517
rect 1334 -2519 1336 -2517
rect 1350 -2519 1352 -2517
rect 1358 -2519 1360 -2517
rect 1368 -2519 1370 -2517
rect 1376 -2519 1378 -2517
rect 1392 -2519 1394 -2517
rect 1400 -2519 1402 -2517
rect -1554 -2595 -1552 -2527
rect -1544 -2595 -1542 -2527
rect -1528 -2595 -1526 -2527
rect -1520 -2595 -1518 -2527
rect -1504 -2595 -1502 -2527
rect -1496 -2595 -1494 -2527
rect -1486 -2595 -1484 -2527
rect -1478 -2595 -1476 -2527
rect -1462 -2595 -1460 -2527
rect -1454 -2560 -1452 -2527
rect -1444 -2560 -1442 -2527
rect -1454 -2562 -1442 -2560
rect -1454 -2595 -1452 -2562
rect -1444 -2595 -1442 -2562
rect -1436 -2595 -1434 -2527
rect -1420 -2595 -1418 -2527
rect -1412 -2595 -1410 -2527
rect -1402 -2595 -1400 -2527
rect -1394 -2595 -1392 -2527
rect -1378 -2595 -1376 -2527
rect -1370 -2595 -1368 -2527
rect -1229 -2595 -1227 -2527
rect -1219 -2595 -1217 -2527
rect -1203 -2595 -1201 -2527
rect -1195 -2595 -1193 -2527
rect -1179 -2595 -1177 -2527
rect -1171 -2595 -1169 -2527
rect -1161 -2595 -1159 -2527
rect -1153 -2595 -1151 -2527
rect -1137 -2595 -1135 -2527
rect -1129 -2560 -1127 -2527
rect -1119 -2560 -1117 -2527
rect -1129 -2562 -1117 -2560
rect -1129 -2595 -1127 -2562
rect -1119 -2595 -1117 -2562
rect -1111 -2595 -1109 -2527
rect -1095 -2595 -1093 -2527
rect -1087 -2595 -1085 -2527
rect -1077 -2595 -1075 -2527
rect -1069 -2595 -1067 -2527
rect -1053 -2595 -1051 -2527
rect -1045 -2595 -1043 -2527
rect -930 -2595 -928 -2527
rect -920 -2595 -918 -2527
rect -904 -2595 -902 -2527
rect -896 -2595 -894 -2527
rect -880 -2595 -878 -2527
rect -872 -2595 -870 -2527
rect -862 -2595 -860 -2527
rect -854 -2595 -852 -2527
rect -838 -2595 -836 -2527
rect -830 -2560 -828 -2527
rect -820 -2560 -818 -2527
rect -830 -2562 -818 -2560
rect -830 -2595 -828 -2562
rect -820 -2595 -818 -2562
rect -812 -2595 -810 -2527
rect -796 -2595 -794 -2527
rect -788 -2595 -786 -2527
rect -778 -2595 -776 -2527
rect -770 -2595 -768 -2527
rect -754 -2595 -752 -2527
rect -746 -2595 -744 -2527
rect -572 -2595 -570 -2527
rect -562 -2595 -560 -2527
rect -546 -2595 -544 -2527
rect -538 -2595 -536 -2527
rect -522 -2595 -520 -2527
rect -514 -2595 -512 -2527
rect -504 -2595 -502 -2527
rect -496 -2595 -494 -2527
rect -480 -2595 -478 -2527
rect -472 -2560 -470 -2527
rect -462 -2560 -460 -2527
rect -472 -2562 -460 -2560
rect -472 -2595 -470 -2562
rect -462 -2595 -460 -2562
rect -454 -2595 -452 -2527
rect -438 -2595 -436 -2527
rect -430 -2595 -428 -2527
rect -420 -2595 -418 -2527
rect -412 -2595 -410 -2527
rect -396 -2595 -394 -2527
rect -388 -2595 -386 -2527
rect -215 -2595 -213 -2527
rect -205 -2595 -203 -2527
rect -189 -2595 -187 -2527
rect -181 -2595 -179 -2527
rect -165 -2595 -163 -2527
rect -157 -2595 -155 -2527
rect -147 -2595 -145 -2527
rect -139 -2595 -137 -2527
rect -123 -2595 -121 -2527
rect -115 -2560 -113 -2527
rect -105 -2560 -103 -2527
rect -115 -2562 -103 -2560
rect -115 -2595 -113 -2562
rect -105 -2595 -103 -2562
rect -97 -2595 -95 -2527
rect -81 -2595 -79 -2527
rect -73 -2595 -71 -2527
rect -63 -2595 -61 -2527
rect -55 -2595 -53 -2527
rect -39 -2595 -37 -2527
rect -31 -2595 -29 -2527
rect 144 -2595 146 -2527
rect 154 -2595 156 -2527
rect 170 -2595 172 -2527
rect 178 -2595 180 -2527
rect 194 -2595 196 -2527
rect 202 -2595 204 -2527
rect 212 -2595 214 -2527
rect 220 -2595 222 -2527
rect 236 -2595 238 -2527
rect 244 -2560 246 -2527
rect 254 -2560 256 -2527
rect 244 -2562 256 -2560
rect 244 -2595 246 -2562
rect 254 -2595 256 -2562
rect 262 -2595 264 -2527
rect 278 -2595 280 -2527
rect 286 -2595 288 -2527
rect 296 -2595 298 -2527
rect 304 -2595 306 -2527
rect 320 -2595 322 -2527
rect 328 -2595 330 -2527
rect 500 -2595 502 -2527
rect 510 -2595 512 -2527
rect 526 -2595 528 -2527
rect 534 -2595 536 -2527
rect 550 -2595 552 -2527
rect 558 -2595 560 -2527
rect 568 -2595 570 -2527
rect 576 -2595 578 -2527
rect 592 -2595 594 -2527
rect 600 -2560 602 -2527
rect 610 -2560 612 -2527
rect 600 -2562 612 -2560
rect 600 -2595 602 -2562
rect 610 -2595 612 -2562
rect 618 -2595 620 -2527
rect 634 -2595 636 -2527
rect 642 -2595 644 -2527
rect 652 -2595 654 -2527
rect 660 -2595 662 -2527
rect 676 -2595 678 -2527
rect 684 -2595 686 -2527
rect 858 -2595 860 -2527
rect 868 -2595 870 -2527
rect 884 -2595 886 -2527
rect 892 -2595 894 -2527
rect 908 -2595 910 -2527
rect 916 -2595 918 -2527
rect 926 -2595 928 -2527
rect 934 -2595 936 -2527
rect 950 -2595 952 -2527
rect 958 -2560 960 -2527
rect 968 -2560 970 -2527
rect 958 -2562 970 -2560
rect 958 -2595 960 -2562
rect 968 -2595 970 -2562
rect 976 -2595 978 -2527
rect 992 -2595 994 -2527
rect 1000 -2595 1002 -2527
rect 1010 -2595 1012 -2527
rect 1018 -2595 1020 -2527
rect 1034 -2595 1036 -2527
rect 1042 -2595 1044 -2527
rect 1216 -2595 1218 -2527
rect 1226 -2595 1228 -2527
rect 1242 -2595 1244 -2527
rect 1250 -2595 1252 -2527
rect 1266 -2595 1268 -2527
rect 1274 -2595 1276 -2527
rect 1284 -2595 1286 -2527
rect 1292 -2595 1294 -2527
rect 1308 -2595 1310 -2527
rect 1316 -2560 1318 -2527
rect 1326 -2560 1328 -2527
rect 1316 -2562 1328 -2560
rect 1316 -2595 1318 -2562
rect 1326 -2595 1328 -2562
rect 1334 -2595 1336 -2527
rect 1350 -2595 1352 -2527
rect 1358 -2595 1360 -2527
rect 1368 -2595 1370 -2527
rect 1376 -2595 1378 -2527
rect 1392 -2595 1394 -2527
rect 1400 -2595 1402 -2527
rect -1554 -2601 -1552 -2599
rect -1544 -2601 -1542 -2599
rect -1528 -2601 -1526 -2599
rect -1520 -2601 -1518 -2599
rect -1504 -2601 -1502 -2599
rect -1496 -2601 -1494 -2599
rect -1486 -2601 -1484 -2599
rect -1478 -2601 -1476 -2599
rect -1462 -2601 -1460 -2599
rect -1454 -2601 -1452 -2599
rect -1444 -2601 -1442 -2599
rect -1436 -2601 -1434 -2599
rect -1420 -2601 -1418 -2599
rect -1412 -2601 -1410 -2599
rect -1402 -2601 -1400 -2599
rect -1394 -2601 -1392 -2599
rect -1378 -2601 -1376 -2599
rect -1370 -2601 -1368 -2599
rect -1229 -2601 -1227 -2599
rect -1219 -2601 -1217 -2599
rect -1203 -2601 -1201 -2599
rect -1195 -2601 -1193 -2599
rect -1179 -2601 -1177 -2599
rect -1171 -2601 -1169 -2599
rect -1161 -2601 -1159 -2599
rect -1153 -2601 -1151 -2599
rect -1137 -2601 -1135 -2599
rect -1129 -2601 -1127 -2599
rect -1119 -2601 -1117 -2599
rect -1111 -2601 -1109 -2599
rect -1095 -2601 -1093 -2599
rect -1087 -2601 -1085 -2599
rect -1077 -2601 -1075 -2599
rect -1069 -2601 -1067 -2599
rect -1053 -2601 -1051 -2599
rect -1045 -2601 -1043 -2599
rect -930 -2601 -928 -2599
rect -920 -2601 -918 -2599
rect -904 -2601 -902 -2599
rect -896 -2601 -894 -2599
rect -880 -2601 -878 -2599
rect -872 -2601 -870 -2599
rect -862 -2601 -860 -2599
rect -854 -2601 -852 -2599
rect -838 -2601 -836 -2599
rect -830 -2601 -828 -2599
rect -820 -2601 -818 -2599
rect -812 -2601 -810 -2599
rect -796 -2601 -794 -2599
rect -788 -2601 -786 -2599
rect -778 -2601 -776 -2599
rect -770 -2601 -768 -2599
rect -754 -2601 -752 -2599
rect -746 -2601 -744 -2599
rect -572 -2601 -570 -2599
rect -562 -2601 -560 -2599
rect -546 -2601 -544 -2599
rect -538 -2601 -536 -2599
rect -522 -2601 -520 -2599
rect -514 -2601 -512 -2599
rect -504 -2601 -502 -2599
rect -496 -2601 -494 -2599
rect -480 -2601 -478 -2599
rect -472 -2601 -470 -2599
rect -462 -2601 -460 -2599
rect -454 -2601 -452 -2599
rect -438 -2601 -436 -2599
rect -430 -2601 -428 -2599
rect -420 -2601 -418 -2599
rect -412 -2601 -410 -2599
rect -396 -2601 -394 -2599
rect -388 -2601 -386 -2599
rect -215 -2601 -213 -2599
rect -205 -2601 -203 -2599
rect -189 -2601 -187 -2599
rect -181 -2601 -179 -2599
rect -165 -2601 -163 -2599
rect -157 -2601 -155 -2599
rect -147 -2601 -145 -2599
rect -139 -2601 -137 -2599
rect -123 -2601 -121 -2599
rect -115 -2601 -113 -2599
rect -105 -2601 -103 -2599
rect -97 -2601 -95 -2599
rect -81 -2601 -79 -2599
rect -73 -2601 -71 -2599
rect -63 -2601 -61 -2599
rect -55 -2601 -53 -2599
rect -39 -2601 -37 -2599
rect -31 -2601 -29 -2599
rect 144 -2601 146 -2599
rect 154 -2601 156 -2599
rect 170 -2601 172 -2599
rect 178 -2601 180 -2599
rect 194 -2601 196 -2599
rect 202 -2601 204 -2599
rect 212 -2601 214 -2599
rect 220 -2601 222 -2599
rect 236 -2601 238 -2599
rect 244 -2601 246 -2599
rect 254 -2601 256 -2599
rect 262 -2601 264 -2599
rect 278 -2601 280 -2599
rect 286 -2601 288 -2599
rect 296 -2601 298 -2599
rect 304 -2601 306 -2599
rect 320 -2601 322 -2599
rect 328 -2601 330 -2599
rect 500 -2601 502 -2599
rect 510 -2601 512 -2599
rect 526 -2601 528 -2599
rect 534 -2601 536 -2599
rect 550 -2601 552 -2599
rect 558 -2601 560 -2599
rect 568 -2601 570 -2599
rect 576 -2601 578 -2599
rect 592 -2601 594 -2599
rect 600 -2601 602 -2599
rect 610 -2601 612 -2599
rect 618 -2601 620 -2599
rect 634 -2601 636 -2599
rect 642 -2601 644 -2599
rect 652 -2601 654 -2599
rect 660 -2601 662 -2599
rect 676 -2601 678 -2599
rect 684 -2601 686 -2599
rect 858 -2601 860 -2599
rect 868 -2601 870 -2599
rect 884 -2601 886 -2599
rect 892 -2601 894 -2599
rect 908 -2601 910 -2599
rect 916 -2601 918 -2599
rect 926 -2601 928 -2599
rect 934 -2601 936 -2599
rect 950 -2601 952 -2599
rect 958 -2601 960 -2599
rect 968 -2601 970 -2599
rect 976 -2601 978 -2599
rect 992 -2601 994 -2599
rect 1000 -2601 1002 -2599
rect 1010 -2601 1012 -2599
rect 1018 -2601 1020 -2599
rect 1034 -2601 1036 -2599
rect 1042 -2601 1044 -2599
rect 1216 -2601 1218 -2599
rect 1226 -2601 1228 -2599
rect 1242 -2601 1244 -2599
rect 1250 -2601 1252 -2599
rect 1266 -2601 1268 -2599
rect 1274 -2601 1276 -2599
rect 1284 -2601 1286 -2599
rect 1292 -2601 1294 -2599
rect 1308 -2601 1310 -2599
rect 1316 -2601 1318 -2599
rect 1326 -2601 1328 -2599
rect 1334 -2601 1336 -2599
rect 1350 -2601 1352 -2599
rect 1358 -2601 1360 -2599
rect 1368 -2601 1370 -2599
rect 1376 -2601 1378 -2599
rect 1392 -2601 1394 -2599
rect 1400 -2601 1402 -2599
rect -1304 -2624 -1302 -2622
rect -1296 -2624 -1294 -2622
rect -1286 -2624 -1284 -2622
rect -930 -2624 -928 -2622
rect -922 -2624 -920 -2622
rect -912 -2624 -910 -2622
rect -572 -2624 -570 -2622
rect -564 -2624 -562 -2622
rect -554 -2624 -552 -2622
rect -214 -2624 -212 -2622
rect -206 -2624 -204 -2622
rect -196 -2624 -194 -2622
rect 144 -2624 146 -2622
rect 152 -2624 154 -2622
rect 162 -2624 164 -2622
rect 500 -2624 502 -2622
rect 508 -2624 510 -2622
rect 518 -2624 520 -2622
rect 858 -2624 860 -2622
rect 866 -2624 868 -2622
rect 876 -2624 878 -2622
rect 1216 -2624 1218 -2622
rect 1224 -2624 1226 -2622
rect 1234 -2624 1236 -2622
rect -1304 -2700 -1302 -2632
rect -1296 -2656 -1294 -2632
rect -1296 -2700 -1294 -2660
rect -1286 -2700 -1284 -2632
rect -930 -2700 -928 -2632
rect -922 -2656 -920 -2632
rect -922 -2700 -920 -2660
rect -912 -2700 -910 -2632
rect -572 -2700 -570 -2632
rect -564 -2656 -562 -2632
rect -564 -2700 -562 -2660
rect -554 -2700 -552 -2632
rect -214 -2700 -212 -2632
rect -206 -2656 -204 -2632
rect -206 -2700 -204 -2660
rect -196 -2700 -194 -2632
rect 144 -2700 146 -2632
rect 152 -2656 154 -2632
rect 152 -2700 154 -2660
rect 162 -2700 164 -2632
rect 500 -2700 502 -2632
rect 508 -2656 510 -2632
rect 508 -2700 510 -2660
rect 518 -2700 520 -2632
rect 858 -2700 860 -2632
rect 866 -2656 868 -2632
rect 866 -2700 868 -2660
rect 876 -2700 878 -2632
rect 1216 -2700 1218 -2632
rect 1224 -2656 1226 -2632
rect 1224 -2700 1226 -2660
rect 1234 -2700 1236 -2632
rect -1304 -2706 -1302 -2704
rect -1296 -2706 -1294 -2704
rect -1286 -2706 -1284 -2704
rect -930 -2706 -928 -2704
rect -922 -2706 -920 -2704
rect -912 -2706 -910 -2704
rect -572 -2706 -570 -2704
rect -564 -2706 -562 -2704
rect -554 -2706 -552 -2704
rect -214 -2706 -212 -2704
rect -206 -2706 -204 -2704
rect -196 -2706 -194 -2704
rect 144 -2706 146 -2704
rect 152 -2706 154 -2704
rect 162 -2706 164 -2704
rect 500 -2706 502 -2704
rect 508 -2706 510 -2704
rect 518 -2706 520 -2704
rect 858 -2706 860 -2704
rect 866 -2706 868 -2704
rect 876 -2706 878 -2704
rect 1216 -2706 1218 -2704
rect 1224 -2706 1226 -2704
rect 1234 -2706 1236 -2704
rect -1229 -2783 -1227 -2781
rect -1219 -2783 -1217 -2781
rect -1203 -2783 -1201 -2781
rect -1193 -2783 -1191 -2781
rect -1185 -2783 -1183 -2781
rect -1175 -2783 -1173 -2781
rect -1159 -2783 -1157 -2781
rect -1151 -2783 -1149 -2781
rect -1141 -2783 -1139 -2781
rect -930 -2783 -928 -2781
rect -920 -2783 -918 -2781
rect -904 -2783 -902 -2781
rect -894 -2783 -892 -2781
rect -878 -2783 -876 -2781
rect -868 -2783 -866 -2781
rect -860 -2783 -858 -2781
rect -850 -2783 -848 -2781
rect -834 -2783 -832 -2781
rect -826 -2783 -824 -2781
rect -816 -2783 -814 -2781
rect -800 -2783 -798 -2781
rect -790 -2783 -788 -2781
rect -782 -2783 -780 -2781
rect -772 -2783 -770 -2781
rect -756 -2783 -754 -2781
rect -748 -2783 -746 -2781
rect -732 -2783 -730 -2781
rect -716 -2783 -714 -2781
rect -708 -2783 -706 -2781
rect -698 -2783 -696 -2781
rect -572 -2783 -570 -2781
rect -562 -2783 -560 -2781
rect -546 -2783 -544 -2781
rect -536 -2783 -534 -2781
rect -520 -2783 -518 -2781
rect -510 -2783 -508 -2781
rect -502 -2783 -500 -2781
rect -492 -2783 -490 -2781
rect -476 -2783 -474 -2781
rect -468 -2783 -466 -2781
rect -458 -2783 -456 -2781
rect -442 -2783 -440 -2781
rect -432 -2783 -430 -2781
rect -424 -2783 -422 -2781
rect -414 -2783 -412 -2781
rect -398 -2783 -396 -2781
rect -390 -2783 -388 -2781
rect -374 -2783 -372 -2781
rect -358 -2783 -356 -2781
rect -350 -2783 -348 -2781
rect -340 -2783 -338 -2781
rect -214 -2783 -212 -2781
rect -204 -2783 -202 -2781
rect -188 -2783 -186 -2781
rect -178 -2783 -176 -2781
rect -162 -2783 -160 -2781
rect -152 -2783 -150 -2781
rect -144 -2783 -142 -2781
rect -134 -2783 -132 -2781
rect -118 -2783 -116 -2781
rect -110 -2783 -108 -2781
rect -100 -2783 -98 -2781
rect -84 -2783 -82 -2781
rect -74 -2783 -72 -2781
rect -66 -2783 -64 -2781
rect -56 -2783 -54 -2781
rect -40 -2783 -38 -2781
rect -32 -2783 -30 -2781
rect -16 -2783 -14 -2781
rect 0 -2783 2 -2781
rect 8 -2783 10 -2781
rect 18 -2783 20 -2781
rect 144 -2783 146 -2781
rect 154 -2783 156 -2781
rect 170 -2783 172 -2781
rect 180 -2783 182 -2781
rect 196 -2783 198 -2781
rect 206 -2783 208 -2781
rect 214 -2783 216 -2781
rect 224 -2783 226 -2781
rect 240 -2783 242 -2781
rect 248 -2783 250 -2781
rect 258 -2783 260 -2781
rect 274 -2783 276 -2781
rect 284 -2783 286 -2781
rect 292 -2783 294 -2781
rect 302 -2783 304 -2781
rect 318 -2783 320 -2781
rect 326 -2783 328 -2781
rect 342 -2783 344 -2781
rect 358 -2783 360 -2781
rect 366 -2783 368 -2781
rect 376 -2783 378 -2781
rect 500 -2783 502 -2781
rect 510 -2783 512 -2781
rect 526 -2783 528 -2781
rect 536 -2783 538 -2781
rect 552 -2783 554 -2781
rect 562 -2783 564 -2781
rect 570 -2783 572 -2781
rect 580 -2783 582 -2781
rect 596 -2783 598 -2781
rect 604 -2783 606 -2781
rect 614 -2783 616 -2781
rect 630 -2783 632 -2781
rect 640 -2783 642 -2781
rect 648 -2783 650 -2781
rect 658 -2783 660 -2781
rect 674 -2783 676 -2781
rect 682 -2783 684 -2781
rect 698 -2783 700 -2781
rect 714 -2783 716 -2781
rect 722 -2783 724 -2781
rect 732 -2783 734 -2781
rect 858 -2783 860 -2781
rect 868 -2783 870 -2781
rect 884 -2783 886 -2781
rect 894 -2783 896 -2781
rect 910 -2783 912 -2781
rect 920 -2783 922 -2781
rect 928 -2783 930 -2781
rect 938 -2783 940 -2781
rect 954 -2783 956 -2781
rect 962 -2783 964 -2781
rect 972 -2783 974 -2781
rect 988 -2783 990 -2781
rect 998 -2783 1000 -2781
rect 1006 -2783 1008 -2781
rect 1016 -2783 1018 -2781
rect 1032 -2783 1034 -2781
rect 1040 -2783 1042 -2781
rect 1056 -2783 1058 -2781
rect 1072 -2783 1074 -2781
rect 1080 -2783 1082 -2781
rect 1090 -2783 1092 -2781
rect 1216 -2783 1218 -2781
rect 1226 -2783 1228 -2781
rect 1242 -2783 1244 -2781
rect 1252 -2783 1254 -2781
rect 1268 -2783 1270 -2781
rect 1278 -2783 1280 -2781
rect 1286 -2783 1288 -2781
rect 1296 -2783 1298 -2781
rect 1312 -2783 1314 -2781
rect 1320 -2783 1322 -2781
rect 1330 -2783 1332 -2781
rect 1346 -2783 1348 -2781
rect 1356 -2783 1358 -2781
rect 1364 -2783 1366 -2781
rect 1374 -2783 1376 -2781
rect 1390 -2783 1392 -2781
rect 1398 -2783 1400 -2781
rect 1414 -2783 1416 -2781
rect 1430 -2783 1432 -2781
rect 1438 -2783 1440 -2781
rect 1448 -2783 1450 -2781
rect -1229 -2859 -1227 -2791
rect -1219 -2859 -1217 -2791
rect -1203 -2859 -1201 -2791
rect -1193 -2859 -1191 -2791
rect -1185 -2859 -1183 -2791
rect -1175 -2859 -1173 -2791
rect -1159 -2859 -1157 -2791
rect -1151 -2859 -1149 -2791
rect -1141 -2859 -1139 -2791
rect -930 -2859 -928 -2791
rect -920 -2859 -918 -2791
rect -904 -2859 -902 -2791
rect -894 -2859 -892 -2791
rect -878 -2859 -876 -2791
rect -868 -2859 -866 -2791
rect -860 -2859 -858 -2791
rect -850 -2859 -848 -2791
rect -834 -2859 -832 -2791
rect -826 -2859 -824 -2791
rect -816 -2859 -814 -2791
rect -800 -2859 -798 -2791
rect -790 -2859 -788 -2791
rect -782 -2859 -780 -2791
rect -772 -2859 -770 -2791
rect -756 -2859 -754 -2791
rect -748 -2859 -746 -2791
rect -732 -2859 -730 -2791
rect -716 -2859 -714 -2791
rect -708 -2859 -706 -2791
rect -698 -2859 -696 -2791
rect -572 -2859 -570 -2791
rect -562 -2859 -560 -2791
rect -546 -2859 -544 -2791
rect -536 -2859 -534 -2791
rect -520 -2859 -518 -2791
rect -510 -2859 -508 -2791
rect -502 -2859 -500 -2791
rect -492 -2859 -490 -2791
rect -476 -2859 -474 -2791
rect -468 -2859 -466 -2791
rect -458 -2859 -456 -2791
rect -442 -2859 -440 -2791
rect -432 -2859 -430 -2791
rect -424 -2859 -422 -2791
rect -414 -2859 -412 -2791
rect -398 -2859 -396 -2791
rect -390 -2859 -388 -2791
rect -374 -2859 -372 -2791
rect -358 -2859 -356 -2791
rect -350 -2859 -348 -2791
rect -340 -2859 -338 -2791
rect -214 -2859 -212 -2791
rect -204 -2859 -202 -2791
rect -188 -2859 -186 -2791
rect -178 -2859 -176 -2791
rect -162 -2859 -160 -2791
rect -152 -2859 -150 -2791
rect -144 -2859 -142 -2791
rect -134 -2859 -132 -2791
rect -118 -2859 -116 -2791
rect -110 -2859 -108 -2791
rect -100 -2859 -98 -2791
rect -84 -2859 -82 -2791
rect -74 -2859 -72 -2791
rect -66 -2859 -64 -2791
rect -56 -2859 -54 -2791
rect -40 -2859 -38 -2791
rect -32 -2859 -30 -2791
rect -16 -2859 -14 -2791
rect 0 -2859 2 -2791
rect 8 -2859 10 -2791
rect 18 -2859 20 -2791
rect 144 -2859 146 -2791
rect 154 -2859 156 -2791
rect 170 -2859 172 -2791
rect 180 -2859 182 -2791
rect 196 -2859 198 -2791
rect 206 -2859 208 -2791
rect 214 -2859 216 -2791
rect 224 -2859 226 -2791
rect 240 -2859 242 -2791
rect 248 -2859 250 -2791
rect 258 -2859 260 -2791
rect 274 -2859 276 -2791
rect 284 -2859 286 -2791
rect 292 -2859 294 -2791
rect 302 -2859 304 -2791
rect 318 -2859 320 -2791
rect 326 -2859 328 -2791
rect 342 -2859 344 -2791
rect 358 -2859 360 -2791
rect 366 -2859 368 -2791
rect 376 -2859 378 -2791
rect 500 -2859 502 -2791
rect 510 -2859 512 -2791
rect 526 -2859 528 -2791
rect 536 -2859 538 -2791
rect 552 -2859 554 -2791
rect 562 -2859 564 -2791
rect 570 -2859 572 -2791
rect 580 -2859 582 -2791
rect 596 -2859 598 -2791
rect 604 -2859 606 -2791
rect 614 -2859 616 -2791
rect 630 -2859 632 -2791
rect 640 -2859 642 -2791
rect 648 -2859 650 -2791
rect 658 -2859 660 -2791
rect 674 -2859 676 -2791
rect 682 -2859 684 -2791
rect 698 -2859 700 -2791
rect 714 -2859 716 -2791
rect 722 -2859 724 -2791
rect 732 -2859 734 -2791
rect 858 -2859 860 -2791
rect 868 -2859 870 -2791
rect 884 -2859 886 -2791
rect 894 -2859 896 -2791
rect 910 -2859 912 -2791
rect 920 -2859 922 -2791
rect 928 -2859 930 -2791
rect 938 -2859 940 -2791
rect 954 -2859 956 -2791
rect 962 -2859 964 -2791
rect 972 -2859 974 -2791
rect 988 -2859 990 -2791
rect 998 -2859 1000 -2791
rect 1006 -2859 1008 -2791
rect 1016 -2859 1018 -2791
rect 1032 -2859 1034 -2791
rect 1040 -2859 1042 -2791
rect 1056 -2859 1058 -2791
rect 1072 -2859 1074 -2791
rect 1080 -2859 1082 -2791
rect 1090 -2859 1092 -2791
rect 1216 -2859 1218 -2791
rect 1226 -2859 1228 -2791
rect 1242 -2859 1244 -2791
rect 1252 -2859 1254 -2791
rect 1268 -2859 1270 -2791
rect 1278 -2859 1280 -2791
rect 1286 -2859 1288 -2791
rect 1296 -2859 1298 -2791
rect 1312 -2859 1314 -2791
rect 1320 -2859 1322 -2791
rect 1330 -2859 1332 -2791
rect 1346 -2859 1348 -2791
rect 1356 -2859 1358 -2791
rect 1364 -2859 1366 -2791
rect 1374 -2859 1376 -2791
rect 1390 -2859 1392 -2791
rect 1398 -2859 1400 -2791
rect 1414 -2859 1416 -2791
rect 1430 -2859 1432 -2791
rect 1438 -2859 1440 -2791
rect 1448 -2859 1450 -2791
rect -1229 -2865 -1227 -2863
rect -1219 -2865 -1217 -2863
rect -1203 -2865 -1201 -2863
rect -1193 -2865 -1191 -2863
rect -1185 -2865 -1183 -2863
rect -1175 -2865 -1173 -2863
rect -1159 -2865 -1157 -2863
rect -1151 -2865 -1149 -2863
rect -1141 -2865 -1139 -2863
rect -930 -2865 -928 -2863
rect -920 -2865 -918 -2863
rect -904 -2865 -902 -2863
rect -894 -2865 -892 -2863
rect -878 -2865 -876 -2863
rect -868 -2865 -866 -2863
rect -860 -2865 -858 -2863
rect -850 -2865 -848 -2863
rect -834 -2865 -832 -2863
rect -826 -2865 -824 -2863
rect -816 -2865 -814 -2863
rect -800 -2865 -798 -2863
rect -790 -2865 -788 -2863
rect -782 -2865 -780 -2863
rect -772 -2865 -770 -2863
rect -756 -2865 -754 -2863
rect -748 -2865 -746 -2863
rect -732 -2865 -730 -2863
rect -716 -2865 -714 -2863
rect -708 -2865 -706 -2863
rect -698 -2865 -696 -2863
rect -572 -2865 -570 -2863
rect -562 -2865 -560 -2863
rect -546 -2865 -544 -2863
rect -536 -2865 -534 -2863
rect -520 -2865 -518 -2863
rect -510 -2865 -508 -2863
rect -502 -2865 -500 -2863
rect -492 -2865 -490 -2863
rect -476 -2865 -474 -2863
rect -468 -2865 -466 -2863
rect -458 -2865 -456 -2863
rect -442 -2865 -440 -2863
rect -432 -2865 -430 -2863
rect -424 -2865 -422 -2863
rect -414 -2865 -412 -2863
rect -398 -2865 -396 -2863
rect -390 -2865 -388 -2863
rect -374 -2865 -372 -2863
rect -358 -2865 -356 -2863
rect -350 -2865 -348 -2863
rect -340 -2865 -338 -2863
rect -214 -2865 -212 -2863
rect -204 -2865 -202 -2863
rect -188 -2865 -186 -2863
rect -178 -2865 -176 -2863
rect -162 -2865 -160 -2863
rect -152 -2865 -150 -2863
rect -144 -2865 -142 -2863
rect -134 -2865 -132 -2863
rect -118 -2865 -116 -2863
rect -110 -2865 -108 -2863
rect -100 -2865 -98 -2863
rect -84 -2865 -82 -2863
rect -74 -2865 -72 -2863
rect -66 -2865 -64 -2863
rect -56 -2865 -54 -2863
rect -40 -2865 -38 -2863
rect -32 -2865 -30 -2863
rect -16 -2865 -14 -2863
rect 0 -2865 2 -2863
rect 8 -2865 10 -2863
rect 18 -2865 20 -2863
rect 144 -2865 146 -2863
rect 154 -2865 156 -2863
rect 170 -2865 172 -2863
rect 180 -2865 182 -2863
rect 196 -2865 198 -2863
rect 206 -2865 208 -2863
rect 214 -2865 216 -2863
rect 224 -2865 226 -2863
rect 240 -2865 242 -2863
rect 248 -2865 250 -2863
rect 258 -2865 260 -2863
rect 274 -2865 276 -2863
rect 284 -2865 286 -2863
rect 292 -2865 294 -2863
rect 302 -2865 304 -2863
rect 318 -2865 320 -2863
rect 326 -2865 328 -2863
rect 342 -2865 344 -2863
rect 358 -2865 360 -2863
rect 366 -2865 368 -2863
rect 376 -2865 378 -2863
rect 500 -2865 502 -2863
rect 510 -2865 512 -2863
rect 526 -2865 528 -2863
rect 536 -2865 538 -2863
rect 552 -2865 554 -2863
rect 562 -2865 564 -2863
rect 570 -2865 572 -2863
rect 580 -2865 582 -2863
rect 596 -2865 598 -2863
rect 604 -2865 606 -2863
rect 614 -2865 616 -2863
rect 630 -2865 632 -2863
rect 640 -2865 642 -2863
rect 648 -2865 650 -2863
rect 658 -2865 660 -2863
rect 674 -2865 676 -2863
rect 682 -2865 684 -2863
rect 698 -2865 700 -2863
rect 714 -2865 716 -2863
rect 722 -2865 724 -2863
rect 732 -2865 734 -2863
rect 858 -2865 860 -2863
rect 868 -2865 870 -2863
rect 884 -2865 886 -2863
rect 894 -2865 896 -2863
rect 910 -2865 912 -2863
rect 920 -2865 922 -2863
rect 928 -2865 930 -2863
rect 938 -2865 940 -2863
rect 954 -2865 956 -2863
rect 962 -2865 964 -2863
rect 972 -2865 974 -2863
rect 988 -2865 990 -2863
rect 998 -2865 1000 -2863
rect 1006 -2865 1008 -2863
rect 1016 -2865 1018 -2863
rect 1032 -2865 1034 -2863
rect 1040 -2865 1042 -2863
rect 1056 -2865 1058 -2863
rect 1072 -2865 1074 -2863
rect 1080 -2865 1082 -2863
rect 1090 -2865 1092 -2863
rect 1216 -2865 1218 -2863
rect 1226 -2865 1228 -2863
rect 1242 -2865 1244 -2863
rect 1252 -2865 1254 -2863
rect 1268 -2865 1270 -2863
rect 1278 -2865 1280 -2863
rect 1286 -2865 1288 -2863
rect 1296 -2865 1298 -2863
rect 1312 -2865 1314 -2863
rect 1320 -2865 1322 -2863
rect 1330 -2865 1332 -2863
rect 1346 -2865 1348 -2863
rect 1356 -2865 1358 -2863
rect 1364 -2865 1366 -2863
rect 1374 -2865 1376 -2863
rect 1390 -2865 1392 -2863
rect 1398 -2865 1400 -2863
rect 1414 -2865 1416 -2863
rect 1430 -2865 1432 -2863
rect 1438 -2865 1440 -2863
rect 1448 -2865 1450 -2863
rect -1554 -2902 -1552 -2900
rect -1544 -2902 -1542 -2900
rect -1528 -2902 -1526 -2900
rect -1520 -2902 -1518 -2900
rect -1504 -2902 -1502 -2900
rect -1496 -2902 -1494 -2900
rect -1486 -2902 -1484 -2900
rect -1478 -2902 -1476 -2900
rect -1462 -2902 -1460 -2900
rect -1454 -2902 -1452 -2900
rect -1444 -2902 -1442 -2900
rect -1436 -2902 -1434 -2900
rect -1420 -2902 -1418 -2900
rect -1412 -2902 -1410 -2900
rect -1402 -2902 -1400 -2900
rect -1394 -2902 -1392 -2900
rect -1378 -2902 -1376 -2900
rect -1370 -2902 -1368 -2900
rect -1229 -2902 -1227 -2900
rect -1219 -2902 -1217 -2900
rect -1203 -2902 -1201 -2900
rect -1195 -2902 -1193 -2900
rect -1179 -2902 -1177 -2900
rect -1171 -2902 -1169 -2900
rect -1161 -2902 -1159 -2900
rect -1153 -2902 -1151 -2900
rect -1137 -2902 -1135 -2900
rect -1129 -2902 -1127 -2900
rect -1119 -2902 -1117 -2900
rect -1111 -2902 -1109 -2900
rect -1095 -2902 -1093 -2900
rect -1087 -2902 -1085 -2900
rect -1077 -2902 -1075 -2900
rect -1069 -2902 -1067 -2900
rect -1053 -2902 -1051 -2900
rect -1045 -2902 -1043 -2900
rect -930 -2902 -928 -2900
rect -920 -2902 -918 -2900
rect -904 -2902 -902 -2900
rect -896 -2902 -894 -2900
rect -880 -2902 -878 -2900
rect -872 -2902 -870 -2900
rect -862 -2902 -860 -2900
rect -854 -2902 -852 -2900
rect -838 -2902 -836 -2900
rect -830 -2902 -828 -2900
rect -820 -2902 -818 -2900
rect -812 -2902 -810 -2900
rect -796 -2902 -794 -2900
rect -788 -2902 -786 -2900
rect -778 -2902 -776 -2900
rect -770 -2902 -768 -2900
rect -754 -2902 -752 -2900
rect -746 -2902 -744 -2900
rect -572 -2902 -570 -2900
rect -562 -2902 -560 -2900
rect -546 -2902 -544 -2900
rect -538 -2902 -536 -2900
rect -522 -2902 -520 -2900
rect -514 -2902 -512 -2900
rect -504 -2902 -502 -2900
rect -496 -2902 -494 -2900
rect -480 -2902 -478 -2900
rect -472 -2902 -470 -2900
rect -462 -2902 -460 -2900
rect -454 -2902 -452 -2900
rect -438 -2902 -436 -2900
rect -430 -2902 -428 -2900
rect -420 -2902 -418 -2900
rect -412 -2902 -410 -2900
rect -396 -2902 -394 -2900
rect -388 -2902 -386 -2900
rect -214 -2902 -212 -2900
rect -204 -2902 -202 -2900
rect -188 -2902 -186 -2900
rect -180 -2902 -178 -2900
rect -164 -2902 -162 -2900
rect -156 -2902 -154 -2900
rect -146 -2902 -144 -2900
rect -138 -2902 -136 -2900
rect -122 -2902 -120 -2900
rect -114 -2902 -112 -2900
rect -104 -2902 -102 -2900
rect -96 -2902 -94 -2900
rect -80 -2902 -78 -2900
rect -72 -2902 -70 -2900
rect -62 -2902 -60 -2900
rect -54 -2902 -52 -2900
rect -38 -2902 -36 -2900
rect -30 -2902 -28 -2900
rect 144 -2902 146 -2900
rect 154 -2902 156 -2900
rect 170 -2902 172 -2900
rect 178 -2902 180 -2900
rect 194 -2902 196 -2900
rect 202 -2902 204 -2900
rect 212 -2902 214 -2900
rect 220 -2902 222 -2900
rect 236 -2902 238 -2900
rect 244 -2902 246 -2900
rect 254 -2902 256 -2900
rect 262 -2902 264 -2900
rect 278 -2902 280 -2900
rect 286 -2902 288 -2900
rect 296 -2902 298 -2900
rect 304 -2902 306 -2900
rect 320 -2902 322 -2900
rect 328 -2902 330 -2900
rect -1554 -2978 -1552 -2910
rect -1544 -2978 -1542 -2910
rect -1528 -2978 -1526 -2910
rect -1520 -2978 -1518 -2910
rect -1504 -2978 -1502 -2910
rect -1496 -2978 -1494 -2910
rect -1486 -2978 -1484 -2910
rect -1478 -2978 -1476 -2910
rect -1462 -2978 -1460 -2910
rect -1454 -2943 -1452 -2910
rect -1444 -2943 -1442 -2910
rect -1454 -2945 -1442 -2943
rect -1454 -2978 -1452 -2945
rect -1444 -2978 -1442 -2945
rect -1436 -2978 -1434 -2910
rect -1420 -2978 -1418 -2910
rect -1412 -2978 -1410 -2910
rect -1402 -2978 -1400 -2910
rect -1394 -2978 -1392 -2910
rect -1378 -2978 -1376 -2910
rect -1370 -2978 -1368 -2910
rect -1229 -2978 -1227 -2910
rect -1219 -2978 -1217 -2910
rect -1203 -2978 -1201 -2910
rect -1195 -2978 -1193 -2910
rect -1179 -2978 -1177 -2910
rect -1171 -2978 -1169 -2910
rect -1161 -2978 -1159 -2910
rect -1153 -2978 -1151 -2910
rect -1137 -2978 -1135 -2910
rect -1129 -2943 -1127 -2910
rect -1119 -2943 -1117 -2910
rect -1129 -2945 -1117 -2943
rect -1129 -2978 -1127 -2945
rect -1119 -2978 -1117 -2945
rect -1111 -2978 -1109 -2910
rect -1095 -2978 -1093 -2910
rect -1087 -2978 -1085 -2910
rect -1077 -2978 -1075 -2910
rect -1069 -2978 -1067 -2910
rect -1053 -2978 -1051 -2910
rect -1045 -2978 -1043 -2910
rect -930 -2978 -928 -2910
rect -920 -2978 -918 -2910
rect -904 -2978 -902 -2910
rect -896 -2978 -894 -2910
rect -880 -2978 -878 -2910
rect -872 -2978 -870 -2910
rect -862 -2978 -860 -2910
rect -854 -2978 -852 -2910
rect -838 -2978 -836 -2910
rect -830 -2943 -828 -2910
rect -820 -2943 -818 -2910
rect -830 -2945 -818 -2943
rect -830 -2978 -828 -2945
rect -820 -2978 -818 -2945
rect -812 -2978 -810 -2910
rect -796 -2978 -794 -2910
rect -788 -2978 -786 -2910
rect -778 -2978 -776 -2910
rect -770 -2978 -768 -2910
rect -754 -2978 -752 -2910
rect -746 -2978 -744 -2910
rect -572 -2978 -570 -2910
rect -562 -2978 -560 -2910
rect -546 -2978 -544 -2910
rect -538 -2978 -536 -2910
rect -522 -2978 -520 -2910
rect -514 -2978 -512 -2910
rect -504 -2978 -502 -2910
rect -496 -2978 -494 -2910
rect -480 -2978 -478 -2910
rect -472 -2943 -470 -2910
rect -462 -2943 -460 -2910
rect -472 -2945 -460 -2943
rect -472 -2978 -470 -2945
rect -462 -2978 -460 -2945
rect -454 -2978 -452 -2910
rect -438 -2978 -436 -2910
rect -430 -2978 -428 -2910
rect -420 -2978 -418 -2910
rect -412 -2978 -410 -2910
rect -396 -2978 -394 -2910
rect -388 -2978 -386 -2910
rect -214 -2978 -212 -2910
rect -204 -2978 -202 -2910
rect -188 -2978 -186 -2910
rect -180 -2978 -178 -2910
rect -164 -2978 -162 -2910
rect -156 -2978 -154 -2910
rect -146 -2978 -144 -2910
rect -138 -2978 -136 -2910
rect -122 -2978 -120 -2910
rect -114 -2943 -112 -2910
rect -104 -2943 -102 -2910
rect -114 -2945 -102 -2943
rect -114 -2978 -112 -2945
rect -104 -2978 -102 -2945
rect -96 -2978 -94 -2910
rect -80 -2978 -78 -2910
rect -72 -2978 -70 -2910
rect -62 -2978 -60 -2910
rect -54 -2978 -52 -2910
rect -38 -2978 -36 -2910
rect -30 -2978 -28 -2910
rect 144 -2978 146 -2910
rect 154 -2978 156 -2910
rect 170 -2978 172 -2910
rect 178 -2978 180 -2910
rect 194 -2978 196 -2910
rect 202 -2978 204 -2910
rect 212 -2978 214 -2910
rect 220 -2978 222 -2910
rect 236 -2978 238 -2910
rect 244 -2943 246 -2910
rect 254 -2943 256 -2910
rect 244 -2945 256 -2943
rect 244 -2978 246 -2945
rect 254 -2978 256 -2945
rect 262 -2978 264 -2910
rect 278 -2978 280 -2910
rect 286 -2978 288 -2910
rect 296 -2978 298 -2910
rect 304 -2978 306 -2910
rect 320 -2978 322 -2910
rect 328 -2978 330 -2910
rect -1554 -2984 -1552 -2982
rect -1544 -2984 -1542 -2982
rect -1528 -2984 -1526 -2982
rect -1520 -2984 -1518 -2982
rect -1504 -2984 -1502 -2982
rect -1496 -2984 -1494 -2982
rect -1486 -2984 -1484 -2982
rect -1478 -2984 -1476 -2982
rect -1462 -2984 -1460 -2982
rect -1454 -2984 -1452 -2982
rect -1444 -2984 -1442 -2982
rect -1436 -2984 -1434 -2982
rect -1420 -2984 -1418 -2982
rect -1412 -2984 -1410 -2982
rect -1402 -2984 -1400 -2982
rect -1394 -2984 -1392 -2982
rect -1378 -2984 -1376 -2982
rect -1370 -2984 -1368 -2982
rect -1229 -2984 -1227 -2982
rect -1219 -2984 -1217 -2982
rect -1203 -2984 -1201 -2982
rect -1195 -2984 -1193 -2982
rect -1179 -2984 -1177 -2982
rect -1171 -2984 -1169 -2982
rect -1161 -2984 -1159 -2982
rect -1153 -2984 -1151 -2982
rect -1137 -2984 -1135 -2982
rect -1129 -2984 -1127 -2982
rect -1119 -2984 -1117 -2982
rect -1111 -2984 -1109 -2982
rect -1095 -2984 -1093 -2982
rect -1087 -2984 -1085 -2982
rect -1077 -2984 -1075 -2982
rect -1069 -2984 -1067 -2982
rect -1053 -2984 -1051 -2982
rect -1045 -2984 -1043 -2982
rect -930 -2984 -928 -2982
rect -920 -2984 -918 -2982
rect -904 -2984 -902 -2982
rect -896 -2984 -894 -2982
rect -880 -2984 -878 -2982
rect -872 -2984 -870 -2982
rect -862 -2984 -860 -2982
rect -854 -2984 -852 -2982
rect -838 -2984 -836 -2982
rect -830 -2984 -828 -2982
rect -820 -2984 -818 -2982
rect -812 -2984 -810 -2982
rect -796 -2984 -794 -2982
rect -788 -2984 -786 -2982
rect -778 -2984 -776 -2982
rect -770 -2984 -768 -2982
rect -754 -2984 -752 -2982
rect -746 -2984 -744 -2982
rect -572 -2984 -570 -2982
rect -562 -2984 -560 -2982
rect -546 -2984 -544 -2982
rect -538 -2984 -536 -2982
rect -522 -2984 -520 -2982
rect -514 -2984 -512 -2982
rect -504 -2984 -502 -2982
rect -496 -2984 -494 -2982
rect -480 -2984 -478 -2982
rect -472 -2984 -470 -2982
rect -462 -2984 -460 -2982
rect -454 -2984 -452 -2982
rect -438 -2984 -436 -2982
rect -430 -2984 -428 -2982
rect -420 -2984 -418 -2982
rect -412 -2984 -410 -2982
rect -396 -2984 -394 -2982
rect -388 -2984 -386 -2982
rect -214 -2984 -212 -2982
rect -204 -2984 -202 -2982
rect -188 -2984 -186 -2982
rect -180 -2984 -178 -2982
rect -164 -2984 -162 -2982
rect -156 -2984 -154 -2982
rect -146 -2984 -144 -2982
rect -138 -2984 -136 -2982
rect -122 -2984 -120 -2982
rect -114 -2984 -112 -2982
rect -104 -2984 -102 -2982
rect -96 -2984 -94 -2982
rect -80 -2984 -78 -2982
rect -72 -2984 -70 -2982
rect -62 -2984 -60 -2982
rect -54 -2984 -52 -2982
rect -38 -2984 -36 -2982
rect -30 -2984 -28 -2982
rect 144 -2984 146 -2982
rect 154 -2984 156 -2982
rect 170 -2984 172 -2982
rect 178 -2984 180 -2982
rect 194 -2984 196 -2982
rect 202 -2984 204 -2982
rect 212 -2984 214 -2982
rect 220 -2984 222 -2982
rect 236 -2984 238 -2982
rect 244 -2984 246 -2982
rect 254 -2984 256 -2982
rect 262 -2984 264 -2982
rect 278 -2984 280 -2982
rect 286 -2984 288 -2982
rect 296 -2984 298 -2982
rect 304 -2984 306 -2982
rect 320 -2984 322 -2982
rect 328 -2984 330 -2982
rect -1554 -3073 -1552 -3071
rect -1544 -3073 -1542 -3071
rect -1528 -3073 -1526 -3071
rect -1520 -3073 -1518 -3071
rect -1504 -3073 -1502 -3071
rect -1496 -3073 -1494 -3071
rect -1486 -3073 -1484 -3071
rect -1478 -3073 -1476 -3071
rect -1462 -3073 -1460 -3071
rect -1454 -3073 -1452 -3071
rect -1444 -3073 -1442 -3071
rect -1436 -3073 -1434 -3071
rect -1420 -3073 -1418 -3071
rect -1412 -3073 -1410 -3071
rect -1402 -3073 -1400 -3071
rect -1394 -3073 -1392 -3071
rect -1378 -3073 -1376 -3071
rect -1370 -3073 -1368 -3071
rect -1229 -3073 -1227 -3071
rect -1219 -3073 -1217 -3071
rect -1203 -3073 -1201 -3071
rect -1195 -3073 -1193 -3071
rect -1179 -3073 -1177 -3071
rect -1171 -3073 -1169 -3071
rect -1161 -3073 -1159 -3071
rect -1153 -3073 -1151 -3071
rect -1137 -3073 -1135 -3071
rect -1129 -3073 -1127 -3071
rect -1119 -3073 -1117 -3071
rect -1111 -3073 -1109 -3071
rect -1095 -3073 -1093 -3071
rect -1087 -3073 -1085 -3071
rect -1077 -3073 -1075 -3071
rect -1069 -3073 -1067 -3071
rect -1053 -3073 -1051 -3071
rect -1045 -3073 -1043 -3071
rect -930 -3073 -928 -3071
rect -920 -3073 -918 -3071
rect -904 -3073 -902 -3071
rect -896 -3073 -894 -3071
rect -880 -3073 -878 -3071
rect -872 -3073 -870 -3071
rect -862 -3073 -860 -3071
rect -854 -3073 -852 -3071
rect -838 -3073 -836 -3071
rect -830 -3073 -828 -3071
rect -820 -3073 -818 -3071
rect -812 -3073 -810 -3071
rect -796 -3073 -794 -3071
rect -788 -3073 -786 -3071
rect -778 -3073 -776 -3071
rect -770 -3073 -768 -3071
rect -754 -3073 -752 -3071
rect -746 -3073 -744 -3071
rect -572 -3073 -570 -3071
rect -562 -3073 -560 -3071
rect -546 -3073 -544 -3071
rect -538 -3073 -536 -3071
rect -522 -3073 -520 -3071
rect -514 -3073 -512 -3071
rect -504 -3073 -502 -3071
rect -496 -3073 -494 -3071
rect -480 -3073 -478 -3071
rect -472 -3073 -470 -3071
rect -462 -3073 -460 -3071
rect -454 -3073 -452 -3071
rect -438 -3073 -436 -3071
rect -430 -3073 -428 -3071
rect -420 -3073 -418 -3071
rect -412 -3073 -410 -3071
rect -396 -3073 -394 -3071
rect -388 -3073 -386 -3071
rect -214 -3073 -212 -3071
rect -204 -3073 -202 -3071
rect -188 -3073 -186 -3071
rect -180 -3073 -178 -3071
rect -164 -3073 -162 -3071
rect -156 -3073 -154 -3071
rect -146 -3073 -144 -3071
rect -138 -3073 -136 -3071
rect -122 -3073 -120 -3071
rect -114 -3073 -112 -3071
rect -104 -3073 -102 -3071
rect -96 -3073 -94 -3071
rect -80 -3073 -78 -3071
rect -72 -3073 -70 -3071
rect -62 -3073 -60 -3071
rect -54 -3073 -52 -3071
rect -38 -3073 -36 -3071
rect -30 -3073 -28 -3071
rect 144 -3073 146 -3071
rect 154 -3073 156 -3071
rect 170 -3073 172 -3071
rect 178 -3073 180 -3071
rect 194 -3073 196 -3071
rect 202 -3073 204 -3071
rect 212 -3073 214 -3071
rect 220 -3073 222 -3071
rect 236 -3073 238 -3071
rect 244 -3073 246 -3071
rect 254 -3073 256 -3071
rect 262 -3073 264 -3071
rect 278 -3073 280 -3071
rect 286 -3073 288 -3071
rect 296 -3073 298 -3071
rect 304 -3073 306 -3071
rect 320 -3073 322 -3071
rect 328 -3073 330 -3071
rect 500 -3073 502 -3071
rect 510 -3073 512 -3071
rect 526 -3073 528 -3071
rect 534 -3073 536 -3071
rect 550 -3073 552 -3071
rect 558 -3073 560 -3071
rect 568 -3073 570 -3071
rect 576 -3073 578 -3071
rect 592 -3073 594 -3071
rect 600 -3073 602 -3071
rect 610 -3073 612 -3071
rect 618 -3073 620 -3071
rect 634 -3073 636 -3071
rect 642 -3073 644 -3071
rect 652 -3073 654 -3071
rect 660 -3073 662 -3071
rect 676 -3073 678 -3071
rect 684 -3073 686 -3071
rect 858 -3073 860 -3071
rect 868 -3073 870 -3071
rect 884 -3073 886 -3071
rect 892 -3073 894 -3071
rect 908 -3073 910 -3071
rect 916 -3073 918 -3071
rect 926 -3073 928 -3071
rect 934 -3073 936 -3071
rect 950 -3073 952 -3071
rect 958 -3073 960 -3071
rect 968 -3073 970 -3071
rect 976 -3073 978 -3071
rect 992 -3073 994 -3071
rect 1000 -3073 1002 -3071
rect 1010 -3073 1012 -3071
rect 1018 -3073 1020 -3071
rect 1034 -3073 1036 -3071
rect 1042 -3073 1044 -3071
rect 1216 -3073 1218 -3071
rect 1226 -3073 1228 -3071
rect 1242 -3073 1244 -3071
rect 1250 -3073 1252 -3071
rect 1266 -3073 1268 -3071
rect 1274 -3073 1276 -3071
rect 1284 -3073 1286 -3071
rect 1292 -3073 1294 -3071
rect 1308 -3073 1310 -3071
rect 1316 -3073 1318 -3071
rect 1326 -3073 1328 -3071
rect 1334 -3073 1336 -3071
rect 1350 -3073 1352 -3071
rect 1358 -3073 1360 -3071
rect 1368 -3073 1370 -3071
rect 1376 -3073 1378 -3071
rect 1392 -3073 1394 -3071
rect 1400 -3073 1402 -3071
rect -1554 -3149 -1552 -3081
rect -1544 -3149 -1542 -3081
rect -1528 -3149 -1526 -3081
rect -1520 -3149 -1518 -3081
rect -1504 -3149 -1502 -3081
rect -1496 -3149 -1494 -3081
rect -1486 -3149 -1484 -3081
rect -1478 -3149 -1476 -3081
rect -1462 -3149 -1460 -3081
rect -1454 -3114 -1452 -3081
rect -1444 -3114 -1442 -3081
rect -1454 -3116 -1442 -3114
rect -1454 -3149 -1452 -3116
rect -1444 -3149 -1442 -3116
rect -1436 -3149 -1434 -3081
rect -1420 -3149 -1418 -3081
rect -1412 -3149 -1410 -3081
rect -1402 -3149 -1400 -3081
rect -1394 -3149 -1392 -3081
rect -1378 -3149 -1376 -3081
rect -1370 -3149 -1368 -3081
rect -1229 -3149 -1227 -3081
rect -1219 -3149 -1217 -3081
rect -1203 -3149 -1201 -3081
rect -1195 -3149 -1193 -3081
rect -1179 -3149 -1177 -3081
rect -1171 -3149 -1169 -3081
rect -1161 -3149 -1159 -3081
rect -1153 -3149 -1151 -3081
rect -1137 -3149 -1135 -3081
rect -1129 -3114 -1127 -3081
rect -1119 -3114 -1117 -3081
rect -1129 -3116 -1117 -3114
rect -1129 -3149 -1127 -3116
rect -1119 -3149 -1117 -3116
rect -1111 -3149 -1109 -3081
rect -1095 -3149 -1093 -3081
rect -1087 -3149 -1085 -3081
rect -1077 -3149 -1075 -3081
rect -1069 -3149 -1067 -3081
rect -1053 -3149 -1051 -3081
rect -1045 -3149 -1043 -3081
rect -930 -3149 -928 -3081
rect -920 -3149 -918 -3081
rect -904 -3149 -902 -3081
rect -896 -3149 -894 -3081
rect -880 -3149 -878 -3081
rect -872 -3149 -870 -3081
rect -862 -3149 -860 -3081
rect -854 -3149 -852 -3081
rect -838 -3149 -836 -3081
rect -830 -3114 -828 -3081
rect -820 -3114 -818 -3081
rect -830 -3116 -818 -3114
rect -830 -3149 -828 -3116
rect -820 -3149 -818 -3116
rect -812 -3149 -810 -3081
rect -796 -3149 -794 -3081
rect -788 -3149 -786 -3081
rect -778 -3149 -776 -3081
rect -770 -3149 -768 -3081
rect -754 -3149 -752 -3081
rect -746 -3149 -744 -3081
rect -572 -3149 -570 -3081
rect -562 -3149 -560 -3081
rect -546 -3149 -544 -3081
rect -538 -3149 -536 -3081
rect -522 -3149 -520 -3081
rect -514 -3149 -512 -3081
rect -504 -3149 -502 -3081
rect -496 -3149 -494 -3081
rect -480 -3149 -478 -3081
rect -472 -3114 -470 -3081
rect -462 -3114 -460 -3081
rect -472 -3116 -460 -3114
rect -472 -3149 -470 -3116
rect -462 -3149 -460 -3116
rect -454 -3149 -452 -3081
rect -438 -3149 -436 -3081
rect -430 -3149 -428 -3081
rect -420 -3149 -418 -3081
rect -412 -3149 -410 -3081
rect -396 -3149 -394 -3081
rect -388 -3149 -386 -3081
rect -214 -3149 -212 -3081
rect -204 -3149 -202 -3081
rect -188 -3149 -186 -3081
rect -180 -3149 -178 -3081
rect -164 -3149 -162 -3081
rect -156 -3149 -154 -3081
rect -146 -3149 -144 -3081
rect -138 -3149 -136 -3081
rect -122 -3149 -120 -3081
rect -114 -3114 -112 -3081
rect -104 -3114 -102 -3081
rect -114 -3116 -102 -3114
rect -114 -3149 -112 -3116
rect -104 -3149 -102 -3116
rect -96 -3149 -94 -3081
rect -80 -3149 -78 -3081
rect -72 -3149 -70 -3081
rect -62 -3149 -60 -3081
rect -54 -3149 -52 -3081
rect -38 -3149 -36 -3081
rect -30 -3149 -28 -3081
rect 144 -3149 146 -3081
rect 154 -3149 156 -3081
rect 170 -3149 172 -3081
rect 178 -3149 180 -3081
rect 194 -3149 196 -3081
rect 202 -3149 204 -3081
rect 212 -3149 214 -3081
rect 220 -3149 222 -3081
rect 236 -3149 238 -3081
rect 244 -3114 246 -3081
rect 254 -3114 256 -3081
rect 244 -3116 256 -3114
rect 244 -3149 246 -3116
rect 254 -3149 256 -3116
rect 262 -3149 264 -3081
rect 278 -3149 280 -3081
rect 286 -3149 288 -3081
rect 296 -3149 298 -3081
rect 304 -3149 306 -3081
rect 320 -3149 322 -3081
rect 328 -3149 330 -3081
rect 500 -3149 502 -3081
rect 510 -3149 512 -3081
rect 526 -3149 528 -3081
rect 534 -3149 536 -3081
rect 550 -3149 552 -3081
rect 558 -3149 560 -3081
rect 568 -3149 570 -3081
rect 576 -3149 578 -3081
rect 592 -3149 594 -3081
rect 600 -3114 602 -3081
rect 610 -3114 612 -3081
rect 600 -3116 612 -3114
rect 600 -3149 602 -3116
rect 610 -3149 612 -3116
rect 618 -3149 620 -3081
rect 634 -3149 636 -3081
rect 642 -3149 644 -3081
rect 652 -3149 654 -3081
rect 660 -3149 662 -3081
rect 676 -3149 678 -3081
rect 684 -3149 686 -3081
rect 858 -3149 860 -3081
rect 868 -3149 870 -3081
rect 884 -3149 886 -3081
rect 892 -3149 894 -3081
rect 908 -3149 910 -3081
rect 916 -3149 918 -3081
rect 926 -3149 928 -3081
rect 934 -3149 936 -3081
rect 950 -3149 952 -3081
rect 958 -3114 960 -3081
rect 968 -3114 970 -3081
rect 958 -3116 970 -3114
rect 958 -3149 960 -3116
rect 968 -3149 970 -3116
rect 976 -3149 978 -3081
rect 992 -3149 994 -3081
rect 1000 -3149 1002 -3081
rect 1010 -3149 1012 -3081
rect 1018 -3149 1020 -3081
rect 1034 -3149 1036 -3081
rect 1042 -3149 1044 -3081
rect 1216 -3149 1218 -3081
rect 1226 -3149 1228 -3081
rect 1242 -3149 1244 -3081
rect 1250 -3149 1252 -3081
rect 1266 -3149 1268 -3081
rect 1274 -3149 1276 -3081
rect 1284 -3149 1286 -3081
rect 1292 -3149 1294 -3081
rect 1308 -3149 1310 -3081
rect 1316 -3114 1318 -3081
rect 1326 -3114 1328 -3081
rect 1316 -3116 1328 -3114
rect 1316 -3149 1318 -3116
rect 1326 -3149 1328 -3116
rect 1334 -3149 1336 -3081
rect 1350 -3149 1352 -3081
rect 1358 -3149 1360 -3081
rect 1368 -3149 1370 -3081
rect 1376 -3149 1378 -3081
rect 1392 -3149 1394 -3081
rect 1400 -3149 1402 -3081
rect -1554 -3155 -1552 -3153
rect -1544 -3155 -1542 -3153
rect -1528 -3155 -1526 -3153
rect -1520 -3155 -1518 -3153
rect -1504 -3155 -1502 -3153
rect -1496 -3155 -1494 -3153
rect -1486 -3155 -1484 -3153
rect -1478 -3155 -1476 -3153
rect -1462 -3155 -1460 -3153
rect -1454 -3155 -1452 -3153
rect -1444 -3155 -1442 -3153
rect -1436 -3155 -1434 -3153
rect -1420 -3155 -1418 -3153
rect -1412 -3155 -1410 -3153
rect -1402 -3155 -1400 -3153
rect -1394 -3155 -1392 -3153
rect -1378 -3155 -1376 -3153
rect -1370 -3155 -1368 -3153
rect -1229 -3155 -1227 -3153
rect -1219 -3155 -1217 -3153
rect -1203 -3155 -1201 -3153
rect -1195 -3155 -1193 -3153
rect -1179 -3155 -1177 -3153
rect -1171 -3155 -1169 -3153
rect -1161 -3155 -1159 -3153
rect -1153 -3155 -1151 -3153
rect -1137 -3155 -1135 -3153
rect -1129 -3155 -1127 -3153
rect -1119 -3155 -1117 -3153
rect -1111 -3155 -1109 -3153
rect -1095 -3155 -1093 -3153
rect -1087 -3155 -1085 -3153
rect -1077 -3155 -1075 -3153
rect -1069 -3155 -1067 -3153
rect -1053 -3155 -1051 -3153
rect -1045 -3155 -1043 -3153
rect -930 -3155 -928 -3153
rect -920 -3155 -918 -3153
rect -904 -3155 -902 -3153
rect -896 -3155 -894 -3153
rect -880 -3155 -878 -3153
rect -872 -3155 -870 -3153
rect -862 -3155 -860 -3153
rect -854 -3155 -852 -3153
rect -838 -3155 -836 -3153
rect -830 -3155 -828 -3153
rect -820 -3155 -818 -3153
rect -812 -3155 -810 -3153
rect -796 -3155 -794 -3153
rect -788 -3155 -786 -3153
rect -778 -3155 -776 -3153
rect -770 -3155 -768 -3153
rect -754 -3155 -752 -3153
rect -746 -3155 -744 -3153
rect -572 -3155 -570 -3153
rect -562 -3155 -560 -3153
rect -546 -3155 -544 -3153
rect -538 -3155 -536 -3153
rect -522 -3155 -520 -3153
rect -514 -3155 -512 -3153
rect -504 -3155 -502 -3153
rect -496 -3155 -494 -3153
rect -480 -3155 -478 -3153
rect -472 -3155 -470 -3153
rect -462 -3155 -460 -3153
rect -454 -3155 -452 -3153
rect -438 -3155 -436 -3153
rect -430 -3155 -428 -3153
rect -420 -3155 -418 -3153
rect -412 -3155 -410 -3153
rect -396 -3155 -394 -3153
rect -388 -3155 -386 -3153
rect -214 -3155 -212 -3153
rect -204 -3155 -202 -3153
rect -188 -3155 -186 -3153
rect -180 -3155 -178 -3153
rect -164 -3155 -162 -3153
rect -156 -3155 -154 -3153
rect -146 -3155 -144 -3153
rect -138 -3155 -136 -3153
rect -122 -3155 -120 -3153
rect -114 -3155 -112 -3153
rect -104 -3155 -102 -3153
rect -96 -3155 -94 -3153
rect -80 -3155 -78 -3153
rect -72 -3155 -70 -3153
rect -62 -3155 -60 -3153
rect -54 -3155 -52 -3153
rect -38 -3155 -36 -3153
rect -30 -3155 -28 -3153
rect 144 -3155 146 -3153
rect 154 -3155 156 -3153
rect 170 -3155 172 -3153
rect 178 -3155 180 -3153
rect 194 -3155 196 -3153
rect 202 -3155 204 -3153
rect 212 -3155 214 -3153
rect 220 -3155 222 -3153
rect 236 -3155 238 -3153
rect 244 -3155 246 -3153
rect 254 -3155 256 -3153
rect 262 -3155 264 -3153
rect 278 -3155 280 -3153
rect 286 -3155 288 -3153
rect 296 -3155 298 -3153
rect 304 -3155 306 -3153
rect 320 -3155 322 -3153
rect 328 -3155 330 -3153
rect 500 -3155 502 -3153
rect 510 -3155 512 -3153
rect 526 -3155 528 -3153
rect 534 -3155 536 -3153
rect 550 -3155 552 -3153
rect 558 -3155 560 -3153
rect 568 -3155 570 -3153
rect 576 -3155 578 -3153
rect 592 -3155 594 -3153
rect 600 -3155 602 -3153
rect 610 -3155 612 -3153
rect 618 -3155 620 -3153
rect 634 -3155 636 -3153
rect 642 -3155 644 -3153
rect 652 -3155 654 -3153
rect 660 -3155 662 -3153
rect 676 -3155 678 -3153
rect 684 -3155 686 -3153
rect 858 -3155 860 -3153
rect 868 -3155 870 -3153
rect 884 -3155 886 -3153
rect 892 -3155 894 -3153
rect 908 -3155 910 -3153
rect 916 -3155 918 -3153
rect 926 -3155 928 -3153
rect 934 -3155 936 -3153
rect 950 -3155 952 -3153
rect 958 -3155 960 -3153
rect 968 -3155 970 -3153
rect 976 -3155 978 -3153
rect 992 -3155 994 -3153
rect 1000 -3155 1002 -3153
rect 1010 -3155 1012 -3153
rect 1018 -3155 1020 -3153
rect 1034 -3155 1036 -3153
rect 1042 -3155 1044 -3153
rect 1216 -3155 1218 -3153
rect 1226 -3155 1228 -3153
rect 1242 -3155 1244 -3153
rect 1250 -3155 1252 -3153
rect 1266 -3155 1268 -3153
rect 1274 -3155 1276 -3153
rect 1284 -3155 1286 -3153
rect 1292 -3155 1294 -3153
rect 1308 -3155 1310 -3153
rect 1316 -3155 1318 -3153
rect 1326 -3155 1328 -3153
rect 1334 -3155 1336 -3153
rect 1350 -3155 1352 -3153
rect 1358 -3155 1360 -3153
rect 1368 -3155 1370 -3153
rect 1376 -3155 1378 -3153
rect 1392 -3155 1394 -3153
rect 1400 -3155 1402 -3153
rect -1554 -3244 -1552 -3242
rect -1544 -3244 -1542 -3242
rect -1528 -3244 -1526 -3242
rect -1520 -3244 -1518 -3242
rect -1504 -3244 -1502 -3242
rect -1496 -3244 -1494 -3242
rect -1486 -3244 -1484 -3242
rect -1478 -3244 -1476 -3242
rect -1462 -3244 -1460 -3242
rect -1454 -3244 -1452 -3242
rect -1444 -3244 -1442 -3242
rect -1436 -3244 -1434 -3242
rect -1420 -3244 -1418 -3242
rect -1412 -3244 -1410 -3242
rect -1402 -3244 -1400 -3242
rect -1394 -3244 -1392 -3242
rect -1378 -3244 -1376 -3242
rect -1370 -3244 -1368 -3242
rect -1229 -3244 -1227 -3242
rect -1219 -3244 -1217 -3242
rect -1203 -3244 -1201 -3242
rect -1195 -3244 -1193 -3242
rect -1179 -3244 -1177 -3242
rect -1171 -3244 -1169 -3242
rect -1161 -3244 -1159 -3242
rect -1153 -3244 -1151 -3242
rect -1137 -3244 -1135 -3242
rect -1129 -3244 -1127 -3242
rect -1119 -3244 -1117 -3242
rect -1111 -3244 -1109 -3242
rect -1095 -3244 -1093 -3242
rect -1087 -3244 -1085 -3242
rect -1077 -3244 -1075 -3242
rect -1069 -3244 -1067 -3242
rect -1053 -3244 -1051 -3242
rect -1045 -3244 -1043 -3242
rect -930 -3244 -928 -3242
rect -920 -3244 -918 -3242
rect -904 -3244 -902 -3242
rect -896 -3244 -894 -3242
rect -880 -3244 -878 -3242
rect -872 -3244 -870 -3242
rect -862 -3244 -860 -3242
rect -854 -3244 -852 -3242
rect -838 -3244 -836 -3242
rect -830 -3244 -828 -3242
rect -820 -3244 -818 -3242
rect -812 -3244 -810 -3242
rect -796 -3244 -794 -3242
rect -788 -3244 -786 -3242
rect -778 -3244 -776 -3242
rect -770 -3244 -768 -3242
rect -754 -3244 -752 -3242
rect -746 -3244 -744 -3242
rect -572 -3244 -570 -3242
rect -562 -3244 -560 -3242
rect -546 -3244 -544 -3242
rect -538 -3244 -536 -3242
rect -522 -3244 -520 -3242
rect -514 -3244 -512 -3242
rect -504 -3244 -502 -3242
rect -496 -3244 -494 -3242
rect -480 -3244 -478 -3242
rect -472 -3244 -470 -3242
rect -462 -3244 -460 -3242
rect -454 -3244 -452 -3242
rect -438 -3244 -436 -3242
rect -430 -3244 -428 -3242
rect -420 -3244 -418 -3242
rect -412 -3244 -410 -3242
rect -396 -3244 -394 -3242
rect -388 -3244 -386 -3242
rect -214 -3244 -212 -3242
rect -204 -3244 -202 -3242
rect -188 -3244 -186 -3242
rect -180 -3244 -178 -3242
rect -164 -3244 -162 -3242
rect -156 -3244 -154 -3242
rect -146 -3244 -144 -3242
rect -138 -3244 -136 -3242
rect -122 -3244 -120 -3242
rect -114 -3244 -112 -3242
rect -104 -3244 -102 -3242
rect -96 -3244 -94 -3242
rect -80 -3244 -78 -3242
rect -72 -3244 -70 -3242
rect -62 -3244 -60 -3242
rect -54 -3244 -52 -3242
rect -38 -3244 -36 -3242
rect -30 -3244 -28 -3242
rect 144 -3244 146 -3242
rect 154 -3244 156 -3242
rect 170 -3244 172 -3242
rect 178 -3244 180 -3242
rect 194 -3244 196 -3242
rect 202 -3244 204 -3242
rect 212 -3244 214 -3242
rect 220 -3244 222 -3242
rect 236 -3244 238 -3242
rect 244 -3244 246 -3242
rect 254 -3244 256 -3242
rect 262 -3244 264 -3242
rect 278 -3244 280 -3242
rect 286 -3244 288 -3242
rect 296 -3244 298 -3242
rect 304 -3244 306 -3242
rect 320 -3244 322 -3242
rect 328 -3244 330 -3242
rect 500 -3244 502 -3242
rect 510 -3244 512 -3242
rect 526 -3244 528 -3242
rect 534 -3244 536 -3242
rect 550 -3244 552 -3242
rect 558 -3244 560 -3242
rect 568 -3244 570 -3242
rect 576 -3244 578 -3242
rect 592 -3244 594 -3242
rect 600 -3244 602 -3242
rect 610 -3244 612 -3242
rect 618 -3244 620 -3242
rect 634 -3244 636 -3242
rect 642 -3244 644 -3242
rect 652 -3244 654 -3242
rect 660 -3244 662 -3242
rect 676 -3244 678 -3242
rect 684 -3244 686 -3242
rect 858 -3244 860 -3242
rect 868 -3244 870 -3242
rect 884 -3244 886 -3242
rect 892 -3244 894 -3242
rect 908 -3244 910 -3242
rect 916 -3244 918 -3242
rect 926 -3244 928 -3242
rect 934 -3244 936 -3242
rect 950 -3244 952 -3242
rect 958 -3244 960 -3242
rect 968 -3244 970 -3242
rect 976 -3244 978 -3242
rect 992 -3244 994 -3242
rect 1000 -3244 1002 -3242
rect 1010 -3244 1012 -3242
rect 1018 -3244 1020 -3242
rect 1034 -3244 1036 -3242
rect 1042 -3244 1044 -3242
rect 1216 -3244 1218 -3242
rect 1226 -3244 1228 -3242
rect 1242 -3244 1244 -3242
rect 1250 -3244 1252 -3242
rect 1266 -3244 1268 -3242
rect 1274 -3244 1276 -3242
rect 1284 -3244 1286 -3242
rect 1292 -3244 1294 -3242
rect 1308 -3244 1310 -3242
rect 1316 -3244 1318 -3242
rect 1326 -3244 1328 -3242
rect 1334 -3244 1336 -3242
rect 1350 -3244 1352 -3242
rect 1358 -3244 1360 -3242
rect 1368 -3244 1370 -3242
rect 1376 -3244 1378 -3242
rect 1392 -3244 1394 -3242
rect 1400 -3244 1402 -3242
rect -1554 -3320 -1552 -3252
rect -1544 -3320 -1542 -3252
rect -1528 -3320 -1526 -3252
rect -1520 -3320 -1518 -3252
rect -1504 -3320 -1502 -3252
rect -1496 -3320 -1494 -3252
rect -1486 -3320 -1484 -3252
rect -1478 -3320 -1476 -3252
rect -1462 -3320 -1460 -3252
rect -1454 -3285 -1452 -3252
rect -1444 -3285 -1442 -3252
rect -1454 -3287 -1442 -3285
rect -1454 -3320 -1452 -3287
rect -1444 -3320 -1442 -3287
rect -1436 -3320 -1434 -3252
rect -1420 -3320 -1418 -3252
rect -1412 -3320 -1410 -3252
rect -1402 -3320 -1400 -3252
rect -1394 -3320 -1392 -3252
rect -1378 -3320 -1376 -3252
rect -1370 -3320 -1368 -3252
rect -1229 -3320 -1227 -3252
rect -1219 -3320 -1217 -3252
rect -1203 -3320 -1201 -3252
rect -1195 -3320 -1193 -3252
rect -1179 -3320 -1177 -3252
rect -1171 -3320 -1169 -3252
rect -1161 -3320 -1159 -3252
rect -1153 -3320 -1151 -3252
rect -1137 -3320 -1135 -3252
rect -1129 -3285 -1127 -3252
rect -1119 -3285 -1117 -3252
rect -1129 -3287 -1117 -3285
rect -1129 -3320 -1127 -3287
rect -1119 -3320 -1117 -3287
rect -1111 -3320 -1109 -3252
rect -1095 -3320 -1093 -3252
rect -1087 -3320 -1085 -3252
rect -1077 -3320 -1075 -3252
rect -1069 -3320 -1067 -3252
rect -1053 -3320 -1051 -3252
rect -1045 -3320 -1043 -3252
rect -930 -3320 -928 -3252
rect -920 -3320 -918 -3252
rect -904 -3320 -902 -3252
rect -896 -3320 -894 -3252
rect -880 -3320 -878 -3252
rect -872 -3320 -870 -3252
rect -862 -3320 -860 -3252
rect -854 -3320 -852 -3252
rect -838 -3320 -836 -3252
rect -830 -3285 -828 -3252
rect -820 -3285 -818 -3252
rect -830 -3287 -818 -3285
rect -830 -3320 -828 -3287
rect -820 -3320 -818 -3287
rect -812 -3320 -810 -3252
rect -796 -3320 -794 -3252
rect -788 -3320 -786 -3252
rect -778 -3320 -776 -3252
rect -770 -3320 -768 -3252
rect -754 -3320 -752 -3252
rect -746 -3320 -744 -3252
rect -572 -3320 -570 -3252
rect -562 -3320 -560 -3252
rect -546 -3320 -544 -3252
rect -538 -3320 -536 -3252
rect -522 -3320 -520 -3252
rect -514 -3320 -512 -3252
rect -504 -3320 -502 -3252
rect -496 -3320 -494 -3252
rect -480 -3320 -478 -3252
rect -472 -3285 -470 -3252
rect -462 -3285 -460 -3252
rect -472 -3287 -460 -3285
rect -472 -3320 -470 -3287
rect -462 -3320 -460 -3287
rect -454 -3320 -452 -3252
rect -438 -3320 -436 -3252
rect -430 -3320 -428 -3252
rect -420 -3320 -418 -3252
rect -412 -3320 -410 -3252
rect -396 -3320 -394 -3252
rect -388 -3320 -386 -3252
rect -214 -3320 -212 -3252
rect -204 -3320 -202 -3252
rect -188 -3320 -186 -3252
rect -180 -3320 -178 -3252
rect -164 -3320 -162 -3252
rect -156 -3320 -154 -3252
rect -146 -3320 -144 -3252
rect -138 -3320 -136 -3252
rect -122 -3320 -120 -3252
rect -114 -3285 -112 -3252
rect -104 -3285 -102 -3252
rect -114 -3287 -102 -3285
rect -114 -3320 -112 -3287
rect -104 -3320 -102 -3287
rect -96 -3320 -94 -3252
rect -80 -3320 -78 -3252
rect -72 -3320 -70 -3252
rect -62 -3320 -60 -3252
rect -54 -3320 -52 -3252
rect -38 -3320 -36 -3252
rect -30 -3320 -28 -3252
rect 144 -3320 146 -3252
rect 154 -3320 156 -3252
rect 170 -3320 172 -3252
rect 178 -3320 180 -3252
rect 194 -3320 196 -3252
rect 202 -3320 204 -3252
rect 212 -3320 214 -3252
rect 220 -3320 222 -3252
rect 236 -3320 238 -3252
rect 244 -3285 246 -3252
rect 254 -3285 256 -3252
rect 244 -3287 256 -3285
rect 244 -3320 246 -3287
rect 254 -3320 256 -3287
rect 262 -3320 264 -3252
rect 278 -3320 280 -3252
rect 286 -3320 288 -3252
rect 296 -3320 298 -3252
rect 304 -3320 306 -3252
rect 320 -3320 322 -3252
rect 328 -3320 330 -3252
rect 500 -3320 502 -3252
rect 510 -3320 512 -3252
rect 526 -3320 528 -3252
rect 534 -3320 536 -3252
rect 550 -3320 552 -3252
rect 558 -3320 560 -3252
rect 568 -3320 570 -3252
rect 576 -3320 578 -3252
rect 592 -3320 594 -3252
rect 600 -3285 602 -3252
rect 610 -3285 612 -3252
rect 600 -3287 612 -3285
rect 600 -3320 602 -3287
rect 610 -3320 612 -3287
rect 618 -3320 620 -3252
rect 634 -3320 636 -3252
rect 642 -3320 644 -3252
rect 652 -3320 654 -3252
rect 660 -3320 662 -3252
rect 676 -3320 678 -3252
rect 684 -3320 686 -3252
rect 858 -3320 860 -3252
rect 868 -3320 870 -3252
rect 884 -3320 886 -3252
rect 892 -3320 894 -3252
rect 908 -3320 910 -3252
rect 916 -3320 918 -3252
rect 926 -3320 928 -3252
rect 934 -3320 936 -3252
rect 950 -3320 952 -3252
rect 958 -3285 960 -3252
rect 968 -3285 970 -3252
rect 958 -3287 970 -3285
rect 958 -3320 960 -3287
rect 968 -3320 970 -3287
rect 976 -3320 978 -3252
rect 992 -3320 994 -3252
rect 1000 -3320 1002 -3252
rect 1010 -3320 1012 -3252
rect 1018 -3320 1020 -3252
rect 1034 -3320 1036 -3252
rect 1042 -3320 1044 -3252
rect 1216 -3320 1218 -3252
rect 1226 -3320 1228 -3252
rect 1242 -3320 1244 -3252
rect 1250 -3320 1252 -3252
rect 1266 -3320 1268 -3252
rect 1274 -3320 1276 -3252
rect 1284 -3320 1286 -3252
rect 1292 -3320 1294 -3252
rect 1308 -3320 1310 -3252
rect 1316 -3285 1318 -3252
rect 1326 -3285 1328 -3252
rect 1316 -3287 1328 -3285
rect 1316 -3320 1318 -3287
rect 1326 -3320 1328 -3287
rect 1334 -3320 1336 -3252
rect 1350 -3320 1352 -3252
rect 1358 -3320 1360 -3252
rect 1368 -3320 1370 -3252
rect 1376 -3320 1378 -3252
rect 1392 -3320 1394 -3252
rect 1400 -3320 1402 -3252
rect -1554 -3326 -1552 -3324
rect -1544 -3326 -1542 -3324
rect -1528 -3326 -1526 -3324
rect -1520 -3326 -1518 -3324
rect -1504 -3326 -1502 -3324
rect -1496 -3326 -1494 -3324
rect -1486 -3326 -1484 -3324
rect -1478 -3326 -1476 -3324
rect -1462 -3326 -1460 -3324
rect -1454 -3326 -1452 -3324
rect -1444 -3326 -1442 -3324
rect -1436 -3326 -1434 -3324
rect -1420 -3326 -1418 -3324
rect -1412 -3326 -1410 -3324
rect -1402 -3326 -1400 -3324
rect -1394 -3326 -1392 -3324
rect -1378 -3326 -1376 -3324
rect -1370 -3326 -1368 -3324
rect -1229 -3326 -1227 -3324
rect -1219 -3326 -1217 -3324
rect -1203 -3326 -1201 -3324
rect -1195 -3326 -1193 -3324
rect -1179 -3326 -1177 -3324
rect -1171 -3326 -1169 -3324
rect -1161 -3326 -1159 -3324
rect -1153 -3326 -1151 -3324
rect -1137 -3326 -1135 -3324
rect -1129 -3326 -1127 -3324
rect -1119 -3326 -1117 -3324
rect -1111 -3326 -1109 -3324
rect -1095 -3326 -1093 -3324
rect -1087 -3326 -1085 -3324
rect -1077 -3326 -1075 -3324
rect -1069 -3326 -1067 -3324
rect -1053 -3326 -1051 -3324
rect -1045 -3326 -1043 -3324
rect -930 -3326 -928 -3324
rect -920 -3326 -918 -3324
rect -904 -3326 -902 -3324
rect -896 -3326 -894 -3324
rect -880 -3326 -878 -3324
rect -872 -3326 -870 -3324
rect -862 -3326 -860 -3324
rect -854 -3326 -852 -3324
rect -838 -3326 -836 -3324
rect -830 -3326 -828 -3324
rect -820 -3326 -818 -3324
rect -812 -3326 -810 -3324
rect -796 -3326 -794 -3324
rect -788 -3326 -786 -3324
rect -778 -3326 -776 -3324
rect -770 -3326 -768 -3324
rect -754 -3326 -752 -3324
rect -746 -3326 -744 -3324
rect -572 -3326 -570 -3324
rect -562 -3326 -560 -3324
rect -546 -3326 -544 -3324
rect -538 -3326 -536 -3324
rect -522 -3326 -520 -3324
rect -514 -3326 -512 -3324
rect -504 -3326 -502 -3324
rect -496 -3326 -494 -3324
rect -480 -3326 -478 -3324
rect -472 -3326 -470 -3324
rect -462 -3326 -460 -3324
rect -454 -3326 -452 -3324
rect -438 -3326 -436 -3324
rect -430 -3326 -428 -3324
rect -420 -3326 -418 -3324
rect -412 -3326 -410 -3324
rect -396 -3326 -394 -3324
rect -388 -3326 -386 -3324
rect -214 -3326 -212 -3324
rect -204 -3326 -202 -3324
rect -188 -3326 -186 -3324
rect -180 -3326 -178 -3324
rect -164 -3326 -162 -3324
rect -156 -3326 -154 -3324
rect -146 -3326 -144 -3324
rect -138 -3326 -136 -3324
rect -122 -3326 -120 -3324
rect -114 -3326 -112 -3324
rect -104 -3326 -102 -3324
rect -96 -3326 -94 -3324
rect -80 -3326 -78 -3324
rect -72 -3326 -70 -3324
rect -62 -3326 -60 -3324
rect -54 -3326 -52 -3324
rect -38 -3326 -36 -3324
rect -30 -3326 -28 -3324
rect 144 -3326 146 -3324
rect 154 -3326 156 -3324
rect 170 -3326 172 -3324
rect 178 -3326 180 -3324
rect 194 -3326 196 -3324
rect 202 -3326 204 -3324
rect 212 -3326 214 -3324
rect 220 -3326 222 -3324
rect 236 -3326 238 -3324
rect 244 -3326 246 -3324
rect 254 -3326 256 -3324
rect 262 -3326 264 -3324
rect 278 -3326 280 -3324
rect 286 -3326 288 -3324
rect 296 -3326 298 -3324
rect 304 -3326 306 -3324
rect 320 -3326 322 -3324
rect 328 -3326 330 -3324
rect 500 -3326 502 -3324
rect 510 -3326 512 -3324
rect 526 -3326 528 -3324
rect 534 -3326 536 -3324
rect 550 -3326 552 -3324
rect 558 -3326 560 -3324
rect 568 -3326 570 -3324
rect 576 -3326 578 -3324
rect 592 -3326 594 -3324
rect 600 -3326 602 -3324
rect 610 -3326 612 -3324
rect 618 -3326 620 -3324
rect 634 -3326 636 -3324
rect 642 -3326 644 -3324
rect 652 -3326 654 -3324
rect 660 -3326 662 -3324
rect 676 -3326 678 -3324
rect 684 -3326 686 -3324
rect 858 -3326 860 -3324
rect 868 -3326 870 -3324
rect 884 -3326 886 -3324
rect 892 -3326 894 -3324
rect 908 -3326 910 -3324
rect 916 -3326 918 -3324
rect 926 -3326 928 -3324
rect 934 -3326 936 -3324
rect 950 -3326 952 -3324
rect 958 -3326 960 -3324
rect 968 -3326 970 -3324
rect 976 -3326 978 -3324
rect 992 -3326 994 -3324
rect 1000 -3326 1002 -3324
rect 1010 -3326 1012 -3324
rect 1018 -3326 1020 -3324
rect 1034 -3326 1036 -3324
rect 1042 -3326 1044 -3324
rect 1216 -3326 1218 -3324
rect 1226 -3326 1228 -3324
rect 1242 -3326 1244 -3324
rect 1250 -3326 1252 -3324
rect 1266 -3326 1268 -3324
rect 1274 -3326 1276 -3324
rect 1284 -3326 1286 -3324
rect 1292 -3326 1294 -3324
rect 1308 -3326 1310 -3324
rect 1316 -3326 1318 -3324
rect 1326 -3326 1328 -3324
rect 1334 -3326 1336 -3324
rect 1350 -3326 1352 -3324
rect 1358 -3326 1360 -3324
rect 1368 -3326 1370 -3324
rect 1376 -3326 1378 -3324
rect 1392 -3326 1394 -3324
rect 1400 -3326 1402 -3324
rect -1304 -3355 -1302 -3353
rect -1296 -3355 -1294 -3353
rect -1286 -3355 -1284 -3353
rect -930 -3355 -928 -3353
rect -922 -3355 -920 -3353
rect -912 -3355 -910 -3353
rect -572 -3355 -570 -3353
rect -564 -3355 -562 -3353
rect -554 -3355 -552 -3353
rect -214 -3355 -212 -3353
rect -206 -3355 -204 -3353
rect -196 -3355 -194 -3353
rect 144 -3355 146 -3353
rect 152 -3355 154 -3353
rect 162 -3355 164 -3353
rect 500 -3355 502 -3353
rect 508 -3355 510 -3353
rect 518 -3355 520 -3353
rect 858 -3355 860 -3353
rect 866 -3355 868 -3353
rect 876 -3355 878 -3353
rect 1216 -3355 1218 -3353
rect 1224 -3355 1226 -3353
rect 1234 -3355 1236 -3353
rect -1304 -3431 -1302 -3363
rect -1296 -3387 -1294 -3363
rect -1296 -3431 -1294 -3391
rect -1286 -3431 -1284 -3363
rect -930 -3431 -928 -3363
rect -922 -3387 -920 -3363
rect -922 -3431 -920 -3391
rect -912 -3431 -910 -3363
rect -572 -3431 -570 -3363
rect -564 -3387 -562 -3363
rect -564 -3431 -562 -3391
rect -554 -3431 -552 -3363
rect -214 -3431 -212 -3363
rect -206 -3387 -204 -3363
rect -206 -3431 -204 -3391
rect -196 -3431 -194 -3363
rect 144 -3431 146 -3363
rect 152 -3387 154 -3363
rect 152 -3431 154 -3391
rect 162 -3431 164 -3363
rect 500 -3431 502 -3363
rect 508 -3387 510 -3363
rect 508 -3431 510 -3391
rect 518 -3431 520 -3363
rect 858 -3431 860 -3363
rect 866 -3387 868 -3363
rect 866 -3431 868 -3391
rect 876 -3431 878 -3363
rect 1216 -3431 1218 -3363
rect 1224 -3387 1226 -3363
rect 1224 -3431 1226 -3391
rect 1234 -3431 1236 -3363
rect -1304 -3437 -1302 -3435
rect -1296 -3437 -1294 -3435
rect -1286 -3437 -1284 -3435
rect -930 -3437 -928 -3435
rect -922 -3437 -920 -3435
rect -912 -3437 -910 -3435
rect -572 -3437 -570 -3435
rect -564 -3437 -562 -3435
rect -554 -3437 -552 -3435
rect -214 -3437 -212 -3435
rect -206 -3437 -204 -3435
rect -196 -3437 -194 -3435
rect 144 -3437 146 -3435
rect 152 -3437 154 -3435
rect 162 -3437 164 -3435
rect 500 -3437 502 -3435
rect 508 -3437 510 -3435
rect 518 -3437 520 -3435
rect 858 -3437 860 -3435
rect 866 -3437 868 -3435
rect 876 -3437 878 -3435
rect 1216 -3437 1218 -3435
rect 1224 -3437 1226 -3435
rect 1234 -3437 1236 -3435
rect -1229 -3514 -1227 -3512
rect -1219 -3514 -1217 -3512
rect -1203 -3514 -1201 -3512
rect -1193 -3514 -1191 -3512
rect -1185 -3514 -1183 -3512
rect -1175 -3514 -1173 -3512
rect -1159 -3514 -1157 -3512
rect -1151 -3514 -1149 -3512
rect -1141 -3514 -1139 -3512
rect -930 -3514 -928 -3512
rect -920 -3514 -918 -3512
rect -904 -3514 -902 -3512
rect -894 -3514 -892 -3512
rect -878 -3514 -876 -3512
rect -868 -3514 -866 -3512
rect -860 -3514 -858 -3512
rect -850 -3514 -848 -3512
rect -834 -3514 -832 -3512
rect -826 -3514 -824 -3512
rect -816 -3514 -814 -3512
rect -800 -3514 -798 -3512
rect -790 -3514 -788 -3512
rect -782 -3514 -780 -3512
rect -772 -3514 -770 -3512
rect -756 -3514 -754 -3512
rect -748 -3514 -746 -3512
rect -732 -3514 -730 -3512
rect -716 -3514 -714 -3512
rect -708 -3514 -706 -3512
rect -698 -3514 -696 -3512
rect -572 -3514 -570 -3512
rect -562 -3514 -560 -3512
rect -546 -3514 -544 -3512
rect -536 -3514 -534 -3512
rect -520 -3514 -518 -3512
rect -510 -3514 -508 -3512
rect -502 -3514 -500 -3512
rect -492 -3514 -490 -3512
rect -476 -3514 -474 -3512
rect -468 -3514 -466 -3512
rect -458 -3514 -456 -3512
rect -442 -3514 -440 -3512
rect -432 -3514 -430 -3512
rect -424 -3514 -422 -3512
rect -414 -3514 -412 -3512
rect -398 -3514 -396 -3512
rect -390 -3514 -388 -3512
rect -374 -3514 -372 -3512
rect -358 -3514 -356 -3512
rect -350 -3514 -348 -3512
rect -340 -3514 -338 -3512
rect -214 -3514 -212 -3512
rect -204 -3514 -202 -3512
rect -188 -3514 -186 -3512
rect -178 -3514 -176 -3512
rect -162 -3514 -160 -3512
rect -152 -3514 -150 -3512
rect -144 -3514 -142 -3512
rect -134 -3514 -132 -3512
rect -118 -3514 -116 -3512
rect -110 -3514 -108 -3512
rect -100 -3514 -98 -3512
rect -84 -3514 -82 -3512
rect -74 -3514 -72 -3512
rect -66 -3514 -64 -3512
rect -56 -3514 -54 -3512
rect -40 -3514 -38 -3512
rect -32 -3514 -30 -3512
rect -16 -3514 -14 -3512
rect 0 -3514 2 -3512
rect 8 -3514 10 -3512
rect 18 -3514 20 -3512
rect 144 -3514 146 -3512
rect 154 -3514 156 -3512
rect 170 -3514 172 -3512
rect 180 -3514 182 -3512
rect 196 -3514 198 -3512
rect 206 -3514 208 -3512
rect 214 -3514 216 -3512
rect 224 -3514 226 -3512
rect 240 -3514 242 -3512
rect 248 -3514 250 -3512
rect 258 -3514 260 -3512
rect 274 -3514 276 -3512
rect 284 -3514 286 -3512
rect 292 -3514 294 -3512
rect 302 -3514 304 -3512
rect 318 -3514 320 -3512
rect 326 -3514 328 -3512
rect 342 -3514 344 -3512
rect 358 -3514 360 -3512
rect 366 -3514 368 -3512
rect 376 -3514 378 -3512
rect 500 -3514 502 -3512
rect 510 -3514 512 -3512
rect 526 -3514 528 -3512
rect 536 -3514 538 -3512
rect 552 -3514 554 -3512
rect 562 -3514 564 -3512
rect 570 -3514 572 -3512
rect 580 -3514 582 -3512
rect 596 -3514 598 -3512
rect 604 -3514 606 -3512
rect 614 -3514 616 -3512
rect 630 -3514 632 -3512
rect 640 -3514 642 -3512
rect 648 -3514 650 -3512
rect 658 -3514 660 -3512
rect 674 -3514 676 -3512
rect 682 -3514 684 -3512
rect 698 -3514 700 -3512
rect 714 -3514 716 -3512
rect 722 -3514 724 -3512
rect 732 -3514 734 -3512
rect 858 -3514 860 -3512
rect 868 -3514 870 -3512
rect 884 -3514 886 -3512
rect 894 -3514 896 -3512
rect 910 -3514 912 -3512
rect 920 -3514 922 -3512
rect 928 -3514 930 -3512
rect 938 -3514 940 -3512
rect 954 -3514 956 -3512
rect 962 -3514 964 -3512
rect 972 -3514 974 -3512
rect 988 -3514 990 -3512
rect 998 -3514 1000 -3512
rect 1006 -3514 1008 -3512
rect 1016 -3514 1018 -3512
rect 1032 -3514 1034 -3512
rect 1040 -3514 1042 -3512
rect 1056 -3514 1058 -3512
rect 1072 -3514 1074 -3512
rect 1080 -3514 1082 -3512
rect 1090 -3514 1092 -3512
rect 1216 -3514 1218 -3512
rect 1226 -3514 1228 -3512
rect 1242 -3514 1244 -3512
rect 1252 -3514 1254 -3512
rect 1268 -3514 1270 -3512
rect 1278 -3514 1280 -3512
rect 1286 -3514 1288 -3512
rect 1296 -3514 1298 -3512
rect 1312 -3514 1314 -3512
rect 1320 -3514 1322 -3512
rect 1330 -3514 1332 -3512
rect 1346 -3514 1348 -3512
rect 1356 -3514 1358 -3512
rect 1364 -3514 1366 -3512
rect 1374 -3514 1376 -3512
rect 1390 -3514 1392 -3512
rect 1398 -3514 1400 -3512
rect 1414 -3514 1416 -3512
rect 1430 -3514 1432 -3512
rect 1438 -3514 1440 -3512
rect 1448 -3514 1450 -3512
rect -1229 -3590 -1227 -3522
rect -1219 -3590 -1217 -3522
rect -1203 -3590 -1201 -3522
rect -1193 -3590 -1191 -3522
rect -1185 -3590 -1183 -3522
rect -1175 -3590 -1173 -3522
rect -1159 -3590 -1157 -3522
rect -1151 -3590 -1149 -3522
rect -1141 -3590 -1139 -3522
rect -930 -3590 -928 -3522
rect -920 -3590 -918 -3522
rect -904 -3590 -902 -3522
rect -894 -3590 -892 -3522
rect -878 -3590 -876 -3522
rect -868 -3590 -866 -3522
rect -860 -3590 -858 -3522
rect -850 -3590 -848 -3522
rect -834 -3590 -832 -3522
rect -826 -3590 -824 -3522
rect -816 -3590 -814 -3522
rect -800 -3590 -798 -3522
rect -790 -3590 -788 -3522
rect -782 -3590 -780 -3522
rect -772 -3590 -770 -3522
rect -756 -3590 -754 -3522
rect -748 -3590 -746 -3522
rect -732 -3590 -730 -3522
rect -716 -3590 -714 -3522
rect -708 -3590 -706 -3522
rect -698 -3590 -696 -3522
rect -572 -3590 -570 -3522
rect -562 -3590 -560 -3522
rect -546 -3590 -544 -3522
rect -536 -3590 -534 -3522
rect -520 -3590 -518 -3522
rect -510 -3590 -508 -3522
rect -502 -3590 -500 -3522
rect -492 -3590 -490 -3522
rect -476 -3590 -474 -3522
rect -468 -3590 -466 -3522
rect -458 -3590 -456 -3522
rect -442 -3590 -440 -3522
rect -432 -3590 -430 -3522
rect -424 -3590 -422 -3522
rect -414 -3590 -412 -3522
rect -398 -3590 -396 -3522
rect -390 -3590 -388 -3522
rect -374 -3590 -372 -3522
rect -358 -3590 -356 -3522
rect -350 -3590 -348 -3522
rect -340 -3590 -338 -3522
rect -214 -3590 -212 -3522
rect -204 -3590 -202 -3522
rect -188 -3590 -186 -3522
rect -178 -3590 -176 -3522
rect -162 -3590 -160 -3522
rect -152 -3590 -150 -3522
rect -144 -3590 -142 -3522
rect -134 -3590 -132 -3522
rect -118 -3590 -116 -3522
rect -110 -3590 -108 -3522
rect -100 -3590 -98 -3522
rect -84 -3590 -82 -3522
rect -74 -3590 -72 -3522
rect -66 -3590 -64 -3522
rect -56 -3590 -54 -3522
rect -40 -3590 -38 -3522
rect -32 -3590 -30 -3522
rect -16 -3590 -14 -3522
rect 0 -3590 2 -3522
rect 8 -3590 10 -3522
rect 18 -3590 20 -3522
rect 144 -3590 146 -3522
rect 154 -3590 156 -3522
rect 170 -3590 172 -3522
rect 180 -3590 182 -3522
rect 196 -3590 198 -3522
rect 206 -3590 208 -3522
rect 214 -3590 216 -3522
rect 224 -3590 226 -3522
rect 240 -3590 242 -3522
rect 248 -3590 250 -3522
rect 258 -3590 260 -3522
rect 274 -3590 276 -3522
rect 284 -3590 286 -3522
rect 292 -3590 294 -3522
rect 302 -3590 304 -3522
rect 318 -3590 320 -3522
rect 326 -3590 328 -3522
rect 342 -3590 344 -3522
rect 358 -3590 360 -3522
rect 366 -3590 368 -3522
rect 376 -3590 378 -3522
rect 500 -3590 502 -3522
rect 510 -3590 512 -3522
rect 526 -3590 528 -3522
rect 536 -3590 538 -3522
rect 552 -3590 554 -3522
rect 562 -3590 564 -3522
rect 570 -3590 572 -3522
rect 580 -3590 582 -3522
rect 596 -3590 598 -3522
rect 604 -3590 606 -3522
rect 614 -3590 616 -3522
rect 630 -3590 632 -3522
rect 640 -3590 642 -3522
rect 648 -3590 650 -3522
rect 658 -3590 660 -3522
rect 674 -3590 676 -3522
rect 682 -3590 684 -3522
rect 698 -3590 700 -3522
rect 714 -3590 716 -3522
rect 722 -3590 724 -3522
rect 732 -3590 734 -3522
rect 858 -3590 860 -3522
rect 868 -3590 870 -3522
rect 884 -3590 886 -3522
rect 894 -3590 896 -3522
rect 910 -3590 912 -3522
rect 920 -3590 922 -3522
rect 928 -3590 930 -3522
rect 938 -3590 940 -3522
rect 954 -3590 956 -3522
rect 962 -3590 964 -3522
rect 972 -3590 974 -3522
rect 988 -3590 990 -3522
rect 998 -3590 1000 -3522
rect 1006 -3590 1008 -3522
rect 1016 -3590 1018 -3522
rect 1032 -3590 1034 -3522
rect 1040 -3590 1042 -3522
rect 1056 -3590 1058 -3522
rect 1072 -3590 1074 -3522
rect 1080 -3590 1082 -3522
rect 1090 -3590 1092 -3522
rect 1216 -3590 1218 -3522
rect 1226 -3590 1228 -3522
rect 1242 -3590 1244 -3522
rect 1252 -3590 1254 -3522
rect 1268 -3590 1270 -3522
rect 1278 -3590 1280 -3522
rect 1286 -3590 1288 -3522
rect 1296 -3590 1298 -3522
rect 1312 -3590 1314 -3522
rect 1320 -3590 1322 -3522
rect 1330 -3590 1332 -3522
rect 1346 -3590 1348 -3522
rect 1356 -3590 1358 -3522
rect 1364 -3590 1366 -3522
rect 1374 -3590 1376 -3522
rect 1390 -3590 1392 -3522
rect 1398 -3590 1400 -3522
rect 1414 -3590 1416 -3522
rect 1430 -3590 1432 -3522
rect 1438 -3590 1440 -3522
rect 1448 -3590 1450 -3522
rect -1229 -3596 -1227 -3594
rect -1219 -3596 -1217 -3594
rect -1203 -3596 -1201 -3594
rect -1193 -3596 -1191 -3594
rect -1185 -3596 -1183 -3594
rect -1175 -3596 -1173 -3594
rect -1159 -3596 -1157 -3594
rect -1151 -3596 -1149 -3594
rect -1141 -3596 -1139 -3594
rect -930 -3596 -928 -3594
rect -920 -3596 -918 -3594
rect -904 -3596 -902 -3594
rect -894 -3596 -892 -3594
rect -878 -3596 -876 -3594
rect -868 -3596 -866 -3594
rect -860 -3596 -858 -3594
rect -850 -3596 -848 -3594
rect -834 -3596 -832 -3594
rect -826 -3596 -824 -3594
rect -816 -3596 -814 -3594
rect -800 -3596 -798 -3594
rect -790 -3596 -788 -3594
rect -782 -3596 -780 -3594
rect -772 -3596 -770 -3594
rect -756 -3596 -754 -3594
rect -748 -3596 -746 -3594
rect -732 -3596 -730 -3594
rect -716 -3596 -714 -3594
rect -708 -3596 -706 -3594
rect -698 -3596 -696 -3594
rect -572 -3596 -570 -3594
rect -562 -3596 -560 -3594
rect -546 -3596 -544 -3594
rect -536 -3596 -534 -3594
rect -520 -3596 -518 -3594
rect -510 -3596 -508 -3594
rect -502 -3596 -500 -3594
rect -492 -3596 -490 -3594
rect -476 -3596 -474 -3594
rect -468 -3596 -466 -3594
rect -458 -3596 -456 -3594
rect -442 -3596 -440 -3594
rect -432 -3596 -430 -3594
rect -424 -3596 -422 -3594
rect -414 -3596 -412 -3594
rect -398 -3596 -396 -3594
rect -390 -3596 -388 -3594
rect -374 -3596 -372 -3594
rect -358 -3596 -356 -3594
rect -350 -3596 -348 -3594
rect -340 -3596 -338 -3594
rect -214 -3596 -212 -3594
rect -204 -3596 -202 -3594
rect -188 -3596 -186 -3594
rect -178 -3596 -176 -3594
rect -162 -3596 -160 -3594
rect -152 -3596 -150 -3594
rect -144 -3596 -142 -3594
rect -134 -3596 -132 -3594
rect -118 -3596 -116 -3594
rect -110 -3596 -108 -3594
rect -100 -3596 -98 -3594
rect -84 -3596 -82 -3594
rect -74 -3596 -72 -3594
rect -66 -3596 -64 -3594
rect -56 -3596 -54 -3594
rect -40 -3596 -38 -3594
rect -32 -3596 -30 -3594
rect -16 -3596 -14 -3594
rect 0 -3596 2 -3594
rect 8 -3596 10 -3594
rect 18 -3596 20 -3594
rect 144 -3596 146 -3594
rect 154 -3596 156 -3594
rect 170 -3596 172 -3594
rect 180 -3596 182 -3594
rect 196 -3596 198 -3594
rect 206 -3596 208 -3594
rect 214 -3596 216 -3594
rect 224 -3596 226 -3594
rect 240 -3596 242 -3594
rect 248 -3596 250 -3594
rect 258 -3596 260 -3594
rect 274 -3596 276 -3594
rect 284 -3596 286 -3594
rect 292 -3596 294 -3594
rect 302 -3596 304 -3594
rect 318 -3596 320 -3594
rect 326 -3596 328 -3594
rect 342 -3596 344 -3594
rect 358 -3596 360 -3594
rect 366 -3596 368 -3594
rect 376 -3596 378 -3594
rect 500 -3596 502 -3594
rect 510 -3596 512 -3594
rect 526 -3596 528 -3594
rect 536 -3596 538 -3594
rect 552 -3596 554 -3594
rect 562 -3596 564 -3594
rect 570 -3596 572 -3594
rect 580 -3596 582 -3594
rect 596 -3596 598 -3594
rect 604 -3596 606 -3594
rect 614 -3596 616 -3594
rect 630 -3596 632 -3594
rect 640 -3596 642 -3594
rect 648 -3596 650 -3594
rect 658 -3596 660 -3594
rect 674 -3596 676 -3594
rect 682 -3596 684 -3594
rect 698 -3596 700 -3594
rect 714 -3596 716 -3594
rect 722 -3596 724 -3594
rect 732 -3596 734 -3594
rect 858 -3596 860 -3594
rect 868 -3596 870 -3594
rect 884 -3596 886 -3594
rect 894 -3596 896 -3594
rect 910 -3596 912 -3594
rect 920 -3596 922 -3594
rect 928 -3596 930 -3594
rect 938 -3596 940 -3594
rect 954 -3596 956 -3594
rect 962 -3596 964 -3594
rect 972 -3596 974 -3594
rect 988 -3596 990 -3594
rect 998 -3596 1000 -3594
rect 1006 -3596 1008 -3594
rect 1016 -3596 1018 -3594
rect 1032 -3596 1034 -3594
rect 1040 -3596 1042 -3594
rect 1056 -3596 1058 -3594
rect 1072 -3596 1074 -3594
rect 1080 -3596 1082 -3594
rect 1090 -3596 1092 -3594
rect 1216 -3596 1218 -3594
rect 1226 -3596 1228 -3594
rect 1242 -3596 1244 -3594
rect 1252 -3596 1254 -3594
rect 1268 -3596 1270 -3594
rect 1278 -3596 1280 -3594
rect 1286 -3596 1288 -3594
rect 1296 -3596 1298 -3594
rect 1312 -3596 1314 -3594
rect 1320 -3596 1322 -3594
rect 1330 -3596 1332 -3594
rect 1346 -3596 1348 -3594
rect 1356 -3596 1358 -3594
rect 1364 -3596 1366 -3594
rect 1374 -3596 1376 -3594
rect 1390 -3596 1392 -3594
rect 1398 -3596 1400 -3594
rect 1414 -3596 1416 -3594
rect 1430 -3596 1432 -3594
rect 1438 -3596 1440 -3594
rect 1448 -3596 1450 -3594
rect -1817 -3644 -1815 -3642
rect -1807 -3644 -1805 -3642
rect -1791 -3644 -1789 -3642
rect -1783 -3644 -1781 -3642
rect -1767 -3644 -1765 -3642
rect -1759 -3644 -1757 -3642
rect -1749 -3644 -1747 -3642
rect -1741 -3644 -1739 -3642
rect -1725 -3644 -1723 -3642
rect -1717 -3644 -1715 -3642
rect -1707 -3644 -1705 -3642
rect -1699 -3644 -1697 -3642
rect -1683 -3644 -1681 -3642
rect -1675 -3644 -1673 -3642
rect -1665 -3644 -1663 -3642
rect -1657 -3644 -1655 -3642
rect -1641 -3644 -1639 -3642
rect -1633 -3644 -1631 -3642
rect -1554 -3644 -1552 -3642
rect -1544 -3644 -1542 -3642
rect -1528 -3644 -1526 -3642
rect -1520 -3644 -1518 -3642
rect -1504 -3644 -1502 -3642
rect -1496 -3644 -1494 -3642
rect -1486 -3644 -1484 -3642
rect -1478 -3644 -1476 -3642
rect -1462 -3644 -1460 -3642
rect -1454 -3644 -1452 -3642
rect -1444 -3644 -1442 -3642
rect -1436 -3644 -1434 -3642
rect -1420 -3644 -1418 -3642
rect -1412 -3644 -1410 -3642
rect -1402 -3644 -1400 -3642
rect -1394 -3644 -1392 -3642
rect -1378 -3644 -1376 -3642
rect -1370 -3644 -1368 -3642
rect -1229 -3644 -1227 -3642
rect -1219 -3644 -1217 -3642
rect -1203 -3644 -1201 -3642
rect -1195 -3644 -1193 -3642
rect -1179 -3644 -1177 -3642
rect -1171 -3644 -1169 -3642
rect -1161 -3644 -1159 -3642
rect -1153 -3644 -1151 -3642
rect -1137 -3644 -1135 -3642
rect -1129 -3644 -1127 -3642
rect -1119 -3644 -1117 -3642
rect -1111 -3644 -1109 -3642
rect -1095 -3644 -1093 -3642
rect -1087 -3644 -1085 -3642
rect -1077 -3644 -1075 -3642
rect -1069 -3644 -1067 -3642
rect -1053 -3644 -1051 -3642
rect -1045 -3644 -1043 -3642
rect -929 -3644 -927 -3642
rect -919 -3644 -917 -3642
rect -903 -3644 -901 -3642
rect -895 -3644 -893 -3642
rect -879 -3644 -877 -3642
rect -871 -3644 -869 -3642
rect -861 -3644 -859 -3642
rect -853 -3644 -851 -3642
rect -837 -3644 -835 -3642
rect -829 -3644 -827 -3642
rect -819 -3644 -817 -3642
rect -811 -3644 -809 -3642
rect -795 -3644 -793 -3642
rect -787 -3644 -785 -3642
rect -777 -3644 -775 -3642
rect -769 -3644 -767 -3642
rect -753 -3644 -751 -3642
rect -745 -3644 -743 -3642
rect -572 -3644 -570 -3642
rect -562 -3644 -560 -3642
rect -546 -3644 -544 -3642
rect -538 -3644 -536 -3642
rect -522 -3644 -520 -3642
rect -514 -3644 -512 -3642
rect -504 -3644 -502 -3642
rect -496 -3644 -494 -3642
rect -480 -3644 -478 -3642
rect -472 -3644 -470 -3642
rect -462 -3644 -460 -3642
rect -454 -3644 -452 -3642
rect -438 -3644 -436 -3642
rect -430 -3644 -428 -3642
rect -420 -3644 -418 -3642
rect -412 -3644 -410 -3642
rect -396 -3644 -394 -3642
rect -388 -3644 -386 -3642
rect -214 -3644 -212 -3642
rect -204 -3644 -202 -3642
rect -188 -3644 -186 -3642
rect -180 -3644 -178 -3642
rect -164 -3644 -162 -3642
rect -156 -3644 -154 -3642
rect -146 -3644 -144 -3642
rect -138 -3644 -136 -3642
rect -122 -3644 -120 -3642
rect -114 -3644 -112 -3642
rect -104 -3644 -102 -3642
rect -96 -3644 -94 -3642
rect -80 -3644 -78 -3642
rect -72 -3644 -70 -3642
rect -62 -3644 -60 -3642
rect -54 -3644 -52 -3642
rect -38 -3644 -36 -3642
rect -30 -3644 -28 -3642
rect -1817 -3720 -1815 -3652
rect -1807 -3720 -1805 -3652
rect -1791 -3720 -1789 -3652
rect -1783 -3720 -1781 -3652
rect -1767 -3720 -1765 -3652
rect -1759 -3720 -1757 -3652
rect -1749 -3720 -1747 -3652
rect -1741 -3720 -1739 -3652
rect -1725 -3720 -1723 -3652
rect -1717 -3685 -1715 -3652
rect -1707 -3685 -1705 -3652
rect -1717 -3687 -1705 -3685
rect -1717 -3720 -1715 -3687
rect -1707 -3720 -1705 -3687
rect -1699 -3720 -1697 -3652
rect -1683 -3720 -1681 -3652
rect -1675 -3720 -1673 -3652
rect -1665 -3720 -1663 -3652
rect -1657 -3720 -1655 -3652
rect -1641 -3720 -1639 -3652
rect -1633 -3720 -1631 -3652
rect -1554 -3720 -1552 -3652
rect -1544 -3720 -1542 -3652
rect -1528 -3720 -1526 -3652
rect -1520 -3720 -1518 -3652
rect -1504 -3720 -1502 -3652
rect -1496 -3720 -1494 -3652
rect -1486 -3720 -1484 -3652
rect -1478 -3720 -1476 -3652
rect -1462 -3720 -1460 -3652
rect -1454 -3685 -1452 -3652
rect -1444 -3685 -1442 -3652
rect -1454 -3687 -1442 -3685
rect -1454 -3720 -1452 -3687
rect -1444 -3720 -1442 -3687
rect -1436 -3720 -1434 -3652
rect -1420 -3720 -1418 -3652
rect -1412 -3720 -1410 -3652
rect -1402 -3720 -1400 -3652
rect -1394 -3720 -1392 -3652
rect -1378 -3720 -1376 -3652
rect -1370 -3720 -1368 -3652
rect -1229 -3720 -1227 -3652
rect -1219 -3720 -1217 -3652
rect -1203 -3720 -1201 -3652
rect -1195 -3720 -1193 -3652
rect -1179 -3720 -1177 -3652
rect -1171 -3720 -1169 -3652
rect -1161 -3720 -1159 -3652
rect -1153 -3720 -1151 -3652
rect -1137 -3720 -1135 -3652
rect -1129 -3685 -1127 -3652
rect -1119 -3685 -1117 -3652
rect -1129 -3687 -1117 -3685
rect -1129 -3720 -1127 -3687
rect -1119 -3720 -1117 -3687
rect -1111 -3720 -1109 -3652
rect -1095 -3720 -1093 -3652
rect -1087 -3720 -1085 -3652
rect -1077 -3720 -1075 -3652
rect -1069 -3720 -1067 -3652
rect -1053 -3720 -1051 -3652
rect -1045 -3720 -1043 -3652
rect -929 -3720 -927 -3652
rect -919 -3720 -917 -3652
rect -903 -3720 -901 -3652
rect -895 -3720 -893 -3652
rect -879 -3720 -877 -3652
rect -871 -3720 -869 -3652
rect -861 -3720 -859 -3652
rect -853 -3720 -851 -3652
rect -837 -3720 -835 -3652
rect -829 -3685 -827 -3652
rect -819 -3685 -817 -3652
rect -829 -3687 -817 -3685
rect -829 -3720 -827 -3687
rect -819 -3720 -817 -3687
rect -811 -3720 -809 -3652
rect -795 -3720 -793 -3652
rect -787 -3720 -785 -3652
rect -777 -3720 -775 -3652
rect -769 -3720 -767 -3652
rect -753 -3720 -751 -3652
rect -745 -3720 -743 -3652
rect -572 -3720 -570 -3652
rect -562 -3720 -560 -3652
rect -546 -3720 -544 -3652
rect -538 -3720 -536 -3652
rect -522 -3720 -520 -3652
rect -514 -3720 -512 -3652
rect -504 -3720 -502 -3652
rect -496 -3720 -494 -3652
rect -480 -3720 -478 -3652
rect -472 -3685 -470 -3652
rect -462 -3685 -460 -3652
rect -472 -3687 -460 -3685
rect -472 -3720 -470 -3687
rect -462 -3720 -460 -3687
rect -454 -3720 -452 -3652
rect -438 -3720 -436 -3652
rect -430 -3720 -428 -3652
rect -420 -3720 -418 -3652
rect -412 -3720 -410 -3652
rect -396 -3720 -394 -3652
rect -388 -3720 -386 -3652
rect -214 -3720 -212 -3652
rect -204 -3720 -202 -3652
rect -188 -3720 -186 -3652
rect -180 -3720 -178 -3652
rect -164 -3720 -162 -3652
rect -156 -3720 -154 -3652
rect -146 -3720 -144 -3652
rect -138 -3720 -136 -3652
rect -122 -3720 -120 -3652
rect -114 -3685 -112 -3652
rect -104 -3685 -102 -3652
rect -114 -3687 -102 -3685
rect -114 -3720 -112 -3687
rect -104 -3720 -102 -3687
rect -96 -3720 -94 -3652
rect -80 -3720 -78 -3652
rect -72 -3720 -70 -3652
rect -62 -3720 -60 -3652
rect -54 -3720 -52 -3652
rect -38 -3720 -36 -3652
rect -30 -3720 -28 -3652
rect -1817 -3726 -1815 -3724
rect -1807 -3726 -1805 -3724
rect -1791 -3726 -1789 -3724
rect -1783 -3726 -1781 -3724
rect -1767 -3726 -1765 -3724
rect -1759 -3726 -1757 -3724
rect -1749 -3726 -1747 -3724
rect -1741 -3726 -1739 -3724
rect -1725 -3726 -1723 -3724
rect -1717 -3726 -1715 -3724
rect -1707 -3726 -1705 -3724
rect -1699 -3726 -1697 -3724
rect -1683 -3726 -1681 -3724
rect -1675 -3726 -1673 -3724
rect -1665 -3726 -1663 -3724
rect -1657 -3726 -1655 -3724
rect -1641 -3726 -1639 -3724
rect -1633 -3726 -1631 -3724
rect -1554 -3726 -1552 -3724
rect -1544 -3726 -1542 -3724
rect -1528 -3726 -1526 -3724
rect -1520 -3726 -1518 -3724
rect -1504 -3726 -1502 -3724
rect -1496 -3726 -1494 -3724
rect -1486 -3726 -1484 -3724
rect -1478 -3726 -1476 -3724
rect -1462 -3726 -1460 -3724
rect -1454 -3726 -1452 -3724
rect -1444 -3726 -1442 -3724
rect -1436 -3726 -1434 -3724
rect -1420 -3726 -1418 -3724
rect -1412 -3726 -1410 -3724
rect -1402 -3726 -1400 -3724
rect -1394 -3726 -1392 -3724
rect -1378 -3726 -1376 -3724
rect -1370 -3726 -1368 -3724
rect -1229 -3726 -1227 -3724
rect -1219 -3726 -1217 -3724
rect -1203 -3726 -1201 -3724
rect -1195 -3726 -1193 -3724
rect -1179 -3726 -1177 -3724
rect -1171 -3726 -1169 -3724
rect -1161 -3726 -1159 -3724
rect -1153 -3726 -1151 -3724
rect -1137 -3726 -1135 -3724
rect -1129 -3726 -1127 -3724
rect -1119 -3726 -1117 -3724
rect -1111 -3726 -1109 -3724
rect -1095 -3726 -1093 -3724
rect -1087 -3726 -1085 -3724
rect -1077 -3726 -1075 -3724
rect -1069 -3726 -1067 -3724
rect -1053 -3726 -1051 -3724
rect -1045 -3726 -1043 -3724
rect -929 -3726 -927 -3724
rect -919 -3726 -917 -3724
rect -903 -3726 -901 -3724
rect -895 -3726 -893 -3724
rect -879 -3726 -877 -3724
rect -871 -3726 -869 -3724
rect -861 -3726 -859 -3724
rect -853 -3726 -851 -3724
rect -837 -3726 -835 -3724
rect -829 -3726 -827 -3724
rect -819 -3726 -817 -3724
rect -811 -3726 -809 -3724
rect -795 -3726 -793 -3724
rect -787 -3726 -785 -3724
rect -777 -3726 -775 -3724
rect -769 -3726 -767 -3724
rect -753 -3726 -751 -3724
rect -745 -3726 -743 -3724
rect -572 -3726 -570 -3724
rect -562 -3726 -560 -3724
rect -546 -3726 -544 -3724
rect -538 -3726 -536 -3724
rect -522 -3726 -520 -3724
rect -514 -3726 -512 -3724
rect -504 -3726 -502 -3724
rect -496 -3726 -494 -3724
rect -480 -3726 -478 -3724
rect -472 -3726 -470 -3724
rect -462 -3726 -460 -3724
rect -454 -3726 -452 -3724
rect -438 -3726 -436 -3724
rect -430 -3726 -428 -3724
rect -420 -3726 -418 -3724
rect -412 -3726 -410 -3724
rect -396 -3726 -394 -3724
rect -388 -3726 -386 -3724
rect -214 -3726 -212 -3724
rect -204 -3726 -202 -3724
rect -188 -3726 -186 -3724
rect -180 -3726 -178 -3724
rect -164 -3726 -162 -3724
rect -156 -3726 -154 -3724
rect -146 -3726 -144 -3724
rect -138 -3726 -136 -3724
rect -122 -3726 -120 -3724
rect -114 -3726 -112 -3724
rect -104 -3726 -102 -3724
rect -96 -3726 -94 -3724
rect -80 -3726 -78 -3724
rect -72 -3726 -70 -3724
rect -62 -3726 -60 -3724
rect -54 -3726 -52 -3724
rect -38 -3726 -36 -3724
rect -30 -3726 -28 -3724
rect -1554 -3815 -1552 -3813
rect -1544 -3815 -1542 -3813
rect -1528 -3815 -1526 -3813
rect -1520 -3815 -1518 -3813
rect -1504 -3815 -1502 -3813
rect -1496 -3815 -1494 -3813
rect -1486 -3815 -1484 -3813
rect -1478 -3815 -1476 -3813
rect -1462 -3815 -1460 -3813
rect -1454 -3815 -1452 -3813
rect -1444 -3815 -1442 -3813
rect -1436 -3815 -1434 -3813
rect -1420 -3815 -1418 -3813
rect -1412 -3815 -1410 -3813
rect -1402 -3815 -1400 -3813
rect -1394 -3815 -1392 -3813
rect -1378 -3815 -1376 -3813
rect -1370 -3815 -1368 -3813
rect -1229 -3815 -1227 -3813
rect -1219 -3815 -1217 -3813
rect -1203 -3815 -1201 -3813
rect -1195 -3815 -1193 -3813
rect -1179 -3815 -1177 -3813
rect -1171 -3815 -1169 -3813
rect -1161 -3815 -1159 -3813
rect -1153 -3815 -1151 -3813
rect -1137 -3815 -1135 -3813
rect -1129 -3815 -1127 -3813
rect -1119 -3815 -1117 -3813
rect -1111 -3815 -1109 -3813
rect -1095 -3815 -1093 -3813
rect -1087 -3815 -1085 -3813
rect -1077 -3815 -1075 -3813
rect -1069 -3815 -1067 -3813
rect -1053 -3815 -1051 -3813
rect -1045 -3815 -1043 -3813
rect -929 -3815 -927 -3813
rect -919 -3815 -917 -3813
rect -903 -3815 -901 -3813
rect -895 -3815 -893 -3813
rect -879 -3815 -877 -3813
rect -871 -3815 -869 -3813
rect -861 -3815 -859 -3813
rect -853 -3815 -851 -3813
rect -837 -3815 -835 -3813
rect -829 -3815 -827 -3813
rect -819 -3815 -817 -3813
rect -811 -3815 -809 -3813
rect -795 -3815 -793 -3813
rect -787 -3815 -785 -3813
rect -777 -3815 -775 -3813
rect -769 -3815 -767 -3813
rect -753 -3815 -751 -3813
rect -745 -3815 -743 -3813
rect -572 -3815 -570 -3813
rect -562 -3815 -560 -3813
rect -546 -3815 -544 -3813
rect -538 -3815 -536 -3813
rect -522 -3815 -520 -3813
rect -514 -3815 -512 -3813
rect -504 -3815 -502 -3813
rect -496 -3815 -494 -3813
rect -480 -3815 -478 -3813
rect -472 -3815 -470 -3813
rect -462 -3815 -460 -3813
rect -454 -3815 -452 -3813
rect -438 -3815 -436 -3813
rect -430 -3815 -428 -3813
rect -420 -3815 -418 -3813
rect -412 -3815 -410 -3813
rect -396 -3815 -394 -3813
rect -388 -3815 -386 -3813
rect -214 -3815 -212 -3813
rect -204 -3815 -202 -3813
rect -188 -3815 -186 -3813
rect -180 -3815 -178 -3813
rect -164 -3815 -162 -3813
rect -156 -3815 -154 -3813
rect -146 -3815 -144 -3813
rect -138 -3815 -136 -3813
rect -122 -3815 -120 -3813
rect -114 -3815 -112 -3813
rect -104 -3815 -102 -3813
rect -96 -3815 -94 -3813
rect -80 -3815 -78 -3813
rect -72 -3815 -70 -3813
rect -62 -3815 -60 -3813
rect -54 -3815 -52 -3813
rect -38 -3815 -36 -3813
rect -30 -3815 -28 -3813
rect 144 -3815 146 -3813
rect 154 -3815 156 -3813
rect 170 -3815 172 -3813
rect 178 -3815 180 -3813
rect 194 -3815 196 -3813
rect 202 -3815 204 -3813
rect 212 -3815 214 -3813
rect 220 -3815 222 -3813
rect 236 -3815 238 -3813
rect 244 -3815 246 -3813
rect 254 -3815 256 -3813
rect 262 -3815 264 -3813
rect 278 -3815 280 -3813
rect 286 -3815 288 -3813
rect 296 -3815 298 -3813
rect 304 -3815 306 -3813
rect 320 -3815 322 -3813
rect 328 -3815 330 -3813
rect 500 -3815 502 -3813
rect 510 -3815 512 -3813
rect 526 -3815 528 -3813
rect 534 -3815 536 -3813
rect 550 -3815 552 -3813
rect 558 -3815 560 -3813
rect 568 -3815 570 -3813
rect 576 -3815 578 -3813
rect 592 -3815 594 -3813
rect 600 -3815 602 -3813
rect 610 -3815 612 -3813
rect 618 -3815 620 -3813
rect 634 -3815 636 -3813
rect 642 -3815 644 -3813
rect 652 -3815 654 -3813
rect 660 -3815 662 -3813
rect 676 -3815 678 -3813
rect 684 -3815 686 -3813
rect 858 -3815 860 -3813
rect 868 -3815 870 -3813
rect 884 -3815 886 -3813
rect 892 -3815 894 -3813
rect 908 -3815 910 -3813
rect 916 -3815 918 -3813
rect 926 -3815 928 -3813
rect 934 -3815 936 -3813
rect 950 -3815 952 -3813
rect 958 -3815 960 -3813
rect 968 -3815 970 -3813
rect 976 -3815 978 -3813
rect 992 -3815 994 -3813
rect 1000 -3815 1002 -3813
rect 1010 -3815 1012 -3813
rect 1018 -3815 1020 -3813
rect 1034 -3815 1036 -3813
rect 1042 -3815 1044 -3813
rect 1216 -3815 1218 -3813
rect 1226 -3815 1228 -3813
rect 1242 -3815 1244 -3813
rect 1250 -3815 1252 -3813
rect 1266 -3815 1268 -3813
rect 1274 -3815 1276 -3813
rect 1284 -3815 1286 -3813
rect 1292 -3815 1294 -3813
rect 1308 -3815 1310 -3813
rect 1316 -3815 1318 -3813
rect 1326 -3815 1328 -3813
rect 1334 -3815 1336 -3813
rect 1350 -3815 1352 -3813
rect 1358 -3815 1360 -3813
rect 1368 -3815 1370 -3813
rect 1376 -3815 1378 -3813
rect 1392 -3815 1394 -3813
rect 1400 -3815 1402 -3813
rect -1554 -3891 -1552 -3823
rect -1544 -3891 -1542 -3823
rect -1528 -3891 -1526 -3823
rect -1520 -3891 -1518 -3823
rect -1504 -3891 -1502 -3823
rect -1496 -3891 -1494 -3823
rect -1486 -3891 -1484 -3823
rect -1478 -3891 -1476 -3823
rect -1462 -3891 -1460 -3823
rect -1454 -3856 -1452 -3823
rect -1444 -3856 -1442 -3823
rect -1454 -3858 -1442 -3856
rect -1454 -3891 -1452 -3858
rect -1444 -3891 -1442 -3858
rect -1436 -3891 -1434 -3823
rect -1420 -3891 -1418 -3823
rect -1412 -3891 -1410 -3823
rect -1402 -3891 -1400 -3823
rect -1394 -3891 -1392 -3823
rect -1378 -3891 -1376 -3823
rect -1370 -3891 -1368 -3823
rect -1229 -3891 -1227 -3823
rect -1219 -3891 -1217 -3823
rect -1203 -3891 -1201 -3823
rect -1195 -3891 -1193 -3823
rect -1179 -3891 -1177 -3823
rect -1171 -3891 -1169 -3823
rect -1161 -3891 -1159 -3823
rect -1153 -3891 -1151 -3823
rect -1137 -3891 -1135 -3823
rect -1129 -3856 -1127 -3823
rect -1119 -3856 -1117 -3823
rect -1129 -3858 -1117 -3856
rect -1129 -3891 -1127 -3858
rect -1119 -3891 -1117 -3858
rect -1111 -3891 -1109 -3823
rect -1095 -3891 -1093 -3823
rect -1087 -3891 -1085 -3823
rect -1077 -3891 -1075 -3823
rect -1069 -3891 -1067 -3823
rect -1053 -3891 -1051 -3823
rect -1045 -3891 -1043 -3823
rect -929 -3891 -927 -3823
rect -919 -3891 -917 -3823
rect -903 -3891 -901 -3823
rect -895 -3891 -893 -3823
rect -879 -3891 -877 -3823
rect -871 -3891 -869 -3823
rect -861 -3891 -859 -3823
rect -853 -3891 -851 -3823
rect -837 -3891 -835 -3823
rect -829 -3856 -827 -3823
rect -819 -3856 -817 -3823
rect -829 -3858 -817 -3856
rect -829 -3891 -827 -3858
rect -819 -3891 -817 -3858
rect -811 -3891 -809 -3823
rect -795 -3891 -793 -3823
rect -787 -3891 -785 -3823
rect -777 -3891 -775 -3823
rect -769 -3891 -767 -3823
rect -753 -3891 -751 -3823
rect -745 -3891 -743 -3823
rect -572 -3891 -570 -3823
rect -562 -3891 -560 -3823
rect -546 -3891 -544 -3823
rect -538 -3891 -536 -3823
rect -522 -3891 -520 -3823
rect -514 -3891 -512 -3823
rect -504 -3891 -502 -3823
rect -496 -3891 -494 -3823
rect -480 -3891 -478 -3823
rect -472 -3856 -470 -3823
rect -462 -3856 -460 -3823
rect -472 -3858 -460 -3856
rect -472 -3891 -470 -3858
rect -462 -3891 -460 -3858
rect -454 -3891 -452 -3823
rect -438 -3891 -436 -3823
rect -430 -3891 -428 -3823
rect -420 -3891 -418 -3823
rect -412 -3891 -410 -3823
rect -396 -3891 -394 -3823
rect -388 -3891 -386 -3823
rect -214 -3891 -212 -3823
rect -204 -3891 -202 -3823
rect -188 -3891 -186 -3823
rect -180 -3891 -178 -3823
rect -164 -3891 -162 -3823
rect -156 -3891 -154 -3823
rect -146 -3891 -144 -3823
rect -138 -3891 -136 -3823
rect -122 -3891 -120 -3823
rect -114 -3856 -112 -3823
rect -104 -3856 -102 -3823
rect -114 -3858 -102 -3856
rect -114 -3891 -112 -3858
rect -104 -3891 -102 -3858
rect -96 -3891 -94 -3823
rect -80 -3891 -78 -3823
rect -72 -3891 -70 -3823
rect -62 -3891 -60 -3823
rect -54 -3891 -52 -3823
rect -38 -3891 -36 -3823
rect -30 -3891 -28 -3823
rect 144 -3891 146 -3823
rect 154 -3891 156 -3823
rect 170 -3891 172 -3823
rect 178 -3891 180 -3823
rect 194 -3891 196 -3823
rect 202 -3891 204 -3823
rect 212 -3891 214 -3823
rect 220 -3891 222 -3823
rect 236 -3891 238 -3823
rect 244 -3856 246 -3823
rect 254 -3856 256 -3823
rect 244 -3858 256 -3856
rect 244 -3891 246 -3858
rect 254 -3891 256 -3858
rect 262 -3891 264 -3823
rect 278 -3891 280 -3823
rect 286 -3891 288 -3823
rect 296 -3891 298 -3823
rect 304 -3891 306 -3823
rect 320 -3891 322 -3823
rect 328 -3891 330 -3823
rect 500 -3891 502 -3823
rect 510 -3891 512 -3823
rect 526 -3891 528 -3823
rect 534 -3891 536 -3823
rect 550 -3891 552 -3823
rect 558 -3891 560 -3823
rect 568 -3891 570 -3823
rect 576 -3891 578 -3823
rect 592 -3891 594 -3823
rect 600 -3856 602 -3823
rect 610 -3856 612 -3823
rect 600 -3858 612 -3856
rect 600 -3891 602 -3858
rect 610 -3891 612 -3858
rect 618 -3891 620 -3823
rect 634 -3891 636 -3823
rect 642 -3891 644 -3823
rect 652 -3891 654 -3823
rect 660 -3891 662 -3823
rect 676 -3891 678 -3823
rect 684 -3891 686 -3823
rect 858 -3891 860 -3823
rect 868 -3891 870 -3823
rect 884 -3891 886 -3823
rect 892 -3891 894 -3823
rect 908 -3891 910 -3823
rect 916 -3891 918 -3823
rect 926 -3891 928 -3823
rect 934 -3891 936 -3823
rect 950 -3891 952 -3823
rect 958 -3856 960 -3823
rect 968 -3856 970 -3823
rect 958 -3858 970 -3856
rect 958 -3891 960 -3858
rect 968 -3891 970 -3858
rect 976 -3891 978 -3823
rect 992 -3891 994 -3823
rect 1000 -3891 1002 -3823
rect 1010 -3891 1012 -3823
rect 1018 -3891 1020 -3823
rect 1034 -3891 1036 -3823
rect 1042 -3891 1044 -3823
rect 1216 -3891 1218 -3823
rect 1226 -3891 1228 -3823
rect 1242 -3891 1244 -3823
rect 1250 -3891 1252 -3823
rect 1266 -3891 1268 -3823
rect 1274 -3891 1276 -3823
rect 1284 -3891 1286 -3823
rect 1292 -3891 1294 -3823
rect 1308 -3891 1310 -3823
rect 1316 -3856 1318 -3823
rect 1326 -3856 1328 -3823
rect 1316 -3858 1328 -3856
rect 1316 -3891 1318 -3858
rect 1326 -3891 1328 -3858
rect 1334 -3891 1336 -3823
rect 1350 -3891 1352 -3823
rect 1358 -3891 1360 -3823
rect 1368 -3891 1370 -3823
rect 1376 -3891 1378 -3823
rect 1392 -3891 1394 -3823
rect 1400 -3891 1402 -3823
rect -1554 -3897 -1552 -3895
rect -1544 -3897 -1542 -3895
rect -1528 -3897 -1526 -3895
rect -1520 -3897 -1518 -3895
rect -1504 -3897 -1502 -3895
rect -1496 -3897 -1494 -3895
rect -1486 -3897 -1484 -3895
rect -1478 -3897 -1476 -3895
rect -1462 -3897 -1460 -3895
rect -1454 -3897 -1452 -3895
rect -1444 -3897 -1442 -3895
rect -1436 -3897 -1434 -3895
rect -1420 -3897 -1418 -3895
rect -1412 -3897 -1410 -3895
rect -1402 -3897 -1400 -3895
rect -1394 -3897 -1392 -3895
rect -1378 -3897 -1376 -3895
rect -1370 -3897 -1368 -3895
rect -1229 -3897 -1227 -3895
rect -1219 -3897 -1217 -3895
rect -1203 -3897 -1201 -3895
rect -1195 -3897 -1193 -3895
rect -1179 -3897 -1177 -3895
rect -1171 -3897 -1169 -3895
rect -1161 -3897 -1159 -3895
rect -1153 -3897 -1151 -3895
rect -1137 -3897 -1135 -3895
rect -1129 -3897 -1127 -3895
rect -1119 -3897 -1117 -3895
rect -1111 -3897 -1109 -3895
rect -1095 -3897 -1093 -3895
rect -1087 -3897 -1085 -3895
rect -1077 -3897 -1075 -3895
rect -1069 -3897 -1067 -3895
rect -1053 -3897 -1051 -3895
rect -1045 -3897 -1043 -3895
rect -929 -3897 -927 -3895
rect -919 -3897 -917 -3895
rect -903 -3897 -901 -3895
rect -895 -3897 -893 -3895
rect -879 -3897 -877 -3895
rect -871 -3897 -869 -3895
rect -861 -3897 -859 -3895
rect -853 -3897 -851 -3895
rect -837 -3897 -835 -3895
rect -829 -3897 -827 -3895
rect -819 -3897 -817 -3895
rect -811 -3897 -809 -3895
rect -795 -3897 -793 -3895
rect -787 -3897 -785 -3895
rect -777 -3897 -775 -3895
rect -769 -3897 -767 -3895
rect -753 -3897 -751 -3895
rect -745 -3897 -743 -3895
rect -572 -3897 -570 -3895
rect -562 -3897 -560 -3895
rect -546 -3897 -544 -3895
rect -538 -3897 -536 -3895
rect -522 -3897 -520 -3895
rect -514 -3897 -512 -3895
rect -504 -3897 -502 -3895
rect -496 -3897 -494 -3895
rect -480 -3897 -478 -3895
rect -472 -3897 -470 -3895
rect -462 -3897 -460 -3895
rect -454 -3897 -452 -3895
rect -438 -3897 -436 -3895
rect -430 -3897 -428 -3895
rect -420 -3897 -418 -3895
rect -412 -3897 -410 -3895
rect -396 -3897 -394 -3895
rect -388 -3897 -386 -3895
rect -214 -3897 -212 -3895
rect -204 -3897 -202 -3895
rect -188 -3897 -186 -3895
rect -180 -3897 -178 -3895
rect -164 -3897 -162 -3895
rect -156 -3897 -154 -3895
rect -146 -3897 -144 -3895
rect -138 -3897 -136 -3895
rect -122 -3897 -120 -3895
rect -114 -3897 -112 -3895
rect -104 -3897 -102 -3895
rect -96 -3897 -94 -3895
rect -80 -3897 -78 -3895
rect -72 -3897 -70 -3895
rect -62 -3897 -60 -3895
rect -54 -3897 -52 -3895
rect -38 -3897 -36 -3895
rect -30 -3897 -28 -3895
rect 144 -3897 146 -3895
rect 154 -3897 156 -3895
rect 170 -3897 172 -3895
rect 178 -3897 180 -3895
rect 194 -3897 196 -3895
rect 202 -3897 204 -3895
rect 212 -3897 214 -3895
rect 220 -3897 222 -3895
rect 236 -3897 238 -3895
rect 244 -3897 246 -3895
rect 254 -3897 256 -3895
rect 262 -3897 264 -3895
rect 278 -3897 280 -3895
rect 286 -3897 288 -3895
rect 296 -3897 298 -3895
rect 304 -3897 306 -3895
rect 320 -3897 322 -3895
rect 328 -3897 330 -3895
rect 500 -3897 502 -3895
rect 510 -3897 512 -3895
rect 526 -3897 528 -3895
rect 534 -3897 536 -3895
rect 550 -3897 552 -3895
rect 558 -3897 560 -3895
rect 568 -3897 570 -3895
rect 576 -3897 578 -3895
rect 592 -3897 594 -3895
rect 600 -3897 602 -3895
rect 610 -3897 612 -3895
rect 618 -3897 620 -3895
rect 634 -3897 636 -3895
rect 642 -3897 644 -3895
rect 652 -3897 654 -3895
rect 660 -3897 662 -3895
rect 676 -3897 678 -3895
rect 684 -3897 686 -3895
rect 858 -3897 860 -3895
rect 868 -3897 870 -3895
rect 884 -3897 886 -3895
rect 892 -3897 894 -3895
rect 908 -3897 910 -3895
rect 916 -3897 918 -3895
rect 926 -3897 928 -3895
rect 934 -3897 936 -3895
rect 950 -3897 952 -3895
rect 958 -3897 960 -3895
rect 968 -3897 970 -3895
rect 976 -3897 978 -3895
rect 992 -3897 994 -3895
rect 1000 -3897 1002 -3895
rect 1010 -3897 1012 -3895
rect 1018 -3897 1020 -3895
rect 1034 -3897 1036 -3895
rect 1042 -3897 1044 -3895
rect 1216 -3897 1218 -3895
rect 1226 -3897 1228 -3895
rect 1242 -3897 1244 -3895
rect 1250 -3897 1252 -3895
rect 1266 -3897 1268 -3895
rect 1274 -3897 1276 -3895
rect 1284 -3897 1286 -3895
rect 1292 -3897 1294 -3895
rect 1308 -3897 1310 -3895
rect 1316 -3897 1318 -3895
rect 1326 -3897 1328 -3895
rect 1334 -3897 1336 -3895
rect 1350 -3897 1352 -3895
rect 1358 -3897 1360 -3895
rect 1368 -3897 1370 -3895
rect 1376 -3897 1378 -3895
rect 1392 -3897 1394 -3895
rect 1400 -3897 1402 -3895
rect -1554 -3990 -1552 -3988
rect -1544 -3990 -1542 -3988
rect -1528 -3990 -1526 -3988
rect -1520 -3990 -1518 -3988
rect -1504 -3990 -1502 -3988
rect -1496 -3990 -1494 -3988
rect -1486 -3990 -1484 -3988
rect -1478 -3990 -1476 -3988
rect -1462 -3990 -1460 -3988
rect -1454 -3990 -1452 -3988
rect -1444 -3990 -1442 -3988
rect -1436 -3990 -1434 -3988
rect -1420 -3990 -1418 -3988
rect -1412 -3990 -1410 -3988
rect -1402 -3990 -1400 -3988
rect -1394 -3990 -1392 -3988
rect -1378 -3990 -1376 -3988
rect -1370 -3990 -1368 -3988
rect -1229 -3990 -1227 -3988
rect -1219 -3990 -1217 -3988
rect -1203 -3990 -1201 -3988
rect -1195 -3990 -1193 -3988
rect -1179 -3990 -1177 -3988
rect -1171 -3990 -1169 -3988
rect -1161 -3990 -1159 -3988
rect -1153 -3990 -1151 -3988
rect -1137 -3990 -1135 -3988
rect -1129 -3990 -1127 -3988
rect -1119 -3990 -1117 -3988
rect -1111 -3990 -1109 -3988
rect -1095 -3990 -1093 -3988
rect -1087 -3990 -1085 -3988
rect -1077 -3990 -1075 -3988
rect -1069 -3990 -1067 -3988
rect -1053 -3990 -1051 -3988
rect -1045 -3990 -1043 -3988
rect -930 -3990 -928 -3988
rect -920 -3990 -918 -3988
rect -904 -3990 -902 -3988
rect -896 -3990 -894 -3988
rect -880 -3990 -878 -3988
rect -872 -3990 -870 -3988
rect -862 -3990 -860 -3988
rect -854 -3990 -852 -3988
rect -838 -3990 -836 -3988
rect -830 -3990 -828 -3988
rect -820 -3990 -818 -3988
rect -812 -3990 -810 -3988
rect -796 -3990 -794 -3988
rect -788 -3990 -786 -3988
rect -778 -3990 -776 -3988
rect -770 -3990 -768 -3988
rect -754 -3990 -752 -3988
rect -746 -3990 -744 -3988
rect -572 -3990 -570 -3988
rect -562 -3990 -560 -3988
rect -546 -3990 -544 -3988
rect -538 -3990 -536 -3988
rect -522 -3990 -520 -3988
rect -514 -3990 -512 -3988
rect -504 -3990 -502 -3988
rect -496 -3990 -494 -3988
rect -480 -3990 -478 -3988
rect -472 -3990 -470 -3988
rect -462 -3990 -460 -3988
rect -454 -3990 -452 -3988
rect -438 -3990 -436 -3988
rect -430 -3990 -428 -3988
rect -420 -3990 -418 -3988
rect -412 -3990 -410 -3988
rect -396 -3990 -394 -3988
rect -388 -3990 -386 -3988
rect -214 -3990 -212 -3988
rect -204 -3990 -202 -3988
rect -188 -3990 -186 -3988
rect -180 -3990 -178 -3988
rect -164 -3990 -162 -3988
rect -156 -3990 -154 -3988
rect -146 -3990 -144 -3988
rect -138 -3990 -136 -3988
rect -122 -3990 -120 -3988
rect -114 -3990 -112 -3988
rect -104 -3990 -102 -3988
rect -96 -3990 -94 -3988
rect -80 -3990 -78 -3988
rect -72 -3990 -70 -3988
rect -62 -3990 -60 -3988
rect -54 -3990 -52 -3988
rect -38 -3990 -36 -3988
rect -30 -3990 -28 -3988
rect 144 -3990 146 -3988
rect 154 -3990 156 -3988
rect 170 -3990 172 -3988
rect 178 -3990 180 -3988
rect 194 -3990 196 -3988
rect 202 -3990 204 -3988
rect 212 -3990 214 -3988
rect 220 -3990 222 -3988
rect 236 -3990 238 -3988
rect 244 -3990 246 -3988
rect 254 -3990 256 -3988
rect 262 -3990 264 -3988
rect 278 -3990 280 -3988
rect 286 -3990 288 -3988
rect 296 -3990 298 -3988
rect 304 -3990 306 -3988
rect 320 -3990 322 -3988
rect 328 -3990 330 -3988
rect 500 -3990 502 -3988
rect 510 -3990 512 -3988
rect 526 -3990 528 -3988
rect 534 -3990 536 -3988
rect 550 -3990 552 -3988
rect 558 -3990 560 -3988
rect 568 -3990 570 -3988
rect 576 -3990 578 -3988
rect 592 -3990 594 -3988
rect 600 -3990 602 -3988
rect 610 -3990 612 -3988
rect 618 -3990 620 -3988
rect 634 -3990 636 -3988
rect 642 -3990 644 -3988
rect 652 -3990 654 -3988
rect 660 -3990 662 -3988
rect 676 -3990 678 -3988
rect 684 -3990 686 -3988
rect 858 -3990 860 -3988
rect 868 -3990 870 -3988
rect 884 -3990 886 -3988
rect 892 -3990 894 -3988
rect 908 -3990 910 -3988
rect 916 -3990 918 -3988
rect 926 -3990 928 -3988
rect 934 -3990 936 -3988
rect 950 -3990 952 -3988
rect 958 -3990 960 -3988
rect 968 -3990 970 -3988
rect 976 -3990 978 -3988
rect 992 -3990 994 -3988
rect 1000 -3990 1002 -3988
rect 1010 -3990 1012 -3988
rect 1018 -3990 1020 -3988
rect 1034 -3990 1036 -3988
rect 1042 -3990 1044 -3988
rect 1216 -3990 1218 -3988
rect 1226 -3990 1228 -3988
rect 1242 -3990 1244 -3988
rect 1250 -3990 1252 -3988
rect 1266 -3990 1268 -3988
rect 1274 -3990 1276 -3988
rect 1284 -3990 1286 -3988
rect 1292 -3990 1294 -3988
rect 1308 -3990 1310 -3988
rect 1316 -3990 1318 -3988
rect 1326 -3990 1328 -3988
rect 1334 -3990 1336 -3988
rect 1350 -3990 1352 -3988
rect 1358 -3990 1360 -3988
rect 1368 -3990 1370 -3988
rect 1376 -3990 1378 -3988
rect 1392 -3990 1394 -3988
rect 1400 -3990 1402 -3988
rect -1554 -4066 -1552 -3998
rect -1544 -4066 -1542 -3998
rect -1528 -4066 -1526 -3998
rect -1520 -4066 -1518 -3998
rect -1504 -4066 -1502 -3998
rect -1496 -4066 -1494 -3998
rect -1486 -4066 -1484 -3998
rect -1478 -4066 -1476 -3998
rect -1462 -4066 -1460 -3998
rect -1454 -4031 -1452 -3998
rect -1444 -4031 -1442 -3998
rect -1454 -4033 -1442 -4031
rect -1454 -4066 -1452 -4033
rect -1444 -4066 -1442 -4033
rect -1436 -4066 -1434 -3998
rect -1420 -4066 -1418 -3998
rect -1412 -4066 -1410 -3998
rect -1402 -4066 -1400 -3998
rect -1394 -4066 -1392 -3998
rect -1378 -4066 -1376 -3998
rect -1370 -4066 -1368 -3998
rect -1229 -4066 -1227 -3998
rect -1219 -4066 -1217 -3998
rect -1203 -4066 -1201 -3998
rect -1195 -4066 -1193 -3998
rect -1179 -4066 -1177 -3998
rect -1171 -4066 -1169 -3998
rect -1161 -4066 -1159 -3998
rect -1153 -4066 -1151 -3998
rect -1137 -4066 -1135 -3998
rect -1129 -4031 -1127 -3998
rect -1119 -4031 -1117 -3998
rect -1129 -4033 -1117 -4031
rect -1129 -4066 -1127 -4033
rect -1119 -4066 -1117 -4033
rect -1111 -4066 -1109 -3998
rect -1095 -4066 -1093 -3998
rect -1087 -4066 -1085 -3998
rect -1077 -4066 -1075 -3998
rect -1069 -4066 -1067 -3998
rect -1053 -4066 -1051 -3998
rect -1045 -4066 -1043 -3998
rect -930 -4066 -928 -3998
rect -920 -4066 -918 -3998
rect -904 -4066 -902 -3998
rect -896 -4066 -894 -3998
rect -880 -4066 -878 -3998
rect -872 -4066 -870 -3998
rect -862 -4066 -860 -3998
rect -854 -4066 -852 -3998
rect -838 -4066 -836 -3998
rect -830 -4031 -828 -3998
rect -820 -4031 -818 -3998
rect -830 -4033 -818 -4031
rect -830 -4066 -828 -4033
rect -820 -4066 -818 -4033
rect -812 -4066 -810 -3998
rect -796 -4066 -794 -3998
rect -788 -4066 -786 -3998
rect -778 -4066 -776 -3998
rect -770 -4066 -768 -3998
rect -754 -4066 -752 -3998
rect -746 -4066 -744 -3998
rect -572 -4066 -570 -3998
rect -562 -4066 -560 -3998
rect -546 -4066 -544 -3998
rect -538 -4066 -536 -3998
rect -522 -4066 -520 -3998
rect -514 -4066 -512 -3998
rect -504 -4066 -502 -3998
rect -496 -4066 -494 -3998
rect -480 -4066 -478 -3998
rect -472 -4031 -470 -3998
rect -462 -4031 -460 -3998
rect -472 -4033 -460 -4031
rect -472 -4066 -470 -4033
rect -462 -4066 -460 -4033
rect -454 -4066 -452 -3998
rect -438 -4066 -436 -3998
rect -430 -4066 -428 -3998
rect -420 -4066 -418 -3998
rect -412 -4066 -410 -3998
rect -396 -4066 -394 -3998
rect -388 -4066 -386 -3998
rect -214 -4066 -212 -3998
rect -204 -4066 -202 -3998
rect -188 -4066 -186 -3998
rect -180 -4066 -178 -3998
rect -164 -4066 -162 -3998
rect -156 -4066 -154 -3998
rect -146 -4066 -144 -3998
rect -138 -4066 -136 -3998
rect -122 -4066 -120 -3998
rect -114 -4031 -112 -3998
rect -104 -4031 -102 -3998
rect -114 -4033 -102 -4031
rect -114 -4066 -112 -4033
rect -104 -4066 -102 -4033
rect -96 -4066 -94 -3998
rect -80 -4066 -78 -3998
rect -72 -4066 -70 -3998
rect -62 -4066 -60 -3998
rect -54 -4066 -52 -3998
rect -38 -4066 -36 -3998
rect -30 -4066 -28 -3998
rect 144 -4066 146 -3998
rect 154 -4066 156 -3998
rect 170 -4066 172 -3998
rect 178 -4066 180 -3998
rect 194 -4066 196 -3998
rect 202 -4066 204 -3998
rect 212 -4066 214 -3998
rect 220 -4066 222 -3998
rect 236 -4066 238 -3998
rect 244 -4031 246 -3998
rect 254 -4031 256 -3998
rect 244 -4033 256 -4031
rect 244 -4066 246 -4033
rect 254 -4066 256 -4033
rect 262 -4066 264 -3998
rect 278 -4066 280 -3998
rect 286 -4066 288 -3998
rect 296 -4066 298 -3998
rect 304 -4066 306 -3998
rect 320 -4066 322 -3998
rect 328 -4066 330 -3998
rect 500 -4066 502 -3998
rect 510 -4066 512 -3998
rect 526 -4066 528 -3998
rect 534 -4066 536 -3998
rect 550 -4066 552 -3998
rect 558 -4066 560 -3998
rect 568 -4066 570 -3998
rect 576 -4066 578 -3998
rect 592 -4066 594 -3998
rect 600 -4031 602 -3998
rect 610 -4031 612 -3998
rect 600 -4033 612 -4031
rect 600 -4066 602 -4033
rect 610 -4066 612 -4033
rect 618 -4066 620 -3998
rect 634 -4066 636 -3998
rect 642 -4066 644 -3998
rect 652 -4066 654 -3998
rect 660 -4066 662 -3998
rect 676 -4066 678 -3998
rect 684 -4066 686 -3998
rect 858 -4066 860 -3998
rect 868 -4066 870 -3998
rect 884 -4066 886 -3998
rect 892 -4066 894 -3998
rect 908 -4066 910 -3998
rect 916 -4066 918 -3998
rect 926 -4066 928 -3998
rect 934 -4066 936 -3998
rect 950 -4066 952 -3998
rect 958 -4031 960 -3998
rect 968 -4031 970 -3998
rect 958 -4033 970 -4031
rect 958 -4066 960 -4033
rect 968 -4066 970 -4033
rect 976 -4066 978 -3998
rect 992 -4066 994 -3998
rect 1000 -4066 1002 -3998
rect 1010 -4066 1012 -3998
rect 1018 -4066 1020 -3998
rect 1034 -4066 1036 -3998
rect 1042 -4066 1044 -3998
rect 1216 -4066 1218 -3998
rect 1226 -4066 1228 -3998
rect 1242 -4066 1244 -3998
rect 1250 -4066 1252 -3998
rect 1266 -4066 1268 -3998
rect 1274 -4066 1276 -3998
rect 1284 -4066 1286 -3998
rect 1292 -4066 1294 -3998
rect 1308 -4066 1310 -3998
rect 1316 -4031 1318 -3998
rect 1326 -4031 1328 -3998
rect 1316 -4033 1328 -4031
rect 1316 -4066 1318 -4033
rect 1326 -4066 1328 -4033
rect 1334 -4066 1336 -3998
rect 1350 -4066 1352 -3998
rect 1358 -4066 1360 -3998
rect 1368 -4066 1370 -3998
rect 1376 -4066 1378 -3998
rect 1392 -4066 1394 -3998
rect 1400 -4066 1402 -3998
rect -1554 -4072 -1552 -4070
rect -1544 -4072 -1542 -4070
rect -1528 -4072 -1526 -4070
rect -1520 -4072 -1518 -4070
rect -1504 -4072 -1502 -4070
rect -1496 -4072 -1494 -4070
rect -1486 -4072 -1484 -4070
rect -1478 -4072 -1476 -4070
rect -1462 -4072 -1460 -4070
rect -1454 -4072 -1452 -4070
rect -1444 -4072 -1442 -4070
rect -1436 -4072 -1434 -4070
rect -1420 -4072 -1418 -4070
rect -1412 -4072 -1410 -4070
rect -1402 -4072 -1400 -4070
rect -1394 -4072 -1392 -4070
rect -1378 -4072 -1376 -4070
rect -1370 -4072 -1368 -4070
rect -1229 -4072 -1227 -4070
rect -1219 -4072 -1217 -4070
rect -1203 -4072 -1201 -4070
rect -1195 -4072 -1193 -4070
rect -1179 -4072 -1177 -4070
rect -1171 -4072 -1169 -4070
rect -1161 -4072 -1159 -4070
rect -1153 -4072 -1151 -4070
rect -1137 -4072 -1135 -4070
rect -1129 -4072 -1127 -4070
rect -1119 -4072 -1117 -4070
rect -1111 -4072 -1109 -4070
rect -1095 -4072 -1093 -4070
rect -1087 -4072 -1085 -4070
rect -1077 -4072 -1075 -4070
rect -1069 -4072 -1067 -4070
rect -1053 -4072 -1051 -4070
rect -1045 -4072 -1043 -4070
rect -930 -4072 -928 -4070
rect -920 -4072 -918 -4070
rect -904 -4072 -902 -4070
rect -896 -4072 -894 -4070
rect -880 -4072 -878 -4070
rect -872 -4072 -870 -4070
rect -862 -4072 -860 -4070
rect -854 -4072 -852 -4070
rect -838 -4072 -836 -4070
rect -830 -4072 -828 -4070
rect -820 -4072 -818 -4070
rect -812 -4072 -810 -4070
rect -796 -4072 -794 -4070
rect -788 -4072 -786 -4070
rect -778 -4072 -776 -4070
rect -770 -4072 -768 -4070
rect -754 -4072 -752 -4070
rect -746 -4072 -744 -4070
rect -572 -4072 -570 -4070
rect -562 -4072 -560 -4070
rect -546 -4072 -544 -4070
rect -538 -4072 -536 -4070
rect -522 -4072 -520 -4070
rect -514 -4072 -512 -4070
rect -504 -4072 -502 -4070
rect -496 -4072 -494 -4070
rect -480 -4072 -478 -4070
rect -472 -4072 -470 -4070
rect -462 -4072 -460 -4070
rect -454 -4072 -452 -4070
rect -438 -4072 -436 -4070
rect -430 -4072 -428 -4070
rect -420 -4072 -418 -4070
rect -412 -4072 -410 -4070
rect -396 -4072 -394 -4070
rect -388 -4072 -386 -4070
rect -214 -4072 -212 -4070
rect -204 -4072 -202 -4070
rect -188 -4072 -186 -4070
rect -180 -4072 -178 -4070
rect -164 -4072 -162 -4070
rect -156 -4072 -154 -4070
rect -146 -4072 -144 -4070
rect -138 -4072 -136 -4070
rect -122 -4072 -120 -4070
rect -114 -4072 -112 -4070
rect -104 -4072 -102 -4070
rect -96 -4072 -94 -4070
rect -80 -4072 -78 -4070
rect -72 -4072 -70 -4070
rect -62 -4072 -60 -4070
rect -54 -4072 -52 -4070
rect -38 -4072 -36 -4070
rect -30 -4072 -28 -4070
rect 144 -4072 146 -4070
rect 154 -4072 156 -4070
rect 170 -4072 172 -4070
rect 178 -4072 180 -4070
rect 194 -4072 196 -4070
rect 202 -4072 204 -4070
rect 212 -4072 214 -4070
rect 220 -4072 222 -4070
rect 236 -4072 238 -4070
rect 244 -4072 246 -4070
rect 254 -4072 256 -4070
rect 262 -4072 264 -4070
rect 278 -4072 280 -4070
rect 286 -4072 288 -4070
rect 296 -4072 298 -4070
rect 304 -4072 306 -4070
rect 320 -4072 322 -4070
rect 328 -4072 330 -4070
rect 500 -4072 502 -4070
rect 510 -4072 512 -4070
rect 526 -4072 528 -4070
rect 534 -4072 536 -4070
rect 550 -4072 552 -4070
rect 558 -4072 560 -4070
rect 568 -4072 570 -4070
rect 576 -4072 578 -4070
rect 592 -4072 594 -4070
rect 600 -4072 602 -4070
rect 610 -4072 612 -4070
rect 618 -4072 620 -4070
rect 634 -4072 636 -4070
rect 642 -4072 644 -4070
rect 652 -4072 654 -4070
rect 660 -4072 662 -4070
rect 676 -4072 678 -4070
rect 684 -4072 686 -4070
rect 858 -4072 860 -4070
rect 868 -4072 870 -4070
rect 884 -4072 886 -4070
rect 892 -4072 894 -4070
rect 908 -4072 910 -4070
rect 916 -4072 918 -4070
rect 926 -4072 928 -4070
rect 934 -4072 936 -4070
rect 950 -4072 952 -4070
rect 958 -4072 960 -4070
rect 968 -4072 970 -4070
rect 976 -4072 978 -4070
rect 992 -4072 994 -4070
rect 1000 -4072 1002 -4070
rect 1010 -4072 1012 -4070
rect 1018 -4072 1020 -4070
rect 1034 -4072 1036 -4070
rect 1042 -4072 1044 -4070
rect 1216 -4072 1218 -4070
rect 1226 -4072 1228 -4070
rect 1242 -4072 1244 -4070
rect 1250 -4072 1252 -4070
rect 1266 -4072 1268 -4070
rect 1274 -4072 1276 -4070
rect 1284 -4072 1286 -4070
rect 1292 -4072 1294 -4070
rect 1308 -4072 1310 -4070
rect 1316 -4072 1318 -4070
rect 1326 -4072 1328 -4070
rect 1334 -4072 1336 -4070
rect 1350 -4072 1352 -4070
rect 1358 -4072 1360 -4070
rect 1368 -4072 1370 -4070
rect 1376 -4072 1378 -4070
rect 1392 -4072 1394 -4070
rect 1400 -4072 1402 -4070
rect -1304 -4105 -1302 -4103
rect -1296 -4105 -1294 -4103
rect -1286 -4105 -1284 -4103
rect -930 -4105 -928 -4103
rect -922 -4105 -920 -4103
rect -912 -4105 -910 -4103
rect -572 -4105 -570 -4103
rect -564 -4105 -562 -4103
rect -554 -4105 -552 -4103
rect -214 -4105 -212 -4103
rect -206 -4105 -204 -4103
rect -196 -4105 -194 -4103
rect 144 -4105 146 -4103
rect 152 -4105 154 -4103
rect 162 -4105 164 -4103
rect 500 -4105 502 -4103
rect 508 -4105 510 -4103
rect 518 -4105 520 -4103
rect 858 -4105 860 -4103
rect 866 -4105 868 -4103
rect 876 -4105 878 -4103
rect 1216 -4105 1218 -4103
rect 1224 -4105 1226 -4103
rect 1234 -4105 1236 -4103
rect -1304 -4181 -1302 -4113
rect -1296 -4137 -1294 -4113
rect -1296 -4181 -1294 -4141
rect -1286 -4181 -1284 -4113
rect -930 -4181 -928 -4113
rect -922 -4137 -920 -4113
rect -922 -4181 -920 -4141
rect -912 -4181 -910 -4113
rect -572 -4181 -570 -4113
rect -564 -4137 -562 -4113
rect -564 -4181 -562 -4141
rect -554 -4181 -552 -4113
rect -214 -4181 -212 -4113
rect -206 -4137 -204 -4113
rect -206 -4181 -204 -4141
rect -196 -4181 -194 -4113
rect 144 -4181 146 -4113
rect 152 -4137 154 -4113
rect 152 -4181 154 -4141
rect 162 -4181 164 -4113
rect 500 -4181 502 -4113
rect 508 -4137 510 -4113
rect 508 -4181 510 -4141
rect 518 -4181 520 -4113
rect 858 -4181 860 -4113
rect 866 -4137 868 -4113
rect 866 -4181 868 -4141
rect 876 -4181 878 -4113
rect 1216 -4181 1218 -4113
rect 1224 -4137 1226 -4113
rect 1224 -4181 1226 -4141
rect 1234 -4181 1236 -4113
rect -1304 -4187 -1302 -4185
rect -1296 -4187 -1294 -4185
rect -1286 -4187 -1284 -4185
rect -930 -4187 -928 -4185
rect -922 -4187 -920 -4185
rect -912 -4187 -910 -4185
rect -572 -4187 -570 -4185
rect -564 -4187 -562 -4185
rect -554 -4187 -552 -4185
rect -214 -4187 -212 -4185
rect -206 -4187 -204 -4185
rect -196 -4187 -194 -4185
rect 144 -4187 146 -4185
rect 152 -4187 154 -4185
rect 162 -4187 164 -4185
rect 500 -4187 502 -4185
rect 508 -4187 510 -4185
rect 518 -4187 520 -4185
rect 858 -4187 860 -4185
rect 866 -4187 868 -4185
rect 876 -4187 878 -4185
rect 1216 -4187 1218 -4185
rect 1224 -4187 1226 -4185
rect 1234 -4187 1236 -4185
rect -1229 -4264 -1227 -4262
rect -1219 -4264 -1217 -4262
rect -1203 -4264 -1201 -4262
rect -1193 -4264 -1191 -4262
rect -1185 -4264 -1183 -4262
rect -1175 -4264 -1173 -4262
rect -1159 -4264 -1157 -4262
rect -1151 -4264 -1149 -4262
rect -1141 -4264 -1139 -4262
rect -930 -4264 -928 -4262
rect -920 -4264 -918 -4262
rect -904 -4264 -902 -4262
rect -894 -4264 -892 -4262
rect -878 -4264 -876 -4262
rect -868 -4264 -866 -4262
rect -860 -4264 -858 -4262
rect -850 -4264 -848 -4262
rect -834 -4264 -832 -4262
rect -826 -4264 -824 -4262
rect -816 -4264 -814 -4262
rect -800 -4264 -798 -4262
rect -790 -4264 -788 -4262
rect -782 -4264 -780 -4262
rect -772 -4264 -770 -4262
rect -756 -4264 -754 -4262
rect -748 -4264 -746 -4262
rect -732 -4264 -730 -4262
rect -716 -4264 -714 -4262
rect -708 -4264 -706 -4262
rect -698 -4264 -696 -4262
rect -572 -4264 -570 -4262
rect -562 -4264 -560 -4262
rect -546 -4264 -544 -4262
rect -536 -4264 -534 -4262
rect -520 -4264 -518 -4262
rect -510 -4264 -508 -4262
rect -502 -4264 -500 -4262
rect -492 -4264 -490 -4262
rect -476 -4264 -474 -4262
rect -468 -4264 -466 -4262
rect -458 -4264 -456 -4262
rect -442 -4264 -440 -4262
rect -432 -4264 -430 -4262
rect -424 -4264 -422 -4262
rect -414 -4264 -412 -4262
rect -398 -4264 -396 -4262
rect -390 -4264 -388 -4262
rect -374 -4264 -372 -4262
rect -358 -4264 -356 -4262
rect -350 -4264 -348 -4262
rect -340 -4264 -338 -4262
rect -214 -4264 -212 -4262
rect -204 -4264 -202 -4262
rect -188 -4264 -186 -4262
rect -178 -4264 -176 -4262
rect -162 -4264 -160 -4262
rect -152 -4264 -150 -4262
rect -144 -4264 -142 -4262
rect -134 -4264 -132 -4262
rect -118 -4264 -116 -4262
rect -110 -4264 -108 -4262
rect -100 -4264 -98 -4262
rect -84 -4264 -82 -4262
rect -74 -4264 -72 -4262
rect -66 -4264 -64 -4262
rect -56 -4264 -54 -4262
rect -40 -4264 -38 -4262
rect -32 -4264 -30 -4262
rect -16 -4264 -14 -4262
rect 0 -4264 2 -4262
rect 8 -4264 10 -4262
rect 18 -4264 20 -4262
rect 144 -4264 146 -4262
rect 154 -4264 156 -4262
rect 170 -4264 172 -4262
rect 180 -4264 182 -4262
rect 196 -4264 198 -4262
rect 206 -4264 208 -4262
rect 214 -4264 216 -4262
rect 224 -4264 226 -4262
rect 240 -4264 242 -4262
rect 248 -4264 250 -4262
rect 258 -4264 260 -4262
rect 274 -4264 276 -4262
rect 284 -4264 286 -4262
rect 292 -4264 294 -4262
rect 302 -4264 304 -4262
rect 318 -4264 320 -4262
rect 326 -4264 328 -4262
rect 342 -4264 344 -4262
rect 358 -4264 360 -4262
rect 366 -4264 368 -4262
rect 376 -4264 378 -4262
rect 500 -4264 502 -4262
rect 510 -4264 512 -4262
rect 526 -4264 528 -4262
rect 536 -4264 538 -4262
rect 552 -4264 554 -4262
rect 562 -4264 564 -4262
rect 570 -4264 572 -4262
rect 580 -4264 582 -4262
rect 596 -4264 598 -4262
rect 604 -4264 606 -4262
rect 614 -4264 616 -4262
rect 630 -4264 632 -4262
rect 640 -4264 642 -4262
rect 648 -4264 650 -4262
rect 658 -4264 660 -4262
rect 674 -4264 676 -4262
rect 682 -4264 684 -4262
rect 698 -4264 700 -4262
rect 714 -4264 716 -4262
rect 722 -4264 724 -4262
rect 732 -4264 734 -4262
rect 858 -4264 860 -4262
rect 868 -4264 870 -4262
rect 884 -4264 886 -4262
rect 894 -4264 896 -4262
rect 910 -4264 912 -4262
rect 920 -4264 922 -4262
rect 928 -4264 930 -4262
rect 938 -4264 940 -4262
rect 954 -4264 956 -4262
rect 962 -4264 964 -4262
rect 972 -4264 974 -4262
rect 988 -4264 990 -4262
rect 998 -4264 1000 -4262
rect 1006 -4264 1008 -4262
rect 1016 -4264 1018 -4262
rect 1032 -4264 1034 -4262
rect 1040 -4264 1042 -4262
rect 1056 -4264 1058 -4262
rect 1072 -4264 1074 -4262
rect 1080 -4264 1082 -4262
rect 1090 -4264 1092 -4262
rect 1216 -4264 1218 -4262
rect 1226 -4264 1228 -4262
rect 1242 -4264 1244 -4262
rect 1252 -4264 1254 -4262
rect 1268 -4264 1270 -4262
rect 1278 -4264 1280 -4262
rect 1286 -4264 1288 -4262
rect 1296 -4264 1298 -4262
rect 1312 -4264 1314 -4262
rect 1320 -4264 1322 -4262
rect 1330 -4264 1332 -4262
rect 1346 -4264 1348 -4262
rect 1356 -4264 1358 -4262
rect 1364 -4264 1366 -4262
rect 1374 -4264 1376 -4262
rect 1390 -4264 1392 -4262
rect 1398 -4264 1400 -4262
rect 1414 -4264 1416 -4262
rect 1430 -4264 1432 -4262
rect 1438 -4264 1440 -4262
rect 1448 -4264 1450 -4262
rect -1229 -4340 -1227 -4272
rect -1219 -4340 -1217 -4272
rect -1203 -4340 -1201 -4272
rect -1193 -4340 -1191 -4272
rect -1185 -4340 -1183 -4272
rect -1175 -4340 -1173 -4272
rect -1159 -4340 -1157 -4272
rect -1151 -4340 -1149 -4272
rect -1141 -4340 -1139 -4272
rect -930 -4340 -928 -4272
rect -920 -4340 -918 -4272
rect -904 -4340 -902 -4272
rect -894 -4340 -892 -4272
rect -878 -4340 -876 -4272
rect -868 -4340 -866 -4272
rect -860 -4340 -858 -4272
rect -850 -4340 -848 -4272
rect -834 -4340 -832 -4272
rect -826 -4340 -824 -4272
rect -816 -4340 -814 -4272
rect -800 -4340 -798 -4272
rect -790 -4340 -788 -4272
rect -782 -4340 -780 -4272
rect -772 -4340 -770 -4272
rect -756 -4340 -754 -4272
rect -748 -4340 -746 -4272
rect -732 -4340 -730 -4272
rect -716 -4340 -714 -4272
rect -708 -4340 -706 -4272
rect -698 -4340 -696 -4272
rect -572 -4340 -570 -4272
rect -562 -4340 -560 -4272
rect -546 -4340 -544 -4272
rect -536 -4340 -534 -4272
rect -520 -4340 -518 -4272
rect -510 -4340 -508 -4272
rect -502 -4340 -500 -4272
rect -492 -4340 -490 -4272
rect -476 -4340 -474 -4272
rect -468 -4340 -466 -4272
rect -458 -4340 -456 -4272
rect -442 -4340 -440 -4272
rect -432 -4340 -430 -4272
rect -424 -4340 -422 -4272
rect -414 -4340 -412 -4272
rect -398 -4340 -396 -4272
rect -390 -4340 -388 -4272
rect -374 -4340 -372 -4272
rect -358 -4340 -356 -4272
rect -350 -4340 -348 -4272
rect -340 -4340 -338 -4272
rect -214 -4340 -212 -4272
rect -204 -4340 -202 -4272
rect -188 -4340 -186 -4272
rect -178 -4340 -176 -4272
rect -162 -4340 -160 -4272
rect -152 -4340 -150 -4272
rect -144 -4340 -142 -4272
rect -134 -4340 -132 -4272
rect -118 -4340 -116 -4272
rect -110 -4340 -108 -4272
rect -100 -4340 -98 -4272
rect -84 -4340 -82 -4272
rect -74 -4340 -72 -4272
rect -66 -4340 -64 -4272
rect -56 -4340 -54 -4272
rect -40 -4340 -38 -4272
rect -32 -4340 -30 -4272
rect -16 -4340 -14 -4272
rect 0 -4340 2 -4272
rect 8 -4340 10 -4272
rect 18 -4340 20 -4272
rect 144 -4340 146 -4272
rect 154 -4340 156 -4272
rect 170 -4340 172 -4272
rect 180 -4340 182 -4272
rect 196 -4340 198 -4272
rect 206 -4340 208 -4272
rect 214 -4340 216 -4272
rect 224 -4340 226 -4272
rect 240 -4340 242 -4272
rect 248 -4340 250 -4272
rect 258 -4340 260 -4272
rect 274 -4340 276 -4272
rect 284 -4340 286 -4272
rect 292 -4340 294 -4272
rect 302 -4340 304 -4272
rect 318 -4340 320 -4272
rect 326 -4340 328 -4272
rect 342 -4340 344 -4272
rect 358 -4340 360 -4272
rect 366 -4340 368 -4272
rect 376 -4340 378 -4272
rect 500 -4340 502 -4272
rect 510 -4340 512 -4272
rect 526 -4340 528 -4272
rect 536 -4340 538 -4272
rect 552 -4340 554 -4272
rect 562 -4340 564 -4272
rect 570 -4340 572 -4272
rect 580 -4340 582 -4272
rect 596 -4340 598 -4272
rect 604 -4340 606 -4272
rect 614 -4340 616 -4272
rect 630 -4340 632 -4272
rect 640 -4340 642 -4272
rect 648 -4340 650 -4272
rect 658 -4340 660 -4272
rect 674 -4340 676 -4272
rect 682 -4340 684 -4272
rect 698 -4340 700 -4272
rect 714 -4340 716 -4272
rect 722 -4340 724 -4272
rect 732 -4340 734 -4272
rect 858 -4340 860 -4272
rect 868 -4340 870 -4272
rect 884 -4340 886 -4272
rect 894 -4340 896 -4272
rect 910 -4340 912 -4272
rect 920 -4340 922 -4272
rect 928 -4340 930 -4272
rect 938 -4340 940 -4272
rect 954 -4340 956 -4272
rect 962 -4340 964 -4272
rect 972 -4340 974 -4272
rect 988 -4340 990 -4272
rect 998 -4340 1000 -4272
rect 1006 -4340 1008 -4272
rect 1016 -4340 1018 -4272
rect 1032 -4340 1034 -4272
rect 1040 -4340 1042 -4272
rect 1056 -4340 1058 -4272
rect 1072 -4340 1074 -4272
rect 1080 -4340 1082 -4272
rect 1090 -4340 1092 -4272
rect 1216 -4340 1218 -4272
rect 1226 -4340 1228 -4272
rect 1242 -4340 1244 -4272
rect 1252 -4340 1254 -4272
rect 1268 -4340 1270 -4272
rect 1278 -4340 1280 -4272
rect 1286 -4340 1288 -4272
rect 1296 -4340 1298 -4272
rect 1312 -4340 1314 -4272
rect 1320 -4340 1322 -4272
rect 1330 -4340 1332 -4272
rect 1346 -4340 1348 -4272
rect 1356 -4340 1358 -4272
rect 1364 -4340 1366 -4272
rect 1374 -4340 1376 -4272
rect 1390 -4340 1392 -4272
rect 1398 -4340 1400 -4272
rect 1414 -4340 1416 -4272
rect 1430 -4340 1432 -4272
rect 1438 -4340 1440 -4272
rect 1448 -4340 1450 -4272
rect -1229 -4346 -1227 -4344
rect -1219 -4346 -1217 -4344
rect -1203 -4346 -1201 -4344
rect -1193 -4346 -1191 -4344
rect -1185 -4346 -1183 -4344
rect -1175 -4346 -1173 -4344
rect -1159 -4346 -1157 -4344
rect -1151 -4346 -1149 -4344
rect -1141 -4346 -1139 -4344
rect -930 -4346 -928 -4344
rect -920 -4346 -918 -4344
rect -904 -4346 -902 -4344
rect -894 -4346 -892 -4344
rect -878 -4346 -876 -4344
rect -868 -4346 -866 -4344
rect -860 -4346 -858 -4344
rect -850 -4346 -848 -4344
rect -834 -4346 -832 -4344
rect -826 -4346 -824 -4344
rect -816 -4346 -814 -4344
rect -800 -4346 -798 -4344
rect -790 -4346 -788 -4344
rect -782 -4346 -780 -4344
rect -772 -4346 -770 -4344
rect -756 -4346 -754 -4344
rect -748 -4346 -746 -4344
rect -732 -4346 -730 -4344
rect -716 -4346 -714 -4344
rect -708 -4346 -706 -4344
rect -698 -4346 -696 -4344
rect -572 -4346 -570 -4344
rect -562 -4346 -560 -4344
rect -546 -4346 -544 -4344
rect -536 -4346 -534 -4344
rect -520 -4346 -518 -4344
rect -510 -4346 -508 -4344
rect -502 -4346 -500 -4344
rect -492 -4346 -490 -4344
rect -476 -4346 -474 -4344
rect -468 -4346 -466 -4344
rect -458 -4346 -456 -4344
rect -442 -4346 -440 -4344
rect -432 -4346 -430 -4344
rect -424 -4346 -422 -4344
rect -414 -4346 -412 -4344
rect -398 -4346 -396 -4344
rect -390 -4346 -388 -4344
rect -374 -4346 -372 -4344
rect -358 -4346 -356 -4344
rect -350 -4346 -348 -4344
rect -340 -4346 -338 -4344
rect -214 -4346 -212 -4344
rect -204 -4346 -202 -4344
rect -188 -4346 -186 -4344
rect -178 -4346 -176 -4344
rect -162 -4346 -160 -4344
rect -152 -4346 -150 -4344
rect -144 -4346 -142 -4344
rect -134 -4346 -132 -4344
rect -118 -4346 -116 -4344
rect -110 -4346 -108 -4344
rect -100 -4346 -98 -4344
rect -84 -4346 -82 -4344
rect -74 -4346 -72 -4344
rect -66 -4346 -64 -4344
rect -56 -4346 -54 -4344
rect -40 -4346 -38 -4344
rect -32 -4346 -30 -4344
rect -16 -4346 -14 -4344
rect 0 -4346 2 -4344
rect 8 -4346 10 -4344
rect 18 -4346 20 -4344
rect 144 -4346 146 -4344
rect 154 -4346 156 -4344
rect 170 -4346 172 -4344
rect 180 -4346 182 -4344
rect 196 -4346 198 -4344
rect 206 -4346 208 -4344
rect 214 -4346 216 -4344
rect 224 -4346 226 -4344
rect 240 -4346 242 -4344
rect 248 -4346 250 -4344
rect 258 -4346 260 -4344
rect 274 -4346 276 -4344
rect 284 -4346 286 -4344
rect 292 -4346 294 -4344
rect 302 -4346 304 -4344
rect 318 -4346 320 -4344
rect 326 -4346 328 -4344
rect 342 -4346 344 -4344
rect 358 -4346 360 -4344
rect 366 -4346 368 -4344
rect 376 -4346 378 -4344
rect 500 -4346 502 -4344
rect 510 -4346 512 -4344
rect 526 -4346 528 -4344
rect 536 -4346 538 -4344
rect 552 -4346 554 -4344
rect 562 -4346 564 -4344
rect 570 -4346 572 -4344
rect 580 -4346 582 -4344
rect 596 -4346 598 -4344
rect 604 -4346 606 -4344
rect 614 -4346 616 -4344
rect 630 -4346 632 -4344
rect 640 -4346 642 -4344
rect 648 -4346 650 -4344
rect 658 -4346 660 -4344
rect 674 -4346 676 -4344
rect 682 -4346 684 -4344
rect 698 -4346 700 -4344
rect 714 -4346 716 -4344
rect 722 -4346 724 -4344
rect 732 -4346 734 -4344
rect 858 -4346 860 -4344
rect 868 -4346 870 -4344
rect 884 -4346 886 -4344
rect 894 -4346 896 -4344
rect 910 -4346 912 -4344
rect 920 -4346 922 -4344
rect 928 -4346 930 -4344
rect 938 -4346 940 -4344
rect 954 -4346 956 -4344
rect 962 -4346 964 -4344
rect 972 -4346 974 -4344
rect 988 -4346 990 -4344
rect 998 -4346 1000 -4344
rect 1006 -4346 1008 -4344
rect 1016 -4346 1018 -4344
rect 1032 -4346 1034 -4344
rect 1040 -4346 1042 -4344
rect 1056 -4346 1058 -4344
rect 1072 -4346 1074 -4344
rect 1080 -4346 1082 -4344
rect 1090 -4346 1092 -4344
rect 1216 -4346 1218 -4344
rect 1226 -4346 1228 -4344
rect 1242 -4346 1244 -4344
rect 1252 -4346 1254 -4344
rect 1268 -4346 1270 -4344
rect 1278 -4346 1280 -4344
rect 1286 -4346 1288 -4344
rect 1296 -4346 1298 -4344
rect 1312 -4346 1314 -4344
rect 1320 -4346 1322 -4344
rect 1330 -4346 1332 -4344
rect 1346 -4346 1348 -4344
rect 1356 -4346 1358 -4344
rect 1364 -4346 1366 -4344
rect 1374 -4346 1376 -4344
rect 1390 -4346 1392 -4344
rect 1398 -4346 1400 -4344
rect 1414 -4346 1416 -4344
rect 1430 -4346 1432 -4344
rect 1438 -4346 1440 -4344
rect 1448 -4346 1450 -4344
rect -1809 -4387 -1807 -4385
rect -1799 -4387 -1797 -4385
rect -1783 -4387 -1781 -4385
rect -1775 -4387 -1773 -4385
rect -1759 -4387 -1757 -4385
rect -1751 -4387 -1749 -4385
rect -1741 -4387 -1739 -4385
rect -1733 -4387 -1731 -4385
rect -1717 -4387 -1715 -4385
rect -1709 -4387 -1707 -4385
rect -1699 -4387 -1697 -4385
rect -1691 -4387 -1689 -4385
rect -1675 -4387 -1673 -4385
rect -1667 -4387 -1665 -4385
rect -1657 -4387 -1655 -4385
rect -1649 -4387 -1647 -4385
rect -1633 -4387 -1631 -4385
rect -1625 -4387 -1623 -4385
rect -1546 -4387 -1544 -4385
rect -1536 -4387 -1534 -4385
rect -1520 -4387 -1518 -4385
rect -1512 -4387 -1510 -4385
rect -1496 -4387 -1494 -4385
rect -1488 -4387 -1486 -4385
rect -1478 -4387 -1476 -4385
rect -1470 -4387 -1468 -4385
rect -1454 -4387 -1452 -4385
rect -1446 -4387 -1444 -4385
rect -1436 -4387 -1434 -4385
rect -1428 -4387 -1426 -4385
rect -1412 -4387 -1410 -4385
rect -1404 -4387 -1402 -4385
rect -1394 -4387 -1392 -4385
rect -1386 -4387 -1384 -4385
rect -1370 -4387 -1368 -4385
rect -1362 -4387 -1360 -4385
rect -1229 -4387 -1227 -4385
rect -1219 -4387 -1217 -4385
rect -1203 -4387 -1201 -4385
rect -1195 -4387 -1193 -4385
rect -1179 -4387 -1177 -4385
rect -1171 -4387 -1169 -4385
rect -1161 -4387 -1159 -4385
rect -1153 -4387 -1151 -4385
rect -1137 -4387 -1135 -4385
rect -1129 -4387 -1127 -4385
rect -1119 -4387 -1117 -4385
rect -1111 -4387 -1109 -4385
rect -1095 -4387 -1093 -4385
rect -1087 -4387 -1085 -4385
rect -1077 -4387 -1075 -4385
rect -1069 -4387 -1067 -4385
rect -1053 -4387 -1051 -4385
rect -1045 -4387 -1043 -4385
rect -930 -4387 -928 -4385
rect -920 -4387 -918 -4385
rect -904 -4387 -902 -4385
rect -896 -4387 -894 -4385
rect -880 -4387 -878 -4385
rect -872 -4387 -870 -4385
rect -862 -4387 -860 -4385
rect -854 -4387 -852 -4385
rect -838 -4387 -836 -4385
rect -830 -4387 -828 -4385
rect -820 -4387 -818 -4385
rect -812 -4387 -810 -4385
rect -796 -4387 -794 -4385
rect -788 -4387 -786 -4385
rect -778 -4387 -776 -4385
rect -770 -4387 -768 -4385
rect -754 -4387 -752 -4385
rect -746 -4387 -744 -4385
rect -572 -4387 -570 -4385
rect -562 -4387 -560 -4385
rect -546 -4387 -544 -4385
rect -538 -4387 -536 -4385
rect -522 -4387 -520 -4385
rect -514 -4387 -512 -4385
rect -504 -4387 -502 -4385
rect -496 -4387 -494 -4385
rect -480 -4387 -478 -4385
rect -472 -4387 -470 -4385
rect -462 -4387 -460 -4385
rect -454 -4387 -452 -4385
rect -438 -4387 -436 -4385
rect -430 -4387 -428 -4385
rect -420 -4387 -418 -4385
rect -412 -4387 -410 -4385
rect -396 -4387 -394 -4385
rect -388 -4387 -386 -4385
rect -1809 -4463 -1807 -4395
rect -1799 -4463 -1797 -4395
rect -1783 -4463 -1781 -4395
rect -1775 -4463 -1773 -4395
rect -1759 -4463 -1757 -4395
rect -1751 -4463 -1749 -4395
rect -1741 -4463 -1739 -4395
rect -1733 -4463 -1731 -4395
rect -1717 -4463 -1715 -4395
rect -1709 -4428 -1707 -4395
rect -1699 -4428 -1697 -4395
rect -1709 -4430 -1697 -4428
rect -1709 -4463 -1707 -4430
rect -1699 -4463 -1697 -4430
rect -1691 -4463 -1689 -4395
rect -1675 -4463 -1673 -4395
rect -1667 -4463 -1665 -4395
rect -1657 -4463 -1655 -4395
rect -1649 -4463 -1647 -4395
rect -1633 -4463 -1631 -4395
rect -1625 -4463 -1623 -4395
rect -1546 -4463 -1544 -4395
rect -1536 -4463 -1534 -4395
rect -1520 -4463 -1518 -4395
rect -1512 -4463 -1510 -4395
rect -1496 -4463 -1494 -4395
rect -1488 -4463 -1486 -4395
rect -1478 -4463 -1476 -4395
rect -1470 -4463 -1468 -4395
rect -1454 -4463 -1452 -4395
rect -1446 -4428 -1444 -4395
rect -1436 -4428 -1434 -4395
rect -1446 -4430 -1434 -4428
rect -1446 -4463 -1444 -4430
rect -1436 -4463 -1434 -4430
rect -1428 -4463 -1426 -4395
rect -1412 -4463 -1410 -4395
rect -1404 -4463 -1402 -4395
rect -1394 -4463 -1392 -4395
rect -1386 -4463 -1384 -4395
rect -1370 -4463 -1368 -4395
rect -1362 -4463 -1360 -4395
rect -1229 -4463 -1227 -4395
rect -1219 -4463 -1217 -4395
rect -1203 -4463 -1201 -4395
rect -1195 -4463 -1193 -4395
rect -1179 -4463 -1177 -4395
rect -1171 -4463 -1169 -4395
rect -1161 -4463 -1159 -4395
rect -1153 -4463 -1151 -4395
rect -1137 -4463 -1135 -4395
rect -1129 -4428 -1127 -4395
rect -1119 -4428 -1117 -4395
rect -1129 -4430 -1117 -4428
rect -1129 -4463 -1127 -4430
rect -1119 -4463 -1117 -4430
rect -1111 -4463 -1109 -4395
rect -1095 -4463 -1093 -4395
rect -1087 -4463 -1085 -4395
rect -1077 -4463 -1075 -4395
rect -1069 -4463 -1067 -4395
rect -1053 -4463 -1051 -4395
rect -1045 -4463 -1043 -4395
rect -930 -4463 -928 -4395
rect -920 -4463 -918 -4395
rect -904 -4463 -902 -4395
rect -896 -4463 -894 -4395
rect -880 -4463 -878 -4395
rect -872 -4463 -870 -4395
rect -862 -4463 -860 -4395
rect -854 -4463 -852 -4395
rect -838 -4463 -836 -4395
rect -830 -4428 -828 -4395
rect -820 -4428 -818 -4395
rect -830 -4430 -818 -4428
rect -830 -4463 -828 -4430
rect -820 -4463 -818 -4430
rect -812 -4463 -810 -4395
rect -796 -4463 -794 -4395
rect -788 -4463 -786 -4395
rect -778 -4463 -776 -4395
rect -770 -4463 -768 -4395
rect -754 -4463 -752 -4395
rect -746 -4463 -744 -4395
rect -572 -4463 -570 -4395
rect -562 -4463 -560 -4395
rect -546 -4463 -544 -4395
rect -538 -4463 -536 -4395
rect -522 -4463 -520 -4395
rect -514 -4463 -512 -4395
rect -504 -4463 -502 -4395
rect -496 -4463 -494 -4395
rect -480 -4463 -478 -4395
rect -472 -4428 -470 -4395
rect -462 -4428 -460 -4395
rect -472 -4430 -460 -4428
rect -472 -4463 -470 -4430
rect -462 -4463 -460 -4430
rect -454 -4463 -452 -4395
rect -438 -4463 -436 -4395
rect -430 -4463 -428 -4395
rect -420 -4463 -418 -4395
rect -412 -4463 -410 -4395
rect -396 -4463 -394 -4395
rect -388 -4463 -386 -4395
rect -1809 -4469 -1807 -4467
rect -1799 -4469 -1797 -4467
rect -1783 -4469 -1781 -4467
rect -1775 -4469 -1773 -4467
rect -1759 -4469 -1757 -4467
rect -1751 -4469 -1749 -4467
rect -1741 -4469 -1739 -4467
rect -1733 -4469 -1731 -4467
rect -1717 -4469 -1715 -4467
rect -1709 -4469 -1707 -4467
rect -1699 -4469 -1697 -4467
rect -1691 -4469 -1689 -4467
rect -1675 -4469 -1673 -4467
rect -1667 -4469 -1665 -4467
rect -1657 -4469 -1655 -4467
rect -1649 -4469 -1647 -4467
rect -1633 -4469 -1631 -4467
rect -1625 -4469 -1623 -4467
rect -1546 -4469 -1544 -4467
rect -1536 -4469 -1534 -4467
rect -1520 -4469 -1518 -4467
rect -1512 -4469 -1510 -4467
rect -1496 -4469 -1494 -4467
rect -1488 -4469 -1486 -4467
rect -1478 -4469 -1476 -4467
rect -1470 -4469 -1468 -4467
rect -1454 -4469 -1452 -4467
rect -1446 -4469 -1444 -4467
rect -1436 -4469 -1434 -4467
rect -1428 -4469 -1426 -4467
rect -1412 -4469 -1410 -4467
rect -1404 -4469 -1402 -4467
rect -1394 -4469 -1392 -4467
rect -1386 -4469 -1384 -4467
rect -1370 -4469 -1368 -4467
rect -1362 -4469 -1360 -4467
rect -1229 -4469 -1227 -4467
rect -1219 -4469 -1217 -4467
rect -1203 -4469 -1201 -4467
rect -1195 -4469 -1193 -4467
rect -1179 -4469 -1177 -4467
rect -1171 -4469 -1169 -4467
rect -1161 -4469 -1159 -4467
rect -1153 -4469 -1151 -4467
rect -1137 -4469 -1135 -4467
rect -1129 -4469 -1127 -4467
rect -1119 -4469 -1117 -4467
rect -1111 -4469 -1109 -4467
rect -1095 -4469 -1093 -4467
rect -1087 -4469 -1085 -4467
rect -1077 -4469 -1075 -4467
rect -1069 -4469 -1067 -4467
rect -1053 -4469 -1051 -4467
rect -1045 -4469 -1043 -4467
rect -930 -4469 -928 -4467
rect -920 -4469 -918 -4467
rect -904 -4469 -902 -4467
rect -896 -4469 -894 -4467
rect -880 -4469 -878 -4467
rect -872 -4469 -870 -4467
rect -862 -4469 -860 -4467
rect -854 -4469 -852 -4467
rect -838 -4469 -836 -4467
rect -830 -4469 -828 -4467
rect -820 -4469 -818 -4467
rect -812 -4469 -810 -4467
rect -796 -4469 -794 -4467
rect -788 -4469 -786 -4467
rect -778 -4469 -776 -4467
rect -770 -4469 -768 -4467
rect -754 -4469 -752 -4467
rect -746 -4469 -744 -4467
rect -572 -4469 -570 -4467
rect -562 -4469 -560 -4467
rect -546 -4469 -544 -4467
rect -538 -4469 -536 -4467
rect -522 -4469 -520 -4467
rect -514 -4469 -512 -4467
rect -504 -4469 -502 -4467
rect -496 -4469 -494 -4467
rect -480 -4469 -478 -4467
rect -472 -4469 -470 -4467
rect -462 -4469 -460 -4467
rect -454 -4469 -452 -4467
rect -438 -4469 -436 -4467
rect -430 -4469 -428 -4467
rect -420 -4469 -418 -4467
rect -412 -4469 -410 -4467
rect -396 -4469 -394 -4467
rect -388 -4469 -386 -4467
rect -1809 -4558 -1807 -4556
rect -1799 -4558 -1797 -4556
rect -1783 -4558 -1781 -4556
rect -1775 -4558 -1773 -4556
rect -1759 -4558 -1757 -4556
rect -1751 -4558 -1749 -4556
rect -1741 -4558 -1739 -4556
rect -1733 -4558 -1731 -4556
rect -1717 -4558 -1715 -4556
rect -1709 -4558 -1707 -4556
rect -1699 -4558 -1697 -4556
rect -1691 -4558 -1689 -4556
rect -1675 -4558 -1673 -4556
rect -1667 -4558 -1665 -4556
rect -1657 -4558 -1655 -4556
rect -1649 -4558 -1647 -4556
rect -1633 -4558 -1631 -4556
rect -1625 -4558 -1623 -4556
rect -1546 -4558 -1544 -4556
rect -1536 -4558 -1534 -4556
rect -1520 -4558 -1518 -4556
rect -1512 -4558 -1510 -4556
rect -1496 -4558 -1494 -4556
rect -1488 -4558 -1486 -4556
rect -1478 -4558 -1476 -4556
rect -1470 -4558 -1468 -4556
rect -1454 -4558 -1452 -4556
rect -1446 -4558 -1444 -4556
rect -1436 -4558 -1434 -4556
rect -1428 -4558 -1426 -4556
rect -1412 -4558 -1410 -4556
rect -1404 -4558 -1402 -4556
rect -1394 -4558 -1392 -4556
rect -1386 -4558 -1384 -4556
rect -1370 -4558 -1368 -4556
rect -1362 -4558 -1360 -4556
rect -1229 -4558 -1227 -4556
rect -1219 -4558 -1217 -4556
rect -1203 -4558 -1201 -4556
rect -1195 -4558 -1193 -4556
rect -1179 -4558 -1177 -4556
rect -1171 -4558 -1169 -4556
rect -1161 -4558 -1159 -4556
rect -1153 -4558 -1151 -4556
rect -1137 -4558 -1135 -4556
rect -1129 -4558 -1127 -4556
rect -1119 -4558 -1117 -4556
rect -1111 -4558 -1109 -4556
rect -1095 -4558 -1093 -4556
rect -1087 -4558 -1085 -4556
rect -1077 -4558 -1075 -4556
rect -1069 -4558 -1067 -4556
rect -1053 -4558 -1051 -4556
rect -1045 -4558 -1043 -4556
rect -930 -4558 -928 -4556
rect -920 -4558 -918 -4556
rect -904 -4558 -902 -4556
rect -896 -4558 -894 -4556
rect -880 -4558 -878 -4556
rect -872 -4558 -870 -4556
rect -862 -4558 -860 -4556
rect -854 -4558 -852 -4556
rect -838 -4558 -836 -4556
rect -830 -4558 -828 -4556
rect -820 -4558 -818 -4556
rect -812 -4558 -810 -4556
rect -796 -4558 -794 -4556
rect -788 -4558 -786 -4556
rect -778 -4558 -776 -4556
rect -770 -4558 -768 -4556
rect -754 -4558 -752 -4556
rect -746 -4558 -744 -4556
rect -572 -4558 -570 -4556
rect -562 -4558 -560 -4556
rect -546 -4558 -544 -4556
rect -538 -4558 -536 -4556
rect -522 -4558 -520 -4556
rect -514 -4558 -512 -4556
rect -504 -4558 -502 -4556
rect -496 -4558 -494 -4556
rect -480 -4558 -478 -4556
rect -472 -4558 -470 -4556
rect -462 -4558 -460 -4556
rect -454 -4558 -452 -4556
rect -438 -4558 -436 -4556
rect -430 -4558 -428 -4556
rect -420 -4558 -418 -4556
rect -412 -4558 -410 -4556
rect -396 -4558 -394 -4556
rect -388 -4558 -386 -4556
rect -214 -4558 -212 -4556
rect -204 -4558 -202 -4556
rect -188 -4558 -186 -4556
rect -180 -4558 -178 -4556
rect -164 -4558 -162 -4556
rect -156 -4558 -154 -4556
rect -146 -4558 -144 -4556
rect -138 -4558 -136 -4556
rect -122 -4558 -120 -4556
rect -114 -4558 -112 -4556
rect -104 -4558 -102 -4556
rect -96 -4558 -94 -4556
rect -80 -4558 -78 -4556
rect -72 -4558 -70 -4556
rect -62 -4558 -60 -4556
rect -54 -4558 -52 -4556
rect -38 -4558 -36 -4556
rect -30 -4558 -28 -4556
rect 144 -4558 146 -4556
rect 154 -4558 156 -4556
rect 170 -4558 172 -4556
rect 178 -4558 180 -4556
rect 194 -4558 196 -4556
rect 202 -4558 204 -4556
rect 212 -4558 214 -4556
rect 220 -4558 222 -4556
rect 236 -4558 238 -4556
rect 244 -4558 246 -4556
rect 254 -4558 256 -4556
rect 262 -4558 264 -4556
rect 278 -4558 280 -4556
rect 286 -4558 288 -4556
rect 296 -4558 298 -4556
rect 304 -4558 306 -4556
rect 320 -4558 322 -4556
rect 328 -4558 330 -4556
rect 500 -4558 502 -4556
rect 510 -4558 512 -4556
rect 526 -4558 528 -4556
rect 534 -4558 536 -4556
rect 550 -4558 552 -4556
rect 558 -4558 560 -4556
rect 568 -4558 570 -4556
rect 576 -4558 578 -4556
rect 592 -4558 594 -4556
rect 600 -4558 602 -4556
rect 610 -4558 612 -4556
rect 618 -4558 620 -4556
rect 634 -4558 636 -4556
rect 642 -4558 644 -4556
rect 652 -4558 654 -4556
rect 660 -4558 662 -4556
rect 676 -4558 678 -4556
rect 684 -4558 686 -4556
rect 858 -4558 860 -4556
rect 868 -4558 870 -4556
rect 884 -4558 886 -4556
rect 892 -4558 894 -4556
rect 908 -4558 910 -4556
rect 916 -4558 918 -4556
rect 926 -4558 928 -4556
rect 934 -4558 936 -4556
rect 950 -4558 952 -4556
rect 958 -4558 960 -4556
rect 968 -4558 970 -4556
rect 976 -4558 978 -4556
rect 992 -4558 994 -4556
rect 1000 -4558 1002 -4556
rect 1010 -4558 1012 -4556
rect 1018 -4558 1020 -4556
rect 1034 -4558 1036 -4556
rect 1042 -4558 1044 -4556
rect 1216 -4558 1218 -4556
rect 1226 -4558 1228 -4556
rect 1242 -4558 1244 -4556
rect 1250 -4558 1252 -4556
rect 1266 -4558 1268 -4556
rect 1274 -4558 1276 -4556
rect 1284 -4558 1286 -4556
rect 1292 -4558 1294 -4556
rect 1308 -4558 1310 -4556
rect 1316 -4558 1318 -4556
rect 1326 -4558 1328 -4556
rect 1334 -4558 1336 -4556
rect 1350 -4558 1352 -4556
rect 1358 -4558 1360 -4556
rect 1368 -4558 1370 -4556
rect 1376 -4558 1378 -4556
rect 1392 -4558 1394 -4556
rect 1400 -4558 1402 -4556
rect -1809 -4634 -1807 -4566
rect -1799 -4634 -1797 -4566
rect -1783 -4634 -1781 -4566
rect -1775 -4634 -1773 -4566
rect -1759 -4634 -1757 -4566
rect -1751 -4634 -1749 -4566
rect -1741 -4634 -1739 -4566
rect -1733 -4634 -1731 -4566
rect -1717 -4634 -1715 -4566
rect -1709 -4599 -1707 -4566
rect -1699 -4599 -1697 -4566
rect -1709 -4601 -1697 -4599
rect -1709 -4634 -1707 -4601
rect -1699 -4634 -1697 -4601
rect -1691 -4634 -1689 -4566
rect -1675 -4634 -1673 -4566
rect -1667 -4634 -1665 -4566
rect -1657 -4634 -1655 -4566
rect -1649 -4634 -1647 -4566
rect -1633 -4634 -1631 -4566
rect -1625 -4634 -1623 -4566
rect -1546 -4634 -1544 -4566
rect -1536 -4634 -1534 -4566
rect -1520 -4634 -1518 -4566
rect -1512 -4634 -1510 -4566
rect -1496 -4634 -1494 -4566
rect -1488 -4634 -1486 -4566
rect -1478 -4634 -1476 -4566
rect -1470 -4634 -1468 -4566
rect -1454 -4634 -1452 -4566
rect -1446 -4599 -1444 -4566
rect -1436 -4599 -1434 -4566
rect -1446 -4601 -1434 -4599
rect -1446 -4634 -1444 -4601
rect -1436 -4634 -1434 -4601
rect -1428 -4634 -1426 -4566
rect -1412 -4634 -1410 -4566
rect -1404 -4634 -1402 -4566
rect -1394 -4634 -1392 -4566
rect -1386 -4634 -1384 -4566
rect -1370 -4634 -1368 -4566
rect -1362 -4634 -1360 -4566
rect -1229 -4634 -1227 -4566
rect -1219 -4634 -1217 -4566
rect -1203 -4634 -1201 -4566
rect -1195 -4634 -1193 -4566
rect -1179 -4634 -1177 -4566
rect -1171 -4634 -1169 -4566
rect -1161 -4634 -1159 -4566
rect -1153 -4634 -1151 -4566
rect -1137 -4634 -1135 -4566
rect -1129 -4599 -1127 -4566
rect -1119 -4599 -1117 -4566
rect -1129 -4601 -1117 -4599
rect -1129 -4634 -1127 -4601
rect -1119 -4634 -1117 -4601
rect -1111 -4634 -1109 -4566
rect -1095 -4634 -1093 -4566
rect -1087 -4634 -1085 -4566
rect -1077 -4634 -1075 -4566
rect -1069 -4634 -1067 -4566
rect -1053 -4634 -1051 -4566
rect -1045 -4634 -1043 -4566
rect -930 -4634 -928 -4566
rect -920 -4634 -918 -4566
rect -904 -4634 -902 -4566
rect -896 -4634 -894 -4566
rect -880 -4634 -878 -4566
rect -872 -4634 -870 -4566
rect -862 -4634 -860 -4566
rect -854 -4634 -852 -4566
rect -838 -4634 -836 -4566
rect -830 -4599 -828 -4566
rect -820 -4599 -818 -4566
rect -830 -4601 -818 -4599
rect -830 -4634 -828 -4601
rect -820 -4634 -818 -4601
rect -812 -4634 -810 -4566
rect -796 -4634 -794 -4566
rect -788 -4634 -786 -4566
rect -778 -4634 -776 -4566
rect -770 -4634 -768 -4566
rect -754 -4634 -752 -4566
rect -746 -4634 -744 -4566
rect -572 -4634 -570 -4566
rect -562 -4634 -560 -4566
rect -546 -4634 -544 -4566
rect -538 -4634 -536 -4566
rect -522 -4634 -520 -4566
rect -514 -4634 -512 -4566
rect -504 -4634 -502 -4566
rect -496 -4634 -494 -4566
rect -480 -4634 -478 -4566
rect -472 -4599 -470 -4566
rect -462 -4599 -460 -4566
rect -472 -4601 -460 -4599
rect -472 -4634 -470 -4601
rect -462 -4634 -460 -4601
rect -454 -4634 -452 -4566
rect -438 -4634 -436 -4566
rect -430 -4634 -428 -4566
rect -420 -4634 -418 -4566
rect -412 -4634 -410 -4566
rect -396 -4634 -394 -4566
rect -388 -4634 -386 -4566
rect -214 -4634 -212 -4566
rect -204 -4634 -202 -4566
rect -188 -4634 -186 -4566
rect -180 -4634 -178 -4566
rect -164 -4634 -162 -4566
rect -156 -4634 -154 -4566
rect -146 -4634 -144 -4566
rect -138 -4634 -136 -4566
rect -122 -4634 -120 -4566
rect -114 -4599 -112 -4566
rect -104 -4599 -102 -4566
rect -114 -4601 -102 -4599
rect -114 -4634 -112 -4601
rect -104 -4634 -102 -4601
rect -96 -4634 -94 -4566
rect -80 -4634 -78 -4566
rect -72 -4634 -70 -4566
rect -62 -4634 -60 -4566
rect -54 -4634 -52 -4566
rect -38 -4634 -36 -4566
rect -30 -4634 -28 -4566
rect 144 -4634 146 -4566
rect 154 -4634 156 -4566
rect 170 -4634 172 -4566
rect 178 -4634 180 -4566
rect 194 -4634 196 -4566
rect 202 -4634 204 -4566
rect 212 -4634 214 -4566
rect 220 -4634 222 -4566
rect 236 -4634 238 -4566
rect 244 -4599 246 -4566
rect 254 -4599 256 -4566
rect 244 -4601 256 -4599
rect 244 -4634 246 -4601
rect 254 -4634 256 -4601
rect 262 -4634 264 -4566
rect 278 -4634 280 -4566
rect 286 -4634 288 -4566
rect 296 -4634 298 -4566
rect 304 -4634 306 -4566
rect 320 -4634 322 -4566
rect 328 -4634 330 -4566
rect 500 -4634 502 -4566
rect 510 -4634 512 -4566
rect 526 -4634 528 -4566
rect 534 -4634 536 -4566
rect 550 -4634 552 -4566
rect 558 -4634 560 -4566
rect 568 -4634 570 -4566
rect 576 -4634 578 -4566
rect 592 -4634 594 -4566
rect 600 -4599 602 -4566
rect 610 -4599 612 -4566
rect 600 -4601 612 -4599
rect 600 -4634 602 -4601
rect 610 -4634 612 -4601
rect 618 -4634 620 -4566
rect 634 -4634 636 -4566
rect 642 -4634 644 -4566
rect 652 -4634 654 -4566
rect 660 -4634 662 -4566
rect 676 -4634 678 -4566
rect 684 -4634 686 -4566
rect 858 -4634 860 -4566
rect 868 -4634 870 -4566
rect 884 -4634 886 -4566
rect 892 -4634 894 -4566
rect 908 -4634 910 -4566
rect 916 -4634 918 -4566
rect 926 -4634 928 -4566
rect 934 -4634 936 -4566
rect 950 -4634 952 -4566
rect 958 -4599 960 -4566
rect 968 -4599 970 -4566
rect 958 -4601 970 -4599
rect 958 -4634 960 -4601
rect 968 -4634 970 -4601
rect 976 -4634 978 -4566
rect 992 -4634 994 -4566
rect 1000 -4634 1002 -4566
rect 1010 -4634 1012 -4566
rect 1018 -4634 1020 -4566
rect 1034 -4634 1036 -4566
rect 1042 -4634 1044 -4566
rect 1216 -4634 1218 -4566
rect 1226 -4634 1228 -4566
rect 1242 -4634 1244 -4566
rect 1250 -4634 1252 -4566
rect 1266 -4634 1268 -4566
rect 1274 -4634 1276 -4566
rect 1284 -4634 1286 -4566
rect 1292 -4634 1294 -4566
rect 1308 -4634 1310 -4566
rect 1316 -4599 1318 -4566
rect 1326 -4599 1328 -4566
rect 1316 -4601 1328 -4599
rect 1316 -4634 1318 -4601
rect 1326 -4634 1328 -4601
rect 1334 -4634 1336 -4566
rect 1350 -4634 1352 -4566
rect 1358 -4634 1360 -4566
rect 1368 -4634 1370 -4566
rect 1376 -4634 1378 -4566
rect 1392 -4634 1394 -4566
rect 1400 -4634 1402 -4566
rect -1809 -4640 -1807 -4638
rect -1799 -4640 -1797 -4638
rect -1783 -4640 -1781 -4638
rect -1775 -4640 -1773 -4638
rect -1759 -4640 -1757 -4638
rect -1751 -4640 -1749 -4638
rect -1741 -4640 -1739 -4638
rect -1733 -4640 -1731 -4638
rect -1717 -4640 -1715 -4638
rect -1709 -4640 -1707 -4638
rect -1699 -4640 -1697 -4638
rect -1691 -4640 -1689 -4638
rect -1675 -4640 -1673 -4638
rect -1667 -4640 -1665 -4638
rect -1657 -4640 -1655 -4638
rect -1649 -4640 -1647 -4638
rect -1633 -4640 -1631 -4638
rect -1625 -4640 -1623 -4638
rect -1546 -4640 -1544 -4638
rect -1536 -4640 -1534 -4638
rect -1520 -4640 -1518 -4638
rect -1512 -4640 -1510 -4638
rect -1496 -4640 -1494 -4638
rect -1488 -4640 -1486 -4638
rect -1478 -4640 -1476 -4638
rect -1470 -4640 -1468 -4638
rect -1454 -4640 -1452 -4638
rect -1446 -4640 -1444 -4638
rect -1436 -4640 -1434 -4638
rect -1428 -4640 -1426 -4638
rect -1412 -4640 -1410 -4638
rect -1404 -4640 -1402 -4638
rect -1394 -4640 -1392 -4638
rect -1386 -4640 -1384 -4638
rect -1370 -4640 -1368 -4638
rect -1362 -4640 -1360 -4638
rect -1229 -4640 -1227 -4638
rect -1219 -4640 -1217 -4638
rect -1203 -4640 -1201 -4638
rect -1195 -4640 -1193 -4638
rect -1179 -4640 -1177 -4638
rect -1171 -4640 -1169 -4638
rect -1161 -4640 -1159 -4638
rect -1153 -4640 -1151 -4638
rect -1137 -4640 -1135 -4638
rect -1129 -4640 -1127 -4638
rect -1119 -4640 -1117 -4638
rect -1111 -4640 -1109 -4638
rect -1095 -4640 -1093 -4638
rect -1087 -4640 -1085 -4638
rect -1077 -4640 -1075 -4638
rect -1069 -4640 -1067 -4638
rect -1053 -4640 -1051 -4638
rect -1045 -4640 -1043 -4638
rect -930 -4640 -928 -4638
rect -920 -4640 -918 -4638
rect -904 -4640 -902 -4638
rect -896 -4640 -894 -4638
rect -880 -4640 -878 -4638
rect -872 -4640 -870 -4638
rect -862 -4640 -860 -4638
rect -854 -4640 -852 -4638
rect -838 -4640 -836 -4638
rect -830 -4640 -828 -4638
rect -820 -4640 -818 -4638
rect -812 -4640 -810 -4638
rect -796 -4640 -794 -4638
rect -788 -4640 -786 -4638
rect -778 -4640 -776 -4638
rect -770 -4640 -768 -4638
rect -754 -4640 -752 -4638
rect -746 -4640 -744 -4638
rect -572 -4640 -570 -4638
rect -562 -4640 -560 -4638
rect -546 -4640 -544 -4638
rect -538 -4640 -536 -4638
rect -522 -4640 -520 -4638
rect -514 -4640 -512 -4638
rect -504 -4640 -502 -4638
rect -496 -4640 -494 -4638
rect -480 -4640 -478 -4638
rect -472 -4640 -470 -4638
rect -462 -4640 -460 -4638
rect -454 -4640 -452 -4638
rect -438 -4640 -436 -4638
rect -430 -4640 -428 -4638
rect -420 -4640 -418 -4638
rect -412 -4640 -410 -4638
rect -396 -4640 -394 -4638
rect -388 -4640 -386 -4638
rect -214 -4640 -212 -4638
rect -204 -4640 -202 -4638
rect -188 -4640 -186 -4638
rect -180 -4640 -178 -4638
rect -164 -4640 -162 -4638
rect -156 -4640 -154 -4638
rect -146 -4640 -144 -4638
rect -138 -4640 -136 -4638
rect -122 -4640 -120 -4638
rect -114 -4640 -112 -4638
rect -104 -4640 -102 -4638
rect -96 -4640 -94 -4638
rect -80 -4640 -78 -4638
rect -72 -4640 -70 -4638
rect -62 -4640 -60 -4638
rect -54 -4640 -52 -4638
rect -38 -4640 -36 -4638
rect -30 -4640 -28 -4638
rect 144 -4640 146 -4638
rect 154 -4640 156 -4638
rect 170 -4640 172 -4638
rect 178 -4640 180 -4638
rect 194 -4640 196 -4638
rect 202 -4640 204 -4638
rect 212 -4640 214 -4638
rect 220 -4640 222 -4638
rect 236 -4640 238 -4638
rect 244 -4640 246 -4638
rect 254 -4640 256 -4638
rect 262 -4640 264 -4638
rect 278 -4640 280 -4638
rect 286 -4640 288 -4638
rect 296 -4640 298 -4638
rect 304 -4640 306 -4638
rect 320 -4640 322 -4638
rect 328 -4640 330 -4638
rect 500 -4640 502 -4638
rect 510 -4640 512 -4638
rect 526 -4640 528 -4638
rect 534 -4640 536 -4638
rect 550 -4640 552 -4638
rect 558 -4640 560 -4638
rect 568 -4640 570 -4638
rect 576 -4640 578 -4638
rect 592 -4640 594 -4638
rect 600 -4640 602 -4638
rect 610 -4640 612 -4638
rect 618 -4640 620 -4638
rect 634 -4640 636 -4638
rect 642 -4640 644 -4638
rect 652 -4640 654 -4638
rect 660 -4640 662 -4638
rect 676 -4640 678 -4638
rect 684 -4640 686 -4638
rect 858 -4640 860 -4638
rect 868 -4640 870 -4638
rect 884 -4640 886 -4638
rect 892 -4640 894 -4638
rect 908 -4640 910 -4638
rect 916 -4640 918 -4638
rect 926 -4640 928 -4638
rect 934 -4640 936 -4638
rect 950 -4640 952 -4638
rect 958 -4640 960 -4638
rect 968 -4640 970 -4638
rect 976 -4640 978 -4638
rect 992 -4640 994 -4638
rect 1000 -4640 1002 -4638
rect 1010 -4640 1012 -4638
rect 1018 -4640 1020 -4638
rect 1034 -4640 1036 -4638
rect 1042 -4640 1044 -4638
rect 1216 -4640 1218 -4638
rect 1226 -4640 1228 -4638
rect 1242 -4640 1244 -4638
rect 1250 -4640 1252 -4638
rect 1266 -4640 1268 -4638
rect 1274 -4640 1276 -4638
rect 1284 -4640 1286 -4638
rect 1292 -4640 1294 -4638
rect 1308 -4640 1310 -4638
rect 1316 -4640 1318 -4638
rect 1326 -4640 1328 -4638
rect 1334 -4640 1336 -4638
rect 1350 -4640 1352 -4638
rect 1358 -4640 1360 -4638
rect 1368 -4640 1370 -4638
rect 1376 -4640 1378 -4638
rect 1392 -4640 1394 -4638
rect 1400 -4640 1402 -4638
rect -1546 -4729 -1544 -4727
rect -1536 -4729 -1534 -4727
rect -1520 -4729 -1518 -4727
rect -1512 -4729 -1510 -4727
rect -1496 -4729 -1494 -4727
rect -1488 -4729 -1486 -4727
rect -1478 -4729 -1476 -4727
rect -1470 -4729 -1468 -4727
rect -1454 -4729 -1452 -4727
rect -1446 -4729 -1444 -4727
rect -1436 -4729 -1434 -4727
rect -1428 -4729 -1426 -4727
rect -1412 -4729 -1410 -4727
rect -1404 -4729 -1402 -4727
rect -1394 -4729 -1392 -4727
rect -1386 -4729 -1384 -4727
rect -1370 -4729 -1368 -4727
rect -1362 -4729 -1360 -4727
rect -1229 -4729 -1227 -4727
rect -1219 -4729 -1217 -4727
rect -1203 -4729 -1201 -4727
rect -1195 -4729 -1193 -4727
rect -1179 -4729 -1177 -4727
rect -1171 -4729 -1169 -4727
rect -1161 -4729 -1159 -4727
rect -1153 -4729 -1151 -4727
rect -1137 -4729 -1135 -4727
rect -1129 -4729 -1127 -4727
rect -1119 -4729 -1117 -4727
rect -1111 -4729 -1109 -4727
rect -1095 -4729 -1093 -4727
rect -1087 -4729 -1085 -4727
rect -1077 -4729 -1075 -4727
rect -1069 -4729 -1067 -4727
rect -1053 -4729 -1051 -4727
rect -1045 -4729 -1043 -4727
rect -930 -4729 -928 -4727
rect -920 -4729 -918 -4727
rect -904 -4729 -902 -4727
rect -896 -4729 -894 -4727
rect -880 -4729 -878 -4727
rect -872 -4729 -870 -4727
rect -862 -4729 -860 -4727
rect -854 -4729 -852 -4727
rect -838 -4729 -836 -4727
rect -830 -4729 -828 -4727
rect -820 -4729 -818 -4727
rect -812 -4729 -810 -4727
rect -796 -4729 -794 -4727
rect -788 -4729 -786 -4727
rect -778 -4729 -776 -4727
rect -770 -4729 -768 -4727
rect -754 -4729 -752 -4727
rect -746 -4729 -744 -4727
rect -572 -4729 -570 -4727
rect -562 -4729 -560 -4727
rect -546 -4729 -544 -4727
rect -538 -4729 -536 -4727
rect -522 -4729 -520 -4727
rect -514 -4729 -512 -4727
rect -504 -4729 -502 -4727
rect -496 -4729 -494 -4727
rect -480 -4729 -478 -4727
rect -472 -4729 -470 -4727
rect -462 -4729 -460 -4727
rect -454 -4729 -452 -4727
rect -438 -4729 -436 -4727
rect -430 -4729 -428 -4727
rect -420 -4729 -418 -4727
rect -412 -4729 -410 -4727
rect -396 -4729 -394 -4727
rect -388 -4729 -386 -4727
rect -214 -4729 -212 -4727
rect -204 -4729 -202 -4727
rect -188 -4729 -186 -4727
rect -180 -4729 -178 -4727
rect -164 -4729 -162 -4727
rect -156 -4729 -154 -4727
rect -146 -4729 -144 -4727
rect -138 -4729 -136 -4727
rect -122 -4729 -120 -4727
rect -114 -4729 -112 -4727
rect -104 -4729 -102 -4727
rect -96 -4729 -94 -4727
rect -80 -4729 -78 -4727
rect -72 -4729 -70 -4727
rect -62 -4729 -60 -4727
rect -54 -4729 -52 -4727
rect -38 -4729 -36 -4727
rect -30 -4729 -28 -4727
rect 144 -4729 146 -4727
rect 154 -4729 156 -4727
rect 170 -4729 172 -4727
rect 178 -4729 180 -4727
rect 194 -4729 196 -4727
rect 202 -4729 204 -4727
rect 212 -4729 214 -4727
rect 220 -4729 222 -4727
rect 236 -4729 238 -4727
rect 244 -4729 246 -4727
rect 254 -4729 256 -4727
rect 262 -4729 264 -4727
rect 278 -4729 280 -4727
rect 286 -4729 288 -4727
rect 296 -4729 298 -4727
rect 304 -4729 306 -4727
rect 320 -4729 322 -4727
rect 328 -4729 330 -4727
rect 500 -4729 502 -4727
rect 510 -4729 512 -4727
rect 526 -4729 528 -4727
rect 534 -4729 536 -4727
rect 550 -4729 552 -4727
rect 558 -4729 560 -4727
rect 568 -4729 570 -4727
rect 576 -4729 578 -4727
rect 592 -4729 594 -4727
rect 600 -4729 602 -4727
rect 610 -4729 612 -4727
rect 618 -4729 620 -4727
rect 634 -4729 636 -4727
rect 642 -4729 644 -4727
rect 652 -4729 654 -4727
rect 660 -4729 662 -4727
rect 676 -4729 678 -4727
rect 684 -4729 686 -4727
rect 858 -4729 860 -4727
rect 868 -4729 870 -4727
rect 884 -4729 886 -4727
rect 892 -4729 894 -4727
rect 908 -4729 910 -4727
rect 916 -4729 918 -4727
rect 926 -4729 928 -4727
rect 934 -4729 936 -4727
rect 950 -4729 952 -4727
rect 958 -4729 960 -4727
rect 968 -4729 970 -4727
rect 976 -4729 978 -4727
rect 992 -4729 994 -4727
rect 1000 -4729 1002 -4727
rect 1010 -4729 1012 -4727
rect 1018 -4729 1020 -4727
rect 1034 -4729 1036 -4727
rect 1042 -4729 1044 -4727
rect 1216 -4729 1218 -4727
rect 1226 -4729 1228 -4727
rect 1242 -4729 1244 -4727
rect 1250 -4729 1252 -4727
rect 1266 -4729 1268 -4727
rect 1274 -4729 1276 -4727
rect 1284 -4729 1286 -4727
rect 1292 -4729 1294 -4727
rect 1308 -4729 1310 -4727
rect 1316 -4729 1318 -4727
rect 1326 -4729 1328 -4727
rect 1334 -4729 1336 -4727
rect 1350 -4729 1352 -4727
rect 1358 -4729 1360 -4727
rect 1368 -4729 1370 -4727
rect 1376 -4729 1378 -4727
rect 1392 -4729 1394 -4727
rect 1400 -4729 1402 -4727
rect -1546 -4805 -1544 -4737
rect -1536 -4805 -1534 -4737
rect -1520 -4805 -1518 -4737
rect -1512 -4805 -1510 -4737
rect -1496 -4805 -1494 -4737
rect -1488 -4805 -1486 -4737
rect -1478 -4805 -1476 -4737
rect -1470 -4805 -1468 -4737
rect -1454 -4805 -1452 -4737
rect -1446 -4770 -1444 -4737
rect -1436 -4770 -1434 -4737
rect -1446 -4772 -1434 -4770
rect -1446 -4805 -1444 -4772
rect -1436 -4805 -1434 -4772
rect -1428 -4805 -1426 -4737
rect -1412 -4805 -1410 -4737
rect -1404 -4805 -1402 -4737
rect -1394 -4805 -1392 -4737
rect -1386 -4805 -1384 -4737
rect -1370 -4805 -1368 -4737
rect -1362 -4805 -1360 -4737
rect -1229 -4805 -1227 -4737
rect -1219 -4805 -1217 -4737
rect -1203 -4805 -1201 -4737
rect -1195 -4805 -1193 -4737
rect -1179 -4805 -1177 -4737
rect -1171 -4805 -1169 -4737
rect -1161 -4805 -1159 -4737
rect -1153 -4805 -1151 -4737
rect -1137 -4805 -1135 -4737
rect -1129 -4770 -1127 -4737
rect -1119 -4770 -1117 -4737
rect -1129 -4772 -1117 -4770
rect -1129 -4805 -1127 -4772
rect -1119 -4805 -1117 -4772
rect -1111 -4805 -1109 -4737
rect -1095 -4805 -1093 -4737
rect -1087 -4805 -1085 -4737
rect -1077 -4805 -1075 -4737
rect -1069 -4805 -1067 -4737
rect -1053 -4805 -1051 -4737
rect -1045 -4805 -1043 -4737
rect -930 -4805 -928 -4737
rect -920 -4805 -918 -4737
rect -904 -4805 -902 -4737
rect -896 -4805 -894 -4737
rect -880 -4805 -878 -4737
rect -872 -4805 -870 -4737
rect -862 -4805 -860 -4737
rect -854 -4805 -852 -4737
rect -838 -4805 -836 -4737
rect -830 -4770 -828 -4737
rect -820 -4770 -818 -4737
rect -830 -4772 -818 -4770
rect -830 -4805 -828 -4772
rect -820 -4805 -818 -4772
rect -812 -4805 -810 -4737
rect -796 -4805 -794 -4737
rect -788 -4805 -786 -4737
rect -778 -4805 -776 -4737
rect -770 -4805 -768 -4737
rect -754 -4805 -752 -4737
rect -746 -4805 -744 -4737
rect -572 -4805 -570 -4737
rect -562 -4805 -560 -4737
rect -546 -4805 -544 -4737
rect -538 -4805 -536 -4737
rect -522 -4805 -520 -4737
rect -514 -4805 -512 -4737
rect -504 -4805 -502 -4737
rect -496 -4805 -494 -4737
rect -480 -4805 -478 -4737
rect -472 -4770 -470 -4737
rect -462 -4770 -460 -4737
rect -472 -4772 -460 -4770
rect -472 -4805 -470 -4772
rect -462 -4805 -460 -4772
rect -454 -4805 -452 -4737
rect -438 -4805 -436 -4737
rect -430 -4805 -428 -4737
rect -420 -4805 -418 -4737
rect -412 -4805 -410 -4737
rect -396 -4805 -394 -4737
rect -388 -4805 -386 -4737
rect -214 -4805 -212 -4737
rect -204 -4805 -202 -4737
rect -188 -4805 -186 -4737
rect -180 -4805 -178 -4737
rect -164 -4805 -162 -4737
rect -156 -4805 -154 -4737
rect -146 -4805 -144 -4737
rect -138 -4805 -136 -4737
rect -122 -4805 -120 -4737
rect -114 -4770 -112 -4737
rect -104 -4770 -102 -4737
rect -114 -4772 -102 -4770
rect -114 -4805 -112 -4772
rect -104 -4805 -102 -4772
rect -96 -4805 -94 -4737
rect -80 -4805 -78 -4737
rect -72 -4805 -70 -4737
rect -62 -4805 -60 -4737
rect -54 -4805 -52 -4737
rect -38 -4805 -36 -4737
rect -30 -4805 -28 -4737
rect 144 -4805 146 -4737
rect 154 -4805 156 -4737
rect 170 -4805 172 -4737
rect 178 -4805 180 -4737
rect 194 -4805 196 -4737
rect 202 -4805 204 -4737
rect 212 -4805 214 -4737
rect 220 -4805 222 -4737
rect 236 -4805 238 -4737
rect 244 -4770 246 -4737
rect 254 -4770 256 -4737
rect 244 -4772 256 -4770
rect 244 -4805 246 -4772
rect 254 -4805 256 -4772
rect 262 -4805 264 -4737
rect 278 -4805 280 -4737
rect 286 -4805 288 -4737
rect 296 -4805 298 -4737
rect 304 -4805 306 -4737
rect 320 -4805 322 -4737
rect 328 -4805 330 -4737
rect 500 -4805 502 -4737
rect 510 -4805 512 -4737
rect 526 -4805 528 -4737
rect 534 -4805 536 -4737
rect 550 -4805 552 -4737
rect 558 -4805 560 -4737
rect 568 -4805 570 -4737
rect 576 -4805 578 -4737
rect 592 -4805 594 -4737
rect 600 -4770 602 -4737
rect 610 -4770 612 -4737
rect 600 -4772 612 -4770
rect 600 -4805 602 -4772
rect 610 -4805 612 -4772
rect 618 -4805 620 -4737
rect 634 -4805 636 -4737
rect 642 -4805 644 -4737
rect 652 -4805 654 -4737
rect 660 -4805 662 -4737
rect 676 -4805 678 -4737
rect 684 -4805 686 -4737
rect 858 -4805 860 -4737
rect 868 -4805 870 -4737
rect 884 -4805 886 -4737
rect 892 -4805 894 -4737
rect 908 -4805 910 -4737
rect 916 -4805 918 -4737
rect 926 -4805 928 -4737
rect 934 -4805 936 -4737
rect 950 -4805 952 -4737
rect 958 -4770 960 -4737
rect 968 -4770 970 -4737
rect 958 -4772 970 -4770
rect 958 -4805 960 -4772
rect 968 -4805 970 -4772
rect 976 -4805 978 -4737
rect 992 -4805 994 -4737
rect 1000 -4805 1002 -4737
rect 1010 -4805 1012 -4737
rect 1018 -4805 1020 -4737
rect 1034 -4805 1036 -4737
rect 1042 -4805 1044 -4737
rect 1216 -4805 1218 -4737
rect 1226 -4805 1228 -4737
rect 1242 -4805 1244 -4737
rect 1250 -4805 1252 -4737
rect 1266 -4805 1268 -4737
rect 1274 -4805 1276 -4737
rect 1284 -4805 1286 -4737
rect 1292 -4805 1294 -4737
rect 1308 -4805 1310 -4737
rect 1316 -4770 1318 -4737
rect 1326 -4770 1328 -4737
rect 1316 -4772 1328 -4770
rect 1316 -4805 1318 -4772
rect 1326 -4805 1328 -4772
rect 1334 -4805 1336 -4737
rect 1350 -4805 1352 -4737
rect 1358 -4805 1360 -4737
rect 1368 -4805 1370 -4737
rect 1376 -4805 1378 -4737
rect 1392 -4805 1394 -4737
rect 1400 -4805 1402 -4737
rect -1546 -4811 -1544 -4809
rect -1536 -4811 -1534 -4809
rect -1520 -4811 -1518 -4809
rect -1512 -4811 -1510 -4809
rect -1496 -4811 -1494 -4809
rect -1488 -4811 -1486 -4809
rect -1478 -4811 -1476 -4809
rect -1470 -4811 -1468 -4809
rect -1454 -4811 -1452 -4809
rect -1446 -4811 -1444 -4809
rect -1436 -4811 -1434 -4809
rect -1428 -4811 -1426 -4809
rect -1412 -4811 -1410 -4809
rect -1404 -4811 -1402 -4809
rect -1394 -4811 -1392 -4809
rect -1386 -4811 -1384 -4809
rect -1370 -4811 -1368 -4809
rect -1362 -4811 -1360 -4809
rect -1229 -4811 -1227 -4809
rect -1219 -4811 -1217 -4809
rect -1203 -4811 -1201 -4809
rect -1195 -4811 -1193 -4809
rect -1179 -4811 -1177 -4809
rect -1171 -4811 -1169 -4809
rect -1161 -4811 -1159 -4809
rect -1153 -4811 -1151 -4809
rect -1137 -4811 -1135 -4809
rect -1129 -4811 -1127 -4809
rect -1119 -4811 -1117 -4809
rect -1111 -4811 -1109 -4809
rect -1095 -4811 -1093 -4809
rect -1087 -4811 -1085 -4809
rect -1077 -4811 -1075 -4809
rect -1069 -4811 -1067 -4809
rect -1053 -4811 -1051 -4809
rect -1045 -4811 -1043 -4809
rect -930 -4811 -928 -4809
rect -920 -4811 -918 -4809
rect -904 -4811 -902 -4809
rect -896 -4811 -894 -4809
rect -880 -4811 -878 -4809
rect -872 -4811 -870 -4809
rect -862 -4811 -860 -4809
rect -854 -4811 -852 -4809
rect -838 -4811 -836 -4809
rect -830 -4811 -828 -4809
rect -820 -4811 -818 -4809
rect -812 -4811 -810 -4809
rect -796 -4811 -794 -4809
rect -788 -4811 -786 -4809
rect -778 -4811 -776 -4809
rect -770 -4811 -768 -4809
rect -754 -4811 -752 -4809
rect -746 -4811 -744 -4809
rect -572 -4811 -570 -4809
rect -562 -4811 -560 -4809
rect -546 -4811 -544 -4809
rect -538 -4811 -536 -4809
rect -522 -4811 -520 -4809
rect -514 -4811 -512 -4809
rect -504 -4811 -502 -4809
rect -496 -4811 -494 -4809
rect -480 -4811 -478 -4809
rect -472 -4811 -470 -4809
rect -462 -4811 -460 -4809
rect -454 -4811 -452 -4809
rect -438 -4811 -436 -4809
rect -430 -4811 -428 -4809
rect -420 -4811 -418 -4809
rect -412 -4811 -410 -4809
rect -396 -4811 -394 -4809
rect -388 -4811 -386 -4809
rect -214 -4811 -212 -4809
rect -204 -4811 -202 -4809
rect -188 -4811 -186 -4809
rect -180 -4811 -178 -4809
rect -164 -4811 -162 -4809
rect -156 -4811 -154 -4809
rect -146 -4811 -144 -4809
rect -138 -4811 -136 -4809
rect -122 -4811 -120 -4809
rect -114 -4811 -112 -4809
rect -104 -4811 -102 -4809
rect -96 -4811 -94 -4809
rect -80 -4811 -78 -4809
rect -72 -4811 -70 -4809
rect -62 -4811 -60 -4809
rect -54 -4811 -52 -4809
rect -38 -4811 -36 -4809
rect -30 -4811 -28 -4809
rect 144 -4811 146 -4809
rect 154 -4811 156 -4809
rect 170 -4811 172 -4809
rect 178 -4811 180 -4809
rect 194 -4811 196 -4809
rect 202 -4811 204 -4809
rect 212 -4811 214 -4809
rect 220 -4811 222 -4809
rect 236 -4811 238 -4809
rect 244 -4811 246 -4809
rect 254 -4811 256 -4809
rect 262 -4811 264 -4809
rect 278 -4811 280 -4809
rect 286 -4811 288 -4809
rect 296 -4811 298 -4809
rect 304 -4811 306 -4809
rect 320 -4811 322 -4809
rect 328 -4811 330 -4809
rect 500 -4811 502 -4809
rect 510 -4811 512 -4809
rect 526 -4811 528 -4809
rect 534 -4811 536 -4809
rect 550 -4811 552 -4809
rect 558 -4811 560 -4809
rect 568 -4811 570 -4809
rect 576 -4811 578 -4809
rect 592 -4811 594 -4809
rect 600 -4811 602 -4809
rect 610 -4811 612 -4809
rect 618 -4811 620 -4809
rect 634 -4811 636 -4809
rect 642 -4811 644 -4809
rect 652 -4811 654 -4809
rect 660 -4811 662 -4809
rect 676 -4811 678 -4809
rect 684 -4811 686 -4809
rect 858 -4811 860 -4809
rect 868 -4811 870 -4809
rect 884 -4811 886 -4809
rect 892 -4811 894 -4809
rect 908 -4811 910 -4809
rect 916 -4811 918 -4809
rect 926 -4811 928 -4809
rect 934 -4811 936 -4809
rect 950 -4811 952 -4809
rect 958 -4811 960 -4809
rect 968 -4811 970 -4809
rect 976 -4811 978 -4809
rect 992 -4811 994 -4809
rect 1000 -4811 1002 -4809
rect 1010 -4811 1012 -4809
rect 1018 -4811 1020 -4809
rect 1034 -4811 1036 -4809
rect 1042 -4811 1044 -4809
rect 1216 -4811 1218 -4809
rect 1226 -4811 1228 -4809
rect 1242 -4811 1244 -4809
rect 1250 -4811 1252 -4809
rect 1266 -4811 1268 -4809
rect 1274 -4811 1276 -4809
rect 1284 -4811 1286 -4809
rect 1292 -4811 1294 -4809
rect 1308 -4811 1310 -4809
rect 1316 -4811 1318 -4809
rect 1326 -4811 1328 -4809
rect 1334 -4811 1336 -4809
rect 1350 -4811 1352 -4809
rect 1358 -4811 1360 -4809
rect 1368 -4811 1370 -4809
rect 1376 -4811 1378 -4809
rect 1392 -4811 1394 -4809
rect 1400 -4811 1402 -4809
rect -1304 -4844 -1302 -4842
rect -1296 -4844 -1294 -4842
rect -1286 -4844 -1284 -4842
rect -930 -4844 -928 -4842
rect -922 -4844 -920 -4842
rect -912 -4844 -910 -4842
rect -572 -4844 -570 -4842
rect -564 -4844 -562 -4842
rect -554 -4844 -552 -4842
rect -214 -4844 -212 -4842
rect -206 -4844 -204 -4842
rect -196 -4844 -194 -4842
rect 144 -4844 146 -4842
rect 152 -4844 154 -4842
rect 162 -4844 164 -4842
rect 500 -4844 502 -4842
rect 508 -4844 510 -4842
rect 518 -4844 520 -4842
rect 858 -4844 860 -4842
rect 866 -4844 868 -4842
rect 876 -4844 878 -4842
rect 1216 -4844 1218 -4842
rect 1224 -4844 1226 -4842
rect 1234 -4844 1236 -4842
rect -1304 -4920 -1302 -4852
rect -1296 -4876 -1294 -4852
rect -1296 -4920 -1294 -4880
rect -1286 -4920 -1284 -4852
rect -930 -4920 -928 -4852
rect -922 -4876 -920 -4852
rect -922 -4920 -920 -4880
rect -912 -4920 -910 -4852
rect -572 -4920 -570 -4852
rect -564 -4876 -562 -4852
rect -564 -4920 -562 -4880
rect -554 -4920 -552 -4852
rect -214 -4920 -212 -4852
rect -206 -4876 -204 -4852
rect -206 -4920 -204 -4880
rect -196 -4920 -194 -4852
rect 144 -4920 146 -4852
rect 152 -4876 154 -4852
rect 152 -4920 154 -4880
rect 162 -4920 164 -4852
rect 500 -4920 502 -4852
rect 508 -4876 510 -4852
rect 508 -4920 510 -4880
rect 518 -4920 520 -4852
rect 858 -4920 860 -4852
rect 866 -4876 868 -4852
rect 866 -4920 868 -4880
rect 876 -4920 878 -4852
rect 1216 -4920 1218 -4852
rect 1224 -4876 1226 -4852
rect 1224 -4920 1226 -4880
rect 1234 -4920 1236 -4852
rect -1304 -4926 -1302 -4924
rect -1296 -4926 -1294 -4924
rect -1286 -4926 -1284 -4924
rect -930 -4926 -928 -4924
rect -922 -4926 -920 -4924
rect -912 -4926 -910 -4924
rect -572 -4926 -570 -4924
rect -564 -4926 -562 -4924
rect -554 -4926 -552 -4924
rect -214 -4926 -212 -4924
rect -206 -4926 -204 -4924
rect -196 -4926 -194 -4924
rect 144 -4926 146 -4924
rect 152 -4926 154 -4924
rect 162 -4926 164 -4924
rect 500 -4926 502 -4924
rect 508 -4926 510 -4924
rect 518 -4926 520 -4924
rect 858 -4926 860 -4924
rect 866 -4926 868 -4924
rect 876 -4926 878 -4924
rect 1216 -4926 1218 -4924
rect 1224 -4926 1226 -4924
rect 1234 -4926 1236 -4924
rect -1229 -5003 -1227 -5001
rect -1219 -5003 -1217 -5001
rect -1203 -5003 -1201 -5001
rect -1193 -5003 -1191 -5001
rect -1185 -5003 -1183 -5001
rect -1175 -5003 -1173 -5001
rect -1159 -5003 -1157 -5001
rect -1151 -5003 -1149 -5001
rect -1141 -5003 -1139 -5001
rect -930 -5003 -928 -5001
rect -920 -5003 -918 -5001
rect -904 -5003 -902 -5001
rect -894 -5003 -892 -5001
rect -878 -5003 -876 -5001
rect -868 -5003 -866 -5001
rect -860 -5003 -858 -5001
rect -850 -5003 -848 -5001
rect -834 -5003 -832 -5001
rect -826 -5003 -824 -5001
rect -816 -5003 -814 -5001
rect -800 -5003 -798 -5001
rect -790 -5003 -788 -5001
rect -782 -5003 -780 -5001
rect -772 -5003 -770 -5001
rect -756 -5003 -754 -5001
rect -748 -5003 -746 -5001
rect -732 -5003 -730 -5001
rect -716 -5003 -714 -5001
rect -708 -5003 -706 -5001
rect -698 -5003 -696 -5001
rect -572 -5003 -570 -5001
rect -562 -5003 -560 -5001
rect -546 -5003 -544 -5001
rect -536 -5003 -534 -5001
rect -520 -5003 -518 -5001
rect -510 -5003 -508 -5001
rect -502 -5003 -500 -5001
rect -492 -5003 -490 -5001
rect -476 -5003 -474 -5001
rect -468 -5003 -466 -5001
rect -458 -5003 -456 -5001
rect -442 -5003 -440 -5001
rect -432 -5003 -430 -5001
rect -424 -5003 -422 -5001
rect -414 -5003 -412 -5001
rect -398 -5003 -396 -5001
rect -390 -5003 -388 -5001
rect -374 -5003 -372 -5001
rect -358 -5003 -356 -5001
rect -350 -5003 -348 -5001
rect -340 -5003 -338 -5001
rect -214 -5003 -212 -5001
rect -204 -5003 -202 -5001
rect -188 -5003 -186 -5001
rect -178 -5003 -176 -5001
rect -162 -5003 -160 -5001
rect -152 -5003 -150 -5001
rect -144 -5003 -142 -5001
rect -134 -5003 -132 -5001
rect -118 -5003 -116 -5001
rect -110 -5003 -108 -5001
rect -100 -5003 -98 -5001
rect -84 -5003 -82 -5001
rect -74 -5003 -72 -5001
rect -66 -5003 -64 -5001
rect -56 -5003 -54 -5001
rect -40 -5003 -38 -5001
rect -32 -5003 -30 -5001
rect -16 -5003 -14 -5001
rect 0 -5003 2 -5001
rect 8 -5003 10 -5001
rect 18 -5003 20 -5001
rect 144 -5003 146 -5001
rect 154 -5003 156 -5001
rect 170 -5003 172 -5001
rect 180 -5003 182 -5001
rect 196 -5003 198 -5001
rect 206 -5003 208 -5001
rect 214 -5003 216 -5001
rect 224 -5003 226 -5001
rect 240 -5003 242 -5001
rect 248 -5003 250 -5001
rect 258 -5003 260 -5001
rect 274 -5003 276 -5001
rect 284 -5003 286 -5001
rect 292 -5003 294 -5001
rect 302 -5003 304 -5001
rect 318 -5003 320 -5001
rect 326 -5003 328 -5001
rect 342 -5003 344 -5001
rect 358 -5003 360 -5001
rect 366 -5003 368 -5001
rect 376 -5003 378 -5001
rect 500 -5003 502 -5001
rect 510 -5003 512 -5001
rect 526 -5003 528 -5001
rect 536 -5003 538 -5001
rect 552 -5003 554 -5001
rect 562 -5003 564 -5001
rect 570 -5003 572 -5001
rect 580 -5003 582 -5001
rect 596 -5003 598 -5001
rect 604 -5003 606 -5001
rect 614 -5003 616 -5001
rect 630 -5003 632 -5001
rect 640 -5003 642 -5001
rect 648 -5003 650 -5001
rect 658 -5003 660 -5001
rect 674 -5003 676 -5001
rect 682 -5003 684 -5001
rect 698 -5003 700 -5001
rect 714 -5003 716 -5001
rect 722 -5003 724 -5001
rect 732 -5003 734 -5001
rect 858 -5003 860 -5001
rect 868 -5003 870 -5001
rect 884 -5003 886 -5001
rect 894 -5003 896 -5001
rect 910 -5003 912 -5001
rect 920 -5003 922 -5001
rect 928 -5003 930 -5001
rect 938 -5003 940 -5001
rect 954 -5003 956 -5001
rect 962 -5003 964 -5001
rect 972 -5003 974 -5001
rect 988 -5003 990 -5001
rect 998 -5003 1000 -5001
rect 1006 -5003 1008 -5001
rect 1016 -5003 1018 -5001
rect 1032 -5003 1034 -5001
rect 1040 -5003 1042 -5001
rect 1056 -5003 1058 -5001
rect 1072 -5003 1074 -5001
rect 1080 -5003 1082 -5001
rect 1090 -5003 1092 -5001
rect 1216 -5003 1218 -5001
rect 1226 -5003 1228 -5001
rect 1242 -5003 1244 -5001
rect 1252 -5003 1254 -5001
rect 1268 -5003 1270 -5001
rect 1278 -5003 1280 -5001
rect 1286 -5003 1288 -5001
rect 1296 -5003 1298 -5001
rect 1312 -5003 1314 -5001
rect 1320 -5003 1322 -5001
rect 1330 -5003 1332 -5001
rect 1346 -5003 1348 -5001
rect 1356 -5003 1358 -5001
rect 1364 -5003 1366 -5001
rect 1374 -5003 1376 -5001
rect 1390 -5003 1392 -5001
rect 1398 -5003 1400 -5001
rect 1414 -5003 1416 -5001
rect 1430 -5003 1432 -5001
rect 1438 -5003 1440 -5001
rect 1448 -5003 1450 -5001
rect -1229 -5079 -1227 -5011
rect -1219 -5079 -1217 -5011
rect -1203 -5079 -1201 -5011
rect -1193 -5079 -1191 -5011
rect -1185 -5079 -1183 -5011
rect -1175 -5079 -1173 -5011
rect -1159 -5079 -1157 -5011
rect -1151 -5079 -1149 -5011
rect -1141 -5079 -1139 -5011
rect -930 -5079 -928 -5011
rect -920 -5079 -918 -5011
rect -904 -5079 -902 -5011
rect -894 -5079 -892 -5011
rect -878 -5079 -876 -5011
rect -868 -5079 -866 -5011
rect -860 -5079 -858 -5011
rect -850 -5079 -848 -5011
rect -834 -5079 -832 -5011
rect -826 -5079 -824 -5011
rect -816 -5079 -814 -5011
rect -800 -5079 -798 -5011
rect -790 -5079 -788 -5011
rect -782 -5079 -780 -5011
rect -772 -5079 -770 -5011
rect -756 -5079 -754 -5011
rect -748 -5079 -746 -5011
rect -732 -5079 -730 -5011
rect -716 -5079 -714 -5011
rect -708 -5079 -706 -5011
rect -698 -5079 -696 -5011
rect -572 -5079 -570 -5011
rect -562 -5079 -560 -5011
rect -546 -5079 -544 -5011
rect -536 -5079 -534 -5011
rect -520 -5079 -518 -5011
rect -510 -5079 -508 -5011
rect -502 -5079 -500 -5011
rect -492 -5079 -490 -5011
rect -476 -5079 -474 -5011
rect -468 -5079 -466 -5011
rect -458 -5079 -456 -5011
rect -442 -5079 -440 -5011
rect -432 -5079 -430 -5011
rect -424 -5079 -422 -5011
rect -414 -5079 -412 -5011
rect -398 -5079 -396 -5011
rect -390 -5079 -388 -5011
rect -374 -5079 -372 -5011
rect -358 -5079 -356 -5011
rect -350 -5079 -348 -5011
rect -340 -5079 -338 -5011
rect -214 -5079 -212 -5011
rect -204 -5079 -202 -5011
rect -188 -5079 -186 -5011
rect -178 -5079 -176 -5011
rect -162 -5079 -160 -5011
rect -152 -5079 -150 -5011
rect -144 -5079 -142 -5011
rect -134 -5079 -132 -5011
rect -118 -5079 -116 -5011
rect -110 -5079 -108 -5011
rect -100 -5079 -98 -5011
rect -84 -5079 -82 -5011
rect -74 -5079 -72 -5011
rect -66 -5079 -64 -5011
rect -56 -5079 -54 -5011
rect -40 -5079 -38 -5011
rect -32 -5079 -30 -5011
rect -16 -5079 -14 -5011
rect 0 -5079 2 -5011
rect 8 -5079 10 -5011
rect 18 -5079 20 -5011
rect 144 -5079 146 -5011
rect 154 -5079 156 -5011
rect 170 -5079 172 -5011
rect 180 -5079 182 -5011
rect 196 -5079 198 -5011
rect 206 -5079 208 -5011
rect 214 -5079 216 -5011
rect 224 -5079 226 -5011
rect 240 -5079 242 -5011
rect 248 -5079 250 -5011
rect 258 -5079 260 -5011
rect 274 -5079 276 -5011
rect 284 -5079 286 -5011
rect 292 -5079 294 -5011
rect 302 -5079 304 -5011
rect 318 -5079 320 -5011
rect 326 -5079 328 -5011
rect 342 -5079 344 -5011
rect 358 -5079 360 -5011
rect 366 -5079 368 -5011
rect 376 -5079 378 -5011
rect 500 -5079 502 -5011
rect 510 -5079 512 -5011
rect 526 -5079 528 -5011
rect 536 -5079 538 -5011
rect 552 -5079 554 -5011
rect 562 -5079 564 -5011
rect 570 -5079 572 -5011
rect 580 -5079 582 -5011
rect 596 -5079 598 -5011
rect 604 -5079 606 -5011
rect 614 -5079 616 -5011
rect 630 -5079 632 -5011
rect 640 -5079 642 -5011
rect 648 -5079 650 -5011
rect 658 -5079 660 -5011
rect 674 -5079 676 -5011
rect 682 -5079 684 -5011
rect 698 -5079 700 -5011
rect 714 -5079 716 -5011
rect 722 -5079 724 -5011
rect 732 -5079 734 -5011
rect 858 -5079 860 -5011
rect 868 -5079 870 -5011
rect 884 -5079 886 -5011
rect 894 -5079 896 -5011
rect 910 -5079 912 -5011
rect 920 -5079 922 -5011
rect 928 -5079 930 -5011
rect 938 -5079 940 -5011
rect 954 -5079 956 -5011
rect 962 -5079 964 -5011
rect 972 -5079 974 -5011
rect 988 -5079 990 -5011
rect 998 -5079 1000 -5011
rect 1006 -5079 1008 -5011
rect 1016 -5079 1018 -5011
rect 1032 -5079 1034 -5011
rect 1040 -5079 1042 -5011
rect 1056 -5079 1058 -5011
rect 1072 -5079 1074 -5011
rect 1080 -5079 1082 -5011
rect 1090 -5079 1092 -5011
rect 1216 -5079 1218 -5011
rect 1226 -5079 1228 -5011
rect 1242 -5079 1244 -5011
rect 1252 -5079 1254 -5011
rect 1268 -5079 1270 -5011
rect 1278 -5079 1280 -5011
rect 1286 -5079 1288 -5011
rect 1296 -5079 1298 -5011
rect 1312 -5079 1314 -5011
rect 1320 -5079 1322 -5011
rect 1330 -5079 1332 -5011
rect 1346 -5079 1348 -5011
rect 1356 -5079 1358 -5011
rect 1364 -5079 1366 -5011
rect 1374 -5079 1376 -5011
rect 1390 -5079 1392 -5011
rect 1398 -5079 1400 -5011
rect 1414 -5079 1416 -5011
rect 1430 -5079 1432 -5011
rect 1438 -5079 1440 -5011
rect 1448 -5079 1450 -5011
rect -1229 -5085 -1227 -5083
rect -1219 -5085 -1217 -5083
rect -1203 -5085 -1201 -5083
rect -1193 -5085 -1191 -5083
rect -1185 -5085 -1183 -5083
rect -1175 -5085 -1173 -5083
rect -1159 -5085 -1157 -5083
rect -1151 -5085 -1149 -5083
rect -1141 -5085 -1139 -5083
rect -930 -5085 -928 -5083
rect -920 -5085 -918 -5083
rect -904 -5085 -902 -5083
rect -894 -5085 -892 -5083
rect -878 -5085 -876 -5083
rect -868 -5085 -866 -5083
rect -860 -5085 -858 -5083
rect -850 -5085 -848 -5083
rect -834 -5085 -832 -5083
rect -826 -5085 -824 -5083
rect -816 -5085 -814 -5083
rect -800 -5085 -798 -5083
rect -790 -5085 -788 -5083
rect -782 -5085 -780 -5083
rect -772 -5085 -770 -5083
rect -756 -5085 -754 -5083
rect -748 -5085 -746 -5083
rect -732 -5085 -730 -5083
rect -716 -5085 -714 -5083
rect -708 -5085 -706 -5083
rect -698 -5085 -696 -5083
rect -572 -5085 -570 -5083
rect -562 -5085 -560 -5083
rect -546 -5085 -544 -5083
rect -536 -5085 -534 -5083
rect -520 -5085 -518 -5083
rect -510 -5085 -508 -5083
rect -502 -5085 -500 -5083
rect -492 -5085 -490 -5083
rect -476 -5085 -474 -5083
rect -468 -5085 -466 -5083
rect -458 -5085 -456 -5083
rect -442 -5085 -440 -5083
rect -432 -5085 -430 -5083
rect -424 -5085 -422 -5083
rect -414 -5085 -412 -5083
rect -398 -5085 -396 -5083
rect -390 -5085 -388 -5083
rect -374 -5085 -372 -5083
rect -358 -5085 -356 -5083
rect -350 -5085 -348 -5083
rect -340 -5085 -338 -5083
rect -214 -5085 -212 -5083
rect -204 -5085 -202 -5083
rect -188 -5085 -186 -5083
rect -178 -5085 -176 -5083
rect -162 -5085 -160 -5083
rect -152 -5085 -150 -5083
rect -144 -5085 -142 -5083
rect -134 -5085 -132 -5083
rect -118 -5085 -116 -5083
rect -110 -5085 -108 -5083
rect -100 -5085 -98 -5083
rect -84 -5085 -82 -5083
rect -74 -5085 -72 -5083
rect -66 -5085 -64 -5083
rect -56 -5085 -54 -5083
rect -40 -5085 -38 -5083
rect -32 -5085 -30 -5083
rect -16 -5085 -14 -5083
rect 0 -5085 2 -5083
rect 8 -5085 10 -5083
rect 18 -5085 20 -5083
rect 144 -5085 146 -5083
rect 154 -5085 156 -5083
rect 170 -5085 172 -5083
rect 180 -5085 182 -5083
rect 196 -5085 198 -5083
rect 206 -5085 208 -5083
rect 214 -5085 216 -5083
rect 224 -5085 226 -5083
rect 240 -5085 242 -5083
rect 248 -5085 250 -5083
rect 258 -5085 260 -5083
rect 274 -5085 276 -5083
rect 284 -5085 286 -5083
rect 292 -5085 294 -5083
rect 302 -5085 304 -5083
rect 318 -5085 320 -5083
rect 326 -5085 328 -5083
rect 342 -5085 344 -5083
rect 358 -5085 360 -5083
rect 366 -5085 368 -5083
rect 376 -5085 378 -5083
rect 500 -5085 502 -5083
rect 510 -5085 512 -5083
rect 526 -5085 528 -5083
rect 536 -5085 538 -5083
rect 552 -5085 554 -5083
rect 562 -5085 564 -5083
rect 570 -5085 572 -5083
rect 580 -5085 582 -5083
rect 596 -5085 598 -5083
rect 604 -5085 606 -5083
rect 614 -5085 616 -5083
rect 630 -5085 632 -5083
rect 640 -5085 642 -5083
rect 648 -5085 650 -5083
rect 658 -5085 660 -5083
rect 674 -5085 676 -5083
rect 682 -5085 684 -5083
rect 698 -5085 700 -5083
rect 714 -5085 716 -5083
rect 722 -5085 724 -5083
rect 732 -5085 734 -5083
rect 858 -5085 860 -5083
rect 868 -5085 870 -5083
rect 884 -5085 886 -5083
rect 894 -5085 896 -5083
rect 910 -5085 912 -5083
rect 920 -5085 922 -5083
rect 928 -5085 930 -5083
rect 938 -5085 940 -5083
rect 954 -5085 956 -5083
rect 962 -5085 964 -5083
rect 972 -5085 974 -5083
rect 988 -5085 990 -5083
rect 998 -5085 1000 -5083
rect 1006 -5085 1008 -5083
rect 1016 -5085 1018 -5083
rect 1032 -5085 1034 -5083
rect 1040 -5085 1042 -5083
rect 1056 -5085 1058 -5083
rect 1072 -5085 1074 -5083
rect 1080 -5085 1082 -5083
rect 1090 -5085 1092 -5083
rect 1216 -5085 1218 -5083
rect 1226 -5085 1228 -5083
rect 1242 -5085 1244 -5083
rect 1252 -5085 1254 -5083
rect 1268 -5085 1270 -5083
rect 1278 -5085 1280 -5083
rect 1286 -5085 1288 -5083
rect 1296 -5085 1298 -5083
rect 1312 -5085 1314 -5083
rect 1320 -5085 1322 -5083
rect 1330 -5085 1332 -5083
rect 1346 -5085 1348 -5083
rect 1356 -5085 1358 -5083
rect 1364 -5085 1366 -5083
rect 1374 -5085 1376 -5083
rect 1390 -5085 1392 -5083
rect 1398 -5085 1400 -5083
rect 1414 -5085 1416 -5083
rect 1430 -5085 1432 -5083
rect 1438 -5085 1440 -5083
rect 1448 -5085 1450 -5083
rect -1805 -5122 -1803 -5120
rect -1795 -5122 -1793 -5120
rect -1779 -5122 -1777 -5120
rect -1771 -5122 -1769 -5120
rect -1755 -5122 -1753 -5120
rect -1747 -5122 -1745 -5120
rect -1737 -5122 -1735 -5120
rect -1729 -5122 -1727 -5120
rect -1713 -5122 -1711 -5120
rect -1705 -5122 -1703 -5120
rect -1695 -5122 -1693 -5120
rect -1687 -5122 -1685 -5120
rect -1671 -5122 -1669 -5120
rect -1663 -5122 -1661 -5120
rect -1653 -5122 -1651 -5120
rect -1645 -5122 -1643 -5120
rect -1629 -5122 -1627 -5120
rect -1621 -5122 -1619 -5120
rect -1542 -5122 -1540 -5120
rect -1532 -5122 -1530 -5120
rect -1516 -5122 -1514 -5120
rect -1508 -5122 -1506 -5120
rect -1492 -5122 -1490 -5120
rect -1484 -5122 -1482 -5120
rect -1474 -5122 -1472 -5120
rect -1466 -5122 -1464 -5120
rect -1450 -5122 -1448 -5120
rect -1442 -5122 -1440 -5120
rect -1432 -5122 -1430 -5120
rect -1424 -5122 -1422 -5120
rect -1408 -5122 -1406 -5120
rect -1400 -5122 -1398 -5120
rect -1390 -5122 -1388 -5120
rect -1382 -5122 -1380 -5120
rect -1366 -5122 -1364 -5120
rect -1358 -5122 -1356 -5120
rect -1229 -5122 -1227 -5120
rect -1219 -5122 -1217 -5120
rect -1203 -5122 -1201 -5120
rect -1195 -5122 -1193 -5120
rect -1179 -5122 -1177 -5120
rect -1171 -5122 -1169 -5120
rect -1161 -5122 -1159 -5120
rect -1153 -5122 -1151 -5120
rect -1137 -5122 -1135 -5120
rect -1129 -5122 -1127 -5120
rect -1119 -5122 -1117 -5120
rect -1111 -5122 -1109 -5120
rect -1095 -5122 -1093 -5120
rect -1087 -5122 -1085 -5120
rect -1077 -5122 -1075 -5120
rect -1069 -5122 -1067 -5120
rect -1053 -5122 -1051 -5120
rect -1045 -5122 -1043 -5120
rect -930 -5122 -928 -5120
rect -920 -5122 -918 -5120
rect -904 -5122 -902 -5120
rect -896 -5122 -894 -5120
rect -880 -5122 -878 -5120
rect -872 -5122 -870 -5120
rect -862 -5122 -860 -5120
rect -854 -5122 -852 -5120
rect -838 -5122 -836 -5120
rect -830 -5122 -828 -5120
rect -820 -5122 -818 -5120
rect -812 -5122 -810 -5120
rect -796 -5122 -794 -5120
rect -788 -5122 -786 -5120
rect -778 -5122 -776 -5120
rect -770 -5122 -768 -5120
rect -754 -5122 -752 -5120
rect -746 -5122 -744 -5120
rect -1805 -5198 -1803 -5130
rect -1795 -5198 -1793 -5130
rect -1779 -5198 -1777 -5130
rect -1771 -5198 -1769 -5130
rect -1755 -5198 -1753 -5130
rect -1747 -5198 -1745 -5130
rect -1737 -5198 -1735 -5130
rect -1729 -5198 -1727 -5130
rect -1713 -5198 -1711 -5130
rect -1705 -5163 -1703 -5130
rect -1695 -5163 -1693 -5130
rect -1705 -5165 -1693 -5163
rect -1705 -5198 -1703 -5165
rect -1695 -5198 -1693 -5165
rect -1687 -5198 -1685 -5130
rect -1671 -5198 -1669 -5130
rect -1663 -5198 -1661 -5130
rect -1653 -5198 -1651 -5130
rect -1645 -5198 -1643 -5130
rect -1629 -5198 -1627 -5130
rect -1621 -5198 -1619 -5130
rect -1542 -5198 -1540 -5130
rect -1532 -5198 -1530 -5130
rect -1516 -5198 -1514 -5130
rect -1508 -5198 -1506 -5130
rect -1492 -5198 -1490 -5130
rect -1484 -5198 -1482 -5130
rect -1474 -5198 -1472 -5130
rect -1466 -5198 -1464 -5130
rect -1450 -5198 -1448 -5130
rect -1442 -5163 -1440 -5130
rect -1432 -5163 -1430 -5130
rect -1442 -5165 -1430 -5163
rect -1442 -5198 -1440 -5165
rect -1432 -5198 -1430 -5165
rect -1424 -5198 -1422 -5130
rect -1408 -5198 -1406 -5130
rect -1400 -5198 -1398 -5130
rect -1390 -5198 -1388 -5130
rect -1382 -5198 -1380 -5130
rect -1366 -5198 -1364 -5130
rect -1358 -5198 -1356 -5130
rect -1229 -5198 -1227 -5130
rect -1219 -5198 -1217 -5130
rect -1203 -5198 -1201 -5130
rect -1195 -5198 -1193 -5130
rect -1179 -5198 -1177 -5130
rect -1171 -5198 -1169 -5130
rect -1161 -5198 -1159 -5130
rect -1153 -5198 -1151 -5130
rect -1137 -5198 -1135 -5130
rect -1129 -5163 -1127 -5130
rect -1119 -5163 -1117 -5130
rect -1129 -5165 -1117 -5163
rect -1129 -5198 -1127 -5165
rect -1119 -5198 -1117 -5165
rect -1111 -5198 -1109 -5130
rect -1095 -5198 -1093 -5130
rect -1087 -5198 -1085 -5130
rect -1077 -5198 -1075 -5130
rect -1069 -5198 -1067 -5130
rect -1053 -5198 -1051 -5130
rect -1045 -5198 -1043 -5130
rect -930 -5198 -928 -5130
rect -920 -5198 -918 -5130
rect -904 -5198 -902 -5130
rect -896 -5198 -894 -5130
rect -880 -5198 -878 -5130
rect -872 -5198 -870 -5130
rect -862 -5198 -860 -5130
rect -854 -5198 -852 -5130
rect -838 -5198 -836 -5130
rect -830 -5163 -828 -5130
rect -820 -5163 -818 -5130
rect -830 -5165 -818 -5163
rect -830 -5198 -828 -5165
rect -820 -5198 -818 -5165
rect -812 -5198 -810 -5130
rect -796 -5198 -794 -5130
rect -788 -5198 -786 -5130
rect -778 -5198 -776 -5130
rect -770 -5198 -768 -5130
rect -754 -5198 -752 -5130
rect -746 -5198 -744 -5130
rect -1805 -5204 -1803 -5202
rect -1795 -5204 -1793 -5202
rect -1779 -5204 -1777 -5202
rect -1771 -5204 -1769 -5202
rect -1755 -5204 -1753 -5202
rect -1747 -5204 -1745 -5202
rect -1737 -5204 -1735 -5202
rect -1729 -5204 -1727 -5202
rect -1713 -5204 -1711 -5202
rect -1705 -5204 -1703 -5202
rect -1695 -5204 -1693 -5202
rect -1687 -5204 -1685 -5202
rect -1671 -5204 -1669 -5202
rect -1663 -5204 -1661 -5202
rect -1653 -5204 -1651 -5202
rect -1645 -5204 -1643 -5202
rect -1629 -5204 -1627 -5202
rect -1621 -5204 -1619 -5202
rect -1542 -5204 -1540 -5202
rect -1532 -5204 -1530 -5202
rect -1516 -5204 -1514 -5202
rect -1508 -5204 -1506 -5202
rect -1492 -5204 -1490 -5202
rect -1484 -5204 -1482 -5202
rect -1474 -5204 -1472 -5202
rect -1466 -5204 -1464 -5202
rect -1450 -5204 -1448 -5202
rect -1442 -5204 -1440 -5202
rect -1432 -5204 -1430 -5202
rect -1424 -5204 -1422 -5202
rect -1408 -5204 -1406 -5202
rect -1400 -5204 -1398 -5202
rect -1390 -5204 -1388 -5202
rect -1382 -5204 -1380 -5202
rect -1366 -5204 -1364 -5202
rect -1358 -5204 -1356 -5202
rect -1229 -5204 -1227 -5202
rect -1219 -5204 -1217 -5202
rect -1203 -5204 -1201 -5202
rect -1195 -5204 -1193 -5202
rect -1179 -5204 -1177 -5202
rect -1171 -5204 -1169 -5202
rect -1161 -5204 -1159 -5202
rect -1153 -5204 -1151 -5202
rect -1137 -5204 -1135 -5202
rect -1129 -5204 -1127 -5202
rect -1119 -5204 -1117 -5202
rect -1111 -5204 -1109 -5202
rect -1095 -5204 -1093 -5202
rect -1087 -5204 -1085 -5202
rect -1077 -5204 -1075 -5202
rect -1069 -5204 -1067 -5202
rect -1053 -5204 -1051 -5202
rect -1045 -5204 -1043 -5202
rect -930 -5204 -928 -5202
rect -920 -5204 -918 -5202
rect -904 -5204 -902 -5202
rect -896 -5204 -894 -5202
rect -880 -5204 -878 -5202
rect -872 -5204 -870 -5202
rect -862 -5204 -860 -5202
rect -854 -5204 -852 -5202
rect -838 -5204 -836 -5202
rect -830 -5204 -828 -5202
rect -820 -5204 -818 -5202
rect -812 -5204 -810 -5202
rect -796 -5204 -794 -5202
rect -788 -5204 -786 -5202
rect -778 -5204 -776 -5202
rect -770 -5204 -768 -5202
rect -754 -5204 -752 -5202
rect -746 -5204 -744 -5202
rect -1805 -5293 -1803 -5291
rect -1795 -5293 -1793 -5291
rect -1779 -5293 -1777 -5291
rect -1771 -5293 -1769 -5291
rect -1755 -5293 -1753 -5291
rect -1747 -5293 -1745 -5291
rect -1737 -5293 -1735 -5291
rect -1729 -5293 -1727 -5291
rect -1713 -5293 -1711 -5291
rect -1705 -5293 -1703 -5291
rect -1695 -5293 -1693 -5291
rect -1687 -5293 -1685 -5291
rect -1671 -5293 -1669 -5291
rect -1663 -5293 -1661 -5291
rect -1653 -5293 -1651 -5291
rect -1645 -5293 -1643 -5291
rect -1629 -5293 -1627 -5291
rect -1621 -5293 -1619 -5291
rect -1542 -5293 -1540 -5291
rect -1532 -5293 -1530 -5291
rect -1516 -5293 -1514 -5291
rect -1508 -5293 -1506 -5291
rect -1492 -5293 -1490 -5291
rect -1484 -5293 -1482 -5291
rect -1474 -5293 -1472 -5291
rect -1466 -5293 -1464 -5291
rect -1450 -5293 -1448 -5291
rect -1442 -5293 -1440 -5291
rect -1432 -5293 -1430 -5291
rect -1424 -5293 -1422 -5291
rect -1408 -5293 -1406 -5291
rect -1400 -5293 -1398 -5291
rect -1390 -5293 -1388 -5291
rect -1382 -5293 -1380 -5291
rect -1366 -5293 -1364 -5291
rect -1358 -5293 -1356 -5291
rect -1229 -5293 -1227 -5291
rect -1219 -5293 -1217 -5291
rect -1203 -5293 -1201 -5291
rect -1195 -5293 -1193 -5291
rect -1179 -5293 -1177 -5291
rect -1171 -5293 -1169 -5291
rect -1161 -5293 -1159 -5291
rect -1153 -5293 -1151 -5291
rect -1137 -5293 -1135 -5291
rect -1129 -5293 -1127 -5291
rect -1119 -5293 -1117 -5291
rect -1111 -5293 -1109 -5291
rect -1095 -5293 -1093 -5291
rect -1087 -5293 -1085 -5291
rect -1077 -5293 -1075 -5291
rect -1069 -5293 -1067 -5291
rect -1053 -5293 -1051 -5291
rect -1045 -5293 -1043 -5291
rect -930 -5293 -928 -5291
rect -920 -5293 -918 -5291
rect -904 -5293 -902 -5291
rect -896 -5293 -894 -5291
rect -880 -5293 -878 -5291
rect -872 -5293 -870 -5291
rect -862 -5293 -860 -5291
rect -854 -5293 -852 -5291
rect -838 -5293 -836 -5291
rect -830 -5293 -828 -5291
rect -820 -5293 -818 -5291
rect -812 -5293 -810 -5291
rect -796 -5293 -794 -5291
rect -788 -5293 -786 -5291
rect -778 -5293 -776 -5291
rect -770 -5293 -768 -5291
rect -754 -5293 -752 -5291
rect -746 -5293 -744 -5291
rect -572 -5293 -570 -5291
rect -562 -5293 -560 -5291
rect -546 -5293 -544 -5291
rect -538 -5293 -536 -5291
rect -522 -5293 -520 -5291
rect -514 -5293 -512 -5291
rect -504 -5293 -502 -5291
rect -496 -5293 -494 -5291
rect -480 -5293 -478 -5291
rect -472 -5293 -470 -5291
rect -462 -5293 -460 -5291
rect -454 -5293 -452 -5291
rect -438 -5293 -436 -5291
rect -430 -5293 -428 -5291
rect -420 -5293 -418 -5291
rect -412 -5293 -410 -5291
rect -396 -5293 -394 -5291
rect -388 -5293 -386 -5291
rect -214 -5293 -212 -5291
rect -204 -5293 -202 -5291
rect -188 -5293 -186 -5291
rect -180 -5293 -178 -5291
rect -164 -5293 -162 -5291
rect -156 -5293 -154 -5291
rect -146 -5293 -144 -5291
rect -138 -5293 -136 -5291
rect -122 -5293 -120 -5291
rect -114 -5293 -112 -5291
rect -104 -5293 -102 -5291
rect -96 -5293 -94 -5291
rect -80 -5293 -78 -5291
rect -72 -5293 -70 -5291
rect -62 -5293 -60 -5291
rect -54 -5293 -52 -5291
rect -38 -5293 -36 -5291
rect -30 -5293 -28 -5291
rect 144 -5293 146 -5291
rect 154 -5293 156 -5291
rect 170 -5293 172 -5291
rect 178 -5293 180 -5291
rect 194 -5293 196 -5291
rect 202 -5293 204 -5291
rect 212 -5293 214 -5291
rect 220 -5293 222 -5291
rect 236 -5293 238 -5291
rect 244 -5293 246 -5291
rect 254 -5293 256 -5291
rect 262 -5293 264 -5291
rect 278 -5293 280 -5291
rect 286 -5293 288 -5291
rect 296 -5293 298 -5291
rect 304 -5293 306 -5291
rect 320 -5293 322 -5291
rect 328 -5293 330 -5291
rect 500 -5293 502 -5291
rect 510 -5293 512 -5291
rect 526 -5293 528 -5291
rect 534 -5293 536 -5291
rect 550 -5293 552 -5291
rect 558 -5293 560 -5291
rect 568 -5293 570 -5291
rect 576 -5293 578 -5291
rect 592 -5293 594 -5291
rect 600 -5293 602 -5291
rect 610 -5293 612 -5291
rect 618 -5293 620 -5291
rect 634 -5293 636 -5291
rect 642 -5293 644 -5291
rect 652 -5293 654 -5291
rect 660 -5293 662 -5291
rect 676 -5293 678 -5291
rect 684 -5293 686 -5291
rect 858 -5293 860 -5291
rect 868 -5293 870 -5291
rect 884 -5293 886 -5291
rect 892 -5293 894 -5291
rect 908 -5293 910 -5291
rect 916 -5293 918 -5291
rect 926 -5293 928 -5291
rect 934 -5293 936 -5291
rect 950 -5293 952 -5291
rect 958 -5293 960 -5291
rect 968 -5293 970 -5291
rect 976 -5293 978 -5291
rect 992 -5293 994 -5291
rect 1000 -5293 1002 -5291
rect 1010 -5293 1012 -5291
rect 1018 -5293 1020 -5291
rect 1034 -5293 1036 -5291
rect 1042 -5293 1044 -5291
rect 1216 -5293 1218 -5291
rect 1226 -5293 1228 -5291
rect 1242 -5293 1244 -5291
rect 1250 -5293 1252 -5291
rect 1266 -5293 1268 -5291
rect 1274 -5293 1276 -5291
rect 1284 -5293 1286 -5291
rect 1292 -5293 1294 -5291
rect 1308 -5293 1310 -5291
rect 1316 -5293 1318 -5291
rect 1326 -5293 1328 -5291
rect 1334 -5293 1336 -5291
rect 1350 -5293 1352 -5291
rect 1358 -5293 1360 -5291
rect 1368 -5293 1370 -5291
rect 1376 -5293 1378 -5291
rect 1392 -5293 1394 -5291
rect 1400 -5293 1402 -5291
rect -1805 -5369 -1803 -5301
rect -1795 -5369 -1793 -5301
rect -1779 -5369 -1777 -5301
rect -1771 -5369 -1769 -5301
rect -1755 -5369 -1753 -5301
rect -1747 -5369 -1745 -5301
rect -1737 -5369 -1735 -5301
rect -1729 -5369 -1727 -5301
rect -1713 -5369 -1711 -5301
rect -1705 -5334 -1703 -5301
rect -1695 -5334 -1693 -5301
rect -1705 -5336 -1693 -5334
rect -1705 -5369 -1703 -5336
rect -1695 -5369 -1693 -5336
rect -1687 -5369 -1685 -5301
rect -1671 -5369 -1669 -5301
rect -1663 -5369 -1661 -5301
rect -1653 -5369 -1651 -5301
rect -1645 -5369 -1643 -5301
rect -1629 -5369 -1627 -5301
rect -1621 -5369 -1619 -5301
rect -1542 -5369 -1540 -5301
rect -1532 -5369 -1530 -5301
rect -1516 -5369 -1514 -5301
rect -1508 -5369 -1506 -5301
rect -1492 -5369 -1490 -5301
rect -1484 -5369 -1482 -5301
rect -1474 -5369 -1472 -5301
rect -1466 -5369 -1464 -5301
rect -1450 -5369 -1448 -5301
rect -1442 -5334 -1440 -5301
rect -1432 -5334 -1430 -5301
rect -1442 -5336 -1430 -5334
rect -1442 -5369 -1440 -5336
rect -1432 -5369 -1430 -5336
rect -1424 -5369 -1422 -5301
rect -1408 -5369 -1406 -5301
rect -1400 -5369 -1398 -5301
rect -1390 -5369 -1388 -5301
rect -1382 -5369 -1380 -5301
rect -1366 -5369 -1364 -5301
rect -1358 -5369 -1356 -5301
rect -1229 -5369 -1227 -5301
rect -1219 -5369 -1217 -5301
rect -1203 -5369 -1201 -5301
rect -1195 -5369 -1193 -5301
rect -1179 -5369 -1177 -5301
rect -1171 -5369 -1169 -5301
rect -1161 -5369 -1159 -5301
rect -1153 -5369 -1151 -5301
rect -1137 -5369 -1135 -5301
rect -1129 -5334 -1127 -5301
rect -1119 -5334 -1117 -5301
rect -1129 -5336 -1117 -5334
rect -1129 -5369 -1127 -5336
rect -1119 -5369 -1117 -5336
rect -1111 -5369 -1109 -5301
rect -1095 -5369 -1093 -5301
rect -1087 -5369 -1085 -5301
rect -1077 -5369 -1075 -5301
rect -1069 -5369 -1067 -5301
rect -1053 -5369 -1051 -5301
rect -1045 -5369 -1043 -5301
rect -930 -5369 -928 -5301
rect -920 -5369 -918 -5301
rect -904 -5369 -902 -5301
rect -896 -5369 -894 -5301
rect -880 -5369 -878 -5301
rect -872 -5369 -870 -5301
rect -862 -5369 -860 -5301
rect -854 -5369 -852 -5301
rect -838 -5369 -836 -5301
rect -830 -5334 -828 -5301
rect -820 -5334 -818 -5301
rect -830 -5336 -818 -5334
rect -830 -5369 -828 -5336
rect -820 -5369 -818 -5336
rect -812 -5369 -810 -5301
rect -796 -5369 -794 -5301
rect -788 -5369 -786 -5301
rect -778 -5369 -776 -5301
rect -770 -5369 -768 -5301
rect -754 -5369 -752 -5301
rect -746 -5369 -744 -5301
rect -572 -5369 -570 -5301
rect -562 -5369 -560 -5301
rect -546 -5369 -544 -5301
rect -538 -5369 -536 -5301
rect -522 -5369 -520 -5301
rect -514 -5369 -512 -5301
rect -504 -5369 -502 -5301
rect -496 -5369 -494 -5301
rect -480 -5369 -478 -5301
rect -472 -5334 -470 -5301
rect -462 -5334 -460 -5301
rect -472 -5336 -460 -5334
rect -472 -5369 -470 -5336
rect -462 -5369 -460 -5336
rect -454 -5369 -452 -5301
rect -438 -5369 -436 -5301
rect -430 -5369 -428 -5301
rect -420 -5369 -418 -5301
rect -412 -5369 -410 -5301
rect -396 -5369 -394 -5301
rect -388 -5369 -386 -5301
rect -214 -5369 -212 -5301
rect -204 -5369 -202 -5301
rect -188 -5369 -186 -5301
rect -180 -5369 -178 -5301
rect -164 -5369 -162 -5301
rect -156 -5369 -154 -5301
rect -146 -5369 -144 -5301
rect -138 -5369 -136 -5301
rect -122 -5369 -120 -5301
rect -114 -5334 -112 -5301
rect -104 -5334 -102 -5301
rect -114 -5336 -102 -5334
rect -114 -5369 -112 -5336
rect -104 -5369 -102 -5336
rect -96 -5369 -94 -5301
rect -80 -5369 -78 -5301
rect -72 -5369 -70 -5301
rect -62 -5369 -60 -5301
rect -54 -5369 -52 -5301
rect -38 -5369 -36 -5301
rect -30 -5369 -28 -5301
rect 144 -5369 146 -5301
rect 154 -5369 156 -5301
rect 170 -5369 172 -5301
rect 178 -5369 180 -5301
rect 194 -5369 196 -5301
rect 202 -5369 204 -5301
rect 212 -5369 214 -5301
rect 220 -5369 222 -5301
rect 236 -5369 238 -5301
rect 244 -5334 246 -5301
rect 254 -5334 256 -5301
rect 244 -5336 256 -5334
rect 244 -5369 246 -5336
rect 254 -5369 256 -5336
rect 262 -5369 264 -5301
rect 278 -5369 280 -5301
rect 286 -5369 288 -5301
rect 296 -5369 298 -5301
rect 304 -5369 306 -5301
rect 320 -5369 322 -5301
rect 328 -5369 330 -5301
rect 500 -5369 502 -5301
rect 510 -5369 512 -5301
rect 526 -5369 528 -5301
rect 534 -5369 536 -5301
rect 550 -5369 552 -5301
rect 558 -5369 560 -5301
rect 568 -5369 570 -5301
rect 576 -5369 578 -5301
rect 592 -5369 594 -5301
rect 600 -5334 602 -5301
rect 610 -5334 612 -5301
rect 600 -5336 612 -5334
rect 600 -5369 602 -5336
rect 610 -5369 612 -5336
rect 618 -5369 620 -5301
rect 634 -5369 636 -5301
rect 642 -5369 644 -5301
rect 652 -5369 654 -5301
rect 660 -5369 662 -5301
rect 676 -5369 678 -5301
rect 684 -5369 686 -5301
rect 858 -5369 860 -5301
rect 868 -5369 870 -5301
rect 884 -5369 886 -5301
rect 892 -5369 894 -5301
rect 908 -5369 910 -5301
rect 916 -5369 918 -5301
rect 926 -5369 928 -5301
rect 934 -5369 936 -5301
rect 950 -5369 952 -5301
rect 958 -5334 960 -5301
rect 968 -5334 970 -5301
rect 958 -5336 970 -5334
rect 958 -5369 960 -5336
rect 968 -5369 970 -5336
rect 976 -5369 978 -5301
rect 992 -5369 994 -5301
rect 1000 -5369 1002 -5301
rect 1010 -5369 1012 -5301
rect 1018 -5369 1020 -5301
rect 1034 -5369 1036 -5301
rect 1042 -5369 1044 -5301
rect 1216 -5369 1218 -5301
rect 1226 -5369 1228 -5301
rect 1242 -5369 1244 -5301
rect 1250 -5369 1252 -5301
rect 1266 -5369 1268 -5301
rect 1274 -5369 1276 -5301
rect 1284 -5369 1286 -5301
rect 1292 -5369 1294 -5301
rect 1308 -5369 1310 -5301
rect 1316 -5334 1318 -5301
rect 1326 -5334 1328 -5301
rect 1316 -5336 1328 -5334
rect 1316 -5369 1318 -5336
rect 1326 -5369 1328 -5336
rect 1334 -5369 1336 -5301
rect 1350 -5369 1352 -5301
rect 1358 -5369 1360 -5301
rect 1368 -5369 1370 -5301
rect 1376 -5369 1378 -5301
rect 1392 -5369 1394 -5301
rect 1400 -5369 1402 -5301
rect -1805 -5375 -1803 -5373
rect -1795 -5375 -1793 -5373
rect -1779 -5375 -1777 -5373
rect -1771 -5375 -1769 -5373
rect -1755 -5375 -1753 -5373
rect -1747 -5375 -1745 -5373
rect -1737 -5375 -1735 -5373
rect -1729 -5375 -1727 -5373
rect -1713 -5375 -1711 -5373
rect -1705 -5375 -1703 -5373
rect -1695 -5375 -1693 -5373
rect -1687 -5375 -1685 -5373
rect -1671 -5375 -1669 -5373
rect -1663 -5375 -1661 -5373
rect -1653 -5375 -1651 -5373
rect -1645 -5375 -1643 -5373
rect -1629 -5375 -1627 -5373
rect -1621 -5375 -1619 -5373
rect -1542 -5375 -1540 -5373
rect -1532 -5375 -1530 -5373
rect -1516 -5375 -1514 -5373
rect -1508 -5375 -1506 -5373
rect -1492 -5375 -1490 -5373
rect -1484 -5375 -1482 -5373
rect -1474 -5375 -1472 -5373
rect -1466 -5375 -1464 -5373
rect -1450 -5375 -1448 -5373
rect -1442 -5375 -1440 -5373
rect -1432 -5375 -1430 -5373
rect -1424 -5375 -1422 -5373
rect -1408 -5375 -1406 -5373
rect -1400 -5375 -1398 -5373
rect -1390 -5375 -1388 -5373
rect -1382 -5375 -1380 -5373
rect -1366 -5375 -1364 -5373
rect -1358 -5375 -1356 -5373
rect -1229 -5375 -1227 -5373
rect -1219 -5375 -1217 -5373
rect -1203 -5375 -1201 -5373
rect -1195 -5375 -1193 -5373
rect -1179 -5375 -1177 -5373
rect -1171 -5375 -1169 -5373
rect -1161 -5375 -1159 -5373
rect -1153 -5375 -1151 -5373
rect -1137 -5375 -1135 -5373
rect -1129 -5375 -1127 -5373
rect -1119 -5375 -1117 -5373
rect -1111 -5375 -1109 -5373
rect -1095 -5375 -1093 -5373
rect -1087 -5375 -1085 -5373
rect -1077 -5375 -1075 -5373
rect -1069 -5375 -1067 -5373
rect -1053 -5375 -1051 -5373
rect -1045 -5375 -1043 -5373
rect -930 -5375 -928 -5373
rect -920 -5375 -918 -5373
rect -904 -5375 -902 -5373
rect -896 -5375 -894 -5373
rect -880 -5375 -878 -5373
rect -872 -5375 -870 -5373
rect -862 -5375 -860 -5373
rect -854 -5375 -852 -5373
rect -838 -5375 -836 -5373
rect -830 -5375 -828 -5373
rect -820 -5375 -818 -5373
rect -812 -5375 -810 -5373
rect -796 -5375 -794 -5373
rect -788 -5375 -786 -5373
rect -778 -5375 -776 -5373
rect -770 -5375 -768 -5373
rect -754 -5375 -752 -5373
rect -746 -5375 -744 -5373
rect -572 -5375 -570 -5373
rect -562 -5375 -560 -5373
rect -546 -5375 -544 -5373
rect -538 -5375 -536 -5373
rect -522 -5375 -520 -5373
rect -514 -5375 -512 -5373
rect -504 -5375 -502 -5373
rect -496 -5375 -494 -5373
rect -480 -5375 -478 -5373
rect -472 -5375 -470 -5373
rect -462 -5375 -460 -5373
rect -454 -5375 -452 -5373
rect -438 -5375 -436 -5373
rect -430 -5375 -428 -5373
rect -420 -5375 -418 -5373
rect -412 -5375 -410 -5373
rect -396 -5375 -394 -5373
rect -388 -5375 -386 -5373
rect -214 -5375 -212 -5373
rect -204 -5375 -202 -5373
rect -188 -5375 -186 -5373
rect -180 -5375 -178 -5373
rect -164 -5375 -162 -5373
rect -156 -5375 -154 -5373
rect -146 -5375 -144 -5373
rect -138 -5375 -136 -5373
rect -122 -5375 -120 -5373
rect -114 -5375 -112 -5373
rect -104 -5375 -102 -5373
rect -96 -5375 -94 -5373
rect -80 -5375 -78 -5373
rect -72 -5375 -70 -5373
rect -62 -5375 -60 -5373
rect -54 -5375 -52 -5373
rect -38 -5375 -36 -5373
rect -30 -5375 -28 -5373
rect 144 -5375 146 -5373
rect 154 -5375 156 -5373
rect 170 -5375 172 -5373
rect 178 -5375 180 -5373
rect 194 -5375 196 -5373
rect 202 -5375 204 -5373
rect 212 -5375 214 -5373
rect 220 -5375 222 -5373
rect 236 -5375 238 -5373
rect 244 -5375 246 -5373
rect 254 -5375 256 -5373
rect 262 -5375 264 -5373
rect 278 -5375 280 -5373
rect 286 -5375 288 -5373
rect 296 -5375 298 -5373
rect 304 -5375 306 -5373
rect 320 -5375 322 -5373
rect 328 -5375 330 -5373
rect 500 -5375 502 -5373
rect 510 -5375 512 -5373
rect 526 -5375 528 -5373
rect 534 -5375 536 -5373
rect 550 -5375 552 -5373
rect 558 -5375 560 -5373
rect 568 -5375 570 -5373
rect 576 -5375 578 -5373
rect 592 -5375 594 -5373
rect 600 -5375 602 -5373
rect 610 -5375 612 -5373
rect 618 -5375 620 -5373
rect 634 -5375 636 -5373
rect 642 -5375 644 -5373
rect 652 -5375 654 -5373
rect 660 -5375 662 -5373
rect 676 -5375 678 -5373
rect 684 -5375 686 -5373
rect 858 -5375 860 -5373
rect 868 -5375 870 -5373
rect 884 -5375 886 -5373
rect 892 -5375 894 -5373
rect 908 -5375 910 -5373
rect 916 -5375 918 -5373
rect 926 -5375 928 -5373
rect 934 -5375 936 -5373
rect 950 -5375 952 -5373
rect 958 -5375 960 -5373
rect 968 -5375 970 -5373
rect 976 -5375 978 -5373
rect 992 -5375 994 -5373
rect 1000 -5375 1002 -5373
rect 1010 -5375 1012 -5373
rect 1018 -5375 1020 -5373
rect 1034 -5375 1036 -5373
rect 1042 -5375 1044 -5373
rect 1216 -5375 1218 -5373
rect 1226 -5375 1228 -5373
rect 1242 -5375 1244 -5373
rect 1250 -5375 1252 -5373
rect 1266 -5375 1268 -5373
rect 1274 -5375 1276 -5373
rect 1284 -5375 1286 -5373
rect 1292 -5375 1294 -5373
rect 1308 -5375 1310 -5373
rect 1316 -5375 1318 -5373
rect 1326 -5375 1328 -5373
rect 1334 -5375 1336 -5373
rect 1350 -5375 1352 -5373
rect 1358 -5375 1360 -5373
rect 1368 -5375 1370 -5373
rect 1376 -5375 1378 -5373
rect 1392 -5375 1394 -5373
rect 1400 -5375 1402 -5373
rect -1805 -5453 -1803 -5451
rect -1795 -5453 -1793 -5451
rect -1779 -5453 -1777 -5451
rect -1771 -5453 -1769 -5451
rect -1755 -5453 -1753 -5451
rect -1747 -5453 -1745 -5451
rect -1737 -5453 -1735 -5451
rect -1729 -5453 -1727 -5451
rect -1713 -5453 -1711 -5451
rect -1705 -5453 -1703 -5451
rect -1695 -5453 -1693 -5451
rect -1687 -5453 -1685 -5451
rect -1671 -5453 -1669 -5451
rect -1663 -5453 -1661 -5451
rect -1653 -5453 -1651 -5451
rect -1645 -5453 -1643 -5451
rect -1629 -5453 -1627 -5451
rect -1621 -5453 -1619 -5451
rect -1542 -5453 -1540 -5451
rect -1532 -5453 -1530 -5451
rect -1516 -5453 -1514 -5451
rect -1508 -5453 -1506 -5451
rect -1492 -5453 -1490 -5451
rect -1484 -5453 -1482 -5451
rect -1474 -5453 -1472 -5451
rect -1466 -5453 -1464 -5451
rect -1450 -5453 -1448 -5451
rect -1442 -5453 -1440 -5451
rect -1432 -5453 -1430 -5451
rect -1424 -5453 -1422 -5451
rect -1408 -5453 -1406 -5451
rect -1400 -5453 -1398 -5451
rect -1390 -5453 -1388 -5451
rect -1382 -5453 -1380 -5451
rect -1366 -5453 -1364 -5451
rect -1358 -5453 -1356 -5451
rect -1229 -5453 -1227 -5451
rect -1219 -5453 -1217 -5451
rect -1203 -5453 -1201 -5451
rect -1195 -5453 -1193 -5451
rect -1179 -5453 -1177 -5451
rect -1171 -5453 -1169 -5451
rect -1161 -5453 -1159 -5451
rect -1153 -5453 -1151 -5451
rect -1137 -5453 -1135 -5451
rect -1129 -5453 -1127 -5451
rect -1119 -5453 -1117 -5451
rect -1111 -5453 -1109 -5451
rect -1095 -5453 -1093 -5451
rect -1087 -5453 -1085 -5451
rect -1077 -5453 -1075 -5451
rect -1069 -5453 -1067 -5451
rect -1053 -5453 -1051 -5451
rect -1045 -5453 -1043 -5451
rect -930 -5453 -928 -5451
rect -920 -5453 -918 -5451
rect -904 -5453 -902 -5451
rect -896 -5453 -894 -5451
rect -880 -5453 -878 -5451
rect -872 -5453 -870 -5451
rect -862 -5453 -860 -5451
rect -854 -5453 -852 -5451
rect -838 -5453 -836 -5451
rect -830 -5453 -828 -5451
rect -820 -5453 -818 -5451
rect -812 -5453 -810 -5451
rect -796 -5453 -794 -5451
rect -788 -5453 -786 -5451
rect -778 -5453 -776 -5451
rect -770 -5453 -768 -5451
rect -754 -5453 -752 -5451
rect -746 -5453 -744 -5451
rect -572 -5453 -570 -5451
rect -562 -5453 -560 -5451
rect -546 -5453 -544 -5451
rect -538 -5453 -536 -5451
rect -522 -5453 -520 -5451
rect -514 -5453 -512 -5451
rect -504 -5453 -502 -5451
rect -496 -5453 -494 -5451
rect -480 -5453 -478 -5451
rect -472 -5453 -470 -5451
rect -462 -5453 -460 -5451
rect -454 -5453 -452 -5451
rect -438 -5453 -436 -5451
rect -430 -5453 -428 -5451
rect -420 -5453 -418 -5451
rect -412 -5453 -410 -5451
rect -396 -5453 -394 -5451
rect -388 -5453 -386 -5451
rect -214 -5453 -212 -5451
rect -204 -5453 -202 -5451
rect -188 -5453 -186 -5451
rect -180 -5453 -178 -5451
rect -164 -5453 -162 -5451
rect -156 -5453 -154 -5451
rect -146 -5453 -144 -5451
rect -138 -5453 -136 -5451
rect -122 -5453 -120 -5451
rect -114 -5453 -112 -5451
rect -104 -5453 -102 -5451
rect -96 -5453 -94 -5451
rect -80 -5453 -78 -5451
rect -72 -5453 -70 -5451
rect -62 -5453 -60 -5451
rect -54 -5453 -52 -5451
rect -38 -5453 -36 -5451
rect -30 -5453 -28 -5451
rect 144 -5453 146 -5451
rect 154 -5453 156 -5451
rect 170 -5453 172 -5451
rect 178 -5453 180 -5451
rect 194 -5453 196 -5451
rect 202 -5453 204 -5451
rect 212 -5453 214 -5451
rect 220 -5453 222 -5451
rect 236 -5453 238 -5451
rect 244 -5453 246 -5451
rect 254 -5453 256 -5451
rect 262 -5453 264 -5451
rect 278 -5453 280 -5451
rect 286 -5453 288 -5451
rect 296 -5453 298 -5451
rect 304 -5453 306 -5451
rect 320 -5453 322 -5451
rect 328 -5453 330 -5451
rect 500 -5453 502 -5451
rect 510 -5453 512 -5451
rect 526 -5453 528 -5451
rect 534 -5453 536 -5451
rect 550 -5453 552 -5451
rect 558 -5453 560 -5451
rect 568 -5453 570 -5451
rect 576 -5453 578 -5451
rect 592 -5453 594 -5451
rect 600 -5453 602 -5451
rect 610 -5453 612 -5451
rect 618 -5453 620 -5451
rect 634 -5453 636 -5451
rect 642 -5453 644 -5451
rect 652 -5453 654 -5451
rect 660 -5453 662 -5451
rect 676 -5453 678 -5451
rect 684 -5453 686 -5451
rect 858 -5453 860 -5451
rect 868 -5453 870 -5451
rect 884 -5453 886 -5451
rect 892 -5453 894 -5451
rect 908 -5453 910 -5451
rect 916 -5453 918 -5451
rect 926 -5453 928 -5451
rect 934 -5453 936 -5451
rect 950 -5453 952 -5451
rect 958 -5453 960 -5451
rect 968 -5453 970 -5451
rect 976 -5453 978 -5451
rect 992 -5453 994 -5451
rect 1000 -5453 1002 -5451
rect 1010 -5453 1012 -5451
rect 1018 -5453 1020 -5451
rect 1034 -5453 1036 -5451
rect 1042 -5453 1044 -5451
rect 1216 -5453 1218 -5451
rect 1226 -5453 1228 -5451
rect 1242 -5453 1244 -5451
rect 1250 -5453 1252 -5451
rect 1266 -5453 1268 -5451
rect 1274 -5453 1276 -5451
rect 1284 -5453 1286 -5451
rect 1292 -5453 1294 -5451
rect 1308 -5453 1310 -5451
rect 1316 -5453 1318 -5451
rect 1326 -5453 1328 -5451
rect 1334 -5453 1336 -5451
rect 1350 -5453 1352 -5451
rect 1358 -5453 1360 -5451
rect 1368 -5453 1370 -5451
rect 1376 -5453 1378 -5451
rect 1392 -5453 1394 -5451
rect 1400 -5453 1402 -5451
rect -1805 -5529 -1803 -5461
rect -1795 -5529 -1793 -5461
rect -1779 -5529 -1777 -5461
rect -1771 -5529 -1769 -5461
rect -1755 -5529 -1753 -5461
rect -1747 -5529 -1745 -5461
rect -1737 -5529 -1735 -5461
rect -1729 -5529 -1727 -5461
rect -1713 -5529 -1711 -5461
rect -1705 -5494 -1703 -5461
rect -1695 -5494 -1693 -5461
rect -1705 -5496 -1693 -5494
rect -1705 -5529 -1703 -5496
rect -1695 -5529 -1693 -5496
rect -1687 -5529 -1685 -5461
rect -1671 -5529 -1669 -5461
rect -1663 -5529 -1661 -5461
rect -1653 -5529 -1651 -5461
rect -1645 -5529 -1643 -5461
rect -1629 -5529 -1627 -5461
rect -1621 -5529 -1619 -5461
rect -1542 -5529 -1540 -5461
rect -1532 -5529 -1530 -5461
rect -1516 -5529 -1514 -5461
rect -1508 -5529 -1506 -5461
rect -1492 -5529 -1490 -5461
rect -1484 -5529 -1482 -5461
rect -1474 -5529 -1472 -5461
rect -1466 -5529 -1464 -5461
rect -1450 -5529 -1448 -5461
rect -1442 -5494 -1440 -5461
rect -1432 -5494 -1430 -5461
rect -1442 -5496 -1430 -5494
rect -1442 -5529 -1440 -5496
rect -1432 -5529 -1430 -5496
rect -1424 -5529 -1422 -5461
rect -1408 -5529 -1406 -5461
rect -1400 -5529 -1398 -5461
rect -1390 -5529 -1388 -5461
rect -1382 -5529 -1380 -5461
rect -1366 -5529 -1364 -5461
rect -1358 -5529 -1356 -5461
rect -1229 -5529 -1227 -5461
rect -1219 -5529 -1217 -5461
rect -1203 -5529 -1201 -5461
rect -1195 -5529 -1193 -5461
rect -1179 -5529 -1177 -5461
rect -1171 -5529 -1169 -5461
rect -1161 -5529 -1159 -5461
rect -1153 -5529 -1151 -5461
rect -1137 -5529 -1135 -5461
rect -1129 -5494 -1127 -5461
rect -1119 -5494 -1117 -5461
rect -1129 -5496 -1117 -5494
rect -1129 -5529 -1127 -5496
rect -1119 -5529 -1117 -5496
rect -1111 -5529 -1109 -5461
rect -1095 -5529 -1093 -5461
rect -1087 -5529 -1085 -5461
rect -1077 -5529 -1075 -5461
rect -1069 -5529 -1067 -5461
rect -1053 -5529 -1051 -5461
rect -1045 -5529 -1043 -5461
rect -930 -5529 -928 -5461
rect -920 -5529 -918 -5461
rect -904 -5529 -902 -5461
rect -896 -5529 -894 -5461
rect -880 -5529 -878 -5461
rect -872 -5529 -870 -5461
rect -862 -5529 -860 -5461
rect -854 -5529 -852 -5461
rect -838 -5529 -836 -5461
rect -830 -5494 -828 -5461
rect -820 -5494 -818 -5461
rect -830 -5496 -818 -5494
rect -830 -5529 -828 -5496
rect -820 -5529 -818 -5496
rect -812 -5529 -810 -5461
rect -796 -5529 -794 -5461
rect -788 -5529 -786 -5461
rect -778 -5529 -776 -5461
rect -770 -5529 -768 -5461
rect -754 -5529 -752 -5461
rect -746 -5529 -744 -5461
rect -572 -5529 -570 -5461
rect -562 -5529 -560 -5461
rect -546 -5529 -544 -5461
rect -538 -5529 -536 -5461
rect -522 -5529 -520 -5461
rect -514 -5529 -512 -5461
rect -504 -5529 -502 -5461
rect -496 -5529 -494 -5461
rect -480 -5529 -478 -5461
rect -472 -5494 -470 -5461
rect -462 -5494 -460 -5461
rect -472 -5496 -460 -5494
rect -472 -5529 -470 -5496
rect -462 -5529 -460 -5496
rect -454 -5529 -452 -5461
rect -438 -5529 -436 -5461
rect -430 -5529 -428 -5461
rect -420 -5529 -418 -5461
rect -412 -5529 -410 -5461
rect -396 -5529 -394 -5461
rect -388 -5529 -386 -5461
rect -214 -5529 -212 -5461
rect -204 -5529 -202 -5461
rect -188 -5529 -186 -5461
rect -180 -5529 -178 -5461
rect -164 -5529 -162 -5461
rect -156 -5529 -154 -5461
rect -146 -5529 -144 -5461
rect -138 -5529 -136 -5461
rect -122 -5529 -120 -5461
rect -114 -5494 -112 -5461
rect -104 -5494 -102 -5461
rect -114 -5496 -102 -5494
rect -114 -5529 -112 -5496
rect -104 -5529 -102 -5496
rect -96 -5529 -94 -5461
rect -80 -5529 -78 -5461
rect -72 -5529 -70 -5461
rect -62 -5529 -60 -5461
rect -54 -5529 -52 -5461
rect -38 -5529 -36 -5461
rect -30 -5529 -28 -5461
rect 144 -5529 146 -5461
rect 154 -5529 156 -5461
rect 170 -5529 172 -5461
rect 178 -5529 180 -5461
rect 194 -5529 196 -5461
rect 202 -5529 204 -5461
rect 212 -5529 214 -5461
rect 220 -5529 222 -5461
rect 236 -5529 238 -5461
rect 244 -5494 246 -5461
rect 254 -5494 256 -5461
rect 244 -5496 256 -5494
rect 244 -5529 246 -5496
rect 254 -5529 256 -5496
rect 262 -5529 264 -5461
rect 278 -5529 280 -5461
rect 286 -5529 288 -5461
rect 296 -5529 298 -5461
rect 304 -5529 306 -5461
rect 320 -5529 322 -5461
rect 328 -5529 330 -5461
rect 500 -5529 502 -5461
rect 510 -5529 512 -5461
rect 526 -5529 528 -5461
rect 534 -5529 536 -5461
rect 550 -5529 552 -5461
rect 558 -5529 560 -5461
rect 568 -5529 570 -5461
rect 576 -5529 578 -5461
rect 592 -5529 594 -5461
rect 600 -5494 602 -5461
rect 610 -5494 612 -5461
rect 600 -5496 612 -5494
rect 600 -5529 602 -5496
rect 610 -5529 612 -5496
rect 618 -5529 620 -5461
rect 634 -5529 636 -5461
rect 642 -5529 644 -5461
rect 652 -5529 654 -5461
rect 660 -5529 662 -5461
rect 676 -5529 678 -5461
rect 684 -5529 686 -5461
rect 858 -5529 860 -5461
rect 868 -5529 870 -5461
rect 884 -5529 886 -5461
rect 892 -5529 894 -5461
rect 908 -5529 910 -5461
rect 916 -5529 918 -5461
rect 926 -5529 928 -5461
rect 934 -5529 936 -5461
rect 950 -5529 952 -5461
rect 958 -5494 960 -5461
rect 968 -5494 970 -5461
rect 958 -5496 970 -5494
rect 958 -5529 960 -5496
rect 968 -5529 970 -5496
rect 976 -5529 978 -5461
rect 992 -5529 994 -5461
rect 1000 -5529 1002 -5461
rect 1010 -5529 1012 -5461
rect 1018 -5529 1020 -5461
rect 1034 -5529 1036 -5461
rect 1042 -5529 1044 -5461
rect 1216 -5529 1218 -5461
rect 1226 -5529 1228 -5461
rect 1242 -5529 1244 -5461
rect 1250 -5529 1252 -5461
rect 1266 -5529 1268 -5461
rect 1274 -5529 1276 -5461
rect 1284 -5529 1286 -5461
rect 1292 -5529 1294 -5461
rect 1308 -5529 1310 -5461
rect 1316 -5494 1318 -5461
rect 1326 -5494 1328 -5461
rect 1316 -5496 1328 -5494
rect 1316 -5529 1318 -5496
rect 1326 -5529 1328 -5496
rect 1334 -5529 1336 -5461
rect 1350 -5529 1352 -5461
rect 1358 -5529 1360 -5461
rect 1368 -5529 1370 -5461
rect 1376 -5529 1378 -5461
rect 1392 -5529 1394 -5461
rect 1400 -5529 1402 -5461
rect -1805 -5535 -1803 -5533
rect -1795 -5535 -1793 -5533
rect -1779 -5535 -1777 -5533
rect -1771 -5535 -1769 -5533
rect -1755 -5535 -1753 -5533
rect -1747 -5535 -1745 -5533
rect -1737 -5535 -1735 -5533
rect -1729 -5535 -1727 -5533
rect -1713 -5535 -1711 -5533
rect -1705 -5535 -1703 -5533
rect -1695 -5535 -1693 -5533
rect -1687 -5535 -1685 -5533
rect -1671 -5535 -1669 -5533
rect -1663 -5535 -1661 -5533
rect -1653 -5535 -1651 -5533
rect -1645 -5535 -1643 -5533
rect -1629 -5535 -1627 -5533
rect -1621 -5535 -1619 -5533
rect -1542 -5535 -1540 -5533
rect -1532 -5535 -1530 -5533
rect -1516 -5535 -1514 -5533
rect -1508 -5535 -1506 -5533
rect -1492 -5535 -1490 -5533
rect -1484 -5535 -1482 -5533
rect -1474 -5535 -1472 -5533
rect -1466 -5535 -1464 -5533
rect -1450 -5535 -1448 -5533
rect -1442 -5535 -1440 -5533
rect -1432 -5535 -1430 -5533
rect -1424 -5535 -1422 -5533
rect -1408 -5535 -1406 -5533
rect -1400 -5535 -1398 -5533
rect -1390 -5535 -1388 -5533
rect -1382 -5535 -1380 -5533
rect -1366 -5535 -1364 -5533
rect -1358 -5535 -1356 -5533
rect -1229 -5535 -1227 -5533
rect -1219 -5535 -1217 -5533
rect -1203 -5535 -1201 -5533
rect -1195 -5535 -1193 -5533
rect -1179 -5535 -1177 -5533
rect -1171 -5535 -1169 -5533
rect -1161 -5535 -1159 -5533
rect -1153 -5535 -1151 -5533
rect -1137 -5535 -1135 -5533
rect -1129 -5535 -1127 -5533
rect -1119 -5535 -1117 -5533
rect -1111 -5535 -1109 -5533
rect -1095 -5535 -1093 -5533
rect -1087 -5535 -1085 -5533
rect -1077 -5535 -1075 -5533
rect -1069 -5535 -1067 -5533
rect -1053 -5535 -1051 -5533
rect -1045 -5535 -1043 -5533
rect -930 -5535 -928 -5533
rect -920 -5535 -918 -5533
rect -904 -5535 -902 -5533
rect -896 -5535 -894 -5533
rect -880 -5535 -878 -5533
rect -872 -5535 -870 -5533
rect -862 -5535 -860 -5533
rect -854 -5535 -852 -5533
rect -838 -5535 -836 -5533
rect -830 -5535 -828 -5533
rect -820 -5535 -818 -5533
rect -812 -5535 -810 -5533
rect -796 -5535 -794 -5533
rect -788 -5535 -786 -5533
rect -778 -5535 -776 -5533
rect -770 -5535 -768 -5533
rect -754 -5535 -752 -5533
rect -746 -5535 -744 -5533
rect -572 -5535 -570 -5533
rect -562 -5535 -560 -5533
rect -546 -5535 -544 -5533
rect -538 -5535 -536 -5533
rect -522 -5535 -520 -5533
rect -514 -5535 -512 -5533
rect -504 -5535 -502 -5533
rect -496 -5535 -494 -5533
rect -480 -5535 -478 -5533
rect -472 -5535 -470 -5533
rect -462 -5535 -460 -5533
rect -454 -5535 -452 -5533
rect -438 -5535 -436 -5533
rect -430 -5535 -428 -5533
rect -420 -5535 -418 -5533
rect -412 -5535 -410 -5533
rect -396 -5535 -394 -5533
rect -388 -5535 -386 -5533
rect -214 -5535 -212 -5533
rect -204 -5535 -202 -5533
rect -188 -5535 -186 -5533
rect -180 -5535 -178 -5533
rect -164 -5535 -162 -5533
rect -156 -5535 -154 -5533
rect -146 -5535 -144 -5533
rect -138 -5535 -136 -5533
rect -122 -5535 -120 -5533
rect -114 -5535 -112 -5533
rect -104 -5535 -102 -5533
rect -96 -5535 -94 -5533
rect -80 -5535 -78 -5533
rect -72 -5535 -70 -5533
rect -62 -5535 -60 -5533
rect -54 -5535 -52 -5533
rect -38 -5535 -36 -5533
rect -30 -5535 -28 -5533
rect 144 -5535 146 -5533
rect 154 -5535 156 -5533
rect 170 -5535 172 -5533
rect 178 -5535 180 -5533
rect 194 -5535 196 -5533
rect 202 -5535 204 -5533
rect 212 -5535 214 -5533
rect 220 -5535 222 -5533
rect 236 -5535 238 -5533
rect 244 -5535 246 -5533
rect 254 -5535 256 -5533
rect 262 -5535 264 -5533
rect 278 -5535 280 -5533
rect 286 -5535 288 -5533
rect 296 -5535 298 -5533
rect 304 -5535 306 -5533
rect 320 -5535 322 -5533
rect 328 -5535 330 -5533
rect 500 -5535 502 -5533
rect 510 -5535 512 -5533
rect 526 -5535 528 -5533
rect 534 -5535 536 -5533
rect 550 -5535 552 -5533
rect 558 -5535 560 -5533
rect 568 -5535 570 -5533
rect 576 -5535 578 -5533
rect 592 -5535 594 -5533
rect 600 -5535 602 -5533
rect 610 -5535 612 -5533
rect 618 -5535 620 -5533
rect 634 -5535 636 -5533
rect 642 -5535 644 -5533
rect 652 -5535 654 -5533
rect 660 -5535 662 -5533
rect 676 -5535 678 -5533
rect 684 -5535 686 -5533
rect 858 -5535 860 -5533
rect 868 -5535 870 -5533
rect 884 -5535 886 -5533
rect 892 -5535 894 -5533
rect 908 -5535 910 -5533
rect 916 -5535 918 -5533
rect 926 -5535 928 -5533
rect 934 -5535 936 -5533
rect 950 -5535 952 -5533
rect 958 -5535 960 -5533
rect 968 -5535 970 -5533
rect 976 -5535 978 -5533
rect 992 -5535 994 -5533
rect 1000 -5535 1002 -5533
rect 1010 -5535 1012 -5533
rect 1018 -5535 1020 -5533
rect 1034 -5535 1036 -5533
rect 1042 -5535 1044 -5533
rect 1216 -5535 1218 -5533
rect 1226 -5535 1228 -5533
rect 1242 -5535 1244 -5533
rect 1250 -5535 1252 -5533
rect 1266 -5535 1268 -5533
rect 1274 -5535 1276 -5533
rect 1284 -5535 1286 -5533
rect 1292 -5535 1294 -5533
rect 1308 -5535 1310 -5533
rect 1316 -5535 1318 -5533
rect 1326 -5535 1328 -5533
rect 1334 -5535 1336 -5533
rect 1350 -5535 1352 -5533
rect 1358 -5535 1360 -5533
rect 1368 -5535 1370 -5533
rect 1376 -5535 1378 -5533
rect 1392 -5535 1394 -5533
rect 1400 -5535 1402 -5533
rect -1304 -5567 -1302 -5565
rect -1296 -5567 -1294 -5565
rect -1286 -5567 -1284 -5565
rect -930 -5567 -928 -5565
rect -922 -5567 -920 -5565
rect -912 -5567 -910 -5565
rect -572 -5567 -570 -5565
rect -564 -5567 -562 -5565
rect -554 -5567 -552 -5565
rect -214 -5567 -212 -5565
rect -206 -5567 -204 -5565
rect -196 -5567 -194 -5565
rect 144 -5567 146 -5565
rect 152 -5567 154 -5565
rect 162 -5567 164 -5565
rect 500 -5567 502 -5565
rect 508 -5567 510 -5565
rect 518 -5567 520 -5565
rect 858 -5567 860 -5565
rect 866 -5567 868 -5565
rect 876 -5567 878 -5565
rect 1216 -5567 1218 -5565
rect 1224 -5567 1226 -5565
rect 1234 -5567 1236 -5565
rect -1304 -5643 -1302 -5575
rect -1296 -5599 -1294 -5575
rect -1296 -5643 -1294 -5603
rect -1286 -5643 -1284 -5575
rect -930 -5643 -928 -5575
rect -922 -5599 -920 -5575
rect -922 -5643 -920 -5603
rect -912 -5643 -910 -5575
rect -572 -5643 -570 -5575
rect -564 -5599 -562 -5575
rect -564 -5643 -562 -5603
rect -554 -5643 -552 -5575
rect -214 -5643 -212 -5575
rect -206 -5599 -204 -5575
rect -206 -5643 -204 -5603
rect -196 -5643 -194 -5575
rect 144 -5643 146 -5575
rect 152 -5599 154 -5575
rect 152 -5643 154 -5603
rect 162 -5643 164 -5575
rect 500 -5643 502 -5575
rect 508 -5599 510 -5575
rect 508 -5643 510 -5603
rect 518 -5643 520 -5575
rect 858 -5643 860 -5575
rect 866 -5599 868 -5575
rect 866 -5643 868 -5603
rect 876 -5643 878 -5575
rect 1216 -5643 1218 -5575
rect 1224 -5599 1226 -5575
rect 1224 -5643 1226 -5603
rect 1234 -5643 1236 -5575
rect -1304 -5649 -1302 -5647
rect -1296 -5649 -1294 -5647
rect -1286 -5649 -1284 -5647
rect -930 -5649 -928 -5647
rect -922 -5649 -920 -5647
rect -912 -5649 -910 -5647
rect -572 -5649 -570 -5647
rect -564 -5649 -562 -5647
rect -554 -5649 -552 -5647
rect -214 -5649 -212 -5647
rect -206 -5649 -204 -5647
rect -196 -5649 -194 -5647
rect 144 -5649 146 -5647
rect 152 -5649 154 -5647
rect 162 -5649 164 -5647
rect 500 -5649 502 -5647
rect 508 -5649 510 -5647
rect 518 -5649 520 -5647
rect 858 -5649 860 -5647
rect 866 -5649 868 -5647
rect 876 -5649 878 -5647
rect 1216 -5649 1218 -5647
rect 1224 -5649 1226 -5647
rect 1234 -5649 1236 -5647
rect -1229 -5726 -1227 -5724
rect -1219 -5726 -1217 -5724
rect -1203 -5726 -1201 -5724
rect -1193 -5726 -1191 -5724
rect -1185 -5726 -1183 -5724
rect -1175 -5726 -1173 -5724
rect -1159 -5726 -1157 -5724
rect -1151 -5726 -1149 -5724
rect -1141 -5726 -1139 -5724
rect -930 -5726 -928 -5724
rect -920 -5726 -918 -5724
rect -904 -5726 -902 -5724
rect -894 -5726 -892 -5724
rect -878 -5726 -876 -5724
rect -868 -5726 -866 -5724
rect -860 -5726 -858 -5724
rect -850 -5726 -848 -5724
rect -834 -5726 -832 -5724
rect -826 -5726 -824 -5724
rect -816 -5726 -814 -5724
rect -800 -5726 -798 -5724
rect -790 -5726 -788 -5724
rect -782 -5726 -780 -5724
rect -772 -5726 -770 -5724
rect -756 -5726 -754 -5724
rect -748 -5726 -746 -5724
rect -732 -5726 -730 -5724
rect -716 -5726 -714 -5724
rect -708 -5726 -706 -5724
rect -698 -5726 -696 -5724
rect -572 -5726 -570 -5724
rect -562 -5726 -560 -5724
rect -546 -5726 -544 -5724
rect -536 -5726 -534 -5724
rect -520 -5726 -518 -5724
rect -510 -5726 -508 -5724
rect -502 -5726 -500 -5724
rect -492 -5726 -490 -5724
rect -476 -5726 -474 -5724
rect -468 -5726 -466 -5724
rect -458 -5726 -456 -5724
rect -442 -5726 -440 -5724
rect -432 -5726 -430 -5724
rect -424 -5726 -422 -5724
rect -414 -5726 -412 -5724
rect -398 -5726 -396 -5724
rect -390 -5726 -388 -5724
rect -374 -5726 -372 -5724
rect -358 -5726 -356 -5724
rect -350 -5726 -348 -5724
rect -340 -5726 -338 -5724
rect -214 -5726 -212 -5724
rect -204 -5726 -202 -5724
rect -188 -5726 -186 -5724
rect -178 -5726 -176 -5724
rect -162 -5726 -160 -5724
rect -152 -5726 -150 -5724
rect -144 -5726 -142 -5724
rect -134 -5726 -132 -5724
rect -118 -5726 -116 -5724
rect -110 -5726 -108 -5724
rect -100 -5726 -98 -5724
rect -84 -5726 -82 -5724
rect -74 -5726 -72 -5724
rect -66 -5726 -64 -5724
rect -56 -5726 -54 -5724
rect -40 -5726 -38 -5724
rect -32 -5726 -30 -5724
rect -16 -5726 -14 -5724
rect 0 -5726 2 -5724
rect 8 -5726 10 -5724
rect 18 -5726 20 -5724
rect 144 -5726 146 -5724
rect 154 -5726 156 -5724
rect 170 -5726 172 -5724
rect 180 -5726 182 -5724
rect 196 -5726 198 -5724
rect 206 -5726 208 -5724
rect 214 -5726 216 -5724
rect 224 -5726 226 -5724
rect 240 -5726 242 -5724
rect 248 -5726 250 -5724
rect 258 -5726 260 -5724
rect 274 -5726 276 -5724
rect 284 -5726 286 -5724
rect 292 -5726 294 -5724
rect 302 -5726 304 -5724
rect 318 -5726 320 -5724
rect 326 -5726 328 -5724
rect 342 -5726 344 -5724
rect 358 -5726 360 -5724
rect 366 -5726 368 -5724
rect 376 -5726 378 -5724
rect 500 -5726 502 -5724
rect 510 -5726 512 -5724
rect 526 -5726 528 -5724
rect 536 -5726 538 -5724
rect 552 -5726 554 -5724
rect 562 -5726 564 -5724
rect 570 -5726 572 -5724
rect 580 -5726 582 -5724
rect 596 -5726 598 -5724
rect 604 -5726 606 -5724
rect 614 -5726 616 -5724
rect 630 -5726 632 -5724
rect 640 -5726 642 -5724
rect 648 -5726 650 -5724
rect 658 -5726 660 -5724
rect 674 -5726 676 -5724
rect 682 -5726 684 -5724
rect 698 -5726 700 -5724
rect 714 -5726 716 -5724
rect 722 -5726 724 -5724
rect 732 -5726 734 -5724
rect 858 -5726 860 -5724
rect 868 -5726 870 -5724
rect 884 -5726 886 -5724
rect 894 -5726 896 -5724
rect 910 -5726 912 -5724
rect 920 -5726 922 -5724
rect 928 -5726 930 -5724
rect 938 -5726 940 -5724
rect 954 -5726 956 -5724
rect 962 -5726 964 -5724
rect 972 -5726 974 -5724
rect 988 -5726 990 -5724
rect 998 -5726 1000 -5724
rect 1006 -5726 1008 -5724
rect 1016 -5726 1018 -5724
rect 1032 -5726 1034 -5724
rect 1040 -5726 1042 -5724
rect 1056 -5726 1058 -5724
rect 1072 -5726 1074 -5724
rect 1080 -5726 1082 -5724
rect 1090 -5726 1092 -5724
rect 1216 -5726 1218 -5724
rect 1226 -5726 1228 -5724
rect 1242 -5726 1244 -5724
rect 1252 -5726 1254 -5724
rect 1268 -5726 1270 -5724
rect 1278 -5726 1280 -5724
rect 1286 -5726 1288 -5724
rect 1296 -5726 1298 -5724
rect 1312 -5726 1314 -5724
rect 1320 -5726 1322 -5724
rect 1330 -5726 1332 -5724
rect 1346 -5726 1348 -5724
rect 1356 -5726 1358 -5724
rect 1364 -5726 1366 -5724
rect 1374 -5726 1376 -5724
rect 1390 -5726 1392 -5724
rect 1398 -5726 1400 -5724
rect 1414 -5726 1416 -5724
rect 1430 -5726 1432 -5724
rect 1438 -5726 1440 -5724
rect 1448 -5726 1450 -5724
rect -1229 -5802 -1227 -5734
rect -1219 -5802 -1217 -5734
rect -1203 -5802 -1201 -5734
rect -1193 -5802 -1191 -5734
rect -1185 -5802 -1183 -5734
rect -1175 -5802 -1173 -5734
rect -1159 -5802 -1157 -5734
rect -1151 -5802 -1149 -5734
rect -1141 -5802 -1139 -5734
rect -930 -5802 -928 -5734
rect -920 -5802 -918 -5734
rect -904 -5802 -902 -5734
rect -894 -5802 -892 -5734
rect -878 -5802 -876 -5734
rect -868 -5802 -866 -5734
rect -860 -5802 -858 -5734
rect -850 -5802 -848 -5734
rect -834 -5802 -832 -5734
rect -826 -5802 -824 -5734
rect -816 -5802 -814 -5734
rect -800 -5802 -798 -5734
rect -790 -5802 -788 -5734
rect -782 -5802 -780 -5734
rect -772 -5802 -770 -5734
rect -756 -5802 -754 -5734
rect -748 -5802 -746 -5734
rect -732 -5802 -730 -5734
rect -716 -5802 -714 -5734
rect -708 -5802 -706 -5734
rect -698 -5802 -696 -5734
rect -572 -5802 -570 -5734
rect -562 -5802 -560 -5734
rect -546 -5802 -544 -5734
rect -536 -5802 -534 -5734
rect -520 -5802 -518 -5734
rect -510 -5802 -508 -5734
rect -502 -5802 -500 -5734
rect -492 -5802 -490 -5734
rect -476 -5802 -474 -5734
rect -468 -5802 -466 -5734
rect -458 -5802 -456 -5734
rect -442 -5802 -440 -5734
rect -432 -5802 -430 -5734
rect -424 -5802 -422 -5734
rect -414 -5802 -412 -5734
rect -398 -5802 -396 -5734
rect -390 -5802 -388 -5734
rect -374 -5802 -372 -5734
rect -358 -5802 -356 -5734
rect -350 -5802 -348 -5734
rect -340 -5802 -338 -5734
rect -214 -5802 -212 -5734
rect -204 -5802 -202 -5734
rect -188 -5802 -186 -5734
rect -178 -5802 -176 -5734
rect -162 -5802 -160 -5734
rect -152 -5802 -150 -5734
rect -144 -5802 -142 -5734
rect -134 -5802 -132 -5734
rect -118 -5802 -116 -5734
rect -110 -5802 -108 -5734
rect -100 -5802 -98 -5734
rect -84 -5802 -82 -5734
rect -74 -5802 -72 -5734
rect -66 -5802 -64 -5734
rect -56 -5802 -54 -5734
rect -40 -5802 -38 -5734
rect -32 -5802 -30 -5734
rect -16 -5802 -14 -5734
rect 0 -5802 2 -5734
rect 8 -5802 10 -5734
rect 18 -5802 20 -5734
rect 144 -5802 146 -5734
rect 154 -5802 156 -5734
rect 170 -5802 172 -5734
rect 180 -5802 182 -5734
rect 196 -5802 198 -5734
rect 206 -5802 208 -5734
rect 214 -5802 216 -5734
rect 224 -5802 226 -5734
rect 240 -5802 242 -5734
rect 248 -5802 250 -5734
rect 258 -5802 260 -5734
rect 274 -5802 276 -5734
rect 284 -5802 286 -5734
rect 292 -5802 294 -5734
rect 302 -5802 304 -5734
rect 318 -5802 320 -5734
rect 326 -5802 328 -5734
rect 342 -5802 344 -5734
rect 358 -5802 360 -5734
rect 366 -5802 368 -5734
rect 376 -5802 378 -5734
rect 500 -5802 502 -5734
rect 510 -5802 512 -5734
rect 526 -5802 528 -5734
rect 536 -5802 538 -5734
rect 552 -5802 554 -5734
rect 562 -5802 564 -5734
rect 570 -5802 572 -5734
rect 580 -5802 582 -5734
rect 596 -5802 598 -5734
rect 604 -5802 606 -5734
rect 614 -5802 616 -5734
rect 630 -5802 632 -5734
rect 640 -5802 642 -5734
rect 648 -5802 650 -5734
rect 658 -5802 660 -5734
rect 674 -5802 676 -5734
rect 682 -5802 684 -5734
rect 698 -5802 700 -5734
rect 714 -5802 716 -5734
rect 722 -5802 724 -5734
rect 732 -5802 734 -5734
rect 858 -5802 860 -5734
rect 868 -5802 870 -5734
rect 884 -5802 886 -5734
rect 894 -5802 896 -5734
rect 910 -5802 912 -5734
rect 920 -5802 922 -5734
rect 928 -5802 930 -5734
rect 938 -5802 940 -5734
rect 954 -5802 956 -5734
rect 962 -5802 964 -5734
rect 972 -5802 974 -5734
rect 988 -5802 990 -5734
rect 998 -5802 1000 -5734
rect 1006 -5802 1008 -5734
rect 1016 -5802 1018 -5734
rect 1032 -5802 1034 -5734
rect 1040 -5802 1042 -5734
rect 1056 -5802 1058 -5734
rect 1072 -5802 1074 -5734
rect 1080 -5802 1082 -5734
rect 1090 -5802 1092 -5734
rect 1216 -5802 1218 -5734
rect 1226 -5802 1228 -5734
rect 1242 -5802 1244 -5734
rect 1252 -5802 1254 -5734
rect 1268 -5802 1270 -5734
rect 1278 -5802 1280 -5734
rect 1286 -5802 1288 -5734
rect 1296 -5802 1298 -5734
rect 1312 -5802 1314 -5734
rect 1320 -5802 1322 -5734
rect 1330 -5802 1332 -5734
rect 1346 -5802 1348 -5734
rect 1356 -5802 1358 -5734
rect 1364 -5802 1366 -5734
rect 1374 -5802 1376 -5734
rect 1390 -5802 1392 -5734
rect 1398 -5802 1400 -5734
rect 1414 -5802 1416 -5734
rect 1430 -5802 1432 -5734
rect 1438 -5802 1440 -5734
rect 1448 -5802 1450 -5734
rect -1229 -5808 -1227 -5806
rect -1219 -5808 -1217 -5806
rect -1203 -5808 -1201 -5806
rect -1193 -5808 -1191 -5806
rect -1185 -5808 -1183 -5806
rect -1175 -5808 -1173 -5806
rect -1159 -5808 -1157 -5806
rect -1151 -5808 -1149 -5806
rect -1141 -5808 -1139 -5806
rect -930 -5808 -928 -5806
rect -920 -5808 -918 -5806
rect -904 -5808 -902 -5806
rect -894 -5808 -892 -5806
rect -878 -5808 -876 -5806
rect -868 -5808 -866 -5806
rect -860 -5808 -858 -5806
rect -850 -5808 -848 -5806
rect -834 -5808 -832 -5806
rect -826 -5808 -824 -5806
rect -816 -5808 -814 -5806
rect -800 -5808 -798 -5806
rect -790 -5808 -788 -5806
rect -782 -5808 -780 -5806
rect -772 -5808 -770 -5806
rect -756 -5808 -754 -5806
rect -748 -5808 -746 -5806
rect -732 -5808 -730 -5806
rect -716 -5808 -714 -5806
rect -708 -5808 -706 -5806
rect -698 -5808 -696 -5806
rect -572 -5808 -570 -5806
rect -562 -5808 -560 -5806
rect -546 -5808 -544 -5806
rect -536 -5808 -534 -5806
rect -520 -5808 -518 -5806
rect -510 -5808 -508 -5806
rect -502 -5808 -500 -5806
rect -492 -5808 -490 -5806
rect -476 -5808 -474 -5806
rect -468 -5808 -466 -5806
rect -458 -5808 -456 -5806
rect -442 -5808 -440 -5806
rect -432 -5808 -430 -5806
rect -424 -5808 -422 -5806
rect -414 -5808 -412 -5806
rect -398 -5808 -396 -5806
rect -390 -5808 -388 -5806
rect -374 -5808 -372 -5806
rect -358 -5808 -356 -5806
rect -350 -5808 -348 -5806
rect -340 -5808 -338 -5806
rect -214 -5808 -212 -5806
rect -204 -5808 -202 -5806
rect -188 -5808 -186 -5806
rect -178 -5808 -176 -5806
rect -162 -5808 -160 -5806
rect -152 -5808 -150 -5806
rect -144 -5808 -142 -5806
rect -134 -5808 -132 -5806
rect -118 -5808 -116 -5806
rect -110 -5808 -108 -5806
rect -100 -5808 -98 -5806
rect -84 -5808 -82 -5806
rect -74 -5808 -72 -5806
rect -66 -5808 -64 -5806
rect -56 -5808 -54 -5806
rect -40 -5808 -38 -5806
rect -32 -5808 -30 -5806
rect -16 -5808 -14 -5806
rect 0 -5808 2 -5806
rect 8 -5808 10 -5806
rect 18 -5808 20 -5806
rect 144 -5808 146 -5806
rect 154 -5808 156 -5806
rect 170 -5808 172 -5806
rect 180 -5808 182 -5806
rect 196 -5808 198 -5806
rect 206 -5808 208 -5806
rect 214 -5808 216 -5806
rect 224 -5808 226 -5806
rect 240 -5808 242 -5806
rect 248 -5808 250 -5806
rect 258 -5808 260 -5806
rect 274 -5808 276 -5806
rect 284 -5808 286 -5806
rect 292 -5808 294 -5806
rect 302 -5808 304 -5806
rect 318 -5808 320 -5806
rect 326 -5808 328 -5806
rect 342 -5808 344 -5806
rect 358 -5808 360 -5806
rect 366 -5808 368 -5806
rect 376 -5808 378 -5806
rect 500 -5808 502 -5806
rect 510 -5808 512 -5806
rect 526 -5808 528 -5806
rect 536 -5808 538 -5806
rect 552 -5808 554 -5806
rect 562 -5808 564 -5806
rect 570 -5808 572 -5806
rect 580 -5808 582 -5806
rect 596 -5808 598 -5806
rect 604 -5808 606 -5806
rect 614 -5808 616 -5806
rect 630 -5808 632 -5806
rect 640 -5808 642 -5806
rect 648 -5808 650 -5806
rect 658 -5808 660 -5806
rect 674 -5808 676 -5806
rect 682 -5808 684 -5806
rect 698 -5808 700 -5806
rect 714 -5808 716 -5806
rect 722 -5808 724 -5806
rect 732 -5808 734 -5806
rect 858 -5808 860 -5806
rect 868 -5808 870 -5806
rect 884 -5808 886 -5806
rect 894 -5808 896 -5806
rect 910 -5808 912 -5806
rect 920 -5808 922 -5806
rect 928 -5808 930 -5806
rect 938 -5808 940 -5806
rect 954 -5808 956 -5806
rect 962 -5808 964 -5806
rect 972 -5808 974 -5806
rect 988 -5808 990 -5806
rect 998 -5808 1000 -5806
rect 1006 -5808 1008 -5806
rect 1016 -5808 1018 -5806
rect 1032 -5808 1034 -5806
rect 1040 -5808 1042 -5806
rect 1056 -5808 1058 -5806
rect 1072 -5808 1074 -5806
rect 1080 -5808 1082 -5806
rect 1090 -5808 1092 -5806
rect 1216 -5808 1218 -5806
rect 1226 -5808 1228 -5806
rect 1242 -5808 1244 -5806
rect 1252 -5808 1254 -5806
rect 1268 -5808 1270 -5806
rect 1278 -5808 1280 -5806
rect 1286 -5808 1288 -5806
rect 1296 -5808 1298 -5806
rect 1312 -5808 1314 -5806
rect 1320 -5808 1322 -5806
rect 1330 -5808 1332 -5806
rect 1346 -5808 1348 -5806
rect 1356 -5808 1358 -5806
rect 1364 -5808 1366 -5806
rect 1374 -5808 1376 -5806
rect 1390 -5808 1392 -5806
rect 1398 -5808 1400 -5806
rect 1414 -5808 1416 -5806
rect 1430 -5808 1432 -5806
rect 1438 -5808 1440 -5806
rect 1448 -5808 1450 -5806
rect -1229 -5849 -1227 -5847
rect -1219 -5849 -1217 -5847
rect -1203 -5849 -1201 -5847
rect -1195 -5849 -1193 -5847
rect -1179 -5849 -1177 -5847
rect -1171 -5849 -1169 -5847
rect -1161 -5849 -1159 -5847
rect -1153 -5849 -1151 -5847
rect -1137 -5849 -1135 -5847
rect -1129 -5849 -1127 -5847
rect -1119 -5849 -1117 -5847
rect -1111 -5849 -1109 -5847
rect -1095 -5849 -1093 -5847
rect -1087 -5849 -1085 -5847
rect -1077 -5849 -1075 -5847
rect -1069 -5849 -1067 -5847
rect -1053 -5849 -1051 -5847
rect -1045 -5849 -1043 -5847
rect -930 -5849 -928 -5847
rect -920 -5849 -918 -5847
rect -904 -5849 -902 -5847
rect -896 -5849 -894 -5847
rect -880 -5849 -878 -5847
rect -872 -5849 -870 -5847
rect -862 -5849 -860 -5847
rect -854 -5849 -852 -5847
rect -838 -5849 -836 -5847
rect -830 -5849 -828 -5847
rect -820 -5849 -818 -5847
rect -812 -5849 -810 -5847
rect -796 -5849 -794 -5847
rect -788 -5849 -786 -5847
rect -778 -5849 -776 -5847
rect -770 -5849 -768 -5847
rect -754 -5849 -752 -5847
rect -746 -5849 -744 -5847
rect -572 -5849 -570 -5847
rect -562 -5849 -560 -5847
rect -546 -5849 -544 -5847
rect -538 -5849 -536 -5847
rect -522 -5849 -520 -5847
rect -514 -5849 -512 -5847
rect -504 -5849 -502 -5847
rect -496 -5849 -494 -5847
rect -480 -5849 -478 -5847
rect -472 -5849 -470 -5847
rect -462 -5849 -460 -5847
rect -454 -5849 -452 -5847
rect -438 -5849 -436 -5847
rect -430 -5849 -428 -5847
rect -420 -5849 -418 -5847
rect -412 -5849 -410 -5847
rect -396 -5849 -394 -5847
rect -388 -5849 -386 -5847
rect -214 -5849 -212 -5847
rect -204 -5849 -202 -5847
rect -188 -5849 -186 -5847
rect -180 -5849 -178 -5847
rect -164 -5849 -162 -5847
rect -156 -5849 -154 -5847
rect -146 -5849 -144 -5847
rect -138 -5849 -136 -5847
rect -122 -5849 -120 -5847
rect -114 -5849 -112 -5847
rect -104 -5849 -102 -5847
rect -96 -5849 -94 -5847
rect -80 -5849 -78 -5847
rect -72 -5849 -70 -5847
rect -62 -5849 -60 -5847
rect -54 -5849 -52 -5847
rect -38 -5849 -36 -5847
rect -30 -5849 -28 -5847
rect 144 -5849 146 -5847
rect 154 -5849 156 -5847
rect 170 -5849 172 -5847
rect 178 -5849 180 -5847
rect 194 -5849 196 -5847
rect 202 -5849 204 -5847
rect 212 -5849 214 -5847
rect 220 -5849 222 -5847
rect 236 -5849 238 -5847
rect 244 -5849 246 -5847
rect 254 -5849 256 -5847
rect 262 -5849 264 -5847
rect 278 -5849 280 -5847
rect 286 -5849 288 -5847
rect 296 -5849 298 -5847
rect 304 -5849 306 -5847
rect 320 -5849 322 -5847
rect 328 -5849 330 -5847
rect 500 -5849 502 -5847
rect 510 -5849 512 -5847
rect 526 -5849 528 -5847
rect 534 -5849 536 -5847
rect 550 -5849 552 -5847
rect 558 -5849 560 -5847
rect 568 -5849 570 -5847
rect 576 -5849 578 -5847
rect 592 -5849 594 -5847
rect 600 -5849 602 -5847
rect 610 -5849 612 -5847
rect 618 -5849 620 -5847
rect 634 -5849 636 -5847
rect 642 -5849 644 -5847
rect 652 -5849 654 -5847
rect 660 -5849 662 -5847
rect 676 -5849 678 -5847
rect 684 -5849 686 -5847
rect 858 -5849 860 -5847
rect 868 -5849 870 -5847
rect 884 -5849 886 -5847
rect 892 -5849 894 -5847
rect 908 -5849 910 -5847
rect 916 -5849 918 -5847
rect 926 -5849 928 -5847
rect 934 -5849 936 -5847
rect 950 -5849 952 -5847
rect 958 -5849 960 -5847
rect 968 -5849 970 -5847
rect 976 -5849 978 -5847
rect 992 -5849 994 -5847
rect 1000 -5849 1002 -5847
rect 1010 -5849 1012 -5847
rect 1018 -5849 1020 -5847
rect 1034 -5849 1036 -5847
rect 1042 -5849 1044 -5847
rect 1216 -5849 1218 -5847
rect 1226 -5849 1228 -5847
rect 1242 -5849 1244 -5847
rect 1250 -5849 1252 -5847
rect 1266 -5849 1268 -5847
rect 1274 -5849 1276 -5847
rect 1284 -5849 1286 -5847
rect 1292 -5849 1294 -5847
rect 1308 -5849 1310 -5847
rect 1316 -5849 1318 -5847
rect 1326 -5849 1328 -5847
rect 1334 -5849 1336 -5847
rect 1350 -5849 1352 -5847
rect 1358 -5849 1360 -5847
rect 1368 -5849 1370 -5847
rect 1376 -5849 1378 -5847
rect 1392 -5849 1394 -5847
rect 1400 -5849 1402 -5847
rect 1560 -5849 1562 -5847
rect 1570 -5849 1572 -5847
rect 1586 -5849 1588 -5847
rect 1594 -5849 1596 -5847
rect 1610 -5849 1612 -5847
rect 1618 -5849 1620 -5847
rect 1628 -5849 1630 -5847
rect 1636 -5849 1638 -5847
rect 1652 -5849 1654 -5847
rect 1660 -5849 1662 -5847
rect 1670 -5849 1672 -5847
rect 1678 -5849 1680 -5847
rect 1694 -5849 1696 -5847
rect 1702 -5849 1704 -5847
rect 1712 -5849 1714 -5847
rect 1720 -5849 1722 -5847
rect 1736 -5849 1738 -5847
rect 1744 -5849 1746 -5847
rect -1229 -5925 -1227 -5857
rect -1219 -5925 -1217 -5857
rect -1203 -5925 -1201 -5857
rect -1195 -5925 -1193 -5857
rect -1179 -5925 -1177 -5857
rect -1171 -5925 -1169 -5857
rect -1161 -5925 -1159 -5857
rect -1153 -5925 -1151 -5857
rect -1137 -5925 -1135 -5857
rect -1129 -5890 -1127 -5857
rect -1119 -5890 -1117 -5857
rect -1129 -5892 -1117 -5890
rect -1129 -5925 -1127 -5892
rect -1119 -5925 -1117 -5892
rect -1111 -5925 -1109 -5857
rect -1095 -5925 -1093 -5857
rect -1087 -5925 -1085 -5857
rect -1077 -5925 -1075 -5857
rect -1069 -5925 -1067 -5857
rect -1053 -5925 -1051 -5857
rect -1045 -5925 -1043 -5857
rect -930 -5925 -928 -5857
rect -920 -5925 -918 -5857
rect -904 -5925 -902 -5857
rect -896 -5925 -894 -5857
rect -880 -5925 -878 -5857
rect -872 -5925 -870 -5857
rect -862 -5925 -860 -5857
rect -854 -5925 -852 -5857
rect -838 -5925 -836 -5857
rect -830 -5890 -828 -5857
rect -820 -5890 -818 -5857
rect -830 -5892 -818 -5890
rect -830 -5925 -828 -5892
rect -820 -5925 -818 -5892
rect -812 -5925 -810 -5857
rect -796 -5925 -794 -5857
rect -788 -5925 -786 -5857
rect -778 -5925 -776 -5857
rect -770 -5925 -768 -5857
rect -754 -5925 -752 -5857
rect -746 -5925 -744 -5857
rect -572 -5925 -570 -5857
rect -562 -5925 -560 -5857
rect -546 -5925 -544 -5857
rect -538 -5925 -536 -5857
rect -522 -5925 -520 -5857
rect -514 -5925 -512 -5857
rect -504 -5925 -502 -5857
rect -496 -5925 -494 -5857
rect -480 -5925 -478 -5857
rect -472 -5890 -470 -5857
rect -462 -5890 -460 -5857
rect -472 -5892 -460 -5890
rect -472 -5925 -470 -5892
rect -462 -5925 -460 -5892
rect -454 -5925 -452 -5857
rect -438 -5925 -436 -5857
rect -430 -5925 -428 -5857
rect -420 -5925 -418 -5857
rect -412 -5925 -410 -5857
rect -396 -5925 -394 -5857
rect -388 -5925 -386 -5857
rect -214 -5925 -212 -5857
rect -204 -5925 -202 -5857
rect -188 -5925 -186 -5857
rect -180 -5925 -178 -5857
rect -164 -5925 -162 -5857
rect -156 -5925 -154 -5857
rect -146 -5925 -144 -5857
rect -138 -5925 -136 -5857
rect -122 -5925 -120 -5857
rect -114 -5890 -112 -5857
rect -104 -5890 -102 -5857
rect -114 -5892 -102 -5890
rect -114 -5925 -112 -5892
rect -104 -5925 -102 -5892
rect -96 -5925 -94 -5857
rect -80 -5925 -78 -5857
rect -72 -5925 -70 -5857
rect -62 -5925 -60 -5857
rect -54 -5925 -52 -5857
rect -38 -5925 -36 -5857
rect -30 -5925 -28 -5857
rect 144 -5925 146 -5857
rect 154 -5925 156 -5857
rect 170 -5925 172 -5857
rect 178 -5925 180 -5857
rect 194 -5925 196 -5857
rect 202 -5925 204 -5857
rect 212 -5925 214 -5857
rect 220 -5925 222 -5857
rect 236 -5925 238 -5857
rect 244 -5890 246 -5857
rect 254 -5890 256 -5857
rect 244 -5892 256 -5890
rect 244 -5925 246 -5892
rect 254 -5925 256 -5892
rect 262 -5925 264 -5857
rect 278 -5925 280 -5857
rect 286 -5925 288 -5857
rect 296 -5925 298 -5857
rect 304 -5925 306 -5857
rect 320 -5925 322 -5857
rect 328 -5925 330 -5857
rect 500 -5925 502 -5857
rect 510 -5925 512 -5857
rect 526 -5925 528 -5857
rect 534 -5925 536 -5857
rect 550 -5925 552 -5857
rect 558 -5925 560 -5857
rect 568 -5925 570 -5857
rect 576 -5925 578 -5857
rect 592 -5925 594 -5857
rect 600 -5890 602 -5857
rect 610 -5890 612 -5857
rect 600 -5892 612 -5890
rect 600 -5925 602 -5892
rect 610 -5925 612 -5892
rect 618 -5925 620 -5857
rect 634 -5925 636 -5857
rect 642 -5925 644 -5857
rect 652 -5925 654 -5857
rect 660 -5925 662 -5857
rect 676 -5925 678 -5857
rect 684 -5925 686 -5857
rect 858 -5925 860 -5857
rect 868 -5925 870 -5857
rect 884 -5925 886 -5857
rect 892 -5925 894 -5857
rect 908 -5925 910 -5857
rect 916 -5925 918 -5857
rect 926 -5925 928 -5857
rect 934 -5925 936 -5857
rect 950 -5925 952 -5857
rect 958 -5890 960 -5857
rect 968 -5890 970 -5857
rect 958 -5892 970 -5890
rect 958 -5925 960 -5892
rect 968 -5925 970 -5892
rect 976 -5925 978 -5857
rect 992 -5925 994 -5857
rect 1000 -5925 1002 -5857
rect 1010 -5925 1012 -5857
rect 1018 -5925 1020 -5857
rect 1034 -5925 1036 -5857
rect 1042 -5925 1044 -5857
rect 1216 -5925 1218 -5857
rect 1226 -5925 1228 -5857
rect 1242 -5925 1244 -5857
rect 1250 -5925 1252 -5857
rect 1266 -5925 1268 -5857
rect 1274 -5925 1276 -5857
rect 1284 -5925 1286 -5857
rect 1292 -5925 1294 -5857
rect 1308 -5925 1310 -5857
rect 1316 -5890 1318 -5857
rect 1326 -5890 1328 -5857
rect 1316 -5892 1328 -5890
rect 1316 -5925 1318 -5892
rect 1326 -5925 1328 -5892
rect 1334 -5925 1336 -5857
rect 1350 -5925 1352 -5857
rect 1358 -5925 1360 -5857
rect 1368 -5925 1370 -5857
rect 1376 -5925 1378 -5857
rect 1392 -5925 1394 -5857
rect 1400 -5925 1402 -5857
rect 1560 -5925 1562 -5857
rect 1570 -5925 1572 -5857
rect 1586 -5925 1588 -5857
rect 1594 -5925 1596 -5857
rect 1610 -5925 1612 -5857
rect 1618 -5925 1620 -5857
rect 1628 -5925 1630 -5857
rect 1636 -5925 1638 -5857
rect 1652 -5925 1654 -5857
rect 1660 -5890 1662 -5857
rect 1670 -5890 1672 -5857
rect 1660 -5892 1672 -5890
rect 1660 -5925 1662 -5892
rect 1670 -5925 1672 -5892
rect 1678 -5925 1680 -5857
rect 1694 -5925 1696 -5857
rect 1702 -5925 1704 -5857
rect 1712 -5925 1714 -5857
rect 1720 -5925 1722 -5857
rect 1736 -5925 1738 -5857
rect 1744 -5925 1746 -5857
rect -1229 -5931 -1227 -5929
rect -1219 -5931 -1217 -5929
rect -1203 -5931 -1201 -5929
rect -1195 -5931 -1193 -5929
rect -1179 -5931 -1177 -5929
rect -1171 -5931 -1169 -5929
rect -1161 -5931 -1159 -5929
rect -1153 -5931 -1151 -5929
rect -1137 -5931 -1135 -5929
rect -1129 -5931 -1127 -5929
rect -1119 -5931 -1117 -5929
rect -1111 -5931 -1109 -5929
rect -1095 -5931 -1093 -5929
rect -1087 -5931 -1085 -5929
rect -1077 -5931 -1075 -5929
rect -1069 -5931 -1067 -5929
rect -1053 -5931 -1051 -5929
rect -1045 -5931 -1043 -5929
rect -930 -5931 -928 -5929
rect -920 -5931 -918 -5929
rect -904 -5931 -902 -5929
rect -896 -5931 -894 -5929
rect -880 -5931 -878 -5929
rect -872 -5931 -870 -5929
rect -862 -5931 -860 -5929
rect -854 -5931 -852 -5929
rect -838 -5931 -836 -5929
rect -830 -5931 -828 -5929
rect -820 -5931 -818 -5929
rect -812 -5931 -810 -5929
rect -796 -5931 -794 -5929
rect -788 -5931 -786 -5929
rect -778 -5931 -776 -5929
rect -770 -5931 -768 -5929
rect -754 -5931 -752 -5929
rect -746 -5931 -744 -5929
rect -572 -5931 -570 -5929
rect -562 -5931 -560 -5929
rect -546 -5931 -544 -5929
rect -538 -5931 -536 -5929
rect -522 -5931 -520 -5929
rect -514 -5931 -512 -5929
rect -504 -5931 -502 -5929
rect -496 -5931 -494 -5929
rect -480 -5931 -478 -5929
rect -472 -5931 -470 -5929
rect -462 -5931 -460 -5929
rect -454 -5931 -452 -5929
rect -438 -5931 -436 -5929
rect -430 -5931 -428 -5929
rect -420 -5931 -418 -5929
rect -412 -5931 -410 -5929
rect -396 -5931 -394 -5929
rect -388 -5931 -386 -5929
rect -214 -5931 -212 -5929
rect -204 -5931 -202 -5929
rect -188 -5931 -186 -5929
rect -180 -5931 -178 -5929
rect -164 -5931 -162 -5929
rect -156 -5931 -154 -5929
rect -146 -5931 -144 -5929
rect -138 -5931 -136 -5929
rect -122 -5931 -120 -5929
rect -114 -5931 -112 -5929
rect -104 -5931 -102 -5929
rect -96 -5931 -94 -5929
rect -80 -5931 -78 -5929
rect -72 -5931 -70 -5929
rect -62 -5931 -60 -5929
rect -54 -5931 -52 -5929
rect -38 -5931 -36 -5929
rect -30 -5931 -28 -5929
rect 144 -5931 146 -5929
rect 154 -5931 156 -5929
rect 170 -5931 172 -5929
rect 178 -5931 180 -5929
rect 194 -5931 196 -5929
rect 202 -5931 204 -5929
rect 212 -5931 214 -5929
rect 220 -5931 222 -5929
rect 236 -5931 238 -5929
rect 244 -5931 246 -5929
rect 254 -5931 256 -5929
rect 262 -5931 264 -5929
rect 278 -5931 280 -5929
rect 286 -5931 288 -5929
rect 296 -5931 298 -5929
rect 304 -5931 306 -5929
rect 320 -5931 322 -5929
rect 328 -5931 330 -5929
rect 500 -5931 502 -5929
rect 510 -5931 512 -5929
rect 526 -5931 528 -5929
rect 534 -5931 536 -5929
rect 550 -5931 552 -5929
rect 558 -5931 560 -5929
rect 568 -5931 570 -5929
rect 576 -5931 578 -5929
rect 592 -5931 594 -5929
rect 600 -5931 602 -5929
rect 610 -5931 612 -5929
rect 618 -5931 620 -5929
rect 634 -5931 636 -5929
rect 642 -5931 644 -5929
rect 652 -5931 654 -5929
rect 660 -5931 662 -5929
rect 676 -5931 678 -5929
rect 684 -5931 686 -5929
rect 858 -5931 860 -5929
rect 868 -5931 870 -5929
rect 884 -5931 886 -5929
rect 892 -5931 894 -5929
rect 908 -5931 910 -5929
rect 916 -5931 918 -5929
rect 926 -5931 928 -5929
rect 934 -5931 936 -5929
rect 950 -5931 952 -5929
rect 958 -5931 960 -5929
rect 968 -5931 970 -5929
rect 976 -5931 978 -5929
rect 992 -5931 994 -5929
rect 1000 -5931 1002 -5929
rect 1010 -5931 1012 -5929
rect 1018 -5931 1020 -5929
rect 1034 -5931 1036 -5929
rect 1042 -5931 1044 -5929
rect 1216 -5931 1218 -5929
rect 1226 -5931 1228 -5929
rect 1242 -5931 1244 -5929
rect 1250 -5931 1252 -5929
rect 1266 -5931 1268 -5929
rect 1274 -5931 1276 -5929
rect 1284 -5931 1286 -5929
rect 1292 -5931 1294 -5929
rect 1308 -5931 1310 -5929
rect 1316 -5931 1318 -5929
rect 1326 -5931 1328 -5929
rect 1334 -5931 1336 -5929
rect 1350 -5931 1352 -5929
rect 1358 -5931 1360 -5929
rect 1368 -5931 1370 -5929
rect 1376 -5931 1378 -5929
rect 1392 -5931 1394 -5929
rect 1400 -5931 1402 -5929
rect 1560 -5931 1562 -5929
rect 1570 -5931 1572 -5929
rect 1586 -5931 1588 -5929
rect 1594 -5931 1596 -5929
rect 1610 -5931 1612 -5929
rect 1618 -5931 1620 -5929
rect 1628 -5931 1630 -5929
rect 1636 -5931 1638 -5929
rect 1652 -5931 1654 -5929
rect 1660 -5931 1662 -5929
rect 1670 -5931 1672 -5929
rect 1678 -5931 1680 -5929
rect 1694 -5931 1696 -5929
rect 1702 -5931 1704 -5929
rect 1712 -5931 1714 -5929
rect 1720 -5931 1722 -5929
rect 1736 -5931 1738 -5929
rect 1744 -5931 1746 -5929
<< ndiffusion >>
rect -1303 -868 -1302 -864
rect -1300 -868 -1294 -864
rect -1292 -868 -1290 -864
rect -1286 -868 -1284 -864
rect -1282 -868 -1281 -864
rect -932 -868 -931 -864
rect -929 -868 -923 -864
rect -921 -868 -919 -864
rect -915 -868 -913 -864
rect -911 -868 -910 -864
rect -573 -868 -572 -864
rect -570 -868 -564 -864
rect -562 -868 -560 -864
rect -556 -868 -554 -864
rect -552 -868 -551 -864
rect -215 -868 -214 -864
rect -212 -868 -206 -864
rect -204 -868 -202 -864
rect -198 -868 -196 -864
rect -194 -868 -193 -864
rect 142 -868 143 -864
rect 145 -868 151 -864
rect 153 -868 155 -864
rect 159 -868 161 -864
rect 163 -868 164 -864
rect 499 -868 500 -864
rect 502 -868 508 -864
rect 510 -868 512 -864
rect 516 -868 518 -864
rect 520 -868 521 -864
rect 857 -868 858 -864
rect 860 -868 866 -864
rect 868 -868 870 -864
rect 874 -868 876 -864
rect 878 -868 879 -864
rect 1215 -868 1216 -864
rect 1218 -868 1224 -864
rect 1226 -868 1228 -864
rect 1232 -868 1234 -864
rect 1236 -868 1237 -864
rect -1226 -1102 -1225 -1098
rect -1223 -1102 -1221 -1098
rect -1217 -1102 -1215 -1098
rect -1213 -1102 -1212 -1098
rect -1200 -1102 -1199 -1098
rect -1197 -1102 -1191 -1098
rect -1189 -1102 -1188 -1098
rect -1176 -1102 -1175 -1098
rect -1173 -1102 -1167 -1098
rect -1165 -1102 -1163 -1098
rect -1159 -1102 -1157 -1098
rect -1155 -1102 -1149 -1098
rect -1147 -1102 -1146 -1098
rect -1134 -1102 -1133 -1098
rect -1131 -1102 -1125 -1098
rect -1123 -1102 -1121 -1098
rect -1117 -1102 -1115 -1098
rect -1113 -1102 -1107 -1098
rect -1105 -1102 -1104 -1098
rect -1092 -1102 -1091 -1098
rect -1089 -1102 -1083 -1098
rect -1081 -1102 -1079 -1098
rect -1075 -1102 -1073 -1098
rect -1071 -1102 -1065 -1098
rect -1063 -1102 -1062 -1098
rect -1050 -1102 -1049 -1098
rect -1047 -1102 -1041 -1098
rect -1039 -1102 -1038 -1098
rect -931 -1102 -930 -1098
rect -928 -1102 -926 -1098
rect -922 -1102 -920 -1098
rect -918 -1102 -917 -1098
rect -905 -1102 -904 -1098
rect -902 -1102 -896 -1098
rect -894 -1102 -893 -1098
rect -881 -1102 -880 -1098
rect -878 -1102 -872 -1098
rect -870 -1102 -868 -1098
rect -864 -1102 -862 -1098
rect -860 -1102 -854 -1098
rect -852 -1102 -851 -1098
rect -839 -1102 -838 -1098
rect -836 -1102 -830 -1098
rect -828 -1102 -826 -1098
rect -822 -1102 -820 -1098
rect -818 -1102 -812 -1098
rect -810 -1102 -809 -1098
rect -797 -1102 -796 -1098
rect -794 -1102 -788 -1098
rect -786 -1102 -784 -1098
rect -780 -1102 -778 -1098
rect -776 -1102 -770 -1098
rect -768 -1102 -767 -1098
rect -755 -1102 -754 -1098
rect -752 -1102 -746 -1098
rect -744 -1102 -743 -1098
rect -573 -1102 -572 -1098
rect -570 -1102 -568 -1098
rect -564 -1102 -562 -1098
rect -560 -1102 -559 -1098
rect -547 -1102 -546 -1098
rect -544 -1102 -538 -1098
rect -536 -1102 -535 -1098
rect -523 -1102 -522 -1098
rect -520 -1102 -514 -1098
rect -512 -1102 -510 -1098
rect -506 -1102 -504 -1098
rect -502 -1102 -496 -1098
rect -494 -1102 -493 -1098
rect -481 -1102 -480 -1098
rect -478 -1102 -472 -1098
rect -470 -1102 -468 -1098
rect -464 -1102 -462 -1098
rect -460 -1102 -454 -1098
rect -452 -1102 -451 -1098
rect -439 -1102 -438 -1098
rect -436 -1102 -430 -1098
rect -428 -1102 -426 -1098
rect -422 -1102 -420 -1098
rect -418 -1102 -412 -1098
rect -410 -1102 -409 -1098
rect -397 -1102 -396 -1098
rect -394 -1102 -388 -1098
rect -386 -1102 -385 -1098
rect -215 -1102 -214 -1098
rect -212 -1102 -210 -1098
rect -206 -1102 -204 -1098
rect -202 -1102 -201 -1098
rect -189 -1102 -188 -1098
rect -186 -1102 -180 -1098
rect -178 -1102 -177 -1098
rect -165 -1102 -164 -1098
rect -162 -1102 -156 -1098
rect -154 -1102 -152 -1098
rect -148 -1102 -146 -1098
rect -144 -1102 -138 -1098
rect -136 -1102 -135 -1098
rect -123 -1102 -122 -1098
rect -120 -1102 -114 -1098
rect -112 -1102 -110 -1098
rect -106 -1102 -104 -1098
rect -102 -1102 -96 -1098
rect -94 -1102 -93 -1098
rect -81 -1102 -80 -1098
rect -78 -1102 -72 -1098
rect -70 -1102 -68 -1098
rect -64 -1102 -62 -1098
rect -60 -1102 -54 -1098
rect -52 -1102 -51 -1098
rect -39 -1102 -38 -1098
rect -36 -1102 -30 -1098
rect -28 -1102 -27 -1098
rect 143 -1102 144 -1098
rect 146 -1102 148 -1098
rect 152 -1102 154 -1098
rect 156 -1102 157 -1098
rect 169 -1102 170 -1098
rect 172 -1102 178 -1098
rect 180 -1102 181 -1098
rect 193 -1102 194 -1098
rect 196 -1102 202 -1098
rect 204 -1102 206 -1098
rect 210 -1102 212 -1098
rect 214 -1102 220 -1098
rect 222 -1102 223 -1098
rect 235 -1102 236 -1098
rect 238 -1102 244 -1098
rect 246 -1102 248 -1098
rect 252 -1102 254 -1098
rect 256 -1102 262 -1098
rect 264 -1102 265 -1098
rect 277 -1102 278 -1098
rect 280 -1102 286 -1098
rect 288 -1102 290 -1098
rect 294 -1102 296 -1098
rect 298 -1102 304 -1098
rect 306 -1102 307 -1098
rect 319 -1102 320 -1098
rect 322 -1102 328 -1098
rect 330 -1102 331 -1098
rect 499 -1102 500 -1098
rect 502 -1102 504 -1098
rect 508 -1102 510 -1098
rect 512 -1102 513 -1098
rect 525 -1102 526 -1098
rect 528 -1102 534 -1098
rect 536 -1102 537 -1098
rect 549 -1102 550 -1098
rect 552 -1102 558 -1098
rect 560 -1102 562 -1098
rect 566 -1102 568 -1098
rect 570 -1102 576 -1098
rect 578 -1102 579 -1098
rect 591 -1102 592 -1098
rect 594 -1102 600 -1098
rect 602 -1102 604 -1098
rect 608 -1102 610 -1098
rect 612 -1102 618 -1098
rect 620 -1102 621 -1098
rect 633 -1102 634 -1098
rect 636 -1102 642 -1098
rect 644 -1102 646 -1098
rect 650 -1102 652 -1098
rect 654 -1102 660 -1098
rect 662 -1102 663 -1098
rect 675 -1102 676 -1098
rect 678 -1102 684 -1098
rect 686 -1102 687 -1098
rect 857 -1102 858 -1098
rect 860 -1102 862 -1098
rect 866 -1102 868 -1098
rect 870 -1102 871 -1098
rect 883 -1102 884 -1098
rect 886 -1102 892 -1098
rect 894 -1102 895 -1098
rect 907 -1102 908 -1098
rect 910 -1102 916 -1098
rect 918 -1102 920 -1098
rect 924 -1102 926 -1098
rect 928 -1102 934 -1098
rect 936 -1102 937 -1098
rect 949 -1102 950 -1098
rect 952 -1102 958 -1098
rect 960 -1102 962 -1098
rect 966 -1102 968 -1098
rect 970 -1102 976 -1098
rect 978 -1102 979 -1098
rect 991 -1102 992 -1098
rect 994 -1102 1000 -1098
rect 1002 -1102 1004 -1098
rect 1008 -1102 1010 -1098
rect 1012 -1102 1018 -1098
rect 1020 -1102 1021 -1098
rect 1033 -1102 1034 -1098
rect 1036 -1102 1042 -1098
rect 1044 -1102 1045 -1098
rect -1305 -1218 -1304 -1214
rect -1302 -1218 -1296 -1214
rect -1294 -1218 -1292 -1214
rect -1288 -1218 -1286 -1214
rect -1284 -1218 -1283 -1214
rect -931 -1218 -930 -1214
rect -928 -1218 -922 -1214
rect -920 -1218 -918 -1214
rect -914 -1218 -912 -1214
rect -910 -1218 -909 -1214
rect -573 -1218 -572 -1214
rect -570 -1218 -564 -1214
rect -562 -1218 -560 -1214
rect -556 -1218 -554 -1214
rect -552 -1218 -551 -1214
rect -215 -1218 -214 -1214
rect -212 -1218 -206 -1214
rect -204 -1218 -202 -1214
rect -198 -1218 -196 -1214
rect -194 -1218 -193 -1214
rect 143 -1218 144 -1214
rect 146 -1218 152 -1214
rect 154 -1218 156 -1214
rect 160 -1218 162 -1214
rect 164 -1218 165 -1214
rect 499 -1218 500 -1214
rect 502 -1218 508 -1214
rect 510 -1218 512 -1214
rect 516 -1218 518 -1214
rect 520 -1218 521 -1214
rect 857 -1218 858 -1214
rect 860 -1218 866 -1214
rect 868 -1218 870 -1214
rect 874 -1218 876 -1214
rect 878 -1218 879 -1214
rect 1215 -1218 1216 -1214
rect 1218 -1218 1224 -1214
rect 1226 -1218 1228 -1214
rect 1232 -1218 1234 -1214
rect 1236 -1218 1237 -1214
rect -1226 -1382 -1225 -1378
rect -1223 -1382 -1221 -1378
rect -1217 -1382 -1215 -1378
rect -1213 -1382 -1212 -1378
rect -1200 -1382 -1199 -1378
rect -1197 -1382 -1195 -1378
rect -1191 -1382 -1189 -1378
rect -1187 -1382 -1181 -1378
rect -1179 -1382 -1177 -1378
rect -1173 -1382 -1171 -1378
rect -1169 -1382 -1168 -1378
rect -1156 -1382 -1155 -1378
rect -1153 -1382 -1147 -1378
rect -1145 -1382 -1143 -1378
rect -1139 -1382 -1137 -1378
rect -1135 -1382 -1134 -1378
rect -931 -1382 -930 -1378
rect -928 -1382 -926 -1378
rect -922 -1382 -920 -1378
rect -918 -1382 -917 -1378
rect -905 -1382 -904 -1378
rect -902 -1382 -900 -1378
rect -896 -1382 -894 -1378
rect -892 -1382 -891 -1378
rect -879 -1382 -878 -1378
rect -876 -1382 -875 -1378
rect -871 -1382 -868 -1378
rect -866 -1382 -860 -1378
rect -858 -1382 -857 -1378
rect -853 -1382 -850 -1378
rect -848 -1382 -847 -1378
rect -835 -1382 -834 -1378
rect -832 -1382 -826 -1378
rect -824 -1382 -822 -1378
rect -818 -1382 -816 -1378
rect -814 -1382 -813 -1378
rect -801 -1382 -800 -1378
rect -798 -1382 -796 -1378
rect -792 -1382 -790 -1378
rect -788 -1382 -782 -1378
rect -780 -1382 -778 -1378
rect -774 -1382 -772 -1378
rect -770 -1382 -769 -1378
rect -757 -1382 -756 -1378
rect -754 -1382 -748 -1378
rect -746 -1382 -745 -1378
rect -733 -1382 -732 -1378
rect -730 -1382 -725 -1378
rect -721 -1382 -716 -1378
rect -714 -1382 -713 -1378
rect -709 -1382 -708 -1378
rect -706 -1382 -704 -1378
rect -700 -1382 -698 -1378
rect -696 -1382 -695 -1378
rect -573 -1382 -572 -1378
rect -570 -1382 -568 -1378
rect -564 -1382 -562 -1378
rect -560 -1382 -559 -1378
rect -547 -1382 -546 -1378
rect -544 -1382 -542 -1378
rect -538 -1382 -536 -1378
rect -534 -1382 -533 -1378
rect -521 -1382 -520 -1378
rect -518 -1382 -517 -1378
rect -513 -1382 -510 -1378
rect -508 -1382 -502 -1378
rect -500 -1382 -499 -1378
rect -495 -1382 -492 -1378
rect -490 -1382 -489 -1378
rect -477 -1382 -476 -1378
rect -474 -1382 -468 -1378
rect -466 -1382 -464 -1378
rect -460 -1382 -458 -1378
rect -456 -1382 -455 -1378
rect -443 -1382 -442 -1378
rect -440 -1382 -438 -1378
rect -434 -1382 -432 -1378
rect -430 -1382 -424 -1378
rect -422 -1382 -420 -1378
rect -416 -1382 -414 -1378
rect -412 -1382 -411 -1378
rect -399 -1382 -398 -1378
rect -396 -1382 -390 -1378
rect -388 -1382 -387 -1378
rect -375 -1382 -374 -1378
rect -372 -1382 -367 -1378
rect -363 -1382 -358 -1378
rect -356 -1382 -355 -1378
rect -351 -1382 -350 -1378
rect -348 -1382 -346 -1378
rect -342 -1382 -340 -1378
rect -338 -1382 -337 -1378
rect -215 -1382 -214 -1378
rect -212 -1382 -210 -1378
rect -206 -1382 -204 -1378
rect -202 -1382 -201 -1378
rect -189 -1382 -188 -1378
rect -186 -1382 -184 -1378
rect -180 -1382 -178 -1378
rect -176 -1382 -175 -1378
rect -163 -1382 -162 -1378
rect -160 -1382 -159 -1378
rect -155 -1382 -152 -1378
rect -150 -1382 -144 -1378
rect -142 -1382 -141 -1378
rect -137 -1382 -134 -1378
rect -132 -1382 -131 -1378
rect -119 -1382 -118 -1378
rect -116 -1382 -110 -1378
rect -108 -1382 -106 -1378
rect -102 -1382 -100 -1378
rect -98 -1382 -97 -1378
rect -85 -1382 -84 -1378
rect -82 -1382 -80 -1378
rect -76 -1382 -74 -1378
rect -72 -1382 -66 -1378
rect -64 -1382 -62 -1378
rect -58 -1382 -56 -1378
rect -54 -1382 -53 -1378
rect -41 -1382 -40 -1378
rect -38 -1382 -32 -1378
rect -30 -1382 -29 -1378
rect -17 -1382 -16 -1378
rect -14 -1382 -9 -1378
rect -5 -1382 0 -1378
rect 2 -1382 3 -1378
rect 7 -1382 8 -1378
rect 10 -1382 12 -1378
rect 16 -1382 18 -1378
rect 20 -1382 21 -1378
rect 143 -1382 144 -1378
rect 146 -1382 148 -1378
rect 152 -1382 154 -1378
rect 156 -1382 157 -1378
rect 169 -1382 170 -1378
rect 172 -1382 174 -1378
rect 178 -1382 180 -1378
rect 182 -1382 183 -1378
rect 195 -1382 196 -1378
rect 198 -1382 199 -1378
rect 203 -1382 206 -1378
rect 208 -1382 214 -1378
rect 216 -1382 217 -1378
rect 221 -1382 224 -1378
rect 226 -1382 227 -1378
rect 239 -1382 240 -1378
rect 242 -1382 248 -1378
rect 250 -1382 252 -1378
rect 256 -1382 258 -1378
rect 260 -1382 261 -1378
rect 273 -1382 274 -1378
rect 276 -1382 278 -1378
rect 282 -1382 284 -1378
rect 286 -1382 292 -1378
rect 294 -1382 296 -1378
rect 300 -1382 302 -1378
rect 304 -1382 305 -1378
rect 317 -1382 318 -1378
rect 320 -1382 326 -1378
rect 328 -1382 329 -1378
rect 341 -1382 342 -1378
rect 344 -1382 349 -1378
rect 353 -1382 358 -1378
rect 360 -1382 361 -1378
rect 365 -1382 366 -1378
rect 368 -1382 370 -1378
rect 374 -1382 376 -1378
rect 378 -1382 379 -1378
rect 499 -1382 500 -1378
rect 502 -1382 504 -1378
rect 508 -1382 510 -1378
rect 512 -1382 513 -1378
rect 525 -1382 526 -1378
rect 528 -1382 530 -1378
rect 534 -1382 536 -1378
rect 538 -1382 539 -1378
rect 551 -1382 552 -1378
rect 554 -1382 555 -1378
rect 559 -1382 562 -1378
rect 564 -1382 570 -1378
rect 572 -1382 573 -1378
rect 577 -1382 580 -1378
rect 582 -1382 583 -1378
rect 595 -1382 596 -1378
rect 598 -1382 604 -1378
rect 606 -1382 608 -1378
rect 612 -1382 614 -1378
rect 616 -1382 617 -1378
rect 629 -1382 630 -1378
rect 632 -1382 634 -1378
rect 638 -1382 640 -1378
rect 642 -1382 648 -1378
rect 650 -1382 652 -1378
rect 656 -1382 658 -1378
rect 660 -1382 661 -1378
rect 673 -1382 674 -1378
rect 676 -1382 682 -1378
rect 684 -1382 685 -1378
rect 697 -1382 698 -1378
rect 700 -1382 705 -1378
rect 709 -1382 714 -1378
rect 716 -1382 717 -1378
rect 721 -1382 722 -1378
rect 724 -1382 726 -1378
rect 730 -1382 732 -1378
rect 734 -1382 735 -1378
rect 857 -1382 858 -1378
rect 860 -1382 862 -1378
rect 866 -1382 868 -1378
rect 870 -1382 871 -1378
rect 883 -1382 884 -1378
rect 886 -1382 888 -1378
rect 892 -1382 894 -1378
rect 896 -1382 897 -1378
rect 909 -1382 910 -1378
rect 912 -1382 913 -1378
rect 917 -1382 920 -1378
rect 922 -1382 928 -1378
rect 930 -1382 931 -1378
rect 935 -1382 938 -1378
rect 940 -1382 941 -1378
rect 953 -1382 954 -1378
rect 956 -1382 962 -1378
rect 964 -1382 966 -1378
rect 970 -1382 972 -1378
rect 974 -1382 975 -1378
rect 987 -1382 988 -1378
rect 990 -1382 992 -1378
rect 996 -1382 998 -1378
rect 1000 -1382 1006 -1378
rect 1008 -1382 1010 -1378
rect 1014 -1382 1016 -1378
rect 1018 -1382 1019 -1378
rect 1031 -1382 1032 -1378
rect 1034 -1382 1040 -1378
rect 1042 -1382 1043 -1378
rect 1055 -1382 1056 -1378
rect 1058 -1382 1063 -1378
rect 1067 -1382 1072 -1378
rect 1074 -1382 1075 -1378
rect 1079 -1382 1080 -1378
rect 1082 -1382 1084 -1378
rect 1088 -1382 1090 -1378
rect 1092 -1382 1093 -1378
rect 1215 -1382 1216 -1378
rect 1218 -1382 1220 -1378
rect 1224 -1382 1226 -1378
rect 1228 -1382 1229 -1378
rect 1241 -1382 1242 -1378
rect 1244 -1382 1246 -1378
rect 1250 -1382 1252 -1378
rect 1254 -1382 1260 -1378
rect 1262 -1382 1264 -1378
rect 1268 -1382 1270 -1378
rect 1272 -1382 1273 -1378
rect 1285 -1382 1286 -1378
rect 1288 -1382 1294 -1378
rect 1296 -1382 1298 -1378
rect 1302 -1382 1304 -1378
rect 1306 -1382 1307 -1378
rect -1226 -1505 -1225 -1501
rect -1223 -1505 -1221 -1501
rect -1217 -1505 -1215 -1501
rect -1213 -1505 -1212 -1501
rect -1200 -1505 -1199 -1501
rect -1197 -1505 -1191 -1501
rect -1189 -1505 -1188 -1501
rect -1176 -1505 -1175 -1501
rect -1173 -1505 -1167 -1501
rect -1165 -1505 -1163 -1501
rect -1159 -1505 -1157 -1501
rect -1155 -1505 -1149 -1501
rect -1147 -1505 -1146 -1501
rect -1134 -1505 -1133 -1501
rect -1131 -1505 -1125 -1501
rect -1123 -1505 -1121 -1501
rect -1117 -1505 -1115 -1501
rect -1113 -1505 -1107 -1501
rect -1105 -1505 -1104 -1501
rect -1092 -1505 -1091 -1501
rect -1089 -1505 -1083 -1501
rect -1081 -1505 -1079 -1501
rect -1075 -1505 -1073 -1501
rect -1071 -1505 -1065 -1501
rect -1063 -1505 -1062 -1501
rect -1050 -1505 -1049 -1501
rect -1047 -1505 -1041 -1501
rect -1039 -1505 -1038 -1501
rect -931 -1505 -930 -1501
rect -928 -1505 -926 -1501
rect -922 -1505 -920 -1501
rect -918 -1505 -917 -1501
rect -905 -1505 -904 -1501
rect -902 -1505 -896 -1501
rect -894 -1505 -893 -1501
rect -881 -1505 -880 -1501
rect -878 -1505 -872 -1501
rect -870 -1505 -868 -1501
rect -864 -1505 -862 -1501
rect -860 -1505 -854 -1501
rect -852 -1505 -851 -1501
rect -839 -1505 -838 -1501
rect -836 -1505 -830 -1501
rect -828 -1505 -826 -1501
rect -822 -1505 -820 -1501
rect -818 -1505 -812 -1501
rect -810 -1505 -809 -1501
rect -797 -1505 -796 -1501
rect -794 -1505 -788 -1501
rect -786 -1505 -784 -1501
rect -780 -1505 -778 -1501
rect -776 -1505 -770 -1501
rect -768 -1505 -767 -1501
rect -755 -1505 -754 -1501
rect -752 -1505 -746 -1501
rect -744 -1505 -743 -1501
rect -573 -1505 -572 -1501
rect -570 -1505 -568 -1501
rect -564 -1505 -562 -1501
rect -560 -1505 -559 -1501
rect -547 -1505 -546 -1501
rect -544 -1505 -538 -1501
rect -536 -1505 -535 -1501
rect -523 -1505 -522 -1501
rect -520 -1505 -514 -1501
rect -512 -1505 -510 -1501
rect -506 -1505 -504 -1501
rect -502 -1505 -496 -1501
rect -494 -1505 -493 -1501
rect -481 -1505 -480 -1501
rect -478 -1505 -472 -1501
rect -470 -1505 -468 -1501
rect -464 -1505 -462 -1501
rect -460 -1505 -454 -1501
rect -452 -1505 -451 -1501
rect -439 -1505 -438 -1501
rect -436 -1505 -430 -1501
rect -428 -1505 -426 -1501
rect -422 -1505 -420 -1501
rect -418 -1505 -412 -1501
rect -410 -1505 -409 -1501
rect -397 -1505 -396 -1501
rect -394 -1505 -388 -1501
rect -386 -1505 -385 -1501
rect -215 -1505 -214 -1501
rect -212 -1505 -210 -1501
rect -206 -1505 -204 -1501
rect -202 -1505 -201 -1501
rect -189 -1505 -188 -1501
rect -186 -1505 -180 -1501
rect -178 -1505 -177 -1501
rect -165 -1505 -164 -1501
rect -162 -1505 -156 -1501
rect -154 -1505 -152 -1501
rect -148 -1505 -146 -1501
rect -144 -1505 -138 -1501
rect -136 -1505 -135 -1501
rect -123 -1505 -122 -1501
rect -120 -1505 -114 -1501
rect -112 -1505 -110 -1501
rect -106 -1505 -104 -1501
rect -102 -1505 -96 -1501
rect -94 -1505 -93 -1501
rect -81 -1505 -80 -1501
rect -78 -1505 -72 -1501
rect -70 -1505 -68 -1501
rect -64 -1505 -62 -1501
rect -60 -1505 -54 -1501
rect -52 -1505 -51 -1501
rect -39 -1505 -38 -1501
rect -36 -1505 -30 -1501
rect -28 -1505 -27 -1501
rect 143 -1505 144 -1501
rect 146 -1505 148 -1501
rect 152 -1505 154 -1501
rect 156 -1505 157 -1501
rect 169 -1505 170 -1501
rect 172 -1505 178 -1501
rect 180 -1505 181 -1501
rect 193 -1505 194 -1501
rect 196 -1505 202 -1501
rect 204 -1505 206 -1501
rect 210 -1505 212 -1501
rect 214 -1505 220 -1501
rect 222 -1505 223 -1501
rect 235 -1505 236 -1501
rect 238 -1505 244 -1501
rect 246 -1505 248 -1501
rect 252 -1505 254 -1501
rect 256 -1505 262 -1501
rect 264 -1505 265 -1501
rect 277 -1505 278 -1501
rect 280 -1505 286 -1501
rect 288 -1505 290 -1501
rect 294 -1505 296 -1501
rect 298 -1505 304 -1501
rect 306 -1505 307 -1501
rect 319 -1505 320 -1501
rect 322 -1505 328 -1501
rect 330 -1505 331 -1501
rect 499 -1505 500 -1501
rect 502 -1505 504 -1501
rect 508 -1505 510 -1501
rect 512 -1505 513 -1501
rect 525 -1505 526 -1501
rect 528 -1505 534 -1501
rect 536 -1505 537 -1501
rect 549 -1505 550 -1501
rect 552 -1505 558 -1501
rect 560 -1505 562 -1501
rect 566 -1505 568 -1501
rect 570 -1505 576 -1501
rect 578 -1505 579 -1501
rect 591 -1505 592 -1501
rect 594 -1505 600 -1501
rect 602 -1505 604 -1501
rect 608 -1505 610 -1501
rect 612 -1505 618 -1501
rect 620 -1505 621 -1501
rect 633 -1505 634 -1501
rect 636 -1505 642 -1501
rect 644 -1505 646 -1501
rect 650 -1505 652 -1501
rect 654 -1505 660 -1501
rect 662 -1505 663 -1501
rect 675 -1505 676 -1501
rect 678 -1505 684 -1501
rect 686 -1505 687 -1501
rect 857 -1505 858 -1501
rect 860 -1505 862 -1501
rect 866 -1505 868 -1501
rect 870 -1505 871 -1501
rect 883 -1505 884 -1501
rect 886 -1505 892 -1501
rect 894 -1505 895 -1501
rect 907 -1505 908 -1501
rect 910 -1505 916 -1501
rect 918 -1505 920 -1501
rect 924 -1505 926 -1501
rect 928 -1505 934 -1501
rect 936 -1505 937 -1501
rect 949 -1505 950 -1501
rect 952 -1505 958 -1501
rect 960 -1505 962 -1501
rect 966 -1505 968 -1501
rect 970 -1505 976 -1501
rect 978 -1505 979 -1501
rect 991 -1505 992 -1501
rect 994 -1505 1000 -1501
rect 1002 -1505 1004 -1501
rect 1008 -1505 1010 -1501
rect 1012 -1505 1018 -1501
rect 1020 -1505 1021 -1501
rect 1033 -1505 1034 -1501
rect 1036 -1505 1042 -1501
rect 1044 -1505 1045 -1501
rect -1226 -1676 -1225 -1672
rect -1223 -1676 -1221 -1672
rect -1217 -1676 -1215 -1672
rect -1213 -1676 -1212 -1672
rect -1200 -1676 -1199 -1672
rect -1197 -1676 -1191 -1672
rect -1189 -1676 -1188 -1672
rect -1176 -1676 -1175 -1672
rect -1173 -1676 -1167 -1672
rect -1165 -1676 -1163 -1672
rect -1159 -1676 -1157 -1672
rect -1155 -1676 -1149 -1672
rect -1147 -1676 -1146 -1672
rect -1134 -1676 -1133 -1672
rect -1131 -1676 -1125 -1672
rect -1123 -1676 -1121 -1672
rect -1117 -1676 -1115 -1672
rect -1113 -1676 -1107 -1672
rect -1105 -1676 -1104 -1672
rect -1092 -1676 -1091 -1672
rect -1089 -1676 -1083 -1672
rect -1081 -1676 -1079 -1672
rect -1075 -1676 -1073 -1672
rect -1071 -1676 -1065 -1672
rect -1063 -1676 -1062 -1672
rect -1050 -1676 -1049 -1672
rect -1047 -1676 -1041 -1672
rect -1039 -1676 -1038 -1672
rect -931 -1676 -930 -1672
rect -928 -1676 -926 -1672
rect -922 -1676 -920 -1672
rect -918 -1676 -917 -1672
rect -905 -1676 -904 -1672
rect -902 -1676 -896 -1672
rect -894 -1676 -893 -1672
rect -881 -1676 -880 -1672
rect -878 -1676 -872 -1672
rect -870 -1676 -868 -1672
rect -864 -1676 -862 -1672
rect -860 -1676 -854 -1672
rect -852 -1676 -851 -1672
rect -839 -1676 -838 -1672
rect -836 -1676 -830 -1672
rect -828 -1676 -826 -1672
rect -822 -1676 -820 -1672
rect -818 -1676 -812 -1672
rect -810 -1676 -809 -1672
rect -797 -1676 -796 -1672
rect -794 -1676 -788 -1672
rect -786 -1676 -784 -1672
rect -780 -1676 -778 -1672
rect -776 -1676 -770 -1672
rect -768 -1676 -767 -1672
rect -755 -1676 -754 -1672
rect -752 -1676 -746 -1672
rect -744 -1676 -743 -1672
rect -573 -1676 -572 -1672
rect -570 -1676 -568 -1672
rect -564 -1676 -562 -1672
rect -560 -1676 -559 -1672
rect -547 -1676 -546 -1672
rect -544 -1676 -538 -1672
rect -536 -1676 -535 -1672
rect -523 -1676 -522 -1672
rect -520 -1676 -514 -1672
rect -512 -1676 -510 -1672
rect -506 -1676 -504 -1672
rect -502 -1676 -496 -1672
rect -494 -1676 -493 -1672
rect -481 -1676 -480 -1672
rect -478 -1676 -472 -1672
rect -470 -1676 -468 -1672
rect -464 -1676 -462 -1672
rect -460 -1676 -454 -1672
rect -452 -1676 -451 -1672
rect -439 -1676 -438 -1672
rect -436 -1676 -430 -1672
rect -428 -1676 -426 -1672
rect -422 -1676 -420 -1672
rect -418 -1676 -412 -1672
rect -410 -1676 -409 -1672
rect -397 -1676 -396 -1672
rect -394 -1676 -388 -1672
rect -386 -1676 -385 -1672
rect -215 -1676 -214 -1672
rect -212 -1676 -210 -1672
rect -206 -1676 -204 -1672
rect -202 -1676 -201 -1672
rect -189 -1676 -188 -1672
rect -186 -1676 -180 -1672
rect -178 -1676 -177 -1672
rect -165 -1676 -164 -1672
rect -162 -1676 -156 -1672
rect -154 -1676 -152 -1672
rect -148 -1676 -146 -1672
rect -144 -1676 -138 -1672
rect -136 -1676 -135 -1672
rect -123 -1676 -122 -1672
rect -120 -1676 -114 -1672
rect -112 -1676 -110 -1672
rect -106 -1676 -104 -1672
rect -102 -1676 -96 -1672
rect -94 -1676 -93 -1672
rect -81 -1676 -80 -1672
rect -78 -1676 -72 -1672
rect -70 -1676 -68 -1672
rect -64 -1676 -62 -1672
rect -60 -1676 -54 -1672
rect -52 -1676 -51 -1672
rect -39 -1676 -38 -1672
rect -36 -1676 -30 -1672
rect -28 -1676 -27 -1672
rect 143 -1676 144 -1672
rect 146 -1676 148 -1672
rect 152 -1676 154 -1672
rect 156 -1676 157 -1672
rect 169 -1676 170 -1672
rect 172 -1676 178 -1672
rect 180 -1676 181 -1672
rect 193 -1676 194 -1672
rect 196 -1676 202 -1672
rect 204 -1676 206 -1672
rect 210 -1676 212 -1672
rect 214 -1676 220 -1672
rect 222 -1676 223 -1672
rect 235 -1676 236 -1672
rect 238 -1676 244 -1672
rect 246 -1676 248 -1672
rect 252 -1676 254 -1672
rect 256 -1676 262 -1672
rect 264 -1676 265 -1672
rect 277 -1676 278 -1672
rect 280 -1676 286 -1672
rect 288 -1676 290 -1672
rect 294 -1676 296 -1672
rect 298 -1676 304 -1672
rect 306 -1676 307 -1672
rect 319 -1676 320 -1672
rect 322 -1676 328 -1672
rect 330 -1676 331 -1672
rect 499 -1676 500 -1672
rect 502 -1676 504 -1672
rect 508 -1676 510 -1672
rect 512 -1676 513 -1672
rect 525 -1676 526 -1672
rect 528 -1676 534 -1672
rect 536 -1676 537 -1672
rect 549 -1676 550 -1672
rect 552 -1676 558 -1672
rect 560 -1676 562 -1672
rect 566 -1676 568 -1672
rect 570 -1676 576 -1672
rect 578 -1676 579 -1672
rect 591 -1676 592 -1672
rect 594 -1676 600 -1672
rect 602 -1676 604 -1672
rect 608 -1676 610 -1672
rect 612 -1676 618 -1672
rect 620 -1676 621 -1672
rect 633 -1676 634 -1672
rect 636 -1676 642 -1672
rect 644 -1676 646 -1672
rect 650 -1676 652 -1672
rect 654 -1676 660 -1672
rect 662 -1676 663 -1672
rect 675 -1676 676 -1672
rect 678 -1676 684 -1672
rect 686 -1676 687 -1672
rect 857 -1676 858 -1672
rect 860 -1676 862 -1672
rect 866 -1676 868 -1672
rect 870 -1676 871 -1672
rect 883 -1676 884 -1672
rect 886 -1676 892 -1672
rect 894 -1676 895 -1672
rect 907 -1676 908 -1672
rect 910 -1676 916 -1672
rect 918 -1676 920 -1672
rect 924 -1676 926 -1672
rect 928 -1676 934 -1672
rect 936 -1676 937 -1672
rect 949 -1676 950 -1672
rect 952 -1676 958 -1672
rect 960 -1676 962 -1672
rect 966 -1676 968 -1672
rect 970 -1676 976 -1672
rect 978 -1676 979 -1672
rect 991 -1676 992 -1672
rect 994 -1676 1000 -1672
rect 1002 -1676 1004 -1672
rect 1008 -1676 1010 -1672
rect 1012 -1676 1018 -1672
rect 1020 -1676 1021 -1672
rect 1033 -1676 1034 -1672
rect 1036 -1676 1042 -1672
rect 1044 -1676 1045 -1672
rect 1215 -1676 1216 -1672
rect 1218 -1676 1220 -1672
rect 1224 -1676 1226 -1672
rect 1228 -1676 1229 -1672
rect 1241 -1676 1242 -1672
rect 1244 -1676 1250 -1672
rect 1252 -1676 1253 -1672
rect 1265 -1676 1266 -1672
rect 1268 -1676 1274 -1672
rect 1276 -1676 1278 -1672
rect 1282 -1676 1284 -1672
rect 1286 -1676 1292 -1672
rect 1294 -1676 1295 -1672
rect 1307 -1676 1308 -1672
rect 1310 -1676 1316 -1672
rect 1318 -1676 1320 -1672
rect 1324 -1676 1326 -1672
rect 1328 -1676 1334 -1672
rect 1336 -1676 1337 -1672
rect 1349 -1676 1350 -1672
rect 1352 -1676 1358 -1672
rect 1360 -1676 1362 -1672
rect 1366 -1676 1368 -1672
rect 1370 -1676 1376 -1672
rect 1378 -1676 1379 -1672
rect 1391 -1676 1392 -1672
rect 1394 -1676 1400 -1672
rect 1402 -1676 1403 -1672
rect -1555 -1847 -1554 -1843
rect -1552 -1847 -1550 -1843
rect -1546 -1847 -1544 -1843
rect -1542 -1847 -1541 -1843
rect -1529 -1847 -1528 -1843
rect -1526 -1847 -1520 -1843
rect -1518 -1847 -1517 -1843
rect -1505 -1847 -1504 -1843
rect -1502 -1847 -1496 -1843
rect -1494 -1847 -1492 -1843
rect -1488 -1847 -1486 -1843
rect -1484 -1847 -1478 -1843
rect -1476 -1847 -1475 -1843
rect -1463 -1847 -1462 -1843
rect -1460 -1847 -1454 -1843
rect -1452 -1847 -1450 -1843
rect -1446 -1847 -1444 -1843
rect -1442 -1847 -1436 -1843
rect -1434 -1847 -1433 -1843
rect -1421 -1847 -1420 -1843
rect -1418 -1847 -1412 -1843
rect -1410 -1847 -1408 -1843
rect -1404 -1847 -1402 -1843
rect -1400 -1847 -1394 -1843
rect -1392 -1847 -1391 -1843
rect -1379 -1847 -1378 -1843
rect -1376 -1847 -1370 -1843
rect -1368 -1847 -1367 -1843
rect -1226 -1847 -1225 -1843
rect -1223 -1847 -1221 -1843
rect -1217 -1847 -1215 -1843
rect -1213 -1847 -1212 -1843
rect -1200 -1847 -1199 -1843
rect -1197 -1847 -1191 -1843
rect -1189 -1847 -1188 -1843
rect -1176 -1847 -1175 -1843
rect -1173 -1847 -1167 -1843
rect -1165 -1847 -1163 -1843
rect -1159 -1847 -1157 -1843
rect -1155 -1847 -1149 -1843
rect -1147 -1847 -1146 -1843
rect -1134 -1847 -1133 -1843
rect -1131 -1847 -1125 -1843
rect -1123 -1847 -1121 -1843
rect -1117 -1847 -1115 -1843
rect -1113 -1847 -1107 -1843
rect -1105 -1847 -1104 -1843
rect -1092 -1847 -1091 -1843
rect -1089 -1847 -1083 -1843
rect -1081 -1847 -1079 -1843
rect -1075 -1847 -1073 -1843
rect -1071 -1847 -1065 -1843
rect -1063 -1847 -1062 -1843
rect -1050 -1847 -1049 -1843
rect -1047 -1847 -1041 -1843
rect -1039 -1847 -1038 -1843
rect -931 -1847 -930 -1843
rect -928 -1847 -926 -1843
rect -922 -1847 -920 -1843
rect -918 -1847 -917 -1843
rect -905 -1847 -904 -1843
rect -902 -1847 -896 -1843
rect -894 -1847 -893 -1843
rect -881 -1847 -880 -1843
rect -878 -1847 -872 -1843
rect -870 -1847 -868 -1843
rect -864 -1847 -862 -1843
rect -860 -1847 -854 -1843
rect -852 -1847 -851 -1843
rect -839 -1847 -838 -1843
rect -836 -1847 -830 -1843
rect -828 -1847 -826 -1843
rect -822 -1847 -820 -1843
rect -818 -1847 -812 -1843
rect -810 -1847 -809 -1843
rect -797 -1847 -796 -1843
rect -794 -1847 -788 -1843
rect -786 -1847 -784 -1843
rect -780 -1847 -778 -1843
rect -776 -1847 -770 -1843
rect -768 -1847 -767 -1843
rect -755 -1847 -754 -1843
rect -752 -1847 -746 -1843
rect -744 -1847 -743 -1843
rect -573 -1847 -572 -1843
rect -570 -1847 -568 -1843
rect -564 -1847 -562 -1843
rect -560 -1847 -559 -1843
rect -547 -1847 -546 -1843
rect -544 -1847 -538 -1843
rect -536 -1847 -535 -1843
rect -523 -1847 -522 -1843
rect -520 -1847 -514 -1843
rect -512 -1847 -510 -1843
rect -506 -1847 -504 -1843
rect -502 -1847 -496 -1843
rect -494 -1847 -493 -1843
rect -481 -1847 -480 -1843
rect -478 -1847 -472 -1843
rect -470 -1847 -468 -1843
rect -464 -1847 -462 -1843
rect -460 -1847 -454 -1843
rect -452 -1847 -451 -1843
rect -439 -1847 -438 -1843
rect -436 -1847 -430 -1843
rect -428 -1847 -426 -1843
rect -422 -1847 -420 -1843
rect -418 -1847 -412 -1843
rect -410 -1847 -409 -1843
rect -397 -1847 -396 -1843
rect -394 -1847 -388 -1843
rect -386 -1847 -385 -1843
rect -215 -1847 -214 -1843
rect -212 -1847 -210 -1843
rect -206 -1847 -204 -1843
rect -202 -1847 -201 -1843
rect -189 -1847 -188 -1843
rect -186 -1847 -180 -1843
rect -178 -1847 -177 -1843
rect -165 -1847 -164 -1843
rect -162 -1847 -156 -1843
rect -154 -1847 -152 -1843
rect -148 -1847 -146 -1843
rect -144 -1847 -138 -1843
rect -136 -1847 -135 -1843
rect -123 -1847 -122 -1843
rect -120 -1847 -114 -1843
rect -112 -1847 -110 -1843
rect -106 -1847 -104 -1843
rect -102 -1847 -96 -1843
rect -94 -1847 -93 -1843
rect -81 -1847 -80 -1843
rect -78 -1847 -72 -1843
rect -70 -1847 -68 -1843
rect -64 -1847 -62 -1843
rect -60 -1847 -54 -1843
rect -52 -1847 -51 -1843
rect -39 -1847 -38 -1843
rect -36 -1847 -30 -1843
rect -28 -1847 -27 -1843
rect 143 -1847 144 -1843
rect 146 -1847 148 -1843
rect 152 -1847 154 -1843
rect 156 -1847 157 -1843
rect 169 -1847 170 -1843
rect 172 -1847 178 -1843
rect 180 -1847 181 -1843
rect 193 -1847 194 -1843
rect 196 -1847 202 -1843
rect 204 -1847 206 -1843
rect 210 -1847 212 -1843
rect 214 -1847 220 -1843
rect 222 -1847 223 -1843
rect 235 -1847 236 -1843
rect 238 -1847 244 -1843
rect 246 -1847 248 -1843
rect 252 -1847 254 -1843
rect 256 -1847 262 -1843
rect 264 -1847 265 -1843
rect 277 -1847 278 -1843
rect 280 -1847 286 -1843
rect 288 -1847 290 -1843
rect 294 -1847 296 -1843
rect 298 -1847 304 -1843
rect 306 -1847 307 -1843
rect 319 -1847 320 -1843
rect 322 -1847 328 -1843
rect 330 -1847 331 -1843
rect 499 -1847 500 -1843
rect 502 -1847 504 -1843
rect 508 -1847 510 -1843
rect 512 -1847 513 -1843
rect 525 -1847 526 -1843
rect 528 -1847 534 -1843
rect 536 -1847 537 -1843
rect 549 -1847 550 -1843
rect 552 -1847 558 -1843
rect 560 -1847 562 -1843
rect 566 -1847 568 -1843
rect 570 -1847 576 -1843
rect 578 -1847 579 -1843
rect 591 -1847 592 -1843
rect 594 -1847 600 -1843
rect 602 -1847 604 -1843
rect 608 -1847 610 -1843
rect 612 -1847 618 -1843
rect 620 -1847 621 -1843
rect 633 -1847 634 -1843
rect 636 -1847 642 -1843
rect 644 -1847 646 -1843
rect 650 -1847 652 -1843
rect 654 -1847 660 -1843
rect 662 -1847 663 -1843
rect 675 -1847 676 -1843
rect 678 -1847 684 -1843
rect 686 -1847 687 -1843
rect 857 -1847 858 -1843
rect 860 -1847 862 -1843
rect 866 -1847 868 -1843
rect 870 -1847 871 -1843
rect 883 -1847 884 -1843
rect 886 -1847 892 -1843
rect 894 -1847 895 -1843
rect 907 -1847 908 -1843
rect 910 -1847 916 -1843
rect 918 -1847 920 -1843
rect 924 -1847 926 -1843
rect 928 -1847 934 -1843
rect 936 -1847 937 -1843
rect 949 -1847 950 -1843
rect 952 -1847 958 -1843
rect 960 -1847 962 -1843
rect 966 -1847 968 -1843
rect 970 -1847 976 -1843
rect 978 -1847 979 -1843
rect 991 -1847 992 -1843
rect 994 -1847 1000 -1843
rect 1002 -1847 1004 -1843
rect 1008 -1847 1010 -1843
rect 1012 -1847 1018 -1843
rect 1020 -1847 1021 -1843
rect 1033 -1847 1034 -1843
rect 1036 -1847 1042 -1843
rect 1044 -1847 1045 -1843
rect 1215 -1847 1216 -1843
rect 1218 -1847 1220 -1843
rect 1224 -1847 1226 -1843
rect 1228 -1847 1229 -1843
rect 1241 -1847 1242 -1843
rect 1244 -1847 1250 -1843
rect 1252 -1847 1253 -1843
rect 1265 -1847 1266 -1843
rect 1268 -1847 1274 -1843
rect 1276 -1847 1278 -1843
rect 1282 -1847 1284 -1843
rect 1286 -1847 1292 -1843
rect 1294 -1847 1295 -1843
rect 1307 -1847 1308 -1843
rect 1310 -1847 1316 -1843
rect 1318 -1847 1320 -1843
rect 1324 -1847 1326 -1843
rect 1328 -1847 1334 -1843
rect 1336 -1847 1337 -1843
rect 1349 -1847 1350 -1843
rect 1352 -1847 1358 -1843
rect 1360 -1847 1362 -1843
rect 1366 -1847 1368 -1843
rect 1370 -1847 1376 -1843
rect 1378 -1847 1379 -1843
rect 1391 -1847 1392 -1843
rect 1394 -1847 1400 -1843
rect 1402 -1847 1403 -1843
rect -1305 -1954 -1304 -1950
rect -1302 -1954 -1296 -1950
rect -1294 -1954 -1292 -1950
rect -1288 -1954 -1286 -1950
rect -1284 -1954 -1283 -1950
rect -931 -1954 -930 -1950
rect -928 -1954 -922 -1950
rect -920 -1954 -918 -1950
rect -914 -1954 -912 -1950
rect -910 -1954 -909 -1950
rect -573 -1954 -572 -1950
rect -570 -1954 -564 -1950
rect -562 -1954 -560 -1950
rect -556 -1954 -554 -1950
rect -552 -1954 -551 -1950
rect -215 -1954 -214 -1950
rect -212 -1954 -206 -1950
rect -204 -1954 -202 -1950
rect -198 -1954 -196 -1950
rect -194 -1954 -193 -1950
rect 143 -1954 144 -1950
rect 146 -1954 152 -1950
rect 154 -1954 156 -1950
rect 160 -1954 162 -1950
rect 164 -1954 165 -1950
rect 499 -1954 500 -1950
rect 502 -1954 508 -1950
rect 510 -1954 512 -1950
rect 516 -1954 518 -1950
rect 520 -1954 521 -1950
rect 857 -1954 858 -1950
rect 860 -1954 866 -1950
rect 868 -1954 870 -1950
rect 874 -1954 876 -1950
rect 878 -1954 879 -1950
rect 1215 -1954 1216 -1950
rect 1218 -1954 1224 -1950
rect 1226 -1954 1228 -1950
rect 1232 -1954 1234 -1950
rect 1236 -1954 1237 -1950
rect -1230 -2113 -1229 -2109
rect -1227 -2113 -1225 -2109
rect -1221 -2113 -1219 -2109
rect -1217 -2113 -1216 -2109
rect -1204 -2113 -1203 -2109
rect -1201 -2113 -1199 -2109
rect -1195 -2113 -1193 -2109
rect -1191 -2113 -1185 -2109
rect -1183 -2113 -1181 -2109
rect -1177 -2113 -1175 -2109
rect -1173 -2113 -1172 -2109
rect -1160 -2113 -1159 -2109
rect -1157 -2113 -1151 -2109
rect -1149 -2113 -1147 -2109
rect -1143 -2113 -1141 -2109
rect -1139 -2113 -1138 -2109
rect -931 -2113 -930 -2109
rect -928 -2113 -926 -2109
rect -922 -2113 -920 -2109
rect -918 -2113 -917 -2109
rect -905 -2113 -904 -2109
rect -902 -2113 -900 -2109
rect -896 -2113 -894 -2109
rect -892 -2113 -891 -2109
rect -879 -2113 -878 -2109
rect -876 -2113 -875 -2109
rect -871 -2113 -868 -2109
rect -866 -2113 -860 -2109
rect -858 -2113 -857 -2109
rect -853 -2113 -850 -2109
rect -848 -2113 -847 -2109
rect -835 -2113 -834 -2109
rect -832 -2113 -826 -2109
rect -824 -2113 -822 -2109
rect -818 -2113 -816 -2109
rect -814 -2113 -813 -2109
rect -801 -2113 -800 -2109
rect -798 -2113 -796 -2109
rect -792 -2113 -790 -2109
rect -788 -2113 -782 -2109
rect -780 -2113 -778 -2109
rect -774 -2113 -772 -2109
rect -770 -2113 -769 -2109
rect -757 -2113 -756 -2109
rect -754 -2113 -748 -2109
rect -746 -2113 -745 -2109
rect -733 -2113 -732 -2109
rect -730 -2113 -725 -2109
rect -721 -2113 -716 -2109
rect -714 -2113 -713 -2109
rect -709 -2113 -708 -2109
rect -706 -2113 -704 -2109
rect -700 -2113 -698 -2109
rect -696 -2113 -695 -2109
rect -573 -2113 -572 -2109
rect -570 -2113 -568 -2109
rect -564 -2113 -562 -2109
rect -560 -2113 -559 -2109
rect -547 -2113 -546 -2109
rect -544 -2113 -542 -2109
rect -538 -2113 -536 -2109
rect -534 -2113 -533 -2109
rect -521 -2113 -520 -2109
rect -518 -2113 -517 -2109
rect -513 -2113 -510 -2109
rect -508 -2113 -502 -2109
rect -500 -2113 -499 -2109
rect -495 -2113 -492 -2109
rect -490 -2113 -489 -2109
rect -477 -2113 -476 -2109
rect -474 -2113 -468 -2109
rect -466 -2113 -464 -2109
rect -460 -2113 -458 -2109
rect -456 -2113 -455 -2109
rect -443 -2113 -442 -2109
rect -440 -2113 -438 -2109
rect -434 -2113 -432 -2109
rect -430 -2113 -424 -2109
rect -422 -2113 -420 -2109
rect -416 -2113 -414 -2109
rect -412 -2113 -411 -2109
rect -399 -2113 -398 -2109
rect -396 -2113 -390 -2109
rect -388 -2113 -387 -2109
rect -375 -2113 -374 -2109
rect -372 -2113 -367 -2109
rect -363 -2113 -358 -2109
rect -356 -2113 -355 -2109
rect -351 -2113 -350 -2109
rect -348 -2113 -346 -2109
rect -342 -2113 -340 -2109
rect -338 -2113 -337 -2109
rect -215 -2113 -214 -2109
rect -212 -2113 -210 -2109
rect -206 -2113 -204 -2109
rect -202 -2113 -201 -2109
rect -189 -2113 -188 -2109
rect -186 -2113 -184 -2109
rect -180 -2113 -178 -2109
rect -176 -2113 -175 -2109
rect -163 -2113 -162 -2109
rect -160 -2113 -159 -2109
rect -155 -2113 -152 -2109
rect -150 -2113 -144 -2109
rect -142 -2113 -141 -2109
rect -137 -2113 -134 -2109
rect -132 -2113 -131 -2109
rect -119 -2113 -118 -2109
rect -116 -2113 -110 -2109
rect -108 -2113 -106 -2109
rect -102 -2113 -100 -2109
rect -98 -2113 -97 -2109
rect -85 -2113 -84 -2109
rect -82 -2113 -80 -2109
rect -76 -2113 -74 -2109
rect -72 -2113 -66 -2109
rect -64 -2113 -62 -2109
rect -58 -2113 -56 -2109
rect -54 -2113 -53 -2109
rect -41 -2113 -40 -2109
rect -38 -2113 -32 -2109
rect -30 -2113 -29 -2109
rect -17 -2113 -16 -2109
rect -14 -2113 -9 -2109
rect -5 -2113 0 -2109
rect 2 -2113 3 -2109
rect 7 -2113 8 -2109
rect 10 -2113 12 -2109
rect 16 -2113 18 -2109
rect 20 -2113 21 -2109
rect 143 -2113 144 -2109
rect 146 -2113 148 -2109
rect 152 -2113 154 -2109
rect 156 -2113 157 -2109
rect 169 -2113 170 -2109
rect 172 -2113 174 -2109
rect 178 -2113 180 -2109
rect 182 -2113 183 -2109
rect 195 -2113 196 -2109
rect 198 -2113 199 -2109
rect 203 -2113 206 -2109
rect 208 -2113 214 -2109
rect 216 -2113 217 -2109
rect 221 -2113 224 -2109
rect 226 -2113 227 -2109
rect 239 -2113 240 -2109
rect 242 -2113 248 -2109
rect 250 -2113 252 -2109
rect 256 -2113 258 -2109
rect 260 -2113 261 -2109
rect 273 -2113 274 -2109
rect 276 -2113 278 -2109
rect 282 -2113 284 -2109
rect 286 -2113 292 -2109
rect 294 -2113 296 -2109
rect 300 -2113 302 -2109
rect 304 -2113 305 -2109
rect 317 -2113 318 -2109
rect 320 -2113 326 -2109
rect 328 -2113 329 -2109
rect 341 -2113 342 -2109
rect 344 -2113 349 -2109
rect 353 -2113 358 -2109
rect 360 -2113 361 -2109
rect 365 -2113 366 -2109
rect 368 -2113 370 -2109
rect 374 -2113 376 -2109
rect 378 -2113 379 -2109
rect 499 -2113 500 -2109
rect 502 -2113 504 -2109
rect 508 -2113 510 -2109
rect 512 -2113 513 -2109
rect 525 -2113 526 -2109
rect 528 -2113 530 -2109
rect 534 -2113 536 -2109
rect 538 -2113 539 -2109
rect 551 -2113 552 -2109
rect 554 -2113 555 -2109
rect 559 -2113 562 -2109
rect 564 -2113 570 -2109
rect 572 -2113 573 -2109
rect 577 -2113 580 -2109
rect 582 -2113 583 -2109
rect 595 -2113 596 -2109
rect 598 -2113 604 -2109
rect 606 -2113 608 -2109
rect 612 -2113 614 -2109
rect 616 -2113 617 -2109
rect 629 -2113 630 -2109
rect 632 -2113 634 -2109
rect 638 -2113 640 -2109
rect 642 -2113 648 -2109
rect 650 -2113 652 -2109
rect 656 -2113 658 -2109
rect 660 -2113 661 -2109
rect 673 -2113 674 -2109
rect 676 -2113 682 -2109
rect 684 -2113 685 -2109
rect 697 -2113 698 -2109
rect 700 -2113 705 -2109
rect 709 -2113 714 -2109
rect 716 -2113 717 -2109
rect 721 -2113 722 -2109
rect 724 -2113 726 -2109
rect 730 -2113 732 -2109
rect 734 -2113 735 -2109
rect 857 -2113 858 -2109
rect 860 -2113 862 -2109
rect 866 -2113 868 -2109
rect 870 -2113 871 -2109
rect 883 -2113 884 -2109
rect 886 -2113 888 -2109
rect 892 -2113 894 -2109
rect 896 -2113 897 -2109
rect 909 -2113 910 -2109
rect 912 -2113 913 -2109
rect 917 -2113 920 -2109
rect 922 -2113 928 -2109
rect 930 -2113 931 -2109
rect 935 -2113 938 -2109
rect 940 -2113 941 -2109
rect 953 -2113 954 -2109
rect 956 -2113 962 -2109
rect 964 -2113 966 -2109
rect 970 -2113 972 -2109
rect 974 -2113 975 -2109
rect 987 -2113 988 -2109
rect 990 -2113 992 -2109
rect 996 -2113 998 -2109
rect 1000 -2113 1006 -2109
rect 1008 -2113 1010 -2109
rect 1014 -2113 1016 -2109
rect 1018 -2113 1019 -2109
rect 1031 -2113 1032 -2109
rect 1034 -2113 1040 -2109
rect 1042 -2113 1043 -2109
rect 1055 -2113 1056 -2109
rect 1058 -2113 1063 -2109
rect 1067 -2113 1072 -2109
rect 1074 -2113 1075 -2109
rect 1079 -2113 1080 -2109
rect 1082 -2113 1084 -2109
rect 1088 -2113 1090 -2109
rect 1092 -2113 1093 -2109
rect 1215 -2113 1216 -2109
rect 1218 -2113 1220 -2109
rect 1224 -2113 1226 -2109
rect 1228 -2113 1229 -2109
rect 1241 -2113 1242 -2109
rect 1244 -2113 1246 -2109
rect 1250 -2113 1252 -2109
rect 1254 -2113 1255 -2109
rect 1267 -2113 1268 -2109
rect 1270 -2113 1271 -2109
rect 1275 -2113 1278 -2109
rect 1280 -2113 1286 -2109
rect 1288 -2113 1289 -2109
rect 1293 -2113 1296 -2109
rect 1298 -2113 1299 -2109
rect 1311 -2113 1312 -2109
rect 1314 -2113 1320 -2109
rect 1322 -2113 1324 -2109
rect 1328 -2113 1330 -2109
rect 1332 -2113 1333 -2109
rect 1345 -2113 1346 -2109
rect 1348 -2113 1350 -2109
rect 1354 -2113 1356 -2109
rect 1358 -2113 1364 -2109
rect 1366 -2113 1368 -2109
rect 1372 -2113 1374 -2109
rect 1376 -2113 1377 -2109
rect 1389 -2113 1390 -2109
rect 1392 -2113 1398 -2109
rect 1400 -2113 1401 -2109
rect 1413 -2113 1414 -2109
rect 1416 -2113 1421 -2109
rect 1425 -2113 1430 -2109
rect 1432 -2113 1433 -2109
rect 1437 -2113 1438 -2109
rect 1440 -2113 1442 -2109
rect 1446 -2113 1448 -2109
rect 1450 -2113 1451 -2109
rect -1230 -2257 -1229 -2253
rect -1227 -2257 -1225 -2253
rect -1221 -2257 -1219 -2253
rect -1217 -2257 -1216 -2253
rect -1204 -2257 -1203 -2253
rect -1201 -2257 -1195 -2253
rect -1193 -2257 -1192 -2253
rect -1180 -2257 -1179 -2253
rect -1177 -2257 -1171 -2253
rect -1169 -2257 -1167 -2253
rect -1163 -2257 -1161 -2253
rect -1159 -2257 -1153 -2253
rect -1151 -2257 -1150 -2253
rect -1138 -2257 -1137 -2253
rect -1135 -2257 -1129 -2253
rect -1127 -2257 -1125 -2253
rect -1121 -2257 -1119 -2253
rect -1117 -2257 -1111 -2253
rect -1109 -2257 -1108 -2253
rect -1096 -2257 -1095 -2253
rect -1093 -2257 -1087 -2253
rect -1085 -2257 -1083 -2253
rect -1079 -2257 -1077 -2253
rect -1075 -2257 -1069 -2253
rect -1067 -2257 -1066 -2253
rect -1054 -2257 -1053 -2253
rect -1051 -2257 -1045 -2253
rect -1043 -2257 -1042 -2253
rect -931 -2257 -930 -2253
rect -928 -2257 -926 -2253
rect -922 -2257 -920 -2253
rect -918 -2257 -917 -2253
rect -905 -2257 -904 -2253
rect -902 -2257 -896 -2253
rect -894 -2257 -893 -2253
rect -881 -2257 -880 -2253
rect -878 -2257 -872 -2253
rect -870 -2257 -868 -2253
rect -864 -2257 -862 -2253
rect -860 -2257 -854 -2253
rect -852 -2257 -851 -2253
rect -839 -2257 -838 -2253
rect -836 -2257 -830 -2253
rect -828 -2257 -826 -2253
rect -822 -2257 -820 -2253
rect -818 -2257 -812 -2253
rect -810 -2257 -809 -2253
rect -797 -2257 -796 -2253
rect -794 -2257 -788 -2253
rect -786 -2257 -784 -2253
rect -780 -2257 -778 -2253
rect -776 -2257 -770 -2253
rect -768 -2257 -767 -2253
rect -755 -2257 -754 -2253
rect -752 -2257 -746 -2253
rect -744 -2257 -743 -2253
rect -573 -2257 -572 -2253
rect -570 -2257 -568 -2253
rect -564 -2257 -562 -2253
rect -560 -2257 -559 -2253
rect -547 -2257 -546 -2253
rect -544 -2257 -538 -2253
rect -536 -2257 -535 -2253
rect -523 -2257 -522 -2253
rect -520 -2257 -514 -2253
rect -512 -2257 -510 -2253
rect -506 -2257 -504 -2253
rect -502 -2257 -496 -2253
rect -494 -2257 -493 -2253
rect -481 -2257 -480 -2253
rect -478 -2257 -472 -2253
rect -470 -2257 -468 -2253
rect -464 -2257 -462 -2253
rect -460 -2257 -454 -2253
rect -452 -2257 -451 -2253
rect -439 -2257 -438 -2253
rect -436 -2257 -430 -2253
rect -428 -2257 -426 -2253
rect -422 -2257 -420 -2253
rect -418 -2257 -412 -2253
rect -410 -2257 -409 -2253
rect -397 -2257 -396 -2253
rect -394 -2257 -388 -2253
rect -386 -2257 -385 -2253
rect -215 -2257 -214 -2253
rect -212 -2257 -210 -2253
rect -206 -2257 -204 -2253
rect -202 -2257 -201 -2253
rect -189 -2257 -188 -2253
rect -186 -2257 -180 -2253
rect -178 -2257 -177 -2253
rect -165 -2257 -164 -2253
rect -162 -2257 -156 -2253
rect -154 -2257 -152 -2253
rect -148 -2257 -146 -2253
rect -144 -2257 -138 -2253
rect -136 -2257 -135 -2253
rect -123 -2257 -122 -2253
rect -120 -2257 -114 -2253
rect -112 -2257 -110 -2253
rect -106 -2257 -104 -2253
rect -102 -2257 -96 -2253
rect -94 -2257 -93 -2253
rect -81 -2257 -80 -2253
rect -78 -2257 -72 -2253
rect -70 -2257 -68 -2253
rect -64 -2257 -62 -2253
rect -60 -2257 -54 -2253
rect -52 -2257 -51 -2253
rect -39 -2257 -38 -2253
rect -36 -2257 -30 -2253
rect -28 -2257 -27 -2253
rect 143 -2257 144 -2253
rect 146 -2257 148 -2253
rect 152 -2257 154 -2253
rect 156 -2257 157 -2253
rect 169 -2257 170 -2253
rect 172 -2257 178 -2253
rect 180 -2257 181 -2253
rect 193 -2257 194 -2253
rect 196 -2257 202 -2253
rect 204 -2257 206 -2253
rect 210 -2257 212 -2253
rect 214 -2257 220 -2253
rect 222 -2257 223 -2253
rect 235 -2257 236 -2253
rect 238 -2257 244 -2253
rect 246 -2257 248 -2253
rect 252 -2257 254 -2253
rect 256 -2257 262 -2253
rect 264 -2257 265 -2253
rect 277 -2257 278 -2253
rect 280 -2257 286 -2253
rect 288 -2257 290 -2253
rect 294 -2257 296 -2253
rect 298 -2257 304 -2253
rect 306 -2257 307 -2253
rect 319 -2257 320 -2253
rect 322 -2257 328 -2253
rect 330 -2257 331 -2253
rect 499 -2257 500 -2253
rect 502 -2257 504 -2253
rect 508 -2257 510 -2253
rect 512 -2257 513 -2253
rect 525 -2257 526 -2253
rect 528 -2257 534 -2253
rect 536 -2257 537 -2253
rect 549 -2257 550 -2253
rect 552 -2257 558 -2253
rect 560 -2257 562 -2253
rect 566 -2257 568 -2253
rect 570 -2257 576 -2253
rect 578 -2257 579 -2253
rect 591 -2257 592 -2253
rect 594 -2257 600 -2253
rect 602 -2257 604 -2253
rect 608 -2257 610 -2253
rect 612 -2257 618 -2253
rect 620 -2257 621 -2253
rect 633 -2257 634 -2253
rect 636 -2257 642 -2253
rect 644 -2257 646 -2253
rect 650 -2257 652 -2253
rect 654 -2257 660 -2253
rect 662 -2257 663 -2253
rect 675 -2257 676 -2253
rect 678 -2257 684 -2253
rect 686 -2257 687 -2253
rect -1555 -2428 -1554 -2424
rect -1552 -2428 -1550 -2424
rect -1546 -2428 -1544 -2424
rect -1542 -2428 -1541 -2424
rect -1529 -2428 -1528 -2424
rect -1526 -2428 -1520 -2424
rect -1518 -2428 -1517 -2424
rect -1505 -2428 -1504 -2424
rect -1502 -2428 -1496 -2424
rect -1494 -2428 -1492 -2424
rect -1488 -2428 -1486 -2424
rect -1484 -2428 -1478 -2424
rect -1476 -2428 -1475 -2424
rect -1463 -2428 -1462 -2424
rect -1460 -2428 -1454 -2424
rect -1452 -2428 -1450 -2424
rect -1446 -2428 -1444 -2424
rect -1442 -2428 -1436 -2424
rect -1434 -2428 -1433 -2424
rect -1421 -2428 -1420 -2424
rect -1418 -2428 -1412 -2424
rect -1410 -2428 -1408 -2424
rect -1404 -2428 -1402 -2424
rect -1400 -2428 -1394 -2424
rect -1392 -2428 -1391 -2424
rect -1379 -2428 -1378 -2424
rect -1376 -2428 -1370 -2424
rect -1368 -2428 -1367 -2424
rect -1230 -2428 -1229 -2424
rect -1227 -2428 -1225 -2424
rect -1221 -2428 -1219 -2424
rect -1217 -2428 -1216 -2424
rect -1204 -2428 -1203 -2424
rect -1201 -2428 -1195 -2424
rect -1193 -2428 -1192 -2424
rect -1180 -2428 -1179 -2424
rect -1177 -2428 -1171 -2424
rect -1169 -2428 -1167 -2424
rect -1163 -2428 -1161 -2424
rect -1159 -2428 -1153 -2424
rect -1151 -2428 -1150 -2424
rect -1138 -2428 -1137 -2424
rect -1135 -2428 -1129 -2424
rect -1127 -2428 -1125 -2424
rect -1121 -2428 -1119 -2424
rect -1117 -2428 -1111 -2424
rect -1109 -2428 -1108 -2424
rect -1096 -2428 -1095 -2424
rect -1093 -2428 -1087 -2424
rect -1085 -2428 -1083 -2424
rect -1079 -2428 -1077 -2424
rect -1075 -2428 -1069 -2424
rect -1067 -2428 -1066 -2424
rect -1054 -2428 -1053 -2424
rect -1051 -2428 -1045 -2424
rect -1043 -2428 -1042 -2424
rect -931 -2428 -930 -2424
rect -928 -2428 -926 -2424
rect -922 -2428 -920 -2424
rect -918 -2428 -917 -2424
rect -905 -2428 -904 -2424
rect -902 -2428 -896 -2424
rect -894 -2428 -893 -2424
rect -881 -2428 -880 -2424
rect -878 -2428 -872 -2424
rect -870 -2428 -868 -2424
rect -864 -2428 -862 -2424
rect -860 -2428 -854 -2424
rect -852 -2428 -851 -2424
rect -839 -2428 -838 -2424
rect -836 -2428 -830 -2424
rect -828 -2428 -826 -2424
rect -822 -2428 -820 -2424
rect -818 -2428 -812 -2424
rect -810 -2428 -809 -2424
rect -797 -2428 -796 -2424
rect -794 -2428 -788 -2424
rect -786 -2428 -784 -2424
rect -780 -2428 -778 -2424
rect -776 -2428 -770 -2424
rect -768 -2428 -767 -2424
rect -755 -2428 -754 -2424
rect -752 -2428 -746 -2424
rect -744 -2428 -743 -2424
rect -573 -2428 -572 -2424
rect -570 -2428 -568 -2424
rect -564 -2428 -562 -2424
rect -560 -2428 -559 -2424
rect -547 -2428 -546 -2424
rect -544 -2428 -538 -2424
rect -536 -2428 -535 -2424
rect -523 -2428 -522 -2424
rect -520 -2428 -514 -2424
rect -512 -2428 -510 -2424
rect -506 -2428 -504 -2424
rect -502 -2428 -496 -2424
rect -494 -2428 -493 -2424
rect -481 -2428 -480 -2424
rect -478 -2428 -472 -2424
rect -470 -2428 -468 -2424
rect -464 -2428 -462 -2424
rect -460 -2428 -454 -2424
rect -452 -2428 -451 -2424
rect -439 -2428 -438 -2424
rect -436 -2428 -430 -2424
rect -428 -2428 -426 -2424
rect -422 -2428 -420 -2424
rect -418 -2428 -412 -2424
rect -410 -2428 -409 -2424
rect -397 -2428 -396 -2424
rect -394 -2428 -388 -2424
rect -386 -2428 -385 -2424
rect -215 -2428 -214 -2424
rect -212 -2428 -210 -2424
rect -206 -2428 -204 -2424
rect -202 -2428 -201 -2424
rect -189 -2428 -188 -2424
rect -186 -2428 -180 -2424
rect -178 -2428 -177 -2424
rect -165 -2428 -164 -2424
rect -162 -2428 -156 -2424
rect -154 -2428 -152 -2424
rect -148 -2428 -146 -2424
rect -144 -2428 -138 -2424
rect -136 -2428 -135 -2424
rect -123 -2428 -122 -2424
rect -120 -2428 -114 -2424
rect -112 -2428 -110 -2424
rect -106 -2428 -104 -2424
rect -102 -2428 -96 -2424
rect -94 -2428 -93 -2424
rect -81 -2428 -80 -2424
rect -78 -2428 -72 -2424
rect -70 -2428 -68 -2424
rect -64 -2428 -62 -2424
rect -60 -2428 -54 -2424
rect -52 -2428 -51 -2424
rect -39 -2428 -38 -2424
rect -36 -2428 -30 -2424
rect -28 -2428 -27 -2424
rect 143 -2428 144 -2424
rect 146 -2428 148 -2424
rect 152 -2428 154 -2424
rect 156 -2428 157 -2424
rect 169 -2428 170 -2424
rect 172 -2428 178 -2424
rect 180 -2428 181 -2424
rect 193 -2428 194 -2424
rect 196 -2428 202 -2424
rect 204 -2428 206 -2424
rect 210 -2428 212 -2424
rect 214 -2428 220 -2424
rect 222 -2428 223 -2424
rect 235 -2428 236 -2424
rect 238 -2428 244 -2424
rect 246 -2428 248 -2424
rect 252 -2428 254 -2424
rect 256 -2428 262 -2424
rect 264 -2428 265 -2424
rect 277 -2428 278 -2424
rect 280 -2428 286 -2424
rect 288 -2428 290 -2424
rect 294 -2428 296 -2424
rect 298 -2428 304 -2424
rect 306 -2428 307 -2424
rect 319 -2428 320 -2424
rect 322 -2428 328 -2424
rect 330 -2428 331 -2424
rect 499 -2428 500 -2424
rect 502 -2428 504 -2424
rect 508 -2428 510 -2424
rect 512 -2428 513 -2424
rect 525 -2428 526 -2424
rect 528 -2428 534 -2424
rect 536 -2428 537 -2424
rect 549 -2428 550 -2424
rect 552 -2428 558 -2424
rect 560 -2428 562 -2424
rect 566 -2428 568 -2424
rect 570 -2428 576 -2424
rect 578 -2428 579 -2424
rect 591 -2428 592 -2424
rect 594 -2428 600 -2424
rect 602 -2428 604 -2424
rect 608 -2428 610 -2424
rect 612 -2428 618 -2424
rect 620 -2428 621 -2424
rect 633 -2428 634 -2424
rect 636 -2428 642 -2424
rect 644 -2428 646 -2424
rect 650 -2428 652 -2424
rect 654 -2428 660 -2424
rect 662 -2428 663 -2424
rect 675 -2428 676 -2424
rect 678 -2428 684 -2424
rect 686 -2428 687 -2424
rect 857 -2428 858 -2424
rect 860 -2428 862 -2424
rect 866 -2428 868 -2424
rect 870 -2428 871 -2424
rect 883 -2428 884 -2424
rect 886 -2428 892 -2424
rect 894 -2428 895 -2424
rect 907 -2428 908 -2424
rect 910 -2428 916 -2424
rect 918 -2428 920 -2424
rect 924 -2428 926 -2424
rect 928 -2428 934 -2424
rect 936 -2428 937 -2424
rect 949 -2428 950 -2424
rect 952 -2428 958 -2424
rect 960 -2428 962 -2424
rect 966 -2428 968 -2424
rect 970 -2428 976 -2424
rect 978 -2428 979 -2424
rect 991 -2428 992 -2424
rect 994 -2428 1000 -2424
rect 1002 -2428 1004 -2424
rect 1008 -2428 1010 -2424
rect 1012 -2428 1018 -2424
rect 1020 -2428 1021 -2424
rect 1033 -2428 1034 -2424
rect 1036 -2428 1042 -2424
rect 1044 -2428 1045 -2424
rect 1215 -2428 1216 -2424
rect 1218 -2428 1220 -2424
rect 1224 -2428 1226 -2424
rect 1228 -2428 1229 -2424
rect 1241 -2428 1242 -2424
rect 1244 -2428 1250 -2424
rect 1252 -2428 1253 -2424
rect 1265 -2428 1266 -2424
rect 1268 -2428 1274 -2424
rect 1276 -2428 1278 -2424
rect 1282 -2428 1284 -2424
rect 1286 -2428 1292 -2424
rect 1294 -2428 1295 -2424
rect 1307 -2428 1308 -2424
rect 1310 -2428 1316 -2424
rect 1318 -2428 1320 -2424
rect 1324 -2428 1326 -2424
rect 1328 -2428 1334 -2424
rect 1336 -2428 1337 -2424
rect 1349 -2428 1350 -2424
rect 1352 -2428 1358 -2424
rect 1360 -2428 1362 -2424
rect 1366 -2428 1368 -2424
rect 1370 -2428 1376 -2424
rect 1378 -2428 1379 -2424
rect 1391 -2428 1392 -2424
rect 1394 -2428 1400 -2424
rect 1402 -2428 1403 -2424
rect -1555 -2599 -1554 -2595
rect -1552 -2599 -1550 -2595
rect -1546 -2599 -1544 -2595
rect -1542 -2599 -1541 -2595
rect -1529 -2599 -1528 -2595
rect -1526 -2599 -1520 -2595
rect -1518 -2599 -1517 -2595
rect -1505 -2599 -1504 -2595
rect -1502 -2599 -1496 -2595
rect -1494 -2599 -1492 -2595
rect -1488 -2599 -1486 -2595
rect -1484 -2599 -1478 -2595
rect -1476 -2599 -1475 -2595
rect -1463 -2599 -1462 -2595
rect -1460 -2599 -1454 -2595
rect -1452 -2599 -1450 -2595
rect -1446 -2599 -1444 -2595
rect -1442 -2599 -1436 -2595
rect -1434 -2599 -1433 -2595
rect -1421 -2599 -1420 -2595
rect -1418 -2599 -1412 -2595
rect -1410 -2599 -1408 -2595
rect -1404 -2599 -1402 -2595
rect -1400 -2599 -1394 -2595
rect -1392 -2599 -1391 -2595
rect -1379 -2599 -1378 -2595
rect -1376 -2599 -1370 -2595
rect -1368 -2599 -1367 -2595
rect -1230 -2599 -1229 -2595
rect -1227 -2599 -1225 -2595
rect -1221 -2599 -1219 -2595
rect -1217 -2599 -1216 -2595
rect -1204 -2599 -1203 -2595
rect -1201 -2599 -1195 -2595
rect -1193 -2599 -1192 -2595
rect -1180 -2599 -1179 -2595
rect -1177 -2599 -1171 -2595
rect -1169 -2599 -1167 -2595
rect -1163 -2599 -1161 -2595
rect -1159 -2599 -1153 -2595
rect -1151 -2599 -1150 -2595
rect -1138 -2599 -1137 -2595
rect -1135 -2599 -1129 -2595
rect -1127 -2599 -1125 -2595
rect -1121 -2599 -1119 -2595
rect -1117 -2599 -1111 -2595
rect -1109 -2599 -1108 -2595
rect -1096 -2599 -1095 -2595
rect -1093 -2599 -1087 -2595
rect -1085 -2599 -1083 -2595
rect -1079 -2599 -1077 -2595
rect -1075 -2599 -1069 -2595
rect -1067 -2599 -1066 -2595
rect -1054 -2599 -1053 -2595
rect -1051 -2599 -1045 -2595
rect -1043 -2599 -1042 -2595
rect -931 -2599 -930 -2595
rect -928 -2599 -926 -2595
rect -922 -2599 -920 -2595
rect -918 -2599 -917 -2595
rect -905 -2599 -904 -2595
rect -902 -2599 -896 -2595
rect -894 -2599 -893 -2595
rect -881 -2599 -880 -2595
rect -878 -2599 -872 -2595
rect -870 -2599 -868 -2595
rect -864 -2599 -862 -2595
rect -860 -2599 -854 -2595
rect -852 -2599 -851 -2595
rect -839 -2599 -838 -2595
rect -836 -2599 -830 -2595
rect -828 -2599 -826 -2595
rect -822 -2599 -820 -2595
rect -818 -2599 -812 -2595
rect -810 -2599 -809 -2595
rect -797 -2599 -796 -2595
rect -794 -2599 -788 -2595
rect -786 -2599 -784 -2595
rect -780 -2599 -778 -2595
rect -776 -2599 -770 -2595
rect -768 -2599 -767 -2595
rect -755 -2599 -754 -2595
rect -752 -2599 -746 -2595
rect -744 -2599 -743 -2595
rect -573 -2599 -572 -2595
rect -570 -2599 -568 -2595
rect -564 -2599 -562 -2595
rect -560 -2599 -559 -2595
rect -547 -2599 -546 -2595
rect -544 -2599 -538 -2595
rect -536 -2599 -535 -2595
rect -523 -2599 -522 -2595
rect -520 -2599 -514 -2595
rect -512 -2599 -510 -2595
rect -506 -2599 -504 -2595
rect -502 -2599 -496 -2595
rect -494 -2599 -493 -2595
rect -481 -2599 -480 -2595
rect -478 -2599 -472 -2595
rect -470 -2599 -468 -2595
rect -464 -2599 -462 -2595
rect -460 -2599 -454 -2595
rect -452 -2599 -451 -2595
rect -439 -2599 -438 -2595
rect -436 -2599 -430 -2595
rect -428 -2599 -426 -2595
rect -422 -2599 -420 -2595
rect -418 -2599 -412 -2595
rect -410 -2599 -409 -2595
rect -397 -2599 -396 -2595
rect -394 -2599 -388 -2595
rect -386 -2599 -385 -2595
rect -216 -2599 -215 -2595
rect -213 -2599 -211 -2595
rect -207 -2599 -205 -2595
rect -203 -2599 -202 -2595
rect -190 -2599 -189 -2595
rect -187 -2599 -181 -2595
rect -179 -2599 -178 -2595
rect -166 -2599 -165 -2595
rect -163 -2599 -157 -2595
rect -155 -2599 -153 -2595
rect -149 -2599 -147 -2595
rect -145 -2599 -139 -2595
rect -137 -2599 -136 -2595
rect -124 -2599 -123 -2595
rect -121 -2599 -115 -2595
rect -113 -2599 -111 -2595
rect -107 -2599 -105 -2595
rect -103 -2599 -97 -2595
rect -95 -2599 -94 -2595
rect -82 -2599 -81 -2595
rect -79 -2599 -73 -2595
rect -71 -2599 -69 -2595
rect -65 -2599 -63 -2595
rect -61 -2599 -55 -2595
rect -53 -2599 -52 -2595
rect -40 -2599 -39 -2595
rect -37 -2599 -31 -2595
rect -29 -2599 -28 -2595
rect 143 -2599 144 -2595
rect 146 -2599 148 -2595
rect 152 -2599 154 -2595
rect 156 -2599 157 -2595
rect 169 -2599 170 -2595
rect 172 -2599 178 -2595
rect 180 -2599 181 -2595
rect 193 -2599 194 -2595
rect 196 -2599 202 -2595
rect 204 -2599 206 -2595
rect 210 -2599 212 -2595
rect 214 -2599 220 -2595
rect 222 -2599 223 -2595
rect 235 -2599 236 -2595
rect 238 -2599 244 -2595
rect 246 -2599 248 -2595
rect 252 -2599 254 -2595
rect 256 -2599 262 -2595
rect 264 -2599 265 -2595
rect 277 -2599 278 -2595
rect 280 -2599 286 -2595
rect 288 -2599 290 -2595
rect 294 -2599 296 -2595
rect 298 -2599 304 -2595
rect 306 -2599 307 -2595
rect 319 -2599 320 -2595
rect 322 -2599 328 -2595
rect 330 -2599 331 -2595
rect 499 -2599 500 -2595
rect 502 -2599 504 -2595
rect 508 -2599 510 -2595
rect 512 -2599 513 -2595
rect 525 -2599 526 -2595
rect 528 -2599 534 -2595
rect 536 -2599 537 -2595
rect 549 -2599 550 -2595
rect 552 -2599 558 -2595
rect 560 -2599 562 -2595
rect 566 -2599 568 -2595
rect 570 -2599 576 -2595
rect 578 -2599 579 -2595
rect 591 -2599 592 -2595
rect 594 -2599 600 -2595
rect 602 -2599 604 -2595
rect 608 -2599 610 -2595
rect 612 -2599 618 -2595
rect 620 -2599 621 -2595
rect 633 -2599 634 -2595
rect 636 -2599 642 -2595
rect 644 -2599 646 -2595
rect 650 -2599 652 -2595
rect 654 -2599 660 -2595
rect 662 -2599 663 -2595
rect 675 -2599 676 -2595
rect 678 -2599 684 -2595
rect 686 -2599 687 -2595
rect 857 -2599 858 -2595
rect 860 -2599 862 -2595
rect 866 -2599 868 -2595
rect 870 -2599 871 -2595
rect 883 -2599 884 -2595
rect 886 -2599 892 -2595
rect 894 -2599 895 -2595
rect 907 -2599 908 -2595
rect 910 -2599 916 -2595
rect 918 -2599 920 -2595
rect 924 -2599 926 -2595
rect 928 -2599 934 -2595
rect 936 -2599 937 -2595
rect 949 -2599 950 -2595
rect 952 -2599 958 -2595
rect 960 -2599 962 -2595
rect 966 -2599 968 -2595
rect 970 -2599 976 -2595
rect 978 -2599 979 -2595
rect 991 -2599 992 -2595
rect 994 -2599 1000 -2595
rect 1002 -2599 1004 -2595
rect 1008 -2599 1010 -2595
rect 1012 -2599 1018 -2595
rect 1020 -2599 1021 -2595
rect 1033 -2599 1034 -2595
rect 1036 -2599 1042 -2595
rect 1044 -2599 1045 -2595
rect 1215 -2599 1216 -2595
rect 1218 -2599 1220 -2595
rect 1224 -2599 1226 -2595
rect 1228 -2599 1229 -2595
rect 1241 -2599 1242 -2595
rect 1244 -2599 1250 -2595
rect 1252 -2599 1253 -2595
rect 1265 -2599 1266 -2595
rect 1268 -2599 1274 -2595
rect 1276 -2599 1278 -2595
rect 1282 -2599 1284 -2595
rect 1286 -2599 1292 -2595
rect 1294 -2599 1295 -2595
rect 1307 -2599 1308 -2595
rect 1310 -2599 1316 -2595
rect 1318 -2599 1320 -2595
rect 1324 -2599 1326 -2595
rect 1328 -2599 1334 -2595
rect 1336 -2599 1337 -2595
rect 1349 -2599 1350 -2595
rect 1352 -2599 1358 -2595
rect 1360 -2599 1362 -2595
rect 1366 -2599 1368 -2595
rect 1370 -2599 1376 -2595
rect 1378 -2599 1379 -2595
rect 1391 -2599 1392 -2595
rect 1394 -2599 1400 -2595
rect 1402 -2599 1403 -2595
rect -1305 -2704 -1304 -2700
rect -1302 -2704 -1296 -2700
rect -1294 -2704 -1292 -2700
rect -1288 -2704 -1286 -2700
rect -1284 -2704 -1283 -2700
rect -931 -2704 -930 -2700
rect -928 -2704 -922 -2700
rect -920 -2704 -918 -2700
rect -914 -2704 -912 -2700
rect -910 -2704 -909 -2700
rect -573 -2704 -572 -2700
rect -570 -2704 -564 -2700
rect -562 -2704 -560 -2700
rect -556 -2704 -554 -2700
rect -552 -2704 -551 -2700
rect -215 -2704 -214 -2700
rect -212 -2704 -206 -2700
rect -204 -2704 -202 -2700
rect -198 -2704 -196 -2700
rect -194 -2704 -193 -2700
rect 143 -2704 144 -2700
rect 146 -2704 152 -2700
rect 154 -2704 156 -2700
rect 160 -2704 162 -2700
rect 164 -2704 165 -2700
rect 499 -2704 500 -2700
rect 502 -2704 508 -2700
rect 510 -2704 512 -2700
rect 516 -2704 518 -2700
rect 520 -2704 521 -2700
rect 857 -2704 858 -2700
rect 860 -2704 866 -2700
rect 868 -2704 870 -2700
rect 874 -2704 876 -2700
rect 878 -2704 879 -2700
rect 1215 -2704 1216 -2700
rect 1218 -2704 1224 -2700
rect 1226 -2704 1228 -2700
rect 1232 -2704 1234 -2700
rect 1236 -2704 1237 -2700
rect -1230 -2863 -1229 -2859
rect -1227 -2863 -1225 -2859
rect -1221 -2863 -1219 -2859
rect -1217 -2863 -1216 -2859
rect -1204 -2863 -1203 -2859
rect -1201 -2863 -1199 -2859
rect -1195 -2863 -1193 -2859
rect -1191 -2863 -1185 -2859
rect -1183 -2863 -1181 -2859
rect -1177 -2863 -1175 -2859
rect -1173 -2863 -1172 -2859
rect -1160 -2863 -1159 -2859
rect -1157 -2863 -1151 -2859
rect -1149 -2863 -1147 -2859
rect -1143 -2863 -1141 -2859
rect -1139 -2863 -1138 -2859
rect -931 -2863 -930 -2859
rect -928 -2863 -926 -2859
rect -922 -2863 -920 -2859
rect -918 -2863 -917 -2859
rect -905 -2863 -904 -2859
rect -902 -2863 -900 -2859
rect -896 -2863 -894 -2859
rect -892 -2863 -891 -2859
rect -879 -2863 -878 -2859
rect -876 -2863 -875 -2859
rect -871 -2863 -868 -2859
rect -866 -2863 -860 -2859
rect -858 -2863 -857 -2859
rect -853 -2863 -850 -2859
rect -848 -2863 -847 -2859
rect -835 -2863 -834 -2859
rect -832 -2863 -826 -2859
rect -824 -2863 -822 -2859
rect -818 -2863 -816 -2859
rect -814 -2863 -813 -2859
rect -801 -2863 -800 -2859
rect -798 -2863 -796 -2859
rect -792 -2863 -790 -2859
rect -788 -2863 -782 -2859
rect -780 -2863 -778 -2859
rect -774 -2863 -772 -2859
rect -770 -2863 -769 -2859
rect -757 -2863 -756 -2859
rect -754 -2863 -748 -2859
rect -746 -2863 -745 -2859
rect -733 -2863 -732 -2859
rect -730 -2863 -725 -2859
rect -721 -2863 -716 -2859
rect -714 -2863 -713 -2859
rect -709 -2863 -708 -2859
rect -706 -2863 -704 -2859
rect -700 -2863 -698 -2859
rect -696 -2863 -695 -2859
rect -573 -2863 -572 -2859
rect -570 -2863 -568 -2859
rect -564 -2863 -562 -2859
rect -560 -2863 -559 -2859
rect -547 -2863 -546 -2859
rect -544 -2863 -542 -2859
rect -538 -2863 -536 -2859
rect -534 -2863 -533 -2859
rect -521 -2863 -520 -2859
rect -518 -2863 -517 -2859
rect -513 -2863 -510 -2859
rect -508 -2863 -502 -2859
rect -500 -2863 -499 -2859
rect -495 -2863 -492 -2859
rect -490 -2863 -489 -2859
rect -477 -2863 -476 -2859
rect -474 -2863 -468 -2859
rect -466 -2863 -464 -2859
rect -460 -2863 -458 -2859
rect -456 -2863 -455 -2859
rect -443 -2863 -442 -2859
rect -440 -2863 -438 -2859
rect -434 -2863 -432 -2859
rect -430 -2863 -424 -2859
rect -422 -2863 -420 -2859
rect -416 -2863 -414 -2859
rect -412 -2863 -411 -2859
rect -399 -2863 -398 -2859
rect -396 -2863 -390 -2859
rect -388 -2863 -387 -2859
rect -375 -2863 -374 -2859
rect -372 -2863 -367 -2859
rect -363 -2863 -358 -2859
rect -356 -2863 -355 -2859
rect -351 -2863 -350 -2859
rect -348 -2863 -346 -2859
rect -342 -2863 -340 -2859
rect -338 -2863 -337 -2859
rect -215 -2863 -214 -2859
rect -212 -2863 -210 -2859
rect -206 -2863 -204 -2859
rect -202 -2863 -201 -2859
rect -189 -2863 -188 -2859
rect -186 -2863 -184 -2859
rect -180 -2863 -178 -2859
rect -176 -2863 -175 -2859
rect -163 -2863 -162 -2859
rect -160 -2863 -159 -2859
rect -155 -2863 -152 -2859
rect -150 -2863 -144 -2859
rect -142 -2863 -141 -2859
rect -137 -2863 -134 -2859
rect -132 -2863 -131 -2859
rect -119 -2863 -118 -2859
rect -116 -2863 -110 -2859
rect -108 -2863 -106 -2859
rect -102 -2863 -100 -2859
rect -98 -2863 -97 -2859
rect -85 -2863 -84 -2859
rect -82 -2863 -80 -2859
rect -76 -2863 -74 -2859
rect -72 -2863 -66 -2859
rect -64 -2863 -62 -2859
rect -58 -2863 -56 -2859
rect -54 -2863 -53 -2859
rect -41 -2863 -40 -2859
rect -38 -2863 -32 -2859
rect -30 -2863 -29 -2859
rect -17 -2863 -16 -2859
rect -14 -2863 -9 -2859
rect -5 -2863 0 -2859
rect 2 -2863 3 -2859
rect 7 -2863 8 -2859
rect 10 -2863 12 -2859
rect 16 -2863 18 -2859
rect 20 -2863 21 -2859
rect 143 -2863 144 -2859
rect 146 -2863 148 -2859
rect 152 -2863 154 -2859
rect 156 -2863 157 -2859
rect 169 -2863 170 -2859
rect 172 -2863 174 -2859
rect 178 -2863 180 -2859
rect 182 -2863 183 -2859
rect 195 -2863 196 -2859
rect 198 -2863 199 -2859
rect 203 -2863 206 -2859
rect 208 -2863 214 -2859
rect 216 -2863 217 -2859
rect 221 -2863 224 -2859
rect 226 -2863 227 -2859
rect 239 -2863 240 -2859
rect 242 -2863 248 -2859
rect 250 -2863 252 -2859
rect 256 -2863 258 -2859
rect 260 -2863 261 -2859
rect 273 -2863 274 -2859
rect 276 -2863 278 -2859
rect 282 -2863 284 -2859
rect 286 -2863 292 -2859
rect 294 -2863 296 -2859
rect 300 -2863 302 -2859
rect 304 -2863 305 -2859
rect 317 -2863 318 -2859
rect 320 -2863 326 -2859
rect 328 -2863 329 -2859
rect 341 -2863 342 -2859
rect 344 -2863 349 -2859
rect 353 -2863 358 -2859
rect 360 -2863 361 -2859
rect 365 -2863 366 -2859
rect 368 -2863 370 -2859
rect 374 -2863 376 -2859
rect 378 -2863 379 -2859
rect 499 -2863 500 -2859
rect 502 -2863 504 -2859
rect 508 -2863 510 -2859
rect 512 -2863 513 -2859
rect 525 -2863 526 -2859
rect 528 -2863 530 -2859
rect 534 -2863 536 -2859
rect 538 -2863 539 -2859
rect 551 -2863 552 -2859
rect 554 -2863 555 -2859
rect 559 -2863 562 -2859
rect 564 -2863 570 -2859
rect 572 -2863 573 -2859
rect 577 -2863 580 -2859
rect 582 -2863 583 -2859
rect 595 -2863 596 -2859
rect 598 -2863 604 -2859
rect 606 -2863 608 -2859
rect 612 -2863 614 -2859
rect 616 -2863 617 -2859
rect 629 -2863 630 -2859
rect 632 -2863 634 -2859
rect 638 -2863 640 -2859
rect 642 -2863 648 -2859
rect 650 -2863 652 -2859
rect 656 -2863 658 -2859
rect 660 -2863 661 -2859
rect 673 -2863 674 -2859
rect 676 -2863 682 -2859
rect 684 -2863 685 -2859
rect 697 -2863 698 -2859
rect 700 -2863 705 -2859
rect 709 -2863 714 -2859
rect 716 -2863 717 -2859
rect 721 -2863 722 -2859
rect 724 -2863 726 -2859
rect 730 -2863 732 -2859
rect 734 -2863 735 -2859
rect 857 -2863 858 -2859
rect 860 -2863 862 -2859
rect 866 -2863 868 -2859
rect 870 -2863 871 -2859
rect 883 -2863 884 -2859
rect 886 -2863 888 -2859
rect 892 -2863 894 -2859
rect 896 -2863 897 -2859
rect 909 -2863 910 -2859
rect 912 -2863 913 -2859
rect 917 -2863 920 -2859
rect 922 -2863 928 -2859
rect 930 -2863 931 -2859
rect 935 -2863 938 -2859
rect 940 -2863 941 -2859
rect 953 -2863 954 -2859
rect 956 -2863 962 -2859
rect 964 -2863 966 -2859
rect 970 -2863 972 -2859
rect 974 -2863 975 -2859
rect 987 -2863 988 -2859
rect 990 -2863 992 -2859
rect 996 -2863 998 -2859
rect 1000 -2863 1006 -2859
rect 1008 -2863 1010 -2859
rect 1014 -2863 1016 -2859
rect 1018 -2863 1019 -2859
rect 1031 -2863 1032 -2859
rect 1034 -2863 1040 -2859
rect 1042 -2863 1043 -2859
rect 1055 -2863 1056 -2859
rect 1058 -2863 1063 -2859
rect 1067 -2863 1072 -2859
rect 1074 -2863 1075 -2859
rect 1079 -2863 1080 -2859
rect 1082 -2863 1084 -2859
rect 1088 -2863 1090 -2859
rect 1092 -2863 1093 -2859
rect 1215 -2863 1216 -2859
rect 1218 -2863 1220 -2859
rect 1224 -2863 1226 -2859
rect 1228 -2863 1229 -2859
rect 1241 -2863 1242 -2859
rect 1244 -2863 1246 -2859
rect 1250 -2863 1252 -2859
rect 1254 -2863 1255 -2859
rect 1267 -2863 1268 -2859
rect 1270 -2863 1271 -2859
rect 1275 -2863 1278 -2859
rect 1280 -2863 1286 -2859
rect 1288 -2863 1289 -2859
rect 1293 -2863 1296 -2859
rect 1298 -2863 1299 -2859
rect 1311 -2863 1312 -2859
rect 1314 -2863 1320 -2859
rect 1322 -2863 1324 -2859
rect 1328 -2863 1330 -2859
rect 1332 -2863 1333 -2859
rect 1345 -2863 1346 -2859
rect 1348 -2863 1350 -2859
rect 1354 -2863 1356 -2859
rect 1358 -2863 1364 -2859
rect 1366 -2863 1368 -2859
rect 1372 -2863 1374 -2859
rect 1376 -2863 1377 -2859
rect 1389 -2863 1390 -2859
rect 1392 -2863 1398 -2859
rect 1400 -2863 1401 -2859
rect 1413 -2863 1414 -2859
rect 1416 -2863 1421 -2859
rect 1425 -2863 1430 -2859
rect 1432 -2863 1433 -2859
rect 1437 -2863 1438 -2859
rect 1440 -2863 1442 -2859
rect 1446 -2863 1448 -2859
rect 1450 -2863 1451 -2859
rect -1555 -2982 -1554 -2978
rect -1552 -2982 -1550 -2978
rect -1546 -2982 -1544 -2978
rect -1542 -2982 -1541 -2978
rect -1529 -2982 -1528 -2978
rect -1526 -2982 -1520 -2978
rect -1518 -2982 -1517 -2978
rect -1505 -2982 -1504 -2978
rect -1502 -2982 -1496 -2978
rect -1494 -2982 -1492 -2978
rect -1488 -2982 -1486 -2978
rect -1484 -2982 -1478 -2978
rect -1476 -2982 -1475 -2978
rect -1463 -2982 -1462 -2978
rect -1460 -2982 -1454 -2978
rect -1452 -2982 -1450 -2978
rect -1446 -2982 -1444 -2978
rect -1442 -2982 -1436 -2978
rect -1434 -2982 -1433 -2978
rect -1421 -2982 -1420 -2978
rect -1418 -2982 -1412 -2978
rect -1410 -2982 -1408 -2978
rect -1404 -2982 -1402 -2978
rect -1400 -2982 -1394 -2978
rect -1392 -2982 -1391 -2978
rect -1379 -2982 -1378 -2978
rect -1376 -2982 -1370 -2978
rect -1368 -2982 -1367 -2978
rect -1230 -2982 -1229 -2978
rect -1227 -2982 -1225 -2978
rect -1221 -2982 -1219 -2978
rect -1217 -2982 -1216 -2978
rect -1204 -2982 -1203 -2978
rect -1201 -2982 -1195 -2978
rect -1193 -2982 -1192 -2978
rect -1180 -2982 -1179 -2978
rect -1177 -2982 -1171 -2978
rect -1169 -2982 -1167 -2978
rect -1163 -2982 -1161 -2978
rect -1159 -2982 -1153 -2978
rect -1151 -2982 -1150 -2978
rect -1138 -2982 -1137 -2978
rect -1135 -2982 -1129 -2978
rect -1127 -2982 -1125 -2978
rect -1121 -2982 -1119 -2978
rect -1117 -2982 -1111 -2978
rect -1109 -2982 -1108 -2978
rect -1096 -2982 -1095 -2978
rect -1093 -2982 -1087 -2978
rect -1085 -2982 -1083 -2978
rect -1079 -2982 -1077 -2978
rect -1075 -2982 -1069 -2978
rect -1067 -2982 -1066 -2978
rect -1054 -2982 -1053 -2978
rect -1051 -2982 -1045 -2978
rect -1043 -2982 -1042 -2978
rect -931 -2982 -930 -2978
rect -928 -2982 -926 -2978
rect -922 -2982 -920 -2978
rect -918 -2982 -917 -2978
rect -905 -2982 -904 -2978
rect -902 -2982 -896 -2978
rect -894 -2982 -893 -2978
rect -881 -2982 -880 -2978
rect -878 -2982 -872 -2978
rect -870 -2982 -868 -2978
rect -864 -2982 -862 -2978
rect -860 -2982 -854 -2978
rect -852 -2982 -851 -2978
rect -839 -2982 -838 -2978
rect -836 -2982 -830 -2978
rect -828 -2982 -826 -2978
rect -822 -2982 -820 -2978
rect -818 -2982 -812 -2978
rect -810 -2982 -809 -2978
rect -797 -2982 -796 -2978
rect -794 -2982 -788 -2978
rect -786 -2982 -784 -2978
rect -780 -2982 -778 -2978
rect -776 -2982 -770 -2978
rect -768 -2982 -767 -2978
rect -755 -2982 -754 -2978
rect -752 -2982 -746 -2978
rect -744 -2982 -743 -2978
rect -573 -2982 -572 -2978
rect -570 -2982 -568 -2978
rect -564 -2982 -562 -2978
rect -560 -2982 -559 -2978
rect -547 -2982 -546 -2978
rect -544 -2982 -538 -2978
rect -536 -2982 -535 -2978
rect -523 -2982 -522 -2978
rect -520 -2982 -514 -2978
rect -512 -2982 -510 -2978
rect -506 -2982 -504 -2978
rect -502 -2982 -496 -2978
rect -494 -2982 -493 -2978
rect -481 -2982 -480 -2978
rect -478 -2982 -472 -2978
rect -470 -2982 -468 -2978
rect -464 -2982 -462 -2978
rect -460 -2982 -454 -2978
rect -452 -2982 -451 -2978
rect -439 -2982 -438 -2978
rect -436 -2982 -430 -2978
rect -428 -2982 -426 -2978
rect -422 -2982 -420 -2978
rect -418 -2982 -412 -2978
rect -410 -2982 -409 -2978
rect -397 -2982 -396 -2978
rect -394 -2982 -388 -2978
rect -386 -2982 -385 -2978
rect -215 -2982 -214 -2978
rect -212 -2982 -210 -2978
rect -206 -2982 -204 -2978
rect -202 -2982 -201 -2978
rect -189 -2982 -188 -2978
rect -186 -2982 -180 -2978
rect -178 -2982 -177 -2978
rect -165 -2982 -164 -2978
rect -162 -2982 -156 -2978
rect -154 -2982 -152 -2978
rect -148 -2982 -146 -2978
rect -144 -2982 -138 -2978
rect -136 -2982 -135 -2978
rect -123 -2982 -122 -2978
rect -120 -2982 -114 -2978
rect -112 -2982 -110 -2978
rect -106 -2982 -104 -2978
rect -102 -2982 -96 -2978
rect -94 -2982 -93 -2978
rect -81 -2982 -80 -2978
rect -78 -2982 -72 -2978
rect -70 -2982 -68 -2978
rect -64 -2982 -62 -2978
rect -60 -2982 -54 -2978
rect -52 -2982 -51 -2978
rect -39 -2982 -38 -2978
rect -36 -2982 -30 -2978
rect -28 -2982 -27 -2978
rect 143 -2982 144 -2978
rect 146 -2982 148 -2978
rect 152 -2982 154 -2978
rect 156 -2982 157 -2978
rect 169 -2982 170 -2978
rect 172 -2982 178 -2978
rect 180 -2982 181 -2978
rect 193 -2982 194 -2978
rect 196 -2982 202 -2978
rect 204 -2982 206 -2978
rect 210 -2982 212 -2978
rect 214 -2982 220 -2978
rect 222 -2982 223 -2978
rect 235 -2982 236 -2978
rect 238 -2982 244 -2978
rect 246 -2982 248 -2978
rect 252 -2982 254 -2978
rect 256 -2982 262 -2978
rect 264 -2982 265 -2978
rect 277 -2982 278 -2978
rect 280 -2982 286 -2978
rect 288 -2982 290 -2978
rect 294 -2982 296 -2978
rect 298 -2982 304 -2978
rect 306 -2982 307 -2978
rect 319 -2982 320 -2978
rect 322 -2982 328 -2978
rect 330 -2982 331 -2978
rect -1555 -3153 -1554 -3149
rect -1552 -3153 -1550 -3149
rect -1546 -3153 -1544 -3149
rect -1542 -3153 -1541 -3149
rect -1529 -3153 -1528 -3149
rect -1526 -3153 -1520 -3149
rect -1518 -3153 -1517 -3149
rect -1505 -3153 -1504 -3149
rect -1502 -3153 -1496 -3149
rect -1494 -3153 -1492 -3149
rect -1488 -3153 -1486 -3149
rect -1484 -3153 -1478 -3149
rect -1476 -3153 -1475 -3149
rect -1463 -3153 -1462 -3149
rect -1460 -3153 -1454 -3149
rect -1452 -3153 -1450 -3149
rect -1446 -3153 -1444 -3149
rect -1442 -3153 -1436 -3149
rect -1434 -3153 -1433 -3149
rect -1421 -3153 -1420 -3149
rect -1418 -3153 -1412 -3149
rect -1410 -3153 -1408 -3149
rect -1404 -3153 -1402 -3149
rect -1400 -3153 -1394 -3149
rect -1392 -3153 -1391 -3149
rect -1379 -3153 -1378 -3149
rect -1376 -3153 -1370 -3149
rect -1368 -3153 -1367 -3149
rect -1230 -3153 -1229 -3149
rect -1227 -3153 -1225 -3149
rect -1221 -3153 -1219 -3149
rect -1217 -3153 -1216 -3149
rect -1204 -3153 -1203 -3149
rect -1201 -3153 -1195 -3149
rect -1193 -3153 -1192 -3149
rect -1180 -3153 -1179 -3149
rect -1177 -3153 -1171 -3149
rect -1169 -3153 -1167 -3149
rect -1163 -3153 -1161 -3149
rect -1159 -3153 -1153 -3149
rect -1151 -3153 -1150 -3149
rect -1138 -3153 -1137 -3149
rect -1135 -3153 -1129 -3149
rect -1127 -3153 -1125 -3149
rect -1121 -3153 -1119 -3149
rect -1117 -3153 -1111 -3149
rect -1109 -3153 -1108 -3149
rect -1096 -3153 -1095 -3149
rect -1093 -3153 -1087 -3149
rect -1085 -3153 -1083 -3149
rect -1079 -3153 -1077 -3149
rect -1075 -3153 -1069 -3149
rect -1067 -3153 -1066 -3149
rect -1054 -3153 -1053 -3149
rect -1051 -3153 -1045 -3149
rect -1043 -3153 -1042 -3149
rect -931 -3153 -930 -3149
rect -928 -3153 -926 -3149
rect -922 -3153 -920 -3149
rect -918 -3153 -917 -3149
rect -905 -3153 -904 -3149
rect -902 -3153 -896 -3149
rect -894 -3153 -893 -3149
rect -881 -3153 -880 -3149
rect -878 -3153 -872 -3149
rect -870 -3153 -868 -3149
rect -864 -3153 -862 -3149
rect -860 -3153 -854 -3149
rect -852 -3153 -851 -3149
rect -839 -3153 -838 -3149
rect -836 -3153 -830 -3149
rect -828 -3153 -826 -3149
rect -822 -3153 -820 -3149
rect -818 -3153 -812 -3149
rect -810 -3153 -809 -3149
rect -797 -3153 -796 -3149
rect -794 -3153 -788 -3149
rect -786 -3153 -784 -3149
rect -780 -3153 -778 -3149
rect -776 -3153 -770 -3149
rect -768 -3153 -767 -3149
rect -755 -3153 -754 -3149
rect -752 -3153 -746 -3149
rect -744 -3153 -743 -3149
rect -573 -3153 -572 -3149
rect -570 -3153 -568 -3149
rect -564 -3153 -562 -3149
rect -560 -3153 -559 -3149
rect -547 -3153 -546 -3149
rect -544 -3153 -538 -3149
rect -536 -3153 -535 -3149
rect -523 -3153 -522 -3149
rect -520 -3153 -514 -3149
rect -512 -3153 -510 -3149
rect -506 -3153 -504 -3149
rect -502 -3153 -496 -3149
rect -494 -3153 -493 -3149
rect -481 -3153 -480 -3149
rect -478 -3153 -472 -3149
rect -470 -3153 -468 -3149
rect -464 -3153 -462 -3149
rect -460 -3153 -454 -3149
rect -452 -3153 -451 -3149
rect -439 -3153 -438 -3149
rect -436 -3153 -430 -3149
rect -428 -3153 -426 -3149
rect -422 -3153 -420 -3149
rect -418 -3153 -412 -3149
rect -410 -3153 -409 -3149
rect -397 -3153 -396 -3149
rect -394 -3153 -388 -3149
rect -386 -3153 -385 -3149
rect -215 -3153 -214 -3149
rect -212 -3153 -210 -3149
rect -206 -3153 -204 -3149
rect -202 -3153 -201 -3149
rect -189 -3153 -188 -3149
rect -186 -3153 -180 -3149
rect -178 -3153 -177 -3149
rect -165 -3153 -164 -3149
rect -162 -3153 -156 -3149
rect -154 -3153 -152 -3149
rect -148 -3153 -146 -3149
rect -144 -3153 -138 -3149
rect -136 -3153 -135 -3149
rect -123 -3153 -122 -3149
rect -120 -3153 -114 -3149
rect -112 -3153 -110 -3149
rect -106 -3153 -104 -3149
rect -102 -3153 -96 -3149
rect -94 -3153 -93 -3149
rect -81 -3153 -80 -3149
rect -78 -3153 -72 -3149
rect -70 -3153 -68 -3149
rect -64 -3153 -62 -3149
rect -60 -3153 -54 -3149
rect -52 -3153 -51 -3149
rect -39 -3153 -38 -3149
rect -36 -3153 -30 -3149
rect -28 -3153 -27 -3149
rect 143 -3153 144 -3149
rect 146 -3153 148 -3149
rect 152 -3153 154 -3149
rect 156 -3153 157 -3149
rect 169 -3153 170 -3149
rect 172 -3153 178 -3149
rect 180 -3153 181 -3149
rect 193 -3153 194 -3149
rect 196 -3153 202 -3149
rect 204 -3153 206 -3149
rect 210 -3153 212 -3149
rect 214 -3153 220 -3149
rect 222 -3153 223 -3149
rect 235 -3153 236 -3149
rect 238 -3153 244 -3149
rect 246 -3153 248 -3149
rect 252 -3153 254 -3149
rect 256 -3153 262 -3149
rect 264 -3153 265 -3149
rect 277 -3153 278 -3149
rect 280 -3153 286 -3149
rect 288 -3153 290 -3149
rect 294 -3153 296 -3149
rect 298 -3153 304 -3149
rect 306 -3153 307 -3149
rect 319 -3153 320 -3149
rect 322 -3153 328 -3149
rect 330 -3153 331 -3149
rect 499 -3153 500 -3149
rect 502 -3153 504 -3149
rect 508 -3153 510 -3149
rect 512 -3153 513 -3149
rect 525 -3153 526 -3149
rect 528 -3153 534 -3149
rect 536 -3153 537 -3149
rect 549 -3153 550 -3149
rect 552 -3153 558 -3149
rect 560 -3153 562 -3149
rect 566 -3153 568 -3149
rect 570 -3153 576 -3149
rect 578 -3153 579 -3149
rect 591 -3153 592 -3149
rect 594 -3153 600 -3149
rect 602 -3153 604 -3149
rect 608 -3153 610 -3149
rect 612 -3153 618 -3149
rect 620 -3153 621 -3149
rect 633 -3153 634 -3149
rect 636 -3153 642 -3149
rect 644 -3153 646 -3149
rect 650 -3153 652 -3149
rect 654 -3153 660 -3149
rect 662 -3153 663 -3149
rect 675 -3153 676 -3149
rect 678 -3153 684 -3149
rect 686 -3153 687 -3149
rect 857 -3153 858 -3149
rect 860 -3153 862 -3149
rect 866 -3153 868 -3149
rect 870 -3153 871 -3149
rect 883 -3153 884 -3149
rect 886 -3153 892 -3149
rect 894 -3153 895 -3149
rect 907 -3153 908 -3149
rect 910 -3153 916 -3149
rect 918 -3153 920 -3149
rect 924 -3153 926 -3149
rect 928 -3153 934 -3149
rect 936 -3153 937 -3149
rect 949 -3153 950 -3149
rect 952 -3153 958 -3149
rect 960 -3153 962 -3149
rect 966 -3153 968 -3149
rect 970 -3153 976 -3149
rect 978 -3153 979 -3149
rect 991 -3153 992 -3149
rect 994 -3153 1000 -3149
rect 1002 -3153 1004 -3149
rect 1008 -3153 1010 -3149
rect 1012 -3153 1018 -3149
rect 1020 -3153 1021 -3149
rect 1033 -3153 1034 -3149
rect 1036 -3153 1042 -3149
rect 1044 -3153 1045 -3149
rect 1215 -3153 1216 -3149
rect 1218 -3153 1220 -3149
rect 1224 -3153 1226 -3149
rect 1228 -3153 1229 -3149
rect 1241 -3153 1242 -3149
rect 1244 -3153 1250 -3149
rect 1252 -3153 1253 -3149
rect 1265 -3153 1266 -3149
rect 1268 -3153 1274 -3149
rect 1276 -3153 1278 -3149
rect 1282 -3153 1284 -3149
rect 1286 -3153 1292 -3149
rect 1294 -3153 1295 -3149
rect 1307 -3153 1308 -3149
rect 1310 -3153 1316 -3149
rect 1318 -3153 1320 -3149
rect 1324 -3153 1326 -3149
rect 1328 -3153 1334 -3149
rect 1336 -3153 1337 -3149
rect 1349 -3153 1350 -3149
rect 1352 -3153 1358 -3149
rect 1360 -3153 1362 -3149
rect 1366 -3153 1368 -3149
rect 1370 -3153 1376 -3149
rect 1378 -3153 1379 -3149
rect 1391 -3153 1392 -3149
rect 1394 -3153 1400 -3149
rect 1402 -3153 1403 -3149
rect -1555 -3324 -1554 -3320
rect -1552 -3324 -1550 -3320
rect -1546 -3324 -1544 -3320
rect -1542 -3324 -1541 -3320
rect -1529 -3324 -1528 -3320
rect -1526 -3324 -1520 -3320
rect -1518 -3324 -1517 -3320
rect -1505 -3324 -1504 -3320
rect -1502 -3324 -1496 -3320
rect -1494 -3324 -1492 -3320
rect -1488 -3324 -1486 -3320
rect -1484 -3324 -1478 -3320
rect -1476 -3324 -1475 -3320
rect -1463 -3324 -1462 -3320
rect -1460 -3324 -1454 -3320
rect -1452 -3324 -1450 -3320
rect -1446 -3324 -1444 -3320
rect -1442 -3324 -1436 -3320
rect -1434 -3324 -1433 -3320
rect -1421 -3324 -1420 -3320
rect -1418 -3324 -1412 -3320
rect -1410 -3324 -1408 -3320
rect -1404 -3324 -1402 -3320
rect -1400 -3324 -1394 -3320
rect -1392 -3324 -1391 -3320
rect -1379 -3324 -1378 -3320
rect -1376 -3324 -1370 -3320
rect -1368 -3324 -1367 -3320
rect -1230 -3324 -1229 -3320
rect -1227 -3324 -1225 -3320
rect -1221 -3324 -1219 -3320
rect -1217 -3324 -1216 -3320
rect -1204 -3324 -1203 -3320
rect -1201 -3324 -1195 -3320
rect -1193 -3324 -1192 -3320
rect -1180 -3324 -1179 -3320
rect -1177 -3324 -1171 -3320
rect -1169 -3324 -1167 -3320
rect -1163 -3324 -1161 -3320
rect -1159 -3324 -1153 -3320
rect -1151 -3324 -1150 -3320
rect -1138 -3324 -1137 -3320
rect -1135 -3324 -1129 -3320
rect -1127 -3324 -1125 -3320
rect -1121 -3324 -1119 -3320
rect -1117 -3324 -1111 -3320
rect -1109 -3324 -1108 -3320
rect -1096 -3324 -1095 -3320
rect -1093 -3324 -1087 -3320
rect -1085 -3324 -1083 -3320
rect -1079 -3324 -1077 -3320
rect -1075 -3324 -1069 -3320
rect -1067 -3324 -1066 -3320
rect -1054 -3324 -1053 -3320
rect -1051 -3324 -1045 -3320
rect -1043 -3324 -1042 -3320
rect -931 -3324 -930 -3320
rect -928 -3324 -926 -3320
rect -922 -3324 -920 -3320
rect -918 -3324 -917 -3320
rect -905 -3324 -904 -3320
rect -902 -3324 -896 -3320
rect -894 -3324 -893 -3320
rect -881 -3324 -880 -3320
rect -878 -3324 -872 -3320
rect -870 -3324 -868 -3320
rect -864 -3324 -862 -3320
rect -860 -3324 -854 -3320
rect -852 -3324 -851 -3320
rect -839 -3324 -838 -3320
rect -836 -3324 -830 -3320
rect -828 -3324 -826 -3320
rect -822 -3324 -820 -3320
rect -818 -3324 -812 -3320
rect -810 -3324 -809 -3320
rect -797 -3324 -796 -3320
rect -794 -3324 -788 -3320
rect -786 -3324 -784 -3320
rect -780 -3324 -778 -3320
rect -776 -3324 -770 -3320
rect -768 -3324 -767 -3320
rect -755 -3324 -754 -3320
rect -752 -3324 -746 -3320
rect -744 -3324 -743 -3320
rect -573 -3324 -572 -3320
rect -570 -3324 -568 -3320
rect -564 -3324 -562 -3320
rect -560 -3324 -559 -3320
rect -547 -3324 -546 -3320
rect -544 -3324 -538 -3320
rect -536 -3324 -535 -3320
rect -523 -3324 -522 -3320
rect -520 -3324 -514 -3320
rect -512 -3324 -510 -3320
rect -506 -3324 -504 -3320
rect -502 -3324 -496 -3320
rect -494 -3324 -493 -3320
rect -481 -3324 -480 -3320
rect -478 -3324 -472 -3320
rect -470 -3324 -468 -3320
rect -464 -3324 -462 -3320
rect -460 -3324 -454 -3320
rect -452 -3324 -451 -3320
rect -439 -3324 -438 -3320
rect -436 -3324 -430 -3320
rect -428 -3324 -426 -3320
rect -422 -3324 -420 -3320
rect -418 -3324 -412 -3320
rect -410 -3324 -409 -3320
rect -397 -3324 -396 -3320
rect -394 -3324 -388 -3320
rect -386 -3324 -385 -3320
rect -215 -3324 -214 -3320
rect -212 -3324 -210 -3320
rect -206 -3324 -204 -3320
rect -202 -3324 -201 -3320
rect -189 -3324 -188 -3320
rect -186 -3324 -180 -3320
rect -178 -3324 -177 -3320
rect -165 -3324 -164 -3320
rect -162 -3324 -156 -3320
rect -154 -3324 -152 -3320
rect -148 -3324 -146 -3320
rect -144 -3324 -138 -3320
rect -136 -3324 -135 -3320
rect -123 -3324 -122 -3320
rect -120 -3324 -114 -3320
rect -112 -3324 -110 -3320
rect -106 -3324 -104 -3320
rect -102 -3324 -96 -3320
rect -94 -3324 -93 -3320
rect -81 -3324 -80 -3320
rect -78 -3324 -72 -3320
rect -70 -3324 -68 -3320
rect -64 -3324 -62 -3320
rect -60 -3324 -54 -3320
rect -52 -3324 -51 -3320
rect -39 -3324 -38 -3320
rect -36 -3324 -30 -3320
rect -28 -3324 -27 -3320
rect 143 -3324 144 -3320
rect 146 -3324 148 -3320
rect 152 -3324 154 -3320
rect 156 -3324 157 -3320
rect 169 -3324 170 -3320
rect 172 -3324 178 -3320
rect 180 -3324 181 -3320
rect 193 -3324 194 -3320
rect 196 -3324 202 -3320
rect 204 -3324 206 -3320
rect 210 -3324 212 -3320
rect 214 -3324 220 -3320
rect 222 -3324 223 -3320
rect 235 -3324 236 -3320
rect 238 -3324 244 -3320
rect 246 -3324 248 -3320
rect 252 -3324 254 -3320
rect 256 -3324 262 -3320
rect 264 -3324 265 -3320
rect 277 -3324 278 -3320
rect 280 -3324 286 -3320
rect 288 -3324 290 -3320
rect 294 -3324 296 -3320
rect 298 -3324 304 -3320
rect 306 -3324 307 -3320
rect 319 -3324 320 -3320
rect 322 -3324 328 -3320
rect 330 -3324 331 -3320
rect 499 -3324 500 -3320
rect 502 -3324 504 -3320
rect 508 -3324 510 -3320
rect 512 -3324 513 -3320
rect 525 -3324 526 -3320
rect 528 -3324 534 -3320
rect 536 -3324 537 -3320
rect 549 -3324 550 -3320
rect 552 -3324 558 -3320
rect 560 -3324 562 -3320
rect 566 -3324 568 -3320
rect 570 -3324 576 -3320
rect 578 -3324 579 -3320
rect 591 -3324 592 -3320
rect 594 -3324 600 -3320
rect 602 -3324 604 -3320
rect 608 -3324 610 -3320
rect 612 -3324 618 -3320
rect 620 -3324 621 -3320
rect 633 -3324 634 -3320
rect 636 -3324 642 -3320
rect 644 -3324 646 -3320
rect 650 -3324 652 -3320
rect 654 -3324 660 -3320
rect 662 -3324 663 -3320
rect 675 -3324 676 -3320
rect 678 -3324 684 -3320
rect 686 -3324 687 -3320
rect 857 -3324 858 -3320
rect 860 -3324 862 -3320
rect 866 -3324 868 -3320
rect 870 -3324 871 -3320
rect 883 -3324 884 -3320
rect 886 -3324 892 -3320
rect 894 -3324 895 -3320
rect 907 -3324 908 -3320
rect 910 -3324 916 -3320
rect 918 -3324 920 -3320
rect 924 -3324 926 -3320
rect 928 -3324 934 -3320
rect 936 -3324 937 -3320
rect 949 -3324 950 -3320
rect 952 -3324 958 -3320
rect 960 -3324 962 -3320
rect 966 -3324 968 -3320
rect 970 -3324 976 -3320
rect 978 -3324 979 -3320
rect 991 -3324 992 -3320
rect 994 -3324 1000 -3320
rect 1002 -3324 1004 -3320
rect 1008 -3324 1010 -3320
rect 1012 -3324 1018 -3320
rect 1020 -3324 1021 -3320
rect 1033 -3324 1034 -3320
rect 1036 -3324 1042 -3320
rect 1044 -3324 1045 -3320
rect 1215 -3324 1216 -3320
rect 1218 -3324 1220 -3320
rect 1224 -3324 1226 -3320
rect 1228 -3324 1229 -3320
rect 1241 -3324 1242 -3320
rect 1244 -3324 1250 -3320
rect 1252 -3324 1253 -3320
rect 1265 -3324 1266 -3320
rect 1268 -3324 1274 -3320
rect 1276 -3324 1278 -3320
rect 1282 -3324 1284 -3320
rect 1286 -3324 1292 -3320
rect 1294 -3324 1295 -3320
rect 1307 -3324 1308 -3320
rect 1310 -3324 1316 -3320
rect 1318 -3324 1320 -3320
rect 1324 -3324 1326 -3320
rect 1328 -3324 1334 -3320
rect 1336 -3324 1337 -3320
rect 1349 -3324 1350 -3320
rect 1352 -3324 1358 -3320
rect 1360 -3324 1362 -3320
rect 1366 -3324 1368 -3320
rect 1370 -3324 1376 -3320
rect 1378 -3324 1379 -3320
rect 1391 -3324 1392 -3320
rect 1394 -3324 1400 -3320
rect 1402 -3324 1403 -3320
rect -1305 -3435 -1304 -3431
rect -1302 -3435 -1296 -3431
rect -1294 -3435 -1292 -3431
rect -1288 -3435 -1286 -3431
rect -1284 -3435 -1283 -3431
rect -931 -3435 -930 -3431
rect -928 -3435 -922 -3431
rect -920 -3435 -918 -3431
rect -914 -3435 -912 -3431
rect -910 -3435 -909 -3431
rect -573 -3435 -572 -3431
rect -570 -3435 -564 -3431
rect -562 -3435 -560 -3431
rect -556 -3435 -554 -3431
rect -552 -3435 -551 -3431
rect -215 -3435 -214 -3431
rect -212 -3435 -206 -3431
rect -204 -3435 -202 -3431
rect -198 -3435 -196 -3431
rect -194 -3435 -193 -3431
rect 143 -3435 144 -3431
rect 146 -3435 152 -3431
rect 154 -3435 156 -3431
rect 160 -3435 162 -3431
rect 164 -3435 165 -3431
rect 499 -3435 500 -3431
rect 502 -3435 508 -3431
rect 510 -3435 512 -3431
rect 516 -3435 518 -3431
rect 520 -3435 521 -3431
rect 857 -3435 858 -3431
rect 860 -3435 866 -3431
rect 868 -3435 870 -3431
rect 874 -3435 876 -3431
rect 878 -3435 879 -3431
rect 1215 -3435 1216 -3431
rect 1218 -3435 1224 -3431
rect 1226 -3435 1228 -3431
rect 1232 -3435 1234 -3431
rect 1236 -3435 1237 -3431
rect -1230 -3594 -1229 -3590
rect -1227 -3594 -1225 -3590
rect -1221 -3594 -1219 -3590
rect -1217 -3594 -1216 -3590
rect -1204 -3594 -1203 -3590
rect -1201 -3594 -1199 -3590
rect -1195 -3594 -1193 -3590
rect -1191 -3594 -1185 -3590
rect -1183 -3594 -1181 -3590
rect -1177 -3594 -1175 -3590
rect -1173 -3594 -1172 -3590
rect -1160 -3594 -1159 -3590
rect -1157 -3594 -1151 -3590
rect -1149 -3594 -1147 -3590
rect -1143 -3594 -1141 -3590
rect -1139 -3594 -1138 -3590
rect -931 -3594 -930 -3590
rect -928 -3594 -926 -3590
rect -922 -3594 -920 -3590
rect -918 -3594 -917 -3590
rect -905 -3594 -904 -3590
rect -902 -3594 -900 -3590
rect -896 -3594 -894 -3590
rect -892 -3594 -891 -3590
rect -879 -3594 -878 -3590
rect -876 -3594 -875 -3590
rect -871 -3594 -868 -3590
rect -866 -3594 -860 -3590
rect -858 -3594 -857 -3590
rect -853 -3594 -850 -3590
rect -848 -3594 -847 -3590
rect -835 -3594 -834 -3590
rect -832 -3594 -826 -3590
rect -824 -3594 -822 -3590
rect -818 -3594 -816 -3590
rect -814 -3594 -813 -3590
rect -801 -3594 -800 -3590
rect -798 -3594 -796 -3590
rect -792 -3594 -790 -3590
rect -788 -3594 -782 -3590
rect -780 -3594 -778 -3590
rect -774 -3594 -772 -3590
rect -770 -3594 -769 -3590
rect -757 -3594 -756 -3590
rect -754 -3594 -748 -3590
rect -746 -3594 -745 -3590
rect -733 -3594 -732 -3590
rect -730 -3594 -725 -3590
rect -721 -3594 -716 -3590
rect -714 -3594 -713 -3590
rect -709 -3594 -708 -3590
rect -706 -3594 -704 -3590
rect -700 -3594 -698 -3590
rect -696 -3594 -695 -3590
rect -573 -3594 -572 -3590
rect -570 -3594 -568 -3590
rect -564 -3594 -562 -3590
rect -560 -3594 -559 -3590
rect -547 -3594 -546 -3590
rect -544 -3594 -542 -3590
rect -538 -3594 -536 -3590
rect -534 -3594 -533 -3590
rect -521 -3594 -520 -3590
rect -518 -3594 -517 -3590
rect -513 -3594 -510 -3590
rect -508 -3594 -502 -3590
rect -500 -3594 -499 -3590
rect -495 -3594 -492 -3590
rect -490 -3594 -489 -3590
rect -477 -3594 -476 -3590
rect -474 -3594 -468 -3590
rect -466 -3594 -464 -3590
rect -460 -3594 -458 -3590
rect -456 -3594 -455 -3590
rect -443 -3594 -442 -3590
rect -440 -3594 -438 -3590
rect -434 -3594 -432 -3590
rect -430 -3594 -424 -3590
rect -422 -3594 -420 -3590
rect -416 -3594 -414 -3590
rect -412 -3594 -411 -3590
rect -399 -3594 -398 -3590
rect -396 -3594 -390 -3590
rect -388 -3594 -387 -3590
rect -375 -3594 -374 -3590
rect -372 -3594 -367 -3590
rect -363 -3594 -358 -3590
rect -356 -3594 -355 -3590
rect -351 -3594 -350 -3590
rect -348 -3594 -346 -3590
rect -342 -3594 -340 -3590
rect -338 -3594 -337 -3590
rect -215 -3594 -214 -3590
rect -212 -3594 -210 -3590
rect -206 -3594 -204 -3590
rect -202 -3594 -201 -3590
rect -189 -3594 -188 -3590
rect -186 -3594 -184 -3590
rect -180 -3594 -178 -3590
rect -176 -3594 -175 -3590
rect -163 -3594 -162 -3590
rect -160 -3594 -159 -3590
rect -155 -3594 -152 -3590
rect -150 -3594 -144 -3590
rect -142 -3594 -141 -3590
rect -137 -3594 -134 -3590
rect -132 -3594 -131 -3590
rect -119 -3594 -118 -3590
rect -116 -3594 -110 -3590
rect -108 -3594 -106 -3590
rect -102 -3594 -100 -3590
rect -98 -3594 -97 -3590
rect -85 -3594 -84 -3590
rect -82 -3594 -80 -3590
rect -76 -3594 -74 -3590
rect -72 -3594 -66 -3590
rect -64 -3594 -62 -3590
rect -58 -3594 -56 -3590
rect -54 -3594 -53 -3590
rect -41 -3594 -40 -3590
rect -38 -3594 -32 -3590
rect -30 -3594 -29 -3590
rect -17 -3594 -16 -3590
rect -14 -3594 -9 -3590
rect -5 -3594 0 -3590
rect 2 -3594 3 -3590
rect 7 -3594 8 -3590
rect 10 -3594 12 -3590
rect 16 -3594 18 -3590
rect 20 -3594 21 -3590
rect 143 -3594 144 -3590
rect 146 -3594 148 -3590
rect 152 -3594 154 -3590
rect 156 -3594 157 -3590
rect 169 -3594 170 -3590
rect 172 -3594 174 -3590
rect 178 -3594 180 -3590
rect 182 -3594 183 -3590
rect 195 -3594 196 -3590
rect 198 -3594 199 -3590
rect 203 -3594 206 -3590
rect 208 -3594 214 -3590
rect 216 -3594 217 -3590
rect 221 -3594 224 -3590
rect 226 -3594 227 -3590
rect 239 -3594 240 -3590
rect 242 -3594 248 -3590
rect 250 -3594 252 -3590
rect 256 -3594 258 -3590
rect 260 -3594 261 -3590
rect 273 -3594 274 -3590
rect 276 -3594 278 -3590
rect 282 -3594 284 -3590
rect 286 -3594 292 -3590
rect 294 -3594 296 -3590
rect 300 -3594 302 -3590
rect 304 -3594 305 -3590
rect 317 -3594 318 -3590
rect 320 -3594 326 -3590
rect 328 -3594 329 -3590
rect 341 -3594 342 -3590
rect 344 -3594 349 -3590
rect 353 -3594 358 -3590
rect 360 -3594 361 -3590
rect 365 -3594 366 -3590
rect 368 -3594 370 -3590
rect 374 -3594 376 -3590
rect 378 -3594 379 -3590
rect 499 -3594 500 -3590
rect 502 -3594 504 -3590
rect 508 -3594 510 -3590
rect 512 -3594 513 -3590
rect 525 -3594 526 -3590
rect 528 -3594 530 -3590
rect 534 -3594 536 -3590
rect 538 -3594 539 -3590
rect 551 -3594 552 -3590
rect 554 -3594 555 -3590
rect 559 -3594 562 -3590
rect 564 -3594 570 -3590
rect 572 -3594 573 -3590
rect 577 -3594 580 -3590
rect 582 -3594 583 -3590
rect 595 -3594 596 -3590
rect 598 -3594 604 -3590
rect 606 -3594 608 -3590
rect 612 -3594 614 -3590
rect 616 -3594 617 -3590
rect 629 -3594 630 -3590
rect 632 -3594 634 -3590
rect 638 -3594 640 -3590
rect 642 -3594 648 -3590
rect 650 -3594 652 -3590
rect 656 -3594 658 -3590
rect 660 -3594 661 -3590
rect 673 -3594 674 -3590
rect 676 -3594 682 -3590
rect 684 -3594 685 -3590
rect 697 -3594 698 -3590
rect 700 -3594 705 -3590
rect 709 -3594 714 -3590
rect 716 -3594 717 -3590
rect 721 -3594 722 -3590
rect 724 -3594 726 -3590
rect 730 -3594 732 -3590
rect 734 -3594 735 -3590
rect 857 -3594 858 -3590
rect 860 -3594 862 -3590
rect 866 -3594 868 -3590
rect 870 -3594 871 -3590
rect 883 -3594 884 -3590
rect 886 -3594 888 -3590
rect 892 -3594 894 -3590
rect 896 -3594 897 -3590
rect 909 -3594 910 -3590
rect 912 -3594 913 -3590
rect 917 -3594 920 -3590
rect 922 -3594 928 -3590
rect 930 -3594 931 -3590
rect 935 -3594 938 -3590
rect 940 -3594 941 -3590
rect 953 -3594 954 -3590
rect 956 -3594 962 -3590
rect 964 -3594 966 -3590
rect 970 -3594 972 -3590
rect 974 -3594 975 -3590
rect 987 -3594 988 -3590
rect 990 -3594 992 -3590
rect 996 -3594 998 -3590
rect 1000 -3594 1006 -3590
rect 1008 -3594 1010 -3590
rect 1014 -3594 1016 -3590
rect 1018 -3594 1019 -3590
rect 1031 -3594 1032 -3590
rect 1034 -3594 1040 -3590
rect 1042 -3594 1043 -3590
rect 1055 -3594 1056 -3590
rect 1058 -3594 1063 -3590
rect 1067 -3594 1072 -3590
rect 1074 -3594 1075 -3590
rect 1079 -3594 1080 -3590
rect 1082 -3594 1084 -3590
rect 1088 -3594 1090 -3590
rect 1092 -3594 1093 -3590
rect 1215 -3594 1216 -3590
rect 1218 -3594 1220 -3590
rect 1224 -3594 1226 -3590
rect 1228 -3594 1229 -3590
rect 1241 -3594 1242 -3590
rect 1244 -3594 1246 -3590
rect 1250 -3594 1252 -3590
rect 1254 -3594 1255 -3590
rect 1267 -3594 1268 -3590
rect 1270 -3594 1271 -3590
rect 1275 -3594 1278 -3590
rect 1280 -3594 1286 -3590
rect 1288 -3594 1289 -3590
rect 1293 -3594 1296 -3590
rect 1298 -3594 1299 -3590
rect 1311 -3594 1312 -3590
rect 1314 -3594 1320 -3590
rect 1322 -3594 1324 -3590
rect 1328 -3594 1330 -3590
rect 1332 -3594 1333 -3590
rect 1345 -3594 1346 -3590
rect 1348 -3594 1350 -3590
rect 1354 -3594 1356 -3590
rect 1358 -3594 1364 -3590
rect 1366 -3594 1368 -3590
rect 1372 -3594 1374 -3590
rect 1376 -3594 1377 -3590
rect 1389 -3594 1390 -3590
rect 1392 -3594 1398 -3590
rect 1400 -3594 1401 -3590
rect 1413 -3594 1414 -3590
rect 1416 -3594 1421 -3590
rect 1425 -3594 1430 -3590
rect 1432 -3594 1433 -3590
rect 1437 -3594 1438 -3590
rect 1440 -3594 1442 -3590
rect 1446 -3594 1448 -3590
rect 1450 -3594 1451 -3590
rect -1818 -3724 -1817 -3720
rect -1815 -3724 -1813 -3720
rect -1809 -3724 -1807 -3720
rect -1805 -3724 -1804 -3720
rect -1792 -3724 -1791 -3720
rect -1789 -3724 -1783 -3720
rect -1781 -3724 -1780 -3720
rect -1768 -3724 -1767 -3720
rect -1765 -3724 -1759 -3720
rect -1757 -3724 -1755 -3720
rect -1751 -3724 -1749 -3720
rect -1747 -3724 -1741 -3720
rect -1739 -3724 -1738 -3720
rect -1726 -3724 -1725 -3720
rect -1723 -3724 -1717 -3720
rect -1715 -3724 -1713 -3720
rect -1709 -3724 -1707 -3720
rect -1705 -3724 -1699 -3720
rect -1697 -3724 -1696 -3720
rect -1684 -3724 -1683 -3720
rect -1681 -3724 -1675 -3720
rect -1673 -3724 -1671 -3720
rect -1667 -3724 -1665 -3720
rect -1663 -3724 -1657 -3720
rect -1655 -3724 -1654 -3720
rect -1642 -3724 -1641 -3720
rect -1639 -3724 -1633 -3720
rect -1631 -3724 -1630 -3720
rect -1555 -3724 -1554 -3720
rect -1552 -3724 -1550 -3720
rect -1546 -3724 -1544 -3720
rect -1542 -3724 -1541 -3720
rect -1529 -3724 -1528 -3720
rect -1526 -3724 -1520 -3720
rect -1518 -3724 -1517 -3720
rect -1505 -3724 -1504 -3720
rect -1502 -3724 -1496 -3720
rect -1494 -3724 -1492 -3720
rect -1488 -3724 -1486 -3720
rect -1484 -3724 -1478 -3720
rect -1476 -3724 -1475 -3720
rect -1463 -3724 -1462 -3720
rect -1460 -3724 -1454 -3720
rect -1452 -3724 -1450 -3720
rect -1446 -3724 -1444 -3720
rect -1442 -3724 -1436 -3720
rect -1434 -3724 -1433 -3720
rect -1421 -3724 -1420 -3720
rect -1418 -3724 -1412 -3720
rect -1410 -3724 -1408 -3720
rect -1404 -3724 -1402 -3720
rect -1400 -3724 -1394 -3720
rect -1392 -3724 -1391 -3720
rect -1379 -3724 -1378 -3720
rect -1376 -3724 -1370 -3720
rect -1368 -3724 -1367 -3720
rect -1230 -3724 -1229 -3720
rect -1227 -3724 -1225 -3720
rect -1221 -3724 -1219 -3720
rect -1217 -3724 -1216 -3720
rect -1204 -3724 -1203 -3720
rect -1201 -3724 -1195 -3720
rect -1193 -3724 -1192 -3720
rect -1180 -3724 -1179 -3720
rect -1177 -3724 -1171 -3720
rect -1169 -3724 -1167 -3720
rect -1163 -3724 -1161 -3720
rect -1159 -3724 -1153 -3720
rect -1151 -3724 -1150 -3720
rect -1138 -3724 -1137 -3720
rect -1135 -3724 -1129 -3720
rect -1127 -3724 -1125 -3720
rect -1121 -3724 -1119 -3720
rect -1117 -3724 -1111 -3720
rect -1109 -3724 -1108 -3720
rect -1096 -3724 -1095 -3720
rect -1093 -3724 -1087 -3720
rect -1085 -3724 -1083 -3720
rect -1079 -3724 -1077 -3720
rect -1075 -3724 -1069 -3720
rect -1067 -3724 -1066 -3720
rect -1054 -3724 -1053 -3720
rect -1051 -3724 -1045 -3720
rect -1043 -3724 -1042 -3720
rect -930 -3724 -929 -3720
rect -927 -3724 -925 -3720
rect -921 -3724 -919 -3720
rect -917 -3724 -916 -3720
rect -904 -3724 -903 -3720
rect -901 -3724 -895 -3720
rect -893 -3724 -892 -3720
rect -880 -3724 -879 -3720
rect -877 -3724 -871 -3720
rect -869 -3724 -867 -3720
rect -863 -3724 -861 -3720
rect -859 -3724 -853 -3720
rect -851 -3724 -850 -3720
rect -838 -3724 -837 -3720
rect -835 -3724 -829 -3720
rect -827 -3724 -825 -3720
rect -821 -3724 -819 -3720
rect -817 -3724 -811 -3720
rect -809 -3724 -808 -3720
rect -796 -3724 -795 -3720
rect -793 -3724 -787 -3720
rect -785 -3724 -783 -3720
rect -779 -3724 -777 -3720
rect -775 -3724 -769 -3720
rect -767 -3724 -766 -3720
rect -754 -3724 -753 -3720
rect -751 -3724 -745 -3720
rect -743 -3724 -742 -3720
rect -573 -3724 -572 -3720
rect -570 -3724 -568 -3720
rect -564 -3724 -562 -3720
rect -560 -3724 -559 -3720
rect -547 -3724 -546 -3720
rect -544 -3724 -538 -3720
rect -536 -3724 -535 -3720
rect -523 -3724 -522 -3720
rect -520 -3724 -514 -3720
rect -512 -3724 -510 -3720
rect -506 -3724 -504 -3720
rect -502 -3724 -496 -3720
rect -494 -3724 -493 -3720
rect -481 -3724 -480 -3720
rect -478 -3724 -472 -3720
rect -470 -3724 -468 -3720
rect -464 -3724 -462 -3720
rect -460 -3724 -454 -3720
rect -452 -3724 -451 -3720
rect -439 -3724 -438 -3720
rect -436 -3724 -430 -3720
rect -428 -3724 -426 -3720
rect -422 -3724 -420 -3720
rect -418 -3724 -412 -3720
rect -410 -3724 -409 -3720
rect -397 -3724 -396 -3720
rect -394 -3724 -388 -3720
rect -386 -3724 -385 -3720
rect -215 -3724 -214 -3720
rect -212 -3724 -210 -3720
rect -206 -3724 -204 -3720
rect -202 -3724 -201 -3720
rect -189 -3724 -188 -3720
rect -186 -3724 -180 -3720
rect -178 -3724 -177 -3720
rect -165 -3724 -164 -3720
rect -162 -3724 -156 -3720
rect -154 -3724 -152 -3720
rect -148 -3724 -146 -3720
rect -144 -3724 -138 -3720
rect -136 -3724 -135 -3720
rect -123 -3724 -122 -3720
rect -120 -3724 -114 -3720
rect -112 -3724 -110 -3720
rect -106 -3724 -104 -3720
rect -102 -3724 -96 -3720
rect -94 -3724 -93 -3720
rect -81 -3724 -80 -3720
rect -78 -3724 -72 -3720
rect -70 -3724 -68 -3720
rect -64 -3724 -62 -3720
rect -60 -3724 -54 -3720
rect -52 -3724 -51 -3720
rect -39 -3724 -38 -3720
rect -36 -3724 -30 -3720
rect -28 -3724 -27 -3720
rect -1555 -3895 -1554 -3891
rect -1552 -3895 -1550 -3891
rect -1546 -3895 -1544 -3891
rect -1542 -3895 -1541 -3891
rect -1529 -3895 -1528 -3891
rect -1526 -3895 -1520 -3891
rect -1518 -3895 -1517 -3891
rect -1505 -3895 -1504 -3891
rect -1502 -3895 -1496 -3891
rect -1494 -3895 -1492 -3891
rect -1488 -3895 -1486 -3891
rect -1484 -3895 -1478 -3891
rect -1476 -3895 -1475 -3891
rect -1463 -3895 -1462 -3891
rect -1460 -3895 -1454 -3891
rect -1452 -3895 -1450 -3891
rect -1446 -3895 -1444 -3891
rect -1442 -3895 -1436 -3891
rect -1434 -3895 -1433 -3891
rect -1421 -3895 -1420 -3891
rect -1418 -3895 -1412 -3891
rect -1410 -3895 -1408 -3891
rect -1404 -3895 -1402 -3891
rect -1400 -3895 -1394 -3891
rect -1392 -3895 -1391 -3891
rect -1379 -3895 -1378 -3891
rect -1376 -3895 -1370 -3891
rect -1368 -3895 -1367 -3891
rect -1230 -3895 -1229 -3891
rect -1227 -3895 -1225 -3891
rect -1221 -3895 -1219 -3891
rect -1217 -3895 -1216 -3891
rect -1204 -3895 -1203 -3891
rect -1201 -3895 -1195 -3891
rect -1193 -3895 -1192 -3891
rect -1180 -3895 -1179 -3891
rect -1177 -3895 -1171 -3891
rect -1169 -3895 -1167 -3891
rect -1163 -3895 -1161 -3891
rect -1159 -3895 -1153 -3891
rect -1151 -3895 -1150 -3891
rect -1138 -3895 -1137 -3891
rect -1135 -3895 -1129 -3891
rect -1127 -3895 -1125 -3891
rect -1121 -3895 -1119 -3891
rect -1117 -3895 -1111 -3891
rect -1109 -3895 -1108 -3891
rect -1096 -3895 -1095 -3891
rect -1093 -3895 -1087 -3891
rect -1085 -3895 -1083 -3891
rect -1079 -3895 -1077 -3891
rect -1075 -3895 -1069 -3891
rect -1067 -3895 -1066 -3891
rect -1054 -3895 -1053 -3891
rect -1051 -3895 -1045 -3891
rect -1043 -3895 -1042 -3891
rect -930 -3895 -929 -3891
rect -927 -3895 -925 -3891
rect -921 -3895 -919 -3891
rect -917 -3895 -916 -3891
rect -904 -3895 -903 -3891
rect -901 -3895 -895 -3891
rect -893 -3895 -892 -3891
rect -880 -3895 -879 -3891
rect -877 -3895 -871 -3891
rect -869 -3895 -867 -3891
rect -863 -3895 -861 -3891
rect -859 -3895 -853 -3891
rect -851 -3895 -850 -3891
rect -838 -3895 -837 -3891
rect -835 -3895 -829 -3891
rect -827 -3895 -825 -3891
rect -821 -3895 -819 -3891
rect -817 -3895 -811 -3891
rect -809 -3895 -808 -3891
rect -796 -3895 -795 -3891
rect -793 -3895 -787 -3891
rect -785 -3895 -783 -3891
rect -779 -3895 -777 -3891
rect -775 -3895 -769 -3891
rect -767 -3895 -766 -3891
rect -754 -3895 -753 -3891
rect -751 -3895 -745 -3891
rect -743 -3895 -742 -3891
rect -573 -3895 -572 -3891
rect -570 -3895 -568 -3891
rect -564 -3895 -562 -3891
rect -560 -3895 -559 -3891
rect -547 -3895 -546 -3891
rect -544 -3895 -538 -3891
rect -536 -3895 -535 -3891
rect -523 -3895 -522 -3891
rect -520 -3895 -514 -3891
rect -512 -3895 -510 -3891
rect -506 -3895 -504 -3891
rect -502 -3895 -496 -3891
rect -494 -3895 -493 -3891
rect -481 -3895 -480 -3891
rect -478 -3895 -472 -3891
rect -470 -3895 -468 -3891
rect -464 -3895 -462 -3891
rect -460 -3895 -454 -3891
rect -452 -3895 -451 -3891
rect -439 -3895 -438 -3891
rect -436 -3895 -430 -3891
rect -428 -3895 -426 -3891
rect -422 -3895 -420 -3891
rect -418 -3895 -412 -3891
rect -410 -3895 -409 -3891
rect -397 -3895 -396 -3891
rect -394 -3895 -388 -3891
rect -386 -3895 -385 -3891
rect -215 -3895 -214 -3891
rect -212 -3895 -210 -3891
rect -206 -3895 -204 -3891
rect -202 -3895 -201 -3891
rect -189 -3895 -188 -3891
rect -186 -3895 -180 -3891
rect -178 -3895 -177 -3891
rect -165 -3895 -164 -3891
rect -162 -3895 -156 -3891
rect -154 -3895 -152 -3891
rect -148 -3895 -146 -3891
rect -144 -3895 -138 -3891
rect -136 -3895 -135 -3891
rect -123 -3895 -122 -3891
rect -120 -3895 -114 -3891
rect -112 -3895 -110 -3891
rect -106 -3895 -104 -3891
rect -102 -3895 -96 -3891
rect -94 -3895 -93 -3891
rect -81 -3895 -80 -3891
rect -78 -3895 -72 -3891
rect -70 -3895 -68 -3891
rect -64 -3895 -62 -3891
rect -60 -3895 -54 -3891
rect -52 -3895 -51 -3891
rect -39 -3895 -38 -3891
rect -36 -3895 -30 -3891
rect -28 -3895 -27 -3891
rect 143 -3895 144 -3891
rect 146 -3895 148 -3891
rect 152 -3895 154 -3891
rect 156 -3895 157 -3891
rect 169 -3895 170 -3891
rect 172 -3895 178 -3891
rect 180 -3895 181 -3891
rect 193 -3895 194 -3891
rect 196 -3895 202 -3891
rect 204 -3895 206 -3891
rect 210 -3895 212 -3891
rect 214 -3895 220 -3891
rect 222 -3895 223 -3891
rect 235 -3895 236 -3891
rect 238 -3895 244 -3891
rect 246 -3895 248 -3891
rect 252 -3895 254 -3891
rect 256 -3895 262 -3891
rect 264 -3895 265 -3891
rect 277 -3895 278 -3891
rect 280 -3895 286 -3891
rect 288 -3895 290 -3891
rect 294 -3895 296 -3891
rect 298 -3895 304 -3891
rect 306 -3895 307 -3891
rect 319 -3895 320 -3891
rect 322 -3895 328 -3891
rect 330 -3895 331 -3891
rect 499 -3895 500 -3891
rect 502 -3895 504 -3891
rect 508 -3895 510 -3891
rect 512 -3895 513 -3891
rect 525 -3895 526 -3891
rect 528 -3895 534 -3891
rect 536 -3895 537 -3891
rect 549 -3895 550 -3891
rect 552 -3895 558 -3891
rect 560 -3895 562 -3891
rect 566 -3895 568 -3891
rect 570 -3895 576 -3891
rect 578 -3895 579 -3891
rect 591 -3895 592 -3891
rect 594 -3895 600 -3891
rect 602 -3895 604 -3891
rect 608 -3895 610 -3891
rect 612 -3895 618 -3891
rect 620 -3895 621 -3891
rect 633 -3895 634 -3891
rect 636 -3895 642 -3891
rect 644 -3895 646 -3891
rect 650 -3895 652 -3891
rect 654 -3895 660 -3891
rect 662 -3895 663 -3891
rect 675 -3895 676 -3891
rect 678 -3895 684 -3891
rect 686 -3895 687 -3891
rect 857 -3895 858 -3891
rect 860 -3895 862 -3891
rect 866 -3895 868 -3891
rect 870 -3895 871 -3891
rect 883 -3895 884 -3891
rect 886 -3895 892 -3891
rect 894 -3895 895 -3891
rect 907 -3895 908 -3891
rect 910 -3895 916 -3891
rect 918 -3895 920 -3891
rect 924 -3895 926 -3891
rect 928 -3895 934 -3891
rect 936 -3895 937 -3891
rect 949 -3895 950 -3891
rect 952 -3895 958 -3891
rect 960 -3895 962 -3891
rect 966 -3895 968 -3891
rect 970 -3895 976 -3891
rect 978 -3895 979 -3891
rect 991 -3895 992 -3891
rect 994 -3895 1000 -3891
rect 1002 -3895 1004 -3891
rect 1008 -3895 1010 -3891
rect 1012 -3895 1018 -3891
rect 1020 -3895 1021 -3891
rect 1033 -3895 1034 -3891
rect 1036 -3895 1042 -3891
rect 1044 -3895 1045 -3891
rect 1215 -3895 1216 -3891
rect 1218 -3895 1220 -3891
rect 1224 -3895 1226 -3891
rect 1228 -3895 1229 -3891
rect 1241 -3895 1242 -3891
rect 1244 -3895 1250 -3891
rect 1252 -3895 1253 -3891
rect 1265 -3895 1266 -3891
rect 1268 -3895 1274 -3891
rect 1276 -3895 1278 -3891
rect 1282 -3895 1284 -3891
rect 1286 -3895 1292 -3891
rect 1294 -3895 1295 -3891
rect 1307 -3895 1308 -3891
rect 1310 -3895 1316 -3891
rect 1318 -3895 1320 -3891
rect 1324 -3895 1326 -3891
rect 1328 -3895 1334 -3891
rect 1336 -3895 1337 -3891
rect 1349 -3895 1350 -3891
rect 1352 -3895 1358 -3891
rect 1360 -3895 1362 -3891
rect 1366 -3895 1368 -3891
rect 1370 -3895 1376 -3891
rect 1378 -3895 1379 -3891
rect 1391 -3895 1392 -3891
rect 1394 -3895 1400 -3891
rect 1402 -3895 1403 -3891
rect -1555 -4070 -1554 -4066
rect -1552 -4070 -1550 -4066
rect -1546 -4070 -1544 -4066
rect -1542 -4070 -1541 -4066
rect -1529 -4070 -1528 -4066
rect -1526 -4070 -1520 -4066
rect -1518 -4070 -1517 -4066
rect -1505 -4070 -1504 -4066
rect -1502 -4070 -1496 -4066
rect -1494 -4070 -1492 -4066
rect -1488 -4070 -1486 -4066
rect -1484 -4070 -1478 -4066
rect -1476 -4070 -1475 -4066
rect -1463 -4070 -1462 -4066
rect -1460 -4070 -1454 -4066
rect -1452 -4070 -1450 -4066
rect -1446 -4070 -1444 -4066
rect -1442 -4070 -1436 -4066
rect -1434 -4070 -1433 -4066
rect -1421 -4070 -1420 -4066
rect -1418 -4070 -1412 -4066
rect -1410 -4070 -1408 -4066
rect -1404 -4070 -1402 -4066
rect -1400 -4070 -1394 -4066
rect -1392 -4070 -1391 -4066
rect -1379 -4070 -1378 -4066
rect -1376 -4070 -1370 -4066
rect -1368 -4070 -1367 -4066
rect -1230 -4070 -1229 -4066
rect -1227 -4070 -1225 -4066
rect -1221 -4070 -1219 -4066
rect -1217 -4070 -1216 -4066
rect -1204 -4070 -1203 -4066
rect -1201 -4070 -1195 -4066
rect -1193 -4070 -1192 -4066
rect -1180 -4070 -1179 -4066
rect -1177 -4070 -1171 -4066
rect -1169 -4070 -1167 -4066
rect -1163 -4070 -1161 -4066
rect -1159 -4070 -1153 -4066
rect -1151 -4070 -1150 -4066
rect -1138 -4070 -1137 -4066
rect -1135 -4070 -1129 -4066
rect -1127 -4070 -1125 -4066
rect -1121 -4070 -1119 -4066
rect -1117 -4070 -1111 -4066
rect -1109 -4070 -1108 -4066
rect -1096 -4070 -1095 -4066
rect -1093 -4070 -1087 -4066
rect -1085 -4070 -1083 -4066
rect -1079 -4070 -1077 -4066
rect -1075 -4070 -1069 -4066
rect -1067 -4070 -1066 -4066
rect -1054 -4070 -1053 -4066
rect -1051 -4070 -1045 -4066
rect -1043 -4070 -1042 -4066
rect -931 -4070 -930 -4066
rect -928 -4070 -926 -4066
rect -922 -4070 -920 -4066
rect -918 -4070 -917 -4066
rect -905 -4070 -904 -4066
rect -902 -4070 -896 -4066
rect -894 -4070 -893 -4066
rect -881 -4070 -880 -4066
rect -878 -4070 -872 -4066
rect -870 -4070 -868 -4066
rect -864 -4070 -862 -4066
rect -860 -4070 -854 -4066
rect -852 -4070 -851 -4066
rect -839 -4070 -838 -4066
rect -836 -4070 -830 -4066
rect -828 -4070 -826 -4066
rect -822 -4070 -820 -4066
rect -818 -4070 -812 -4066
rect -810 -4070 -809 -4066
rect -797 -4070 -796 -4066
rect -794 -4070 -788 -4066
rect -786 -4070 -784 -4066
rect -780 -4070 -778 -4066
rect -776 -4070 -770 -4066
rect -768 -4070 -767 -4066
rect -755 -4070 -754 -4066
rect -752 -4070 -746 -4066
rect -744 -4070 -743 -4066
rect -573 -4070 -572 -4066
rect -570 -4070 -568 -4066
rect -564 -4070 -562 -4066
rect -560 -4070 -559 -4066
rect -547 -4070 -546 -4066
rect -544 -4070 -538 -4066
rect -536 -4070 -535 -4066
rect -523 -4070 -522 -4066
rect -520 -4070 -514 -4066
rect -512 -4070 -510 -4066
rect -506 -4070 -504 -4066
rect -502 -4070 -496 -4066
rect -494 -4070 -493 -4066
rect -481 -4070 -480 -4066
rect -478 -4070 -472 -4066
rect -470 -4070 -468 -4066
rect -464 -4070 -462 -4066
rect -460 -4070 -454 -4066
rect -452 -4070 -451 -4066
rect -439 -4070 -438 -4066
rect -436 -4070 -430 -4066
rect -428 -4070 -426 -4066
rect -422 -4070 -420 -4066
rect -418 -4070 -412 -4066
rect -410 -4070 -409 -4066
rect -397 -4070 -396 -4066
rect -394 -4070 -388 -4066
rect -386 -4070 -385 -4066
rect -215 -4070 -214 -4066
rect -212 -4070 -210 -4066
rect -206 -4070 -204 -4066
rect -202 -4070 -201 -4066
rect -189 -4070 -188 -4066
rect -186 -4070 -180 -4066
rect -178 -4070 -177 -4066
rect -165 -4070 -164 -4066
rect -162 -4070 -156 -4066
rect -154 -4070 -152 -4066
rect -148 -4070 -146 -4066
rect -144 -4070 -138 -4066
rect -136 -4070 -135 -4066
rect -123 -4070 -122 -4066
rect -120 -4070 -114 -4066
rect -112 -4070 -110 -4066
rect -106 -4070 -104 -4066
rect -102 -4070 -96 -4066
rect -94 -4070 -93 -4066
rect -81 -4070 -80 -4066
rect -78 -4070 -72 -4066
rect -70 -4070 -68 -4066
rect -64 -4070 -62 -4066
rect -60 -4070 -54 -4066
rect -52 -4070 -51 -4066
rect -39 -4070 -38 -4066
rect -36 -4070 -30 -4066
rect -28 -4070 -27 -4066
rect 143 -4070 144 -4066
rect 146 -4070 148 -4066
rect 152 -4070 154 -4066
rect 156 -4070 157 -4066
rect 169 -4070 170 -4066
rect 172 -4070 178 -4066
rect 180 -4070 181 -4066
rect 193 -4070 194 -4066
rect 196 -4070 202 -4066
rect 204 -4070 206 -4066
rect 210 -4070 212 -4066
rect 214 -4070 220 -4066
rect 222 -4070 223 -4066
rect 235 -4070 236 -4066
rect 238 -4070 244 -4066
rect 246 -4070 248 -4066
rect 252 -4070 254 -4066
rect 256 -4070 262 -4066
rect 264 -4070 265 -4066
rect 277 -4070 278 -4066
rect 280 -4070 286 -4066
rect 288 -4070 290 -4066
rect 294 -4070 296 -4066
rect 298 -4070 304 -4066
rect 306 -4070 307 -4066
rect 319 -4070 320 -4066
rect 322 -4070 328 -4066
rect 330 -4070 331 -4066
rect 499 -4070 500 -4066
rect 502 -4070 504 -4066
rect 508 -4070 510 -4066
rect 512 -4070 513 -4066
rect 525 -4070 526 -4066
rect 528 -4070 534 -4066
rect 536 -4070 537 -4066
rect 549 -4070 550 -4066
rect 552 -4070 558 -4066
rect 560 -4070 562 -4066
rect 566 -4070 568 -4066
rect 570 -4070 576 -4066
rect 578 -4070 579 -4066
rect 591 -4070 592 -4066
rect 594 -4070 600 -4066
rect 602 -4070 604 -4066
rect 608 -4070 610 -4066
rect 612 -4070 618 -4066
rect 620 -4070 621 -4066
rect 633 -4070 634 -4066
rect 636 -4070 642 -4066
rect 644 -4070 646 -4066
rect 650 -4070 652 -4066
rect 654 -4070 660 -4066
rect 662 -4070 663 -4066
rect 675 -4070 676 -4066
rect 678 -4070 684 -4066
rect 686 -4070 687 -4066
rect 857 -4070 858 -4066
rect 860 -4070 862 -4066
rect 866 -4070 868 -4066
rect 870 -4070 871 -4066
rect 883 -4070 884 -4066
rect 886 -4070 892 -4066
rect 894 -4070 895 -4066
rect 907 -4070 908 -4066
rect 910 -4070 916 -4066
rect 918 -4070 920 -4066
rect 924 -4070 926 -4066
rect 928 -4070 934 -4066
rect 936 -4070 937 -4066
rect 949 -4070 950 -4066
rect 952 -4070 958 -4066
rect 960 -4070 962 -4066
rect 966 -4070 968 -4066
rect 970 -4070 976 -4066
rect 978 -4070 979 -4066
rect 991 -4070 992 -4066
rect 994 -4070 1000 -4066
rect 1002 -4070 1004 -4066
rect 1008 -4070 1010 -4066
rect 1012 -4070 1018 -4066
rect 1020 -4070 1021 -4066
rect 1033 -4070 1034 -4066
rect 1036 -4070 1042 -4066
rect 1044 -4070 1045 -4066
rect 1215 -4070 1216 -4066
rect 1218 -4070 1220 -4066
rect 1224 -4070 1226 -4066
rect 1228 -4070 1229 -4066
rect 1241 -4070 1242 -4066
rect 1244 -4070 1250 -4066
rect 1252 -4070 1253 -4066
rect 1265 -4070 1266 -4066
rect 1268 -4070 1274 -4066
rect 1276 -4070 1278 -4066
rect 1282 -4070 1284 -4066
rect 1286 -4070 1292 -4066
rect 1294 -4070 1295 -4066
rect 1307 -4070 1308 -4066
rect 1310 -4070 1316 -4066
rect 1318 -4070 1320 -4066
rect 1324 -4070 1326 -4066
rect 1328 -4070 1334 -4066
rect 1336 -4070 1337 -4066
rect 1349 -4070 1350 -4066
rect 1352 -4070 1358 -4066
rect 1360 -4070 1362 -4066
rect 1366 -4070 1368 -4066
rect 1370 -4070 1376 -4066
rect 1378 -4070 1379 -4066
rect 1391 -4070 1392 -4066
rect 1394 -4070 1400 -4066
rect 1402 -4070 1403 -4066
rect -1305 -4185 -1304 -4181
rect -1302 -4185 -1296 -4181
rect -1294 -4185 -1292 -4181
rect -1288 -4185 -1286 -4181
rect -1284 -4185 -1283 -4181
rect -931 -4185 -930 -4181
rect -928 -4185 -922 -4181
rect -920 -4185 -918 -4181
rect -914 -4185 -912 -4181
rect -910 -4185 -909 -4181
rect -573 -4185 -572 -4181
rect -570 -4185 -564 -4181
rect -562 -4185 -560 -4181
rect -556 -4185 -554 -4181
rect -552 -4185 -551 -4181
rect -215 -4185 -214 -4181
rect -212 -4185 -206 -4181
rect -204 -4185 -202 -4181
rect -198 -4185 -196 -4181
rect -194 -4185 -193 -4181
rect 143 -4185 144 -4181
rect 146 -4185 152 -4181
rect 154 -4185 156 -4181
rect 160 -4185 162 -4181
rect 164 -4185 165 -4181
rect 499 -4185 500 -4181
rect 502 -4185 508 -4181
rect 510 -4185 512 -4181
rect 516 -4185 518 -4181
rect 520 -4185 521 -4181
rect 857 -4185 858 -4181
rect 860 -4185 866 -4181
rect 868 -4185 870 -4181
rect 874 -4185 876 -4181
rect 878 -4185 879 -4181
rect 1215 -4185 1216 -4181
rect 1218 -4185 1224 -4181
rect 1226 -4185 1228 -4181
rect 1232 -4185 1234 -4181
rect 1236 -4185 1237 -4181
rect -1230 -4344 -1229 -4340
rect -1227 -4344 -1225 -4340
rect -1221 -4344 -1219 -4340
rect -1217 -4344 -1216 -4340
rect -1204 -4344 -1203 -4340
rect -1201 -4344 -1199 -4340
rect -1195 -4344 -1193 -4340
rect -1191 -4344 -1185 -4340
rect -1183 -4344 -1181 -4340
rect -1177 -4344 -1175 -4340
rect -1173 -4344 -1172 -4340
rect -1160 -4344 -1159 -4340
rect -1157 -4344 -1151 -4340
rect -1149 -4344 -1147 -4340
rect -1143 -4344 -1141 -4340
rect -1139 -4344 -1138 -4340
rect -931 -4344 -930 -4340
rect -928 -4344 -926 -4340
rect -922 -4344 -920 -4340
rect -918 -4344 -917 -4340
rect -905 -4344 -904 -4340
rect -902 -4344 -900 -4340
rect -896 -4344 -894 -4340
rect -892 -4344 -891 -4340
rect -879 -4344 -878 -4340
rect -876 -4344 -875 -4340
rect -871 -4344 -868 -4340
rect -866 -4344 -860 -4340
rect -858 -4344 -857 -4340
rect -853 -4344 -850 -4340
rect -848 -4344 -847 -4340
rect -835 -4344 -834 -4340
rect -832 -4344 -826 -4340
rect -824 -4344 -822 -4340
rect -818 -4344 -816 -4340
rect -814 -4344 -813 -4340
rect -801 -4344 -800 -4340
rect -798 -4344 -796 -4340
rect -792 -4344 -790 -4340
rect -788 -4344 -782 -4340
rect -780 -4344 -778 -4340
rect -774 -4344 -772 -4340
rect -770 -4344 -769 -4340
rect -757 -4344 -756 -4340
rect -754 -4344 -748 -4340
rect -746 -4344 -745 -4340
rect -733 -4344 -732 -4340
rect -730 -4344 -725 -4340
rect -721 -4344 -716 -4340
rect -714 -4344 -713 -4340
rect -709 -4344 -708 -4340
rect -706 -4344 -704 -4340
rect -700 -4344 -698 -4340
rect -696 -4344 -695 -4340
rect -573 -4344 -572 -4340
rect -570 -4344 -568 -4340
rect -564 -4344 -562 -4340
rect -560 -4344 -559 -4340
rect -547 -4344 -546 -4340
rect -544 -4344 -542 -4340
rect -538 -4344 -536 -4340
rect -534 -4344 -533 -4340
rect -521 -4344 -520 -4340
rect -518 -4344 -517 -4340
rect -513 -4344 -510 -4340
rect -508 -4344 -502 -4340
rect -500 -4344 -499 -4340
rect -495 -4344 -492 -4340
rect -490 -4344 -489 -4340
rect -477 -4344 -476 -4340
rect -474 -4344 -468 -4340
rect -466 -4344 -464 -4340
rect -460 -4344 -458 -4340
rect -456 -4344 -455 -4340
rect -443 -4344 -442 -4340
rect -440 -4344 -438 -4340
rect -434 -4344 -432 -4340
rect -430 -4344 -424 -4340
rect -422 -4344 -420 -4340
rect -416 -4344 -414 -4340
rect -412 -4344 -411 -4340
rect -399 -4344 -398 -4340
rect -396 -4344 -390 -4340
rect -388 -4344 -387 -4340
rect -375 -4344 -374 -4340
rect -372 -4344 -367 -4340
rect -363 -4344 -358 -4340
rect -356 -4344 -355 -4340
rect -351 -4344 -350 -4340
rect -348 -4344 -346 -4340
rect -342 -4344 -340 -4340
rect -338 -4344 -337 -4340
rect -215 -4344 -214 -4340
rect -212 -4344 -210 -4340
rect -206 -4344 -204 -4340
rect -202 -4344 -201 -4340
rect -189 -4344 -188 -4340
rect -186 -4344 -184 -4340
rect -180 -4344 -178 -4340
rect -176 -4344 -175 -4340
rect -163 -4344 -162 -4340
rect -160 -4344 -159 -4340
rect -155 -4344 -152 -4340
rect -150 -4344 -144 -4340
rect -142 -4344 -141 -4340
rect -137 -4344 -134 -4340
rect -132 -4344 -131 -4340
rect -119 -4344 -118 -4340
rect -116 -4344 -110 -4340
rect -108 -4344 -106 -4340
rect -102 -4344 -100 -4340
rect -98 -4344 -97 -4340
rect -85 -4344 -84 -4340
rect -82 -4344 -80 -4340
rect -76 -4344 -74 -4340
rect -72 -4344 -66 -4340
rect -64 -4344 -62 -4340
rect -58 -4344 -56 -4340
rect -54 -4344 -53 -4340
rect -41 -4344 -40 -4340
rect -38 -4344 -32 -4340
rect -30 -4344 -29 -4340
rect -17 -4344 -16 -4340
rect -14 -4344 -9 -4340
rect -5 -4344 0 -4340
rect 2 -4344 3 -4340
rect 7 -4344 8 -4340
rect 10 -4344 12 -4340
rect 16 -4344 18 -4340
rect 20 -4344 21 -4340
rect 143 -4344 144 -4340
rect 146 -4344 148 -4340
rect 152 -4344 154 -4340
rect 156 -4344 157 -4340
rect 169 -4344 170 -4340
rect 172 -4344 174 -4340
rect 178 -4344 180 -4340
rect 182 -4344 183 -4340
rect 195 -4344 196 -4340
rect 198 -4344 199 -4340
rect 203 -4344 206 -4340
rect 208 -4344 214 -4340
rect 216 -4344 217 -4340
rect 221 -4344 224 -4340
rect 226 -4344 227 -4340
rect 239 -4344 240 -4340
rect 242 -4344 248 -4340
rect 250 -4344 252 -4340
rect 256 -4344 258 -4340
rect 260 -4344 261 -4340
rect 273 -4344 274 -4340
rect 276 -4344 278 -4340
rect 282 -4344 284 -4340
rect 286 -4344 292 -4340
rect 294 -4344 296 -4340
rect 300 -4344 302 -4340
rect 304 -4344 305 -4340
rect 317 -4344 318 -4340
rect 320 -4344 326 -4340
rect 328 -4344 329 -4340
rect 341 -4344 342 -4340
rect 344 -4344 349 -4340
rect 353 -4344 358 -4340
rect 360 -4344 361 -4340
rect 365 -4344 366 -4340
rect 368 -4344 370 -4340
rect 374 -4344 376 -4340
rect 378 -4344 379 -4340
rect 499 -4344 500 -4340
rect 502 -4344 504 -4340
rect 508 -4344 510 -4340
rect 512 -4344 513 -4340
rect 525 -4344 526 -4340
rect 528 -4344 530 -4340
rect 534 -4344 536 -4340
rect 538 -4344 539 -4340
rect 551 -4344 552 -4340
rect 554 -4344 555 -4340
rect 559 -4344 562 -4340
rect 564 -4344 570 -4340
rect 572 -4344 573 -4340
rect 577 -4344 580 -4340
rect 582 -4344 583 -4340
rect 595 -4344 596 -4340
rect 598 -4344 604 -4340
rect 606 -4344 608 -4340
rect 612 -4344 614 -4340
rect 616 -4344 617 -4340
rect 629 -4344 630 -4340
rect 632 -4344 634 -4340
rect 638 -4344 640 -4340
rect 642 -4344 648 -4340
rect 650 -4344 652 -4340
rect 656 -4344 658 -4340
rect 660 -4344 661 -4340
rect 673 -4344 674 -4340
rect 676 -4344 682 -4340
rect 684 -4344 685 -4340
rect 697 -4344 698 -4340
rect 700 -4344 705 -4340
rect 709 -4344 714 -4340
rect 716 -4344 717 -4340
rect 721 -4344 722 -4340
rect 724 -4344 726 -4340
rect 730 -4344 732 -4340
rect 734 -4344 735 -4340
rect 857 -4344 858 -4340
rect 860 -4344 862 -4340
rect 866 -4344 868 -4340
rect 870 -4344 871 -4340
rect 883 -4344 884 -4340
rect 886 -4344 888 -4340
rect 892 -4344 894 -4340
rect 896 -4344 897 -4340
rect 909 -4344 910 -4340
rect 912 -4344 913 -4340
rect 917 -4344 920 -4340
rect 922 -4344 928 -4340
rect 930 -4344 931 -4340
rect 935 -4344 938 -4340
rect 940 -4344 941 -4340
rect 953 -4344 954 -4340
rect 956 -4344 962 -4340
rect 964 -4344 966 -4340
rect 970 -4344 972 -4340
rect 974 -4344 975 -4340
rect 987 -4344 988 -4340
rect 990 -4344 992 -4340
rect 996 -4344 998 -4340
rect 1000 -4344 1006 -4340
rect 1008 -4344 1010 -4340
rect 1014 -4344 1016 -4340
rect 1018 -4344 1019 -4340
rect 1031 -4344 1032 -4340
rect 1034 -4344 1040 -4340
rect 1042 -4344 1043 -4340
rect 1055 -4344 1056 -4340
rect 1058 -4344 1063 -4340
rect 1067 -4344 1072 -4340
rect 1074 -4344 1075 -4340
rect 1079 -4344 1080 -4340
rect 1082 -4344 1084 -4340
rect 1088 -4344 1090 -4340
rect 1092 -4344 1093 -4340
rect 1215 -4344 1216 -4340
rect 1218 -4344 1220 -4340
rect 1224 -4344 1226 -4340
rect 1228 -4344 1229 -4340
rect 1241 -4344 1242 -4340
rect 1244 -4344 1246 -4340
rect 1250 -4344 1252 -4340
rect 1254 -4344 1255 -4340
rect 1267 -4344 1268 -4340
rect 1270 -4344 1271 -4340
rect 1275 -4344 1278 -4340
rect 1280 -4344 1286 -4340
rect 1288 -4344 1289 -4340
rect 1293 -4344 1296 -4340
rect 1298 -4344 1299 -4340
rect 1311 -4344 1312 -4340
rect 1314 -4344 1320 -4340
rect 1322 -4344 1324 -4340
rect 1328 -4344 1330 -4340
rect 1332 -4344 1333 -4340
rect 1345 -4344 1346 -4340
rect 1348 -4344 1350 -4340
rect 1354 -4344 1356 -4340
rect 1358 -4344 1364 -4340
rect 1366 -4344 1368 -4340
rect 1372 -4344 1374 -4340
rect 1376 -4344 1377 -4340
rect 1389 -4344 1390 -4340
rect 1392 -4344 1398 -4340
rect 1400 -4344 1401 -4340
rect 1413 -4344 1414 -4340
rect 1416 -4344 1421 -4340
rect 1425 -4344 1430 -4340
rect 1432 -4344 1433 -4340
rect 1437 -4344 1438 -4340
rect 1440 -4344 1442 -4340
rect 1446 -4344 1448 -4340
rect 1450 -4344 1451 -4340
rect -1810 -4467 -1809 -4463
rect -1807 -4467 -1805 -4463
rect -1801 -4467 -1799 -4463
rect -1797 -4467 -1796 -4463
rect -1784 -4467 -1783 -4463
rect -1781 -4467 -1775 -4463
rect -1773 -4467 -1772 -4463
rect -1760 -4467 -1759 -4463
rect -1757 -4467 -1751 -4463
rect -1749 -4467 -1747 -4463
rect -1743 -4467 -1741 -4463
rect -1739 -4467 -1733 -4463
rect -1731 -4467 -1730 -4463
rect -1718 -4467 -1717 -4463
rect -1715 -4467 -1709 -4463
rect -1707 -4467 -1705 -4463
rect -1701 -4467 -1699 -4463
rect -1697 -4467 -1691 -4463
rect -1689 -4467 -1688 -4463
rect -1676 -4467 -1675 -4463
rect -1673 -4467 -1667 -4463
rect -1665 -4467 -1663 -4463
rect -1659 -4467 -1657 -4463
rect -1655 -4467 -1649 -4463
rect -1647 -4467 -1646 -4463
rect -1634 -4467 -1633 -4463
rect -1631 -4467 -1625 -4463
rect -1623 -4467 -1622 -4463
rect -1547 -4467 -1546 -4463
rect -1544 -4467 -1542 -4463
rect -1538 -4467 -1536 -4463
rect -1534 -4467 -1533 -4463
rect -1521 -4467 -1520 -4463
rect -1518 -4467 -1512 -4463
rect -1510 -4467 -1509 -4463
rect -1497 -4467 -1496 -4463
rect -1494 -4467 -1488 -4463
rect -1486 -4467 -1484 -4463
rect -1480 -4467 -1478 -4463
rect -1476 -4467 -1470 -4463
rect -1468 -4467 -1467 -4463
rect -1455 -4467 -1454 -4463
rect -1452 -4467 -1446 -4463
rect -1444 -4467 -1442 -4463
rect -1438 -4467 -1436 -4463
rect -1434 -4467 -1428 -4463
rect -1426 -4467 -1425 -4463
rect -1413 -4467 -1412 -4463
rect -1410 -4467 -1404 -4463
rect -1402 -4467 -1400 -4463
rect -1396 -4467 -1394 -4463
rect -1392 -4467 -1386 -4463
rect -1384 -4467 -1383 -4463
rect -1371 -4467 -1370 -4463
rect -1368 -4467 -1362 -4463
rect -1360 -4467 -1359 -4463
rect -1230 -4467 -1229 -4463
rect -1227 -4467 -1225 -4463
rect -1221 -4467 -1219 -4463
rect -1217 -4467 -1216 -4463
rect -1204 -4467 -1203 -4463
rect -1201 -4467 -1195 -4463
rect -1193 -4467 -1192 -4463
rect -1180 -4467 -1179 -4463
rect -1177 -4467 -1171 -4463
rect -1169 -4467 -1167 -4463
rect -1163 -4467 -1161 -4463
rect -1159 -4467 -1153 -4463
rect -1151 -4467 -1150 -4463
rect -1138 -4467 -1137 -4463
rect -1135 -4467 -1129 -4463
rect -1127 -4467 -1125 -4463
rect -1121 -4467 -1119 -4463
rect -1117 -4467 -1111 -4463
rect -1109 -4467 -1108 -4463
rect -1096 -4467 -1095 -4463
rect -1093 -4467 -1087 -4463
rect -1085 -4467 -1083 -4463
rect -1079 -4467 -1077 -4463
rect -1075 -4467 -1069 -4463
rect -1067 -4467 -1066 -4463
rect -1054 -4467 -1053 -4463
rect -1051 -4467 -1045 -4463
rect -1043 -4467 -1042 -4463
rect -931 -4467 -930 -4463
rect -928 -4467 -926 -4463
rect -922 -4467 -920 -4463
rect -918 -4467 -917 -4463
rect -905 -4467 -904 -4463
rect -902 -4467 -896 -4463
rect -894 -4467 -893 -4463
rect -881 -4467 -880 -4463
rect -878 -4467 -872 -4463
rect -870 -4467 -868 -4463
rect -864 -4467 -862 -4463
rect -860 -4467 -854 -4463
rect -852 -4467 -851 -4463
rect -839 -4467 -838 -4463
rect -836 -4467 -830 -4463
rect -828 -4467 -826 -4463
rect -822 -4467 -820 -4463
rect -818 -4467 -812 -4463
rect -810 -4467 -809 -4463
rect -797 -4467 -796 -4463
rect -794 -4467 -788 -4463
rect -786 -4467 -784 -4463
rect -780 -4467 -778 -4463
rect -776 -4467 -770 -4463
rect -768 -4467 -767 -4463
rect -755 -4467 -754 -4463
rect -752 -4467 -746 -4463
rect -744 -4467 -743 -4463
rect -573 -4467 -572 -4463
rect -570 -4467 -568 -4463
rect -564 -4467 -562 -4463
rect -560 -4467 -559 -4463
rect -547 -4467 -546 -4463
rect -544 -4467 -538 -4463
rect -536 -4467 -535 -4463
rect -523 -4467 -522 -4463
rect -520 -4467 -514 -4463
rect -512 -4467 -510 -4463
rect -506 -4467 -504 -4463
rect -502 -4467 -496 -4463
rect -494 -4467 -493 -4463
rect -481 -4467 -480 -4463
rect -478 -4467 -472 -4463
rect -470 -4467 -468 -4463
rect -464 -4467 -462 -4463
rect -460 -4467 -454 -4463
rect -452 -4467 -451 -4463
rect -439 -4467 -438 -4463
rect -436 -4467 -430 -4463
rect -428 -4467 -426 -4463
rect -422 -4467 -420 -4463
rect -418 -4467 -412 -4463
rect -410 -4467 -409 -4463
rect -397 -4467 -396 -4463
rect -394 -4467 -388 -4463
rect -386 -4467 -385 -4463
rect -1810 -4638 -1809 -4634
rect -1807 -4638 -1805 -4634
rect -1801 -4638 -1799 -4634
rect -1797 -4638 -1796 -4634
rect -1784 -4638 -1783 -4634
rect -1781 -4638 -1775 -4634
rect -1773 -4638 -1772 -4634
rect -1760 -4638 -1759 -4634
rect -1757 -4638 -1751 -4634
rect -1749 -4638 -1747 -4634
rect -1743 -4638 -1741 -4634
rect -1739 -4638 -1733 -4634
rect -1731 -4638 -1730 -4634
rect -1718 -4638 -1717 -4634
rect -1715 -4638 -1709 -4634
rect -1707 -4638 -1705 -4634
rect -1701 -4638 -1699 -4634
rect -1697 -4638 -1691 -4634
rect -1689 -4638 -1688 -4634
rect -1676 -4638 -1675 -4634
rect -1673 -4638 -1667 -4634
rect -1665 -4638 -1663 -4634
rect -1659 -4638 -1657 -4634
rect -1655 -4638 -1649 -4634
rect -1647 -4638 -1646 -4634
rect -1634 -4638 -1633 -4634
rect -1631 -4638 -1625 -4634
rect -1623 -4638 -1622 -4634
rect -1547 -4638 -1546 -4634
rect -1544 -4638 -1542 -4634
rect -1538 -4638 -1536 -4634
rect -1534 -4638 -1533 -4634
rect -1521 -4638 -1520 -4634
rect -1518 -4638 -1512 -4634
rect -1510 -4638 -1509 -4634
rect -1497 -4638 -1496 -4634
rect -1494 -4638 -1488 -4634
rect -1486 -4638 -1484 -4634
rect -1480 -4638 -1478 -4634
rect -1476 -4638 -1470 -4634
rect -1468 -4638 -1467 -4634
rect -1455 -4638 -1454 -4634
rect -1452 -4638 -1446 -4634
rect -1444 -4638 -1442 -4634
rect -1438 -4638 -1436 -4634
rect -1434 -4638 -1428 -4634
rect -1426 -4638 -1425 -4634
rect -1413 -4638 -1412 -4634
rect -1410 -4638 -1404 -4634
rect -1402 -4638 -1400 -4634
rect -1396 -4638 -1394 -4634
rect -1392 -4638 -1386 -4634
rect -1384 -4638 -1383 -4634
rect -1371 -4638 -1370 -4634
rect -1368 -4638 -1362 -4634
rect -1360 -4638 -1359 -4634
rect -1230 -4638 -1229 -4634
rect -1227 -4638 -1225 -4634
rect -1221 -4638 -1219 -4634
rect -1217 -4638 -1216 -4634
rect -1204 -4638 -1203 -4634
rect -1201 -4638 -1195 -4634
rect -1193 -4638 -1192 -4634
rect -1180 -4638 -1179 -4634
rect -1177 -4638 -1171 -4634
rect -1169 -4638 -1167 -4634
rect -1163 -4638 -1161 -4634
rect -1159 -4638 -1153 -4634
rect -1151 -4638 -1150 -4634
rect -1138 -4638 -1137 -4634
rect -1135 -4638 -1129 -4634
rect -1127 -4638 -1125 -4634
rect -1121 -4638 -1119 -4634
rect -1117 -4638 -1111 -4634
rect -1109 -4638 -1108 -4634
rect -1096 -4638 -1095 -4634
rect -1093 -4638 -1087 -4634
rect -1085 -4638 -1083 -4634
rect -1079 -4638 -1077 -4634
rect -1075 -4638 -1069 -4634
rect -1067 -4638 -1066 -4634
rect -1054 -4638 -1053 -4634
rect -1051 -4638 -1045 -4634
rect -1043 -4638 -1042 -4634
rect -931 -4638 -930 -4634
rect -928 -4638 -926 -4634
rect -922 -4638 -920 -4634
rect -918 -4638 -917 -4634
rect -905 -4638 -904 -4634
rect -902 -4638 -896 -4634
rect -894 -4638 -893 -4634
rect -881 -4638 -880 -4634
rect -878 -4638 -872 -4634
rect -870 -4638 -868 -4634
rect -864 -4638 -862 -4634
rect -860 -4638 -854 -4634
rect -852 -4638 -851 -4634
rect -839 -4638 -838 -4634
rect -836 -4638 -830 -4634
rect -828 -4638 -826 -4634
rect -822 -4638 -820 -4634
rect -818 -4638 -812 -4634
rect -810 -4638 -809 -4634
rect -797 -4638 -796 -4634
rect -794 -4638 -788 -4634
rect -786 -4638 -784 -4634
rect -780 -4638 -778 -4634
rect -776 -4638 -770 -4634
rect -768 -4638 -767 -4634
rect -755 -4638 -754 -4634
rect -752 -4638 -746 -4634
rect -744 -4638 -743 -4634
rect -573 -4638 -572 -4634
rect -570 -4638 -568 -4634
rect -564 -4638 -562 -4634
rect -560 -4638 -559 -4634
rect -547 -4638 -546 -4634
rect -544 -4638 -538 -4634
rect -536 -4638 -535 -4634
rect -523 -4638 -522 -4634
rect -520 -4638 -514 -4634
rect -512 -4638 -510 -4634
rect -506 -4638 -504 -4634
rect -502 -4638 -496 -4634
rect -494 -4638 -493 -4634
rect -481 -4638 -480 -4634
rect -478 -4638 -472 -4634
rect -470 -4638 -468 -4634
rect -464 -4638 -462 -4634
rect -460 -4638 -454 -4634
rect -452 -4638 -451 -4634
rect -439 -4638 -438 -4634
rect -436 -4638 -430 -4634
rect -428 -4638 -426 -4634
rect -422 -4638 -420 -4634
rect -418 -4638 -412 -4634
rect -410 -4638 -409 -4634
rect -397 -4638 -396 -4634
rect -394 -4638 -388 -4634
rect -386 -4638 -385 -4634
rect -215 -4638 -214 -4634
rect -212 -4638 -210 -4634
rect -206 -4638 -204 -4634
rect -202 -4638 -201 -4634
rect -189 -4638 -188 -4634
rect -186 -4638 -180 -4634
rect -178 -4638 -177 -4634
rect -165 -4638 -164 -4634
rect -162 -4638 -156 -4634
rect -154 -4638 -152 -4634
rect -148 -4638 -146 -4634
rect -144 -4638 -138 -4634
rect -136 -4638 -135 -4634
rect -123 -4638 -122 -4634
rect -120 -4638 -114 -4634
rect -112 -4638 -110 -4634
rect -106 -4638 -104 -4634
rect -102 -4638 -96 -4634
rect -94 -4638 -93 -4634
rect -81 -4638 -80 -4634
rect -78 -4638 -72 -4634
rect -70 -4638 -68 -4634
rect -64 -4638 -62 -4634
rect -60 -4638 -54 -4634
rect -52 -4638 -51 -4634
rect -39 -4638 -38 -4634
rect -36 -4638 -30 -4634
rect -28 -4638 -27 -4634
rect 143 -4638 144 -4634
rect 146 -4638 148 -4634
rect 152 -4638 154 -4634
rect 156 -4638 157 -4634
rect 169 -4638 170 -4634
rect 172 -4638 178 -4634
rect 180 -4638 181 -4634
rect 193 -4638 194 -4634
rect 196 -4638 202 -4634
rect 204 -4638 206 -4634
rect 210 -4638 212 -4634
rect 214 -4638 220 -4634
rect 222 -4638 223 -4634
rect 235 -4638 236 -4634
rect 238 -4638 244 -4634
rect 246 -4638 248 -4634
rect 252 -4638 254 -4634
rect 256 -4638 262 -4634
rect 264 -4638 265 -4634
rect 277 -4638 278 -4634
rect 280 -4638 286 -4634
rect 288 -4638 290 -4634
rect 294 -4638 296 -4634
rect 298 -4638 304 -4634
rect 306 -4638 307 -4634
rect 319 -4638 320 -4634
rect 322 -4638 328 -4634
rect 330 -4638 331 -4634
rect 499 -4638 500 -4634
rect 502 -4638 504 -4634
rect 508 -4638 510 -4634
rect 512 -4638 513 -4634
rect 525 -4638 526 -4634
rect 528 -4638 534 -4634
rect 536 -4638 537 -4634
rect 549 -4638 550 -4634
rect 552 -4638 558 -4634
rect 560 -4638 562 -4634
rect 566 -4638 568 -4634
rect 570 -4638 576 -4634
rect 578 -4638 579 -4634
rect 591 -4638 592 -4634
rect 594 -4638 600 -4634
rect 602 -4638 604 -4634
rect 608 -4638 610 -4634
rect 612 -4638 618 -4634
rect 620 -4638 621 -4634
rect 633 -4638 634 -4634
rect 636 -4638 642 -4634
rect 644 -4638 646 -4634
rect 650 -4638 652 -4634
rect 654 -4638 660 -4634
rect 662 -4638 663 -4634
rect 675 -4638 676 -4634
rect 678 -4638 684 -4634
rect 686 -4638 687 -4634
rect 857 -4638 858 -4634
rect 860 -4638 862 -4634
rect 866 -4638 868 -4634
rect 870 -4638 871 -4634
rect 883 -4638 884 -4634
rect 886 -4638 892 -4634
rect 894 -4638 895 -4634
rect 907 -4638 908 -4634
rect 910 -4638 916 -4634
rect 918 -4638 920 -4634
rect 924 -4638 926 -4634
rect 928 -4638 934 -4634
rect 936 -4638 937 -4634
rect 949 -4638 950 -4634
rect 952 -4638 958 -4634
rect 960 -4638 962 -4634
rect 966 -4638 968 -4634
rect 970 -4638 976 -4634
rect 978 -4638 979 -4634
rect 991 -4638 992 -4634
rect 994 -4638 1000 -4634
rect 1002 -4638 1004 -4634
rect 1008 -4638 1010 -4634
rect 1012 -4638 1018 -4634
rect 1020 -4638 1021 -4634
rect 1033 -4638 1034 -4634
rect 1036 -4638 1042 -4634
rect 1044 -4638 1045 -4634
rect 1215 -4638 1216 -4634
rect 1218 -4638 1220 -4634
rect 1224 -4638 1226 -4634
rect 1228 -4638 1229 -4634
rect 1241 -4638 1242 -4634
rect 1244 -4638 1250 -4634
rect 1252 -4638 1253 -4634
rect 1265 -4638 1266 -4634
rect 1268 -4638 1274 -4634
rect 1276 -4638 1278 -4634
rect 1282 -4638 1284 -4634
rect 1286 -4638 1292 -4634
rect 1294 -4638 1295 -4634
rect 1307 -4638 1308 -4634
rect 1310 -4638 1316 -4634
rect 1318 -4638 1320 -4634
rect 1324 -4638 1326 -4634
rect 1328 -4638 1334 -4634
rect 1336 -4638 1337 -4634
rect 1349 -4638 1350 -4634
rect 1352 -4638 1358 -4634
rect 1360 -4638 1362 -4634
rect 1366 -4638 1368 -4634
rect 1370 -4638 1376 -4634
rect 1378 -4638 1379 -4634
rect 1391 -4638 1392 -4634
rect 1394 -4638 1400 -4634
rect 1402 -4638 1403 -4634
rect -1547 -4809 -1546 -4805
rect -1544 -4809 -1542 -4805
rect -1538 -4809 -1536 -4805
rect -1534 -4809 -1533 -4805
rect -1521 -4809 -1520 -4805
rect -1518 -4809 -1512 -4805
rect -1510 -4809 -1509 -4805
rect -1497 -4809 -1496 -4805
rect -1494 -4809 -1488 -4805
rect -1486 -4809 -1484 -4805
rect -1480 -4809 -1478 -4805
rect -1476 -4809 -1470 -4805
rect -1468 -4809 -1467 -4805
rect -1455 -4809 -1454 -4805
rect -1452 -4809 -1446 -4805
rect -1444 -4809 -1442 -4805
rect -1438 -4809 -1436 -4805
rect -1434 -4809 -1428 -4805
rect -1426 -4809 -1425 -4805
rect -1413 -4809 -1412 -4805
rect -1410 -4809 -1404 -4805
rect -1402 -4809 -1400 -4805
rect -1396 -4809 -1394 -4805
rect -1392 -4809 -1386 -4805
rect -1384 -4809 -1383 -4805
rect -1371 -4809 -1370 -4805
rect -1368 -4809 -1362 -4805
rect -1360 -4809 -1359 -4805
rect -1230 -4809 -1229 -4805
rect -1227 -4809 -1225 -4805
rect -1221 -4809 -1219 -4805
rect -1217 -4809 -1216 -4805
rect -1204 -4809 -1203 -4805
rect -1201 -4809 -1195 -4805
rect -1193 -4809 -1192 -4805
rect -1180 -4809 -1179 -4805
rect -1177 -4809 -1171 -4805
rect -1169 -4809 -1167 -4805
rect -1163 -4809 -1161 -4805
rect -1159 -4809 -1153 -4805
rect -1151 -4809 -1150 -4805
rect -1138 -4809 -1137 -4805
rect -1135 -4809 -1129 -4805
rect -1127 -4809 -1125 -4805
rect -1121 -4809 -1119 -4805
rect -1117 -4809 -1111 -4805
rect -1109 -4809 -1108 -4805
rect -1096 -4809 -1095 -4805
rect -1093 -4809 -1087 -4805
rect -1085 -4809 -1083 -4805
rect -1079 -4809 -1077 -4805
rect -1075 -4809 -1069 -4805
rect -1067 -4809 -1066 -4805
rect -1054 -4809 -1053 -4805
rect -1051 -4809 -1045 -4805
rect -1043 -4809 -1042 -4805
rect -931 -4809 -930 -4805
rect -928 -4809 -926 -4805
rect -922 -4809 -920 -4805
rect -918 -4809 -917 -4805
rect -905 -4809 -904 -4805
rect -902 -4809 -896 -4805
rect -894 -4809 -893 -4805
rect -881 -4809 -880 -4805
rect -878 -4809 -872 -4805
rect -870 -4809 -868 -4805
rect -864 -4809 -862 -4805
rect -860 -4809 -854 -4805
rect -852 -4809 -851 -4805
rect -839 -4809 -838 -4805
rect -836 -4809 -830 -4805
rect -828 -4809 -826 -4805
rect -822 -4809 -820 -4805
rect -818 -4809 -812 -4805
rect -810 -4809 -809 -4805
rect -797 -4809 -796 -4805
rect -794 -4809 -788 -4805
rect -786 -4809 -784 -4805
rect -780 -4809 -778 -4805
rect -776 -4809 -770 -4805
rect -768 -4809 -767 -4805
rect -755 -4809 -754 -4805
rect -752 -4809 -746 -4805
rect -744 -4809 -743 -4805
rect -573 -4809 -572 -4805
rect -570 -4809 -568 -4805
rect -564 -4809 -562 -4805
rect -560 -4809 -559 -4805
rect -547 -4809 -546 -4805
rect -544 -4809 -538 -4805
rect -536 -4809 -535 -4805
rect -523 -4809 -522 -4805
rect -520 -4809 -514 -4805
rect -512 -4809 -510 -4805
rect -506 -4809 -504 -4805
rect -502 -4809 -496 -4805
rect -494 -4809 -493 -4805
rect -481 -4809 -480 -4805
rect -478 -4809 -472 -4805
rect -470 -4809 -468 -4805
rect -464 -4809 -462 -4805
rect -460 -4809 -454 -4805
rect -452 -4809 -451 -4805
rect -439 -4809 -438 -4805
rect -436 -4809 -430 -4805
rect -428 -4809 -426 -4805
rect -422 -4809 -420 -4805
rect -418 -4809 -412 -4805
rect -410 -4809 -409 -4805
rect -397 -4809 -396 -4805
rect -394 -4809 -388 -4805
rect -386 -4809 -385 -4805
rect -215 -4809 -214 -4805
rect -212 -4809 -210 -4805
rect -206 -4809 -204 -4805
rect -202 -4809 -201 -4805
rect -189 -4809 -188 -4805
rect -186 -4809 -180 -4805
rect -178 -4809 -177 -4805
rect -165 -4809 -164 -4805
rect -162 -4809 -156 -4805
rect -154 -4809 -152 -4805
rect -148 -4809 -146 -4805
rect -144 -4809 -138 -4805
rect -136 -4809 -135 -4805
rect -123 -4809 -122 -4805
rect -120 -4809 -114 -4805
rect -112 -4809 -110 -4805
rect -106 -4809 -104 -4805
rect -102 -4809 -96 -4805
rect -94 -4809 -93 -4805
rect -81 -4809 -80 -4805
rect -78 -4809 -72 -4805
rect -70 -4809 -68 -4805
rect -64 -4809 -62 -4805
rect -60 -4809 -54 -4805
rect -52 -4809 -51 -4805
rect -39 -4809 -38 -4805
rect -36 -4809 -30 -4805
rect -28 -4809 -27 -4805
rect 143 -4809 144 -4805
rect 146 -4809 148 -4805
rect 152 -4809 154 -4805
rect 156 -4809 157 -4805
rect 169 -4809 170 -4805
rect 172 -4809 178 -4805
rect 180 -4809 181 -4805
rect 193 -4809 194 -4805
rect 196 -4809 202 -4805
rect 204 -4809 206 -4805
rect 210 -4809 212 -4805
rect 214 -4809 220 -4805
rect 222 -4809 223 -4805
rect 235 -4809 236 -4805
rect 238 -4809 244 -4805
rect 246 -4809 248 -4805
rect 252 -4809 254 -4805
rect 256 -4809 262 -4805
rect 264 -4809 265 -4805
rect 277 -4809 278 -4805
rect 280 -4809 286 -4805
rect 288 -4809 290 -4805
rect 294 -4809 296 -4805
rect 298 -4809 304 -4805
rect 306 -4809 307 -4805
rect 319 -4809 320 -4805
rect 322 -4809 328 -4805
rect 330 -4809 331 -4805
rect 499 -4809 500 -4805
rect 502 -4809 504 -4805
rect 508 -4809 510 -4805
rect 512 -4809 513 -4805
rect 525 -4809 526 -4805
rect 528 -4809 534 -4805
rect 536 -4809 537 -4805
rect 549 -4809 550 -4805
rect 552 -4809 558 -4805
rect 560 -4809 562 -4805
rect 566 -4809 568 -4805
rect 570 -4809 576 -4805
rect 578 -4809 579 -4805
rect 591 -4809 592 -4805
rect 594 -4809 600 -4805
rect 602 -4809 604 -4805
rect 608 -4809 610 -4805
rect 612 -4809 618 -4805
rect 620 -4809 621 -4805
rect 633 -4809 634 -4805
rect 636 -4809 642 -4805
rect 644 -4809 646 -4805
rect 650 -4809 652 -4805
rect 654 -4809 660 -4805
rect 662 -4809 663 -4805
rect 675 -4809 676 -4805
rect 678 -4809 684 -4805
rect 686 -4809 687 -4805
rect 857 -4809 858 -4805
rect 860 -4809 862 -4805
rect 866 -4809 868 -4805
rect 870 -4809 871 -4805
rect 883 -4809 884 -4805
rect 886 -4809 892 -4805
rect 894 -4809 895 -4805
rect 907 -4809 908 -4805
rect 910 -4809 916 -4805
rect 918 -4809 920 -4805
rect 924 -4809 926 -4805
rect 928 -4809 934 -4805
rect 936 -4809 937 -4805
rect 949 -4809 950 -4805
rect 952 -4809 958 -4805
rect 960 -4809 962 -4805
rect 966 -4809 968 -4805
rect 970 -4809 976 -4805
rect 978 -4809 979 -4805
rect 991 -4809 992 -4805
rect 994 -4809 1000 -4805
rect 1002 -4809 1004 -4805
rect 1008 -4809 1010 -4805
rect 1012 -4809 1018 -4805
rect 1020 -4809 1021 -4805
rect 1033 -4809 1034 -4805
rect 1036 -4809 1042 -4805
rect 1044 -4809 1045 -4805
rect 1215 -4809 1216 -4805
rect 1218 -4809 1220 -4805
rect 1224 -4809 1226 -4805
rect 1228 -4809 1229 -4805
rect 1241 -4809 1242 -4805
rect 1244 -4809 1250 -4805
rect 1252 -4809 1253 -4805
rect 1265 -4809 1266 -4805
rect 1268 -4809 1274 -4805
rect 1276 -4809 1278 -4805
rect 1282 -4809 1284 -4805
rect 1286 -4809 1292 -4805
rect 1294 -4809 1295 -4805
rect 1307 -4809 1308 -4805
rect 1310 -4809 1316 -4805
rect 1318 -4809 1320 -4805
rect 1324 -4809 1326 -4805
rect 1328 -4809 1334 -4805
rect 1336 -4809 1337 -4805
rect 1349 -4809 1350 -4805
rect 1352 -4809 1358 -4805
rect 1360 -4809 1362 -4805
rect 1366 -4809 1368 -4805
rect 1370 -4809 1376 -4805
rect 1378 -4809 1379 -4805
rect 1391 -4809 1392 -4805
rect 1394 -4809 1400 -4805
rect 1402 -4809 1403 -4805
rect -1305 -4924 -1304 -4920
rect -1302 -4924 -1296 -4920
rect -1294 -4924 -1292 -4920
rect -1288 -4924 -1286 -4920
rect -1284 -4924 -1283 -4920
rect -931 -4924 -930 -4920
rect -928 -4924 -922 -4920
rect -920 -4924 -918 -4920
rect -914 -4924 -912 -4920
rect -910 -4924 -909 -4920
rect -573 -4924 -572 -4920
rect -570 -4924 -564 -4920
rect -562 -4924 -560 -4920
rect -556 -4924 -554 -4920
rect -552 -4924 -551 -4920
rect -215 -4924 -214 -4920
rect -212 -4924 -206 -4920
rect -204 -4924 -202 -4920
rect -198 -4924 -196 -4920
rect -194 -4924 -193 -4920
rect 143 -4924 144 -4920
rect 146 -4924 152 -4920
rect 154 -4924 156 -4920
rect 160 -4924 162 -4920
rect 164 -4924 165 -4920
rect 499 -4924 500 -4920
rect 502 -4924 508 -4920
rect 510 -4924 512 -4920
rect 516 -4924 518 -4920
rect 520 -4924 521 -4920
rect 857 -4924 858 -4920
rect 860 -4924 866 -4920
rect 868 -4924 870 -4920
rect 874 -4924 876 -4920
rect 878 -4924 879 -4920
rect 1215 -4924 1216 -4920
rect 1218 -4924 1224 -4920
rect 1226 -4924 1228 -4920
rect 1232 -4924 1234 -4920
rect 1236 -4924 1237 -4920
rect -1230 -5083 -1229 -5079
rect -1227 -5083 -1225 -5079
rect -1221 -5083 -1219 -5079
rect -1217 -5083 -1216 -5079
rect -1204 -5083 -1203 -5079
rect -1201 -5083 -1199 -5079
rect -1195 -5083 -1193 -5079
rect -1191 -5083 -1185 -5079
rect -1183 -5083 -1181 -5079
rect -1177 -5083 -1175 -5079
rect -1173 -5083 -1172 -5079
rect -1160 -5083 -1159 -5079
rect -1157 -5083 -1151 -5079
rect -1149 -5083 -1147 -5079
rect -1143 -5083 -1141 -5079
rect -1139 -5083 -1138 -5079
rect -931 -5083 -930 -5079
rect -928 -5083 -926 -5079
rect -922 -5083 -920 -5079
rect -918 -5083 -917 -5079
rect -905 -5083 -904 -5079
rect -902 -5083 -900 -5079
rect -896 -5083 -894 -5079
rect -892 -5083 -891 -5079
rect -879 -5083 -878 -5079
rect -876 -5083 -875 -5079
rect -871 -5083 -868 -5079
rect -866 -5083 -860 -5079
rect -858 -5083 -857 -5079
rect -853 -5083 -850 -5079
rect -848 -5083 -847 -5079
rect -835 -5083 -834 -5079
rect -832 -5083 -826 -5079
rect -824 -5083 -822 -5079
rect -818 -5083 -816 -5079
rect -814 -5083 -813 -5079
rect -801 -5083 -800 -5079
rect -798 -5083 -796 -5079
rect -792 -5083 -790 -5079
rect -788 -5083 -782 -5079
rect -780 -5083 -778 -5079
rect -774 -5083 -772 -5079
rect -770 -5083 -769 -5079
rect -757 -5083 -756 -5079
rect -754 -5083 -748 -5079
rect -746 -5083 -745 -5079
rect -733 -5083 -732 -5079
rect -730 -5083 -725 -5079
rect -721 -5083 -716 -5079
rect -714 -5083 -713 -5079
rect -709 -5083 -708 -5079
rect -706 -5083 -704 -5079
rect -700 -5083 -698 -5079
rect -696 -5083 -695 -5079
rect -573 -5083 -572 -5079
rect -570 -5083 -568 -5079
rect -564 -5083 -562 -5079
rect -560 -5083 -559 -5079
rect -547 -5083 -546 -5079
rect -544 -5083 -542 -5079
rect -538 -5083 -536 -5079
rect -534 -5083 -533 -5079
rect -521 -5083 -520 -5079
rect -518 -5083 -517 -5079
rect -513 -5083 -510 -5079
rect -508 -5083 -502 -5079
rect -500 -5083 -499 -5079
rect -495 -5083 -492 -5079
rect -490 -5083 -489 -5079
rect -477 -5083 -476 -5079
rect -474 -5083 -468 -5079
rect -466 -5083 -464 -5079
rect -460 -5083 -458 -5079
rect -456 -5083 -455 -5079
rect -443 -5083 -442 -5079
rect -440 -5083 -438 -5079
rect -434 -5083 -432 -5079
rect -430 -5083 -424 -5079
rect -422 -5083 -420 -5079
rect -416 -5083 -414 -5079
rect -412 -5083 -411 -5079
rect -399 -5083 -398 -5079
rect -396 -5083 -390 -5079
rect -388 -5083 -387 -5079
rect -375 -5083 -374 -5079
rect -372 -5083 -367 -5079
rect -363 -5083 -358 -5079
rect -356 -5083 -355 -5079
rect -351 -5083 -350 -5079
rect -348 -5083 -346 -5079
rect -342 -5083 -340 -5079
rect -338 -5083 -337 -5079
rect -215 -5083 -214 -5079
rect -212 -5083 -210 -5079
rect -206 -5083 -204 -5079
rect -202 -5083 -201 -5079
rect -189 -5083 -188 -5079
rect -186 -5083 -184 -5079
rect -180 -5083 -178 -5079
rect -176 -5083 -175 -5079
rect -163 -5083 -162 -5079
rect -160 -5083 -159 -5079
rect -155 -5083 -152 -5079
rect -150 -5083 -144 -5079
rect -142 -5083 -141 -5079
rect -137 -5083 -134 -5079
rect -132 -5083 -131 -5079
rect -119 -5083 -118 -5079
rect -116 -5083 -110 -5079
rect -108 -5083 -106 -5079
rect -102 -5083 -100 -5079
rect -98 -5083 -97 -5079
rect -85 -5083 -84 -5079
rect -82 -5083 -80 -5079
rect -76 -5083 -74 -5079
rect -72 -5083 -66 -5079
rect -64 -5083 -62 -5079
rect -58 -5083 -56 -5079
rect -54 -5083 -53 -5079
rect -41 -5083 -40 -5079
rect -38 -5083 -32 -5079
rect -30 -5083 -29 -5079
rect -17 -5083 -16 -5079
rect -14 -5083 -9 -5079
rect -5 -5083 0 -5079
rect 2 -5083 3 -5079
rect 7 -5083 8 -5079
rect 10 -5083 12 -5079
rect 16 -5083 18 -5079
rect 20 -5083 21 -5079
rect 143 -5083 144 -5079
rect 146 -5083 148 -5079
rect 152 -5083 154 -5079
rect 156 -5083 157 -5079
rect 169 -5083 170 -5079
rect 172 -5083 174 -5079
rect 178 -5083 180 -5079
rect 182 -5083 183 -5079
rect 195 -5083 196 -5079
rect 198 -5083 199 -5079
rect 203 -5083 206 -5079
rect 208 -5083 214 -5079
rect 216 -5083 217 -5079
rect 221 -5083 224 -5079
rect 226 -5083 227 -5079
rect 239 -5083 240 -5079
rect 242 -5083 248 -5079
rect 250 -5083 252 -5079
rect 256 -5083 258 -5079
rect 260 -5083 261 -5079
rect 273 -5083 274 -5079
rect 276 -5083 278 -5079
rect 282 -5083 284 -5079
rect 286 -5083 292 -5079
rect 294 -5083 296 -5079
rect 300 -5083 302 -5079
rect 304 -5083 305 -5079
rect 317 -5083 318 -5079
rect 320 -5083 326 -5079
rect 328 -5083 329 -5079
rect 341 -5083 342 -5079
rect 344 -5083 349 -5079
rect 353 -5083 358 -5079
rect 360 -5083 361 -5079
rect 365 -5083 366 -5079
rect 368 -5083 370 -5079
rect 374 -5083 376 -5079
rect 378 -5083 379 -5079
rect 499 -5083 500 -5079
rect 502 -5083 504 -5079
rect 508 -5083 510 -5079
rect 512 -5083 513 -5079
rect 525 -5083 526 -5079
rect 528 -5083 530 -5079
rect 534 -5083 536 -5079
rect 538 -5083 539 -5079
rect 551 -5083 552 -5079
rect 554 -5083 555 -5079
rect 559 -5083 562 -5079
rect 564 -5083 570 -5079
rect 572 -5083 573 -5079
rect 577 -5083 580 -5079
rect 582 -5083 583 -5079
rect 595 -5083 596 -5079
rect 598 -5083 604 -5079
rect 606 -5083 608 -5079
rect 612 -5083 614 -5079
rect 616 -5083 617 -5079
rect 629 -5083 630 -5079
rect 632 -5083 634 -5079
rect 638 -5083 640 -5079
rect 642 -5083 648 -5079
rect 650 -5083 652 -5079
rect 656 -5083 658 -5079
rect 660 -5083 661 -5079
rect 673 -5083 674 -5079
rect 676 -5083 682 -5079
rect 684 -5083 685 -5079
rect 697 -5083 698 -5079
rect 700 -5083 705 -5079
rect 709 -5083 714 -5079
rect 716 -5083 717 -5079
rect 721 -5083 722 -5079
rect 724 -5083 726 -5079
rect 730 -5083 732 -5079
rect 734 -5083 735 -5079
rect 857 -5083 858 -5079
rect 860 -5083 862 -5079
rect 866 -5083 868 -5079
rect 870 -5083 871 -5079
rect 883 -5083 884 -5079
rect 886 -5083 888 -5079
rect 892 -5083 894 -5079
rect 896 -5083 897 -5079
rect 909 -5083 910 -5079
rect 912 -5083 913 -5079
rect 917 -5083 920 -5079
rect 922 -5083 928 -5079
rect 930 -5083 931 -5079
rect 935 -5083 938 -5079
rect 940 -5083 941 -5079
rect 953 -5083 954 -5079
rect 956 -5083 962 -5079
rect 964 -5083 966 -5079
rect 970 -5083 972 -5079
rect 974 -5083 975 -5079
rect 987 -5083 988 -5079
rect 990 -5083 992 -5079
rect 996 -5083 998 -5079
rect 1000 -5083 1006 -5079
rect 1008 -5083 1010 -5079
rect 1014 -5083 1016 -5079
rect 1018 -5083 1019 -5079
rect 1031 -5083 1032 -5079
rect 1034 -5083 1040 -5079
rect 1042 -5083 1043 -5079
rect 1055 -5083 1056 -5079
rect 1058 -5083 1063 -5079
rect 1067 -5083 1072 -5079
rect 1074 -5083 1075 -5079
rect 1079 -5083 1080 -5079
rect 1082 -5083 1084 -5079
rect 1088 -5083 1090 -5079
rect 1092 -5083 1093 -5079
rect 1215 -5083 1216 -5079
rect 1218 -5083 1220 -5079
rect 1224 -5083 1226 -5079
rect 1228 -5083 1229 -5079
rect 1241 -5083 1242 -5079
rect 1244 -5083 1246 -5079
rect 1250 -5083 1252 -5079
rect 1254 -5083 1255 -5079
rect 1267 -5083 1268 -5079
rect 1270 -5083 1271 -5079
rect 1275 -5083 1278 -5079
rect 1280 -5083 1286 -5079
rect 1288 -5083 1289 -5079
rect 1293 -5083 1296 -5079
rect 1298 -5083 1299 -5079
rect 1311 -5083 1312 -5079
rect 1314 -5083 1320 -5079
rect 1322 -5083 1324 -5079
rect 1328 -5083 1330 -5079
rect 1332 -5083 1333 -5079
rect 1345 -5083 1346 -5079
rect 1348 -5083 1350 -5079
rect 1354 -5083 1356 -5079
rect 1358 -5083 1364 -5079
rect 1366 -5083 1368 -5079
rect 1372 -5083 1374 -5079
rect 1376 -5083 1377 -5079
rect 1389 -5083 1390 -5079
rect 1392 -5083 1398 -5079
rect 1400 -5083 1401 -5079
rect 1413 -5083 1414 -5079
rect 1416 -5083 1421 -5079
rect 1425 -5083 1430 -5079
rect 1432 -5083 1433 -5079
rect 1437 -5083 1438 -5079
rect 1440 -5083 1442 -5079
rect 1446 -5083 1448 -5079
rect 1450 -5083 1451 -5079
rect -1806 -5202 -1805 -5198
rect -1803 -5202 -1801 -5198
rect -1797 -5202 -1795 -5198
rect -1793 -5202 -1792 -5198
rect -1780 -5202 -1779 -5198
rect -1777 -5202 -1771 -5198
rect -1769 -5202 -1768 -5198
rect -1756 -5202 -1755 -5198
rect -1753 -5202 -1747 -5198
rect -1745 -5202 -1743 -5198
rect -1739 -5202 -1737 -5198
rect -1735 -5202 -1729 -5198
rect -1727 -5202 -1726 -5198
rect -1714 -5202 -1713 -5198
rect -1711 -5202 -1705 -5198
rect -1703 -5202 -1701 -5198
rect -1697 -5202 -1695 -5198
rect -1693 -5202 -1687 -5198
rect -1685 -5202 -1684 -5198
rect -1672 -5202 -1671 -5198
rect -1669 -5202 -1663 -5198
rect -1661 -5202 -1659 -5198
rect -1655 -5202 -1653 -5198
rect -1651 -5202 -1645 -5198
rect -1643 -5202 -1642 -5198
rect -1630 -5202 -1629 -5198
rect -1627 -5202 -1621 -5198
rect -1619 -5202 -1618 -5198
rect -1543 -5202 -1542 -5198
rect -1540 -5202 -1538 -5198
rect -1534 -5202 -1532 -5198
rect -1530 -5202 -1529 -5198
rect -1517 -5202 -1516 -5198
rect -1514 -5202 -1508 -5198
rect -1506 -5202 -1505 -5198
rect -1493 -5202 -1492 -5198
rect -1490 -5202 -1484 -5198
rect -1482 -5202 -1480 -5198
rect -1476 -5202 -1474 -5198
rect -1472 -5202 -1466 -5198
rect -1464 -5202 -1463 -5198
rect -1451 -5202 -1450 -5198
rect -1448 -5202 -1442 -5198
rect -1440 -5202 -1438 -5198
rect -1434 -5202 -1432 -5198
rect -1430 -5202 -1424 -5198
rect -1422 -5202 -1421 -5198
rect -1409 -5202 -1408 -5198
rect -1406 -5202 -1400 -5198
rect -1398 -5202 -1396 -5198
rect -1392 -5202 -1390 -5198
rect -1388 -5202 -1382 -5198
rect -1380 -5202 -1379 -5198
rect -1367 -5202 -1366 -5198
rect -1364 -5202 -1358 -5198
rect -1356 -5202 -1355 -5198
rect -1230 -5202 -1229 -5198
rect -1227 -5202 -1225 -5198
rect -1221 -5202 -1219 -5198
rect -1217 -5202 -1216 -5198
rect -1204 -5202 -1203 -5198
rect -1201 -5202 -1195 -5198
rect -1193 -5202 -1192 -5198
rect -1180 -5202 -1179 -5198
rect -1177 -5202 -1171 -5198
rect -1169 -5202 -1167 -5198
rect -1163 -5202 -1161 -5198
rect -1159 -5202 -1153 -5198
rect -1151 -5202 -1150 -5198
rect -1138 -5202 -1137 -5198
rect -1135 -5202 -1129 -5198
rect -1127 -5202 -1125 -5198
rect -1121 -5202 -1119 -5198
rect -1117 -5202 -1111 -5198
rect -1109 -5202 -1108 -5198
rect -1096 -5202 -1095 -5198
rect -1093 -5202 -1087 -5198
rect -1085 -5202 -1083 -5198
rect -1079 -5202 -1077 -5198
rect -1075 -5202 -1069 -5198
rect -1067 -5202 -1066 -5198
rect -1054 -5202 -1053 -5198
rect -1051 -5202 -1045 -5198
rect -1043 -5202 -1042 -5198
rect -931 -5202 -930 -5198
rect -928 -5202 -926 -5198
rect -922 -5202 -920 -5198
rect -918 -5202 -917 -5198
rect -905 -5202 -904 -5198
rect -902 -5202 -896 -5198
rect -894 -5202 -893 -5198
rect -881 -5202 -880 -5198
rect -878 -5202 -872 -5198
rect -870 -5202 -868 -5198
rect -864 -5202 -862 -5198
rect -860 -5202 -854 -5198
rect -852 -5202 -851 -5198
rect -839 -5202 -838 -5198
rect -836 -5202 -830 -5198
rect -828 -5202 -826 -5198
rect -822 -5202 -820 -5198
rect -818 -5202 -812 -5198
rect -810 -5202 -809 -5198
rect -797 -5202 -796 -5198
rect -794 -5202 -788 -5198
rect -786 -5202 -784 -5198
rect -780 -5202 -778 -5198
rect -776 -5202 -770 -5198
rect -768 -5202 -767 -5198
rect -755 -5202 -754 -5198
rect -752 -5202 -746 -5198
rect -744 -5202 -743 -5198
rect -1806 -5373 -1805 -5369
rect -1803 -5373 -1801 -5369
rect -1797 -5373 -1795 -5369
rect -1793 -5373 -1792 -5369
rect -1780 -5373 -1779 -5369
rect -1777 -5373 -1771 -5369
rect -1769 -5373 -1768 -5369
rect -1756 -5373 -1755 -5369
rect -1753 -5373 -1747 -5369
rect -1745 -5373 -1743 -5369
rect -1739 -5373 -1737 -5369
rect -1735 -5373 -1729 -5369
rect -1727 -5373 -1726 -5369
rect -1714 -5373 -1713 -5369
rect -1711 -5373 -1705 -5369
rect -1703 -5373 -1701 -5369
rect -1697 -5373 -1695 -5369
rect -1693 -5373 -1687 -5369
rect -1685 -5373 -1684 -5369
rect -1672 -5373 -1671 -5369
rect -1669 -5373 -1663 -5369
rect -1661 -5373 -1659 -5369
rect -1655 -5373 -1653 -5369
rect -1651 -5373 -1645 -5369
rect -1643 -5373 -1642 -5369
rect -1630 -5373 -1629 -5369
rect -1627 -5373 -1621 -5369
rect -1619 -5373 -1618 -5369
rect -1543 -5373 -1542 -5369
rect -1540 -5373 -1538 -5369
rect -1534 -5373 -1532 -5369
rect -1530 -5373 -1529 -5369
rect -1517 -5373 -1516 -5369
rect -1514 -5373 -1508 -5369
rect -1506 -5373 -1505 -5369
rect -1493 -5373 -1492 -5369
rect -1490 -5373 -1484 -5369
rect -1482 -5373 -1480 -5369
rect -1476 -5373 -1474 -5369
rect -1472 -5373 -1466 -5369
rect -1464 -5373 -1463 -5369
rect -1451 -5373 -1450 -5369
rect -1448 -5373 -1442 -5369
rect -1440 -5373 -1438 -5369
rect -1434 -5373 -1432 -5369
rect -1430 -5373 -1424 -5369
rect -1422 -5373 -1421 -5369
rect -1409 -5373 -1408 -5369
rect -1406 -5373 -1400 -5369
rect -1398 -5373 -1396 -5369
rect -1392 -5373 -1390 -5369
rect -1388 -5373 -1382 -5369
rect -1380 -5373 -1379 -5369
rect -1367 -5373 -1366 -5369
rect -1364 -5373 -1358 -5369
rect -1356 -5373 -1355 -5369
rect -1230 -5373 -1229 -5369
rect -1227 -5373 -1225 -5369
rect -1221 -5373 -1219 -5369
rect -1217 -5373 -1216 -5369
rect -1204 -5373 -1203 -5369
rect -1201 -5373 -1195 -5369
rect -1193 -5373 -1192 -5369
rect -1180 -5373 -1179 -5369
rect -1177 -5373 -1171 -5369
rect -1169 -5373 -1167 -5369
rect -1163 -5373 -1161 -5369
rect -1159 -5373 -1153 -5369
rect -1151 -5373 -1150 -5369
rect -1138 -5373 -1137 -5369
rect -1135 -5373 -1129 -5369
rect -1127 -5373 -1125 -5369
rect -1121 -5373 -1119 -5369
rect -1117 -5373 -1111 -5369
rect -1109 -5373 -1108 -5369
rect -1096 -5373 -1095 -5369
rect -1093 -5373 -1087 -5369
rect -1085 -5373 -1083 -5369
rect -1079 -5373 -1077 -5369
rect -1075 -5373 -1069 -5369
rect -1067 -5373 -1066 -5369
rect -1054 -5373 -1053 -5369
rect -1051 -5373 -1045 -5369
rect -1043 -5373 -1042 -5369
rect -931 -5373 -930 -5369
rect -928 -5373 -926 -5369
rect -922 -5373 -920 -5369
rect -918 -5373 -917 -5369
rect -905 -5373 -904 -5369
rect -902 -5373 -896 -5369
rect -894 -5373 -893 -5369
rect -881 -5373 -880 -5369
rect -878 -5373 -872 -5369
rect -870 -5373 -868 -5369
rect -864 -5373 -862 -5369
rect -860 -5373 -854 -5369
rect -852 -5373 -851 -5369
rect -839 -5373 -838 -5369
rect -836 -5373 -830 -5369
rect -828 -5373 -826 -5369
rect -822 -5373 -820 -5369
rect -818 -5373 -812 -5369
rect -810 -5373 -809 -5369
rect -797 -5373 -796 -5369
rect -794 -5373 -788 -5369
rect -786 -5373 -784 -5369
rect -780 -5373 -778 -5369
rect -776 -5373 -770 -5369
rect -768 -5373 -767 -5369
rect -755 -5373 -754 -5369
rect -752 -5373 -746 -5369
rect -744 -5373 -743 -5369
rect -573 -5373 -572 -5369
rect -570 -5373 -568 -5369
rect -564 -5373 -562 -5369
rect -560 -5373 -559 -5369
rect -547 -5373 -546 -5369
rect -544 -5373 -538 -5369
rect -536 -5373 -535 -5369
rect -523 -5373 -522 -5369
rect -520 -5373 -514 -5369
rect -512 -5373 -510 -5369
rect -506 -5373 -504 -5369
rect -502 -5373 -496 -5369
rect -494 -5373 -493 -5369
rect -481 -5373 -480 -5369
rect -478 -5373 -472 -5369
rect -470 -5373 -468 -5369
rect -464 -5373 -462 -5369
rect -460 -5373 -454 -5369
rect -452 -5373 -451 -5369
rect -439 -5373 -438 -5369
rect -436 -5373 -430 -5369
rect -428 -5373 -426 -5369
rect -422 -5373 -420 -5369
rect -418 -5373 -412 -5369
rect -410 -5373 -409 -5369
rect -397 -5373 -396 -5369
rect -394 -5373 -388 -5369
rect -386 -5373 -385 -5369
rect -215 -5373 -214 -5369
rect -212 -5373 -210 -5369
rect -206 -5373 -204 -5369
rect -202 -5373 -201 -5369
rect -189 -5373 -188 -5369
rect -186 -5373 -180 -5369
rect -178 -5373 -177 -5369
rect -165 -5373 -164 -5369
rect -162 -5373 -156 -5369
rect -154 -5373 -152 -5369
rect -148 -5373 -146 -5369
rect -144 -5373 -138 -5369
rect -136 -5373 -135 -5369
rect -123 -5373 -122 -5369
rect -120 -5373 -114 -5369
rect -112 -5373 -110 -5369
rect -106 -5373 -104 -5369
rect -102 -5373 -96 -5369
rect -94 -5373 -93 -5369
rect -81 -5373 -80 -5369
rect -78 -5373 -72 -5369
rect -70 -5373 -68 -5369
rect -64 -5373 -62 -5369
rect -60 -5373 -54 -5369
rect -52 -5373 -51 -5369
rect -39 -5373 -38 -5369
rect -36 -5373 -30 -5369
rect -28 -5373 -27 -5369
rect 143 -5373 144 -5369
rect 146 -5373 148 -5369
rect 152 -5373 154 -5369
rect 156 -5373 157 -5369
rect 169 -5373 170 -5369
rect 172 -5373 178 -5369
rect 180 -5373 181 -5369
rect 193 -5373 194 -5369
rect 196 -5373 202 -5369
rect 204 -5373 206 -5369
rect 210 -5373 212 -5369
rect 214 -5373 220 -5369
rect 222 -5373 223 -5369
rect 235 -5373 236 -5369
rect 238 -5373 244 -5369
rect 246 -5373 248 -5369
rect 252 -5373 254 -5369
rect 256 -5373 262 -5369
rect 264 -5373 265 -5369
rect 277 -5373 278 -5369
rect 280 -5373 286 -5369
rect 288 -5373 290 -5369
rect 294 -5373 296 -5369
rect 298 -5373 304 -5369
rect 306 -5373 307 -5369
rect 319 -5373 320 -5369
rect 322 -5373 328 -5369
rect 330 -5373 331 -5369
rect 499 -5373 500 -5369
rect 502 -5373 504 -5369
rect 508 -5373 510 -5369
rect 512 -5373 513 -5369
rect 525 -5373 526 -5369
rect 528 -5373 534 -5369
rect 536 -5373 537 -5369
rect 549 -5373 550 -5369
rect 552 -5373 558 -5369
rect 560 -5373 562 -5369
rect 566 -5373 568 -5369
rect 570 -5373 576 -5369
rect 578 -5373 579 -5369
rect 591 -5373 592 -5369
rect 594 -5373 600 -5369
rect 602 -5373 604 -5369
rect 608 -5373 610 -5369
rect 612 -5373 618 -5369
rect 620 -5373 621 -5369
rect 633 -5373 634 -5369
rect 636 -5373 642 -5369
rect 644 -5373 646 -5369
rect 650 -5373 652 -5369
rect 654 -5373 660 -5369
rect 662 -5373 663 -5369
rect 675 -5373 676 -5369
rect 678 -5373 684 -5369
rect 686 -5373 687 -5369
rect 857 -5373 858 -5369
rect 860 -5373 862 -5369
rect 866 -5373 868 -5369
rect 870 -5373 871 -5369
rect 883 -5373 884 -5369
rect 886 -5373 892 -5369
rect 894 -5373 895 -5369
rect 907 -5373 908 -5369
rect 910 -5373 916 -5369
rect 918 -5373 920 -5369
rect 924 -5373 926 -5369
rect 928 -5373 934 -5369
rect 936 -5373 937 -5369
rect 949 -5373 950 -5369
rect 952 -5373 958 -5369
rect 960 -5373 962 -5369
rect 966 -5373 968 -5369
rect 970 -5373 976 -5369
rect 978 -5373 979 -5369
rect 991 -5373 992 -5369
rect 994 -5373 1000 -5369
rect 1002 -5373 1004 -5369
rect 1008 -5373 1010 -5369
rect 1012 -5373 1018 -5369
rect 1020 -5373 1021 -5369
rect 1033 -5373 1034 -5369
rect 1036 -5373 1042 -5369
rect 1044 -5373 1045 -5369
rect 1215 -5373 1216 -5369
rect 1218 -5373 1220 -5369
rect 1224 -5373 1226 -5369
rect 1228 -5373 1229 -5369
rect 1241 -5373 1242 -5369
rect 1244 -5373 1250 -5369
rect 1252 -5373 1253 -5369
rect 1265 -5373 1266 -5369
rect 1268 -5373 1274 -5369
rect 1276 -5373 1278 -5369
rect 1282 -5373 1284 -5369
rect 1286 -5373 1292 -5369
rect 1294 -5373 1295 -5369
rect 1307 -5373 1308 -5369
rect 1310 -5373 1316 -5369
rect 1318 -5373 1320 -5369
rect 1324 -5373 1326 -5369
rect 1328 -5373 1334 -5369
rect 1336 -5373 1337 -5369
rect 1349 -5373 1350 -5369
rect 1352 -5373 1358 -5369
rect 1360 -5373 1362 -5369
rect 1366 -5373 1368 -5369
rect 1370 -5373 1376 -5369
rect 1378 -5373 1379 -5369
rect 1391 -5373 1392 -5369
rect 1394 -5373 1400 -5369
rect 1402 -5373 1403 -5369
rect -1806 -5533 -1805 -5529
rect -1803 -5533 -1801 -5529
rect -1797 -5533 -1795 -5529
rect -1793 -5533 -1792 -5529
rect -1780 -5533 -1779 -5529
rect -1777 -5533 -1771 -5529
rect -1769 -5533 -1768 -5529
rect -1756 -5533 -1755 -5529
rect -1753 -5533 -1747 -5529
rect -1745 -5533 -1743 -5529
rect -1739 -5533 -1737 -5529
rect -1735 -5533 -1729 -5529
rect -1727 -5533 -1726 -5529
rect -1714 -5533 -1713 -5529
rect -1711 -5533 -1705 -5529
rect -1703 -5533 -1701 -5529
rect -1697 -5533 -1695 -5529
rect -1693 -5533 -1687 -5529
rect -1685 -5533 -1684 -5529
rect -1672 -5533 -1671 -5529
rect -1669 -5533 -1663 -5529
rect -1661 -5533 -1659 -5529
rect -1655 -5533 -1653 -5529
rect -1651 -5533 -1645 -5529
rect -1643 -5533 -1642 -5529
rect -1630 -5533 -1629 -5529
rect -1627 -5533 -1621 -5529
rect -1619 -5533 -1618 -5529
rect -1543 -5533 -1542 -5529
rect -1540 -5533 -1538 -5529
rect -1534 -5533 -1532 -5529
rect -1530 -5533 -1529 -5529
rect -1517 -5533 -1516 -5529
rect -1514 -5533 -1508 -5529
rect -1506 -5533 -1505 -5529
rect -1493 -5533 -1492 -5529
rect -1490 -5533 -1484 -5529
rect -1482 -5533 -1480 -5529
rect -1476 -5533 -1474 -5529
rect -1472 -5533 -1466 -5529
rect -1464 -5533 -1463 -5529
rect -1451 -5533 -1450 -5529
rect -1448 -5533 -1442 -5529
rect -1440 -5533 -1438 -5529
rect -1434 -5533 -1432 -5529
rect -1430 -5533 -1424 -5529
rect -1422 -5533 -1421 -5529
rect -1409 -5533 -1408 -5529
rect -1406 -5533 -1400 -5529
rect -1398 -5533 -1396 -5529
rect -1392 -5533 -1390 -5529
rect -1388 -5533 -1382 -5529
rect -1380 -5533 -1379 -5529
rect -1367 -5533 -1366 -5529
rect -1364 -5533 -1358 -5529
rect -1356 -5533 -1355 -5529
rect -1230 -5533 -1229 -5529
rect -1227 -5533 -1225 -5529
rect -1221 -5533 -1219 -5529
rect -1217 -5533 -1216 -5529
rect -1204 -5533 -1203 -5529
rect -1201 -5533 -1195 -5529
rect -1193 -5533 -1192 -5529
rect -1180 -5533 -1179 -5529
rect -1177 -5533 -1171 -5529
rect -1169 -5533 -1167 -5529
rect -1163 -5533 -1161 -5529
rect -1159 -5533 -1153 -5529
rect -1151 -5533 -1150 -5529
rect -1138 -5533 -1137 -5529
rect -1135 -5533 -1129 -5529
rect -1127 -5533 -1125 -5529
rect -1121 -5533 -1119 -5529
rect -1117 -5533 -1111 -5529
rect -1109 -5533 -1108 -5529
rect -1096 -5533 -1095 -5529
rect -1093 -5533 -1087 -5529
rect -1085 -5533 -1083 -5529
rect -1079 -5533 -1077 -5529
rect -1075 -5533 -1069 -5529
rect -1067 -5533 -1066 -5529
rect -1054 -5533 -1053 -5529
rect -1051 -5533 -1045 -5529
rect -1043 -5533 -1042 -5529
rect -931 -5533 -930 -5529
rect -928 -5533 -926 -5529
rect -922 -5533 -920 -5529
rect -918 -5533 -917 -5529
rect -905 -5533 -904 -5529
rect -902 -5533 -896 -5529
rect -894 -5533 -893 -5529
rect -881 -5533 -880 -5529
rect -878 -5533 -872 -5529
rect -870 -5533 -868 -5529
rect -864 -5533 -862 -5529
rect -860 -5533 -854 -5529
rect -852 -5533 -851 -5529
rect -839 -5533 -838 -5529
rect -836 -5533 -830 -5529
rect -828 -5533 -826 -5529
rect -822 -5533 -820 -5529
rect -818 -5533 -812 -5529
rect -810 -5533 -809 -5529
rect -797 -5533 -796 -5529
rect -794 -5533 -788 -5529
rect -786 -5533 -784 -5529
rect -780 -5533 -778 -5529
rect -776 -5533 -770 -5529
rect -768 -5533 -767 -5529
rect -755 -5533 -754 -5529
rect -752 -5533 -746 -5529
rect -744 -5533 -743 -5529
rect -573 -5533 -572 -5529
rect -570 -5533 -568 -5529
rect -564 -5533 -562 -5529
rect -560 -5533 -559 -5529
rect -547 -5533 -546 -5529
rect -544 -5533 -538 -5529
rect -536 -5533 -535 -5529
rect -523 -5533 -522 -5529
rect -520 -5533 -514 -5529
rect -512 -5533 -510 -5529
rect -506 -5533 -504 -5529
rect -502 -5533 -496 -5529
rect -494 -5533 -493 -5529
rect -481 -5533 -480 -5529
rect -478 -5533 -472 -5529
rect -470 -5533 -468 -5529
rect -464 -5533 -462 -5529
rect -460 -5533 -454 -5529
rect -452 -5533 -451 -5529
rect -439 -5533 -438 -5529
rect -436 -5533 -430 -5529
rect -428 -5533 -426 -5529
rect -422 -5533 -420 -5529
rect -418 -5533 -412 -5529
rect -410 -5533 -409 -5529
rect -397 -5533 -396 -5529
rect -394 -5533 -388 -5529
rect -386 -5533 -385 -5529
rect -215 -5533 -214 -5529
rect -212 -5533 -210 -5529
rect -206 -5533 -204 -5529
rect -202 -5533 -201 -5529
rect -189 -5533 -188 -5529
rect -186 -5533 -180 -5529
rect -178 -5533 -177 -5529
rect -165 -5533 -164 -5529
rect -162 -5533 -156 -5529
rect -154 -5533 -152 -5529
rect -148 -5533 -146 -5529
rect -144 -5533 -138 -5529
rect -136 -5533 -135 -5529
rect -123 -5533 -122 -5529
rect -120 -5533 -114 -5529
rect -112 -5533 -110 -5529
rect -106 -5533 -104 -5529
rect -102 -5533 -96 -5529
rect -94 -5533 -93 -5529
rect -81 -5533 -80 -5529
rect -78 -5533 -72 -5529
rect -70 -5533 -68 -5529
rect -64 -5533 -62 -5529
rect -60 -5533 -54 -5529
rect -52 -5533 -51 -5529
rect -39 -5533 -38 -5529
rect -36 -5533 -30 -5529
rect -28 -5533 -27 -5529
rect 143 -5533 144 -5529
rect 146 -5533 148 -5529
rect 152 -5533 154 -5529
rect 156 -5533 157 -5529
rect 169 -5533 170 -5529
rect 172 -5533 178 -5529
rect 180 -5533 181 -5529
rect 193 -5533 194 -5529
rect 196 -5533 202 -5529
rect 204 -5533 206 -5529
rect 210 -5533 212 -5529
rect 214 -5533 220 -5529
rect 222 -5533 223 -5529
rect 235 -5533 236 -5529
rect 238 -5533 244 -5529
rect 246 -5533 248 -5529
rect 252 -5533 254 -5529
rect 256 -5533 262 -5529
rect 264 -5533 265 -5529
rect 277 -5533 278 -5529
rect 280 -5533 286 -5529
rect 288 -5533 290 -5529
rect 294 -5533 296 -5529
rect 298 -5533 304 -5529
rect 306 -5533 307 -5529
rect 319 -5533 320 -5529
rect 322 -5533 328 -5529
rect 330 -5533 331 -5529
rect 499 -5533 500 -5529
rect 502 -5533 504 -5529
rect 508 -5533 510 -5529
rect 512 -5533 513 -5529
rect 525 -5533 526 -5529
rect 528 -5533 534 -5529
rect 536 -5533 537 -5529
rect 549 -5533 550 -5529
rect 552 -5533 558 -5529
rect 560 -5533 562 -5529
rect 566 -5533 568 -5529
rect 570 -5533 576 -5529
rect 578 -5533 579 -5529
rect 591 -5533 592 -5529
rect 594 -5533 600 -5529
rect 602 -5533 604 -5529
rect 608 -5533 610 -5529
rect 612 -5533 618 -5529
rect 620 -5533 621 -5529
rect 633 -5533 634 -5529
rect 636 -5533 642 -5529
rect 644 -5533 646 -5529
rect 650 -5533 652 -5529
rect 654 -5533 660 -5529
rect 662 -5533 663 -5529
rect 675 -5533 676 -5529
rect 678 -5533 684 -5529
rect 686 -5533 687 -5529
rect 857 -5533 858 -5529
rect 860 -5533 862 -5529
rect 866 -5533 868 -5529
rect 870 -5533 871 -5529
rect 883 -5533 884 -5529
rect 886 -5533 892 -5529
rect 894 -5533 895 -5529
rect 907 -5533 908 -5529
rect 910 -5533 916 -5529
rect 918 -5533 920 -5529
rect 924 -5533 926 -5529
rect 928 -5533 934 -5529
rect 936 -5533 937 -5529
rect 949 -5533 950 -5529
rect 952 -5533 958 -5529
rect 960 -5533 962 -5529
rect 966 -5533 968 -5529
rect 970 -5533 976 -5529
rect 978 -5533 979 -5529
rect 991 -5533 992 -5529
rect 994 -5533 1000 -5529
rect 1002 -5533 1004 -5529
rect 1008 -5533 1010 -5529
rect 1012 -5533 1018 -5529
rect 1020 -5533 1021 -5529
rect 1033 -5533 1034 -5529
rect 1036 -5533 1042 -5529
rect 1044 -5533 1045 -5529
rect 1215 -5533 1216 -5529
rect 1218 -5533 1220 -5529
rect 1224 -5533 1226 -5529
rect 1228 -5533 1229 -5529
rect 1241 -5533 1242 -5529
rect 1244 -5533 1250 -5529
rect 1252 -5533 1253 -5529
rect 1265 -5533 1266 -5529
rect 1268 -5533 1274 -5529
rect 1276 -5533 1278 -5529
rect 1282 -5533 1284 -5529
rect 1286 -5533 1292 -5529
rect 1294 -5533 1295 -5529
rect 1307 -5533 1308 -5529
rect 1310 -5533 1316 -5529
rect 1318 -5533 1320 -5529
rect 1324 -5533 1326 -5529
rect 1328 -5533 1334 -5529
rect 1336 -5533 1337 -5529
rect 1349 -5533 1350 -5529
rect 1352 -5533 1358 -5529
rect 1360 -5533 1362 -5529
rect 1366 -5533 1368 -5529
rect 1370 -5533 1376 -5529
rect 1378 -5533 1379 -5529
rect 1391 -5533 1392 -5529
rect 1394 -5533 1400 -5529
rect 1402 -5533 1403 -5529
rect -1305 -5647 -1304 -5643
rect -1302 -5647 -1296 -5643
rect -1294 -5647 -1292 -5643
rect -1288 -5647 -1286 -5643
rect -1284 -5647 -1283 -5643
rect -931 -5647 -930 -5643
rect -928 -5647 -922 -5643
rect -920 -5647 -918 -5643
rect -914 -5647 -912 -5643
rect -910 -5647 -909 -5643
rect -573 -5647 -572 -5643
rect -570 -5647 -564 -5643
rect -562 -5647 -560 -5643
rect -556 -5647 -554 -5643
rect -552 -5647 -551 -5643
rect -215 -5647 -214 -5643
rect -212 -5647 -206 -5643
rect -204 -5647 -202 -5643
rect -198 -5647 -196 -5643
rect -194 -5647 -193 -5643
rect 143 -5647 144 -5643
rect 146 -5647 152 -5643
rect 154 -5647 156 -5643
rect 160 -5647 162 -5643
rect 164 -5647 165 -5643
rect 499 -5647 500 -5643
rect 502 -5647 508 -5643
rect 510 -5647 512 -5643
rect 516 -5647 518 -5643
rect 520 -5647 521 -5643
rect 857 -5647 858 -5643
rect 860 -5647 866 -5643
rect 868 -5647 870 -5643
rect 874 -5647 876 -5643
rect 878 -5647 879 -5643
rect 1215 -5647 1216 -5643
rect 1218 -5647 1224 -5643
rect 1226 -5647 1228 -5643
rect 1232 -5647 1234 -5643
rect 1236 -5647 1237 -5643
rect -1230 -5806 -1229 -5802
rect -1227 -5806 -1225 -5802
rect -1221 -5806 -1219 -5802
rect -1217 -5806 -1216 -5802
rect -1204 -5806 -1203 -5802
rect -1201 -5806 -1199 -5802
rect -1195 -5806 -1193 -5802
rect -1191 -5806 -1185 -5802
rect -1183 -5806 -1181 -5802
rect -1177 -5806 -1175 -5802
rect -1173 -5806 -1172 -5802
rect -1160 -5806 -1159 -5802
rect -1157 -5806 -1151 -5802
rect -1149 -5806 -1147 -5802
rect -1143 -5806 -1141 -5802
rect -1139 -5806 -1138 -5802
rect -931 -5806 -930 -5802
rect -928 -5806 -926 -5802
rect -922 -5806 -920 -5802
rect -918 -5806 -917 -5802
rect -905 -5806 -904 -5802
rect -902 -5806 -900 -5802
rect -896 -5806 -894 -5802
rect -892 -5806 -891 -5802
rect -879 -5806 -878 -5802
rect -876 -5806 -875 -5802
rect -871 -5806 -868 -5802
rect -866 -5806 -860 -5802
rect -858 -5806 -857 -5802
rect -853 -5806 -850 -5802
rect -848 -5806 -847 -5802
rect -835 -5806 -834 -5802
rect -832 -5806 -826 -5802
rect -824 -5806 -822 -5802
rect -818 -5806 -816 -5802
rect -814 -5806 -813 -5802
rect -801 -5806 -800 -5802
rect -798 -5806 -796 -5802
rect -792 -5806 -790 -5802
rect -788 -5806 -782 -5802
rect -780 -5806 -778 -5802
rect -774 -5806 -772 -5802
rect -770 -5806 -769 -5802
rect -757 -5806 -756 -5802
rect -754 -5806 -748 -5802
rect -746 -5806 -745 -5802
rect -733 -5806 -732 -5802
rect -730 -5806 -725 -5802
rect -721 -5806 -716 -5802
rect -714 -5806 -713 -5802
rect -709 -5806 -708 -5802
rect -706 -5806 -704 -5802
rect -700 -5806 -698 -5802
rect -696 -5806 -695 -5802
rect -573 -5806 -572 -5802
rect -570 -5806 -568 -5802
rect -564 -5806 -562 -5802
rect -560 -5806 -559 -5802
rect -547 -5806 -546 -5802
rect -544 -5806 -542 -5802
rect -538 -5806 -536 -5802
rect -534 -5806 -533 -5802
rect -521 -5806 -520 -5802
rect -518 -5806 -517 -5802
rect -513 -5806 -510 -5802
rect -508 -5806 -502 -5802
rect -500 -5806 -499 -5802
rect -495 -5806 -492 -5802
rect -490 -5806 -489 -5802
rect -477 -5806 -476 -5802
rect -474 -5806 -468 -5802
rect -466 -5806 -464 -5802
rect -460 -5806 -458 -5802
rect -456 -5806 -455 -5802
rect -443 -5806 -442 -5802
rect -440 -5806 -438 -5802
rect -434 -5806 -432 -5802
rect -430 -5806 -424 -5802
rect -422 -5806 -420 -5802
rect -416 -5806 -414 -5802
rect -412 -5806 -411 -5802
rect -399 -5806 -398 -5802
rect -396 -5806 -390 -5802
rect -388 -5806 -387 -5802
rect -375 -5806 -374 -5802
rect -372 -5806 -367 -5802
rect -363 -5806 -358 -5802
rect -356 -5806 -355 -5802
rect -351 -5806 -350 -5802
rect -348 -5806 -346 -5802
rect -342 -5806 -340 -5802
rect -338 -5806 -337 -5802
rect -215 -5806 -214 -5802
rect -212 -5806 -210 -5802
rect -206 -5806 -204 -5802
rect -202 -5806 -201 -5802
rect -189 -5806 -188 -5802
rect -186 -5806 -184 -5802
rect -180 -5806 -178 -5802
rect -176 -5806 -175 -5802
rect -163 -5806 -162 -5802
rect -160 -5806 -159 -5802
rect -155 -5806 -152 -5802
rect -150 -5806 -144 -5802
rect -142 -5806 -141 -5802
rect -137 -5806 -134 -5802
rect -132 -5806 -131 -5802
rect -119 -5806 -118 -5802
rect -116 -5806 -110 -5802
rect -108 -5806 -106 -5802
rect -102 -5806 -100 -5802
rect -98 -5806 -97 -5802
rect -85 -5806 -84 -5802
rect -82 -5806 -80 -5802
rect -76 -5806 -74 -5802
rect -72 -5806 -66 -5802
rect -64 -5806 -62 -5802
rect -58 -5806 -56 -5802
rect -54 -5806 -53 -5802
rect -41 -5806 -40 -5802
rect -38 -5806 -32 -5802
rect -30 -5806 -29 -5802
rect -17 -5806 -16 -5802
rect -14 -5806 -9 -5802
rect -5 -5806 0 -5802
rect 2 -5806 3 -5802
rect 7 -5806 8 -5802
rect 10 -5806 12 -5802
rect 16 -5806 18 -5802
rect 20 -5806 21 -5802
rect 143 -5806 144 -5802
rect 146 -5806 148 -5802
rect 152 -5806 154 -5802
rect 156 -5806 157 -5802
rect 169 -5806 170 -5802
rect 172 -5806 174 -5802
rect 178 -5806 180 -5802
rect 182 -5806 183 -5802
rect 195 -5806 196 -5802
rect 198 -5806 199 -5802
rect 203 -5806 206 -5802
rect 208 -5806 214 -5802
rect 216 -5806 217 -5802
rect 221 -5806 224 -5802
rect 226 -5806 227 -5802
rect 239 -5806 240 -5802
rect 242 -5806 248 -5802
rect 250 -5806 252 -5802
rect 256 -5806 258 -5802
rect 260 -5806 261 -5802
rect 273 -5806 274 -5802
rect 276 -5806 278 -5802
rect 282 -5806 284 -5802
rect 286 -5806 292 -5802
rect 294 -5806 296 -5802
rect 300 -5806 302 -5802
rect 304 -5806 305 -5802
rect 317 -5806 318 -5802
rect 320 -5806 326 -5802
rect 328 -5806 329 -5802
rect 341 -5806 342 -5802
rect 344 -5806 349 -5802
rect 353 -5806 358 -5802
rect 360 -5806 361 -5802
rect 365 -5806 366 -5802
rect 368 -5806 370 -5802
rect 374 -5806 376 -5802
rect 378 -5806 379 -5802
rect 499 -5806 500 -5802
rect 502 -5806 504 -5802
rect 508 -5806 510 -5802
rect 512 -5806 513 -5802
rect 525 -5806 526 -5802
rect 528 -5806 530 -5802
rect 534 -5806 536 -5802
rect 538 -5806 539 -5802
rect 551 -5806 552 -5802
rect 554 -5806 555 -5802
rect 559 -5806 562 -5802
rect 564 -5806 570 -5802
rect 572 -5806 573 -5802
rect 577 -5806 580 -5802
rect 582 -5806 583 -5802
rect 595 -5806 596 -5802
rect 598 -5806 604 -5802
rect 606 -5806 608 -5802
rect 612 -5806 614 -5802
rect 616 -5806 617 -5802
rect 629 -5806 630 -5802
rect 632 -5806 634 -5802
rect 638 -5806 640 -5802
rect 642 -5806 648 -5802
rect 650 -5806 652 -5802
rect 656 -5806 658 -5802
rect 660 -5806 661 -5802
rect 673 -5806 674 -5802
rect 676 -5806 682 -5802
rect 684 -5806 685 -5802
rect 697 -5806 698 -5802
rect 700 -5806 705 -5802
rect 709 -5806 714 -5802
rect 716 -5806 717 -5802
rect 721 -5806 722 -5802
rect 724 -5806 726 -5802
rect 730 -5806 732 -5802
rect 734 -5806 735 -5802
rect 857 -5806 858 -5802
rect 860 -5806 862 -5802
rect 866 -5806 868 -5802
rect 870 -5806 871 -5802
rect 883 -5806 884 -5802
rect 886 -5806 888 -5802
rect 892 -5806 894 -5802
rect 896 -5806 897 -5802
rect 909 -5806 910 -5802
rect 912 -5806 913 -5802
rect 917 -5806 920 -5802
rect 922 -5806 928 -5802
rect 930 -5806 931 -5802
rect 935 -5806 938 -5802
rect 940 -5806 941 -5802
rect 953 -5806 954 -5802
rect 956 -5806 962 -5802
rect 964 -5806 966 -5802
rect 970 -5806 972 -5802
rect 974 -5806 975 -5802
rect 987 -5806 988 -5802
rect 990 -5806 992 -5802
rect 996 -5806 998 -5802
rect 1000 -5806 1006 -5802
rect 1008 -5806 1010 -5802
rect 1014 -5806 1016 -5802
rect 1018 -5806 1019 -5802
rect 1031 -5806 1032 -5802
rect 1034 -5806 1040 -5802
rect 1042 -5806 1043 -5802
rect 1055 -5806 1056 -5802
rect 1058 -5806 1063 -5802
rect 1067 -5806 1072 -5802
rect 1074 -5806 1075 -5802
rect 1079 -5806 1080 -5802
rect 1082 -5806 1084 -5802
rect 1088 -5806 1090 -5802
rect 1092 -5806 1093 -5802
rect 1215 -5806 1216 -5802
rect 1218 -5806 1220 -5802
rect 1224 -5806 1226 -5802
rect 1228 -5806 1229 -5802
rect 1241 -5806 1242 -5802
rect 1244 -5806 1246 -5802
rect 1250 -5806 1252 -5802
rect 1254 -5806 1255 -5802
rect 1267 -5806 1268 -5802
rect 1270 -5806 1271 -5802
rect 1275 -5806 1278 -5802
rect 1280 -5806 1286 -5802
rect 1288 -5806 1289 -5802
rect 1293 -5806 1296 -5802
rect 1298 -5806 1299 -5802
rect 1311 -5806 1312 -5802
rect 1314 -5806 1320 -5802
rect 1322 -5806 1324 -5802
rect 1328 -5806 1330 -5802
rect 1332 -5806 1333 -5802
rect 1345 -5806 1346 -5802
rect 1348 -5806 1350 -5802
rect 1354 -5806 1356 -5802
rect 1358 -5806 1364 -5802
rect 1366 -5806 1368 -5802
rect 1372 -5806 1374 -5802
rect 1376 -5806 1377 -5802
rect 1389 -5806 1390 -5802
rect 1392 -5806 1398 -5802
rect 1400 -5806 1401 -5802
rect 1413 -5806 1414 -5802
rect 1416 -5806 1421 -5802
rect 1425 -5806 1430 -5802
rect 1432 -5806 1433 -5802
rect 1437 -5806 1438 -5802
rect 1440 -5806 1442 -5802
rect 1446 -5806 1448 -5802
rect 1450 -5806 1451 -5802
rect -1230 -5929 -1229 -5925
rect -1227 -5929 -1225 -5925
rect -1221 -5929 -1219 -5925
rect -1217 -5929 -1216 -5925
rect -1204 -5929 -1203 -5925
rect -1201 -5929 -1195 -5925
rect -1193 -5929 -1192 -5925
rect -1180 -5929 -1179 -5925
rect -1177 -5929 -1171 -5925
rect -1169 -5929 -1167 -5925
rect -1163 -5929 -1161 -5925
rect -1159 -5929 -1153 -5925
rect -1151 -5929 -1150 -5925
rect -1138 -5929 -1137 -5925
rect -1135 -5929 -1129 -5925
rect -1127 -5929 -1125 -5925
rect -1121 -5929 -1119 -5925
rect -1117 -5929 -1111 -5925
rect -1109 -5929 -1108 -5925
rect -1096 -5929 -1095 -5925
rect -1093 -5929 -1087 -5925
rect -1085 -5929 -1083 -5925
rect -1079 -5929 -1077 -5925
rect -1075 -5929 -1069 -5925
rect -1067 -5929 -1066 -5925
rect -1054 -5929 -1053 -5925
rect -1051 -5929 -1045 -5925
rect -1043 -5929 -1042 -5925
rect -931 -5929 -930 -5925
rect -928 -5929 -926 -5925
rect -922 -5929 -920 -5925
rect -918 -5929 -917 -5925
rect -905 -5929 -904 -5925
rect -902 -5929 -896 -5925
rect -894 -5929 -893 -5925
rect -881 -5929 -880 -5925
rect -878 -5929 -872 -5925
rect -870 -5929 -868 -5925
rect -864 -5929 -862 -5925
rect -860 -5929 -854 -5925
rect -852 -5929 -851 -5925
rect -839 -5929 -838 -5925
rect -836 -5929 -830 -5925
rect -828 -5929 -826 -5925
rect -822 -5929 -820 -5925
rect -818 -5929 -812 -5925
rect -810 -5929 -809 -5925
rect -797 -5929 -796 -5925
rect -794 -5929 -788 -5925
rect -786 -5929 -784 -5925
rect -780 -5929 -778 -5925
rect -776 -5929 -770 -5925
rect -768 -5929 -767 -5925
rect -755 -5929 -754 -5925
rect -752 -5929 -746 -5925
rect -744 -5929 -743 -5925
rect -573 -5929 -572 -5925
rect -570 -5929 -568 -5925
rect -564 -5929 -562 -5925
rect -560 -5929 -559 -5925
rect -547 -5929 -546 -5925
rect -544 -5929 -538 -5925
rect -536 -5929 -535 -5925
rect -523 -5929 -522 -5925
rect -520 -5929 -514 -5925
rect -512 -5929 -510 -5925
rect -506 -5929 -504 -5925
rect -502 -5929 -496 -5925
rect -494 -5929 -493 -5925
rect -481 -5929 -480 -5925
rect -478 -5929 -472 -5925
rect -470 -5929 -468 -5925
rect -464 -5929 -462 -5925
rect -460 -5929 -454 -5925
rect -452 -5929 -451 -5925
rect -439 -5929 -438 -5925
rect -436 -5929 -430 -5925
rect -428 -5929 -426 -5925
rect -422 -5929 -420 -5925
rect -418 -5929 -412 -5925
rect -410 -5929 -409 -5925
rect -397 -5929 -396 -5925
rect -394 -5929 -388 -5925
rect -386 -5929 -385 -5925
rect -215 -5929 -214 -5925
rect -212 -5929 -210 -5925
rect -206 -5929 -204 -5925
rect -202 -5929 -201 -5925
rect -189 -5929 -188 -5925
rect -186 -5929 -180 -5925
rect -178 -5929 -177 -5925
rect -165 -5929 -164 -5925
rect -162 -5929 -156 -5925
rect -154 -5929 -152 -5925
rect -148 -5929 -146 -5925
rect -144 -5929 -138 -5925
rect -136 -5929 -135 -5925
rect -123 -5929 -122 -5925
rect -120 -5929 -114 -5925
rect -112 -5929 -110 -5925
rect -106 -5929 -104 -5925
rect -102 -5929 -96 -5925
rect -94 -5929 -93 -5925
rect -81 -5929 -80 -5925
rect -78 -5929 -72 -5925
rect -70 -5929 -68 -5925
rect -64 -5929 -62 -5925
rect -60 -5929 -54 -5925
rect -52 -5929 -51 -5925
rect -39 -5929 -38 -5925
rect -36 -5929 -30 -5925
rect -28 -5929 -27 -5925
rect 143 -5929 144 -5925
rect 146 -5929 148 -5925
rect 152 -5929 154 -5925
rect 156 -5929 157 -5925
rect 169 -5929 170 -5925
rect 172 -5929 178 -5925
rect 180 -5929 181 -5925
rect 193 -5929 194 -5925
rect 196 -5929 202 -5925
rect 204 -5929 206 -5925
rect 210 -5929 212 -5925
rect 214 -5929 220 -5925
rect 222 -5929 223 -5925
rect 235 -5929 236 -5925
rect 238 -5929 244 -5925
rect 246 -5929 248 -5925
rect 252 -5929 254 -5925
rect 256 -5929 262 -5925
rect 264 -5929 265 -5925
rect 277 -5929 278 -5925
rect 280 -5929 286 -5925
rect 288 -5929 290 -5925
rect 294 -5929 296 -5925
rect 298 -5929 304 -5925
rect 306 -5929 307 -5925
rect 319 -5929 320 -5925
rect 322 -5929 328 -5925
rect 330 -5929 331 -5925
rect 499 -5929 500 -5925
rect 502 -5929 504 -5925
rect 508 -5929 510 -5925
rect 512 -5929 513 -5925
rect 525 -5929 526 -5925
rect 528 -5929 534 -5925
rect 536 -5929 537 -5925
rect 549 -5929 550 -5925
rect 552 -5929 558 -5925
rect 560 -5929 562 -5925
rect 566 -5929 568 -5925
rect 570 -5929 576 -5925
rect 578 -5929 579 -5925
rect 591 -5929 592 -5925
rect 594 -5929 600 -5925
rect 602 -5929 604 -5925
rect 608 -5929 610 -5925
rect 612 -5929 618 -5925
rect 620 -5929 621 -5925
rect 633 -5929 634 -5925
rect 636 -5929 642 -5925
rect 644 -5929 646 -5925
rect 650 -5929 652 -5925
rect 654 -5929 660 -5925
rect 662 -5929 663 -5925
rect 675 -5929 676 -5925
rect 678 -5929 684 -5925
rect 686 -5929 687 -5925
rect 857 -5929 858 -5925
rect 860 -5929 862 -5925
rect 866 -5929 868 -5925
rect 870 -5929 871 -5925
rect 883 -5929 884 -5925
rect 886 -5929 892 -5925
rect 894 -5929 895 -5925
rect 907 -5929 908 -5925
rect 910 -5929 916 -5925
rect 918 -5929 920 -5925
rect 924 -5929 926 -5925
rect 928 -5929 934 -5925
rect 936 -5929 937 -5925
rect 949 -5929 950 -5925
rect 952 -5929 958 -5925
rect 960 -5929 962 -5925
rect 966 -5929 968 -5925
rect 970 -5929 976 -5925
rect 978 -5929 979 -5925
rect 991 -5929 992 -5925
rect 994 -5929 1000 -5925
rect 1002 -5929 1004 -5925
rect 1008 -5929 1010 -5925
rect 1012 -5929 1018 -5925
rect 1020 -5929 1021 -5925
rect 1033 -5929 1034 -5925
rect 1036 -5929 1042 -5925
rect 1044 -5929 1045 -5925
rect 1215 -5929 1216 -5925
rect 1218 -5929 1220 -5925
rect 1224 -5929 1226 -5925
rect 1228 -5929 1229 -5925
rect 1241 -5929 1242 -5925
rect 1244 -5929 1250 -5925
rect 1252 -5929 1253 -5925
rect 1265 -5929 1266 -5925
rect 1268 -5929 1274 -5925
rect 1276 -5929 1278 -5925
rect 1282 -5929 1284 -5925
rect 1286 -5929 1292 -5925
rect 1294 -5929 1295 -5925
rect 1307 -5929 1308 -5925
rect 1310 -5929 1316 -5925
rect 1318 -5929 1320 -5925
rect 1324 -5929 1326 -5925
rect 1328 -5929 1334 -5925
rect 1336 -5929 1337 -5925
rect 1349 -5929 1350 -5925
rect 1352 -5929 1358 -5925
rect 1360 -5929 1362 -5925
rect 1366 -5929 1368 -5925
rect 1370 -5929 1376 -5925
rect 1378 -5929 1379 -5925
rect 1391 -5929 1392 -5925
rect 1394 -5929 1400 -5925
rect 1402 -5929 1403 -5925
rect 1559 -5929 1560 -5925
rect 1562 -5929 1564 -5925
rect 1568 -5929 1570 -5925
rect 1572 -5929 1573 -5925
rect 1585 -5929 1586 -5925
rect 1588 -5929 1594 -5925
rect 1596 -5929 1597 -5925
rect 1609 -5929 1610 -5925
rect 1612 -5929 1618 -5925
rect 1620 -5929 1622 -5925
rect 1626 -5929 1628 -5925
rect 1630 -5929 1636 -5925
rect 1638 -5929 1639 -5925
rect 1651 -5929 1652 -5925
rect 1654 -5929 1660 -5925
rect 1662 -5929 1664 -5925
rect 1668 -5929 1670 -5925
rect 1672 -5929 1678 -5925
rect 1680 -5929 1681 -5925
rect 1693 -5929 1694 -5925
rect 1696 -5929 1702 -5925
rect 1704 -5929 1706 -5925
rect 1710 -5929 1712 -5925
rect 1714 -5929 1720 -5925
rect 1722 -5929 1723 -5925
rect 1735 -5929 1736 -5925
rect 1738 -5929 1744 -5925
rect 1746 -5929 1747 -5925
<< pdiffusion >>
rect -1303 -796 -1302 -788
rect -1300 -796 -1299 -788
rect -1295 -796 -1294 -788
rect -1292 -796 -1290 -788
rect -1286 -796 -1284 -788
rect -1282 -796 -1281 -788
rect -932 -796 -931 -788
rect -929 -796 -928 -788
rect -924 -796 -923 -788
rect -921 -796 -919 -788
rect -915 -796 -913 -788
rect -911 -796 -910 -788
rect -573 -796 -572 -788
rect -570 -796 -569 -788
rect -565 -796 -564 -788
rect -562 -796 -560 -788
rect -556 -796 -554 -788
rect -552 -796 -551 -788
rect -215 -796 -214 -788
rect -212 -796 -211 -788
rect -207 -796 -206 -788
rect -204 -796 -202 -788
rect -198 -796 -196 -788
rect -194 -796 -193 -788
rect 142 -796 143 -788
rect 145 -796 146 -788
rect 150 -796 151 -788
rect 153 -796 155 -788
rect 159 -796 161 -788
rect 163 -796 164 -788
rect 499 -796 500 -788
rect 502 -796 503 -788
rect 507 -796 508 -788
rect 510 -796 512 -788
rect 516 -796 518 -788
rect 520 -796 521 -788
rect 857 -796 858 -788
rect 860 -796 861 -788
rect 865 -796 866 -788
rect 868 -796 870 -788
rect 874 -796 876 -788
rect 878 -796 879 -788
rect 1215 -796 1216 -788
rect 1218 -796 1219 -788
rect 1223 -796 1224 -788
rect 1226 -796 1228 -788
rect 1232 -796 1234 -788
rect 1236 -796 1237 -788
rect -1226 -1030 -1225 -1022
rect -1223 -1030 -1221 -1022
rect -1217 -1030 -1215 -1022
rect -1213 -1030 -1212 -1022
rect -1200 -1030 -1199 -1022
rect -1197 -1030 -1196 -1022
rect -1192 -1030 -1191 -1022
rect -1189 -1030 -1184 -1022
rect -1180 -1030 -1175 -1022
rect -1173 -1030 -1172 -1022
rect -1168 -1030 -1167 -1022
rect -1165 -1030 -1163 -1022
rect -1159 -1030 -1157 -1022
rect -1155 -1030 -1154 -1022
rect -1150 -1030 -1149 -1022
rect -1147 -1030 -1142 -1022
rect -1138 -1030 -1133 -1022
rect -1131 -1030 -1130 -1022
rect -1126 -1030 -1125 -1022
rect -1123 -1030 -1121 -1022
rect -1117 -1030 -1115 -1022
rect -1113 -1030 -1112 -1022
rect -1108 -1030 -1107 -1022
rect -1105 -1030 -1100 -1022
rect -1096 -1030 -1091 -1022
rect -1089 -1030 -1088 -1022
rect -1084 -1030 -1083 -1022
rect -1081 -1030 -1079 -1022
rect -1075 -1030 -1073 -1022
rect -1071 -1030 -1070 -1022
rect -1066 -1030 -1065 -1022
rect -1063 -1030 -1058 -1022
rect -1054 -1030 -1049 -1022
rect -1047 -1030 -1046 -1022
rect -1042 -1030 -1041 -1022
rect -1039 -1030 -1038 -1022
rect -931 -1030 -930 -1022
rect -928 -1030 -926 -1022
rect -922 -1030 -920 -1022
rect -918 -1030 -917 -1022
rect -905 -1030 -904 -1022
rect -902 -1030 -901 -1022
rect -897 -1030 -896 -1022
rect -894 -1030 -889 -1022
rect -885 -1030 -880 -1022
rect -878 -1030 -877 -1022
rect -873 -1030 -872 -1022
rect -870 -1030 -868 -1022
rect -864 -1030 -862 -1022
rect -860 -1030 -859 -1022
rect -855 -1030 -854 -1022
rect -852 -1030 -847 -1022
rect -843 -1030 -838 -1022
rect -836 -1030 -835 -1022
rect -831 -1030 -830 -1022
rect -828 -1030 -826 -1022
rect -822 -1030 -820 -1022
rect -818 -1030 -817 -1022
rect -813 -1030 -812 -1022
rect -810 -1030 -805 -1022
rect -801 -1030 -796 -1022
rect -794 -1030 -793 -1022
rect -789 -1030 -788 -1022
rect -786 -1030 -784 -1022
rect -780 -1030 -778 -1022
rect -776 -1030 -775 -1022
rect -771 -1030 -770 -1022
rect -768 -1030 -763 -1022
rect -759 -1030 -754 -1022
rect -752 -1030 -751 -1022
rect -747 -1030 -746 -1022
rect -744 -1030 -743 -1022
rect -573 -1030 -572 -1022
rect -570 -1030 -568 -1022
rect -564 -1030 -562 -1022
rect -560 -1030 -559 -1022
rect -547 -1030 -546 -1022
rect -544 -1030 -543 -1022
rect -539 -1030 -538 -1022
rect -536 -1030 -531 -1022
rect -527 -1030 -522 -1022
rect -520 -1030 -519 -1022
rect -515 -1030 -514 -1022
rect -512 -1030 -510 -1022
rect -506 -1030 -504 -1022
rect -502 -1030 -501 -1022
rect -497 -1030 -496 -1022
rect -494 -1030 -489 -1022
rect -485 -1030 -480 -1022
rect -478 -1030 -477 -1022
rect -473 -1030 -472 -1022
rect -470 -1030 -468 -1022
rect -464 -1030 -462 -1022
rect -460 -1030 -459 -1022
rect -455 -1030 -454 -1022
rect -452 -1030 -447 -1022
rect -443 -1030 -438 -1022
rect -436 -1030 -435 -1022
rect -431 -1030 -430 -1022
rect -428 -1030 -426 -1022
rect -422 -1030 -420 -1022
rect -418 -1030 -417 -1022
rect -413 -1030 -412 -1022
rect -410 -1030 -405 -1022
rect -401 -1030 -396 -1022
rect -394 -1030 -393 -1022
rect -389 -1030 -388 -1022
rect -386 -1030 -385 -1022
rect -215 -1030 -214 -1022
rect -212 -1030 -210 -1022
rect -206 -1030 -204 -1022
rect -202 -1030 -201 -1022
rect -189 -1030 -188 -1022
rect -186 -1030 -185 -1022
rect -181 -1030 -180 -1022
rect -178 -1030 -173 -1022
rect -169 -1030 -164 -1022
rect -162 -1030 -161 -1022
rect -157 -1030 -156 -1022
rect -154 -1030 -152 -1022
rect -148 -1030 -146 -1022
rect -144 -1030 -143 -1022
rect -139 -1030 -138 -1022
rect -136 -1030 -131 -1022
rect -127 -1030 -122 -1022
rect -120 -1030 -119 -1022
rect -115 -1030 -114 -1022
rect -112 -1030 -110 -1022
rect -106 -1030 -104 -1022
rect -102 -1030 -101 -1022
rect -97 -1030 -96 -1022
rect -94 -1030 -89 -1022
rect -85 -1030 -80 -1022
rect -78 -1030 -77 -1022
rect -73 -1030 -72 -1022
rect -70 -1030 -68 -1022
rect -64 -1030 -62 -1022
rect -60 -1030 -59 -1022
rect -55 -1030 -54 -1022
rect -52 -1030 -47 -1022
rect -43 -1030 -38 -1022
rect -36 -1030 -35 -1022
rect -31 -1030 -30 -1022
rect -28 -1030 -27 -1022
rect 143 -1030 144 -1022
rect 146 -1030 148 -1022
rect 152 -1030 154 -1022
rect 156 -1030 157 -1022
rect 169 -1030 170 -1022
rect 172 -1030 173 -1022
rect 177 -1030 178 -1022
rect 180 -1030 185 -1022
rect 189 -1030 194 -1022
rect 196 -1030 197 -1022
rect 201 -1030 202 -1022
rect 204 -1030 206 -1022
rect 210 -1030 212 -1022
rect 214 -1030 215 -1022
rect 219 -1030 220 -1022
rect 222 -1030 227 -1022
rect 231 -1030 236 -1022
rect 238 -1030 239 -1022
rect 243 -1030 244 -1022
rect 246 -1030 248 -1022
rect 252 -1030 254 -1022
rect 256 -1030 257 -1022
rect 261 -1030 262 -1022
rect 264 -1030 269 -1022
rect 273 -1030 278 -1022
rect 280 -1030 281 -1022
rect 285 -1030 286 -1022
rect 288 -1030 290 -1022
rect 294 -1030 296 -1022
rect 298 -1030 299 -1022
rect 303 -1030 304 -1022
rect 306 -1030 311 -1022
rect 315 -1030 320 -1022
rect 322 -1030 323 -1022
rect 327 -1030 328 -1022
rect 330 -1030 331 -1022
rect 499 -1030 500 -1022
rect 502 -1030 504 -1022
rect 508 -1030 510 -1022
rect 512 -1030 513 -1022
rect 525 -1030 526 -1022
rect 528 -1030 529 -1022
rect 533 -1030 534 -1022
rect 536 -1030 541 -1022
rect 545 -1030 550 -1022
rect 552 -1030 553 -1022
rect 557 -1030 558 -1022
rect 560 -1030 562 -1022
rect 566 -1030 568 -1022
rect 570 -1030 571 -1022
rect 575 -1030 576 -1022
rect 578 -1030 583 -1022
rect 587 -1030 592 -1022
rect 594 -1030 595 -1022
rect 599 -1030 600 -1022
rect 602 -1030 604 -1022
rect 608 -1030 610 -1022
rect 612 -1030 613 -1022
rect 617 -1030 618 -1022
rect 620 -1030 625 -1022
rect 629 -1030 634 -1022
rect 636 -1030 637 -1022
rect 641 -1030 642 -1022
rect 644 -1030 646 -1022
rect 650 -1030 652 -1022
rect 654 -1030 655 -1022
rect 659 -1030 660 -1022
rect 662 -1030 667 -1022
rect 671 -1030 676 -1022
rect 678 -1030 679 -1022
rect 683 -1030 684 -1022
rect 686 -1030 687 -1022
rect 857 -1030 858 -1022
rect 860 -1030 862 -1022
rect 866 -1030 868 -1022
rect 870 -1030 871 -1022
rect 883 -1030 884 -1022
rect 886 -1030 887 -1022
rect 891 -1030 892 -1022
rect 894 -1030 899 -1022
rect 903 -1030 908 -1022
rect 910 -1030 911 -1022
rect 915 -1030 916 -1022
rect 918 -1030 920 -1022
rect 924 -1030 926 -1022
rect 928 -1030 929 -1022
rect 933 -1030 934 -1022
rect 936 -1030 941 -1022
rect 945 -1030 950 -1022
rect 952 -1030 953 -1022
rect 957 -1030 958 -1022
rect 960 -1030 962 -1022
rect 966 -1030 968 -1022
rect 970 -1030 971 -1022
rect 975 -1030 976 -1022
rect 978 -1030 983 -1022
rect 987 -1030 992 -1022
rect 994 -1030 995 -1022
rect 999 -1030 1000 -1022
rect 1002 -1030 1004 -1022
rect 1008 -1030 1010 -1022
rect 1012 -1030 1013 -1022
rect 1017 -1030 1018 -1022
rect 1020 -1030 1025 -1022
rect 1029 -1030 1034 -1022
rect 1036 -1030 1037 -1022
rect 1041 -1030 1042 -1022
rect 1044 -1030 1045 -1022
rect -1305 -1146 -1304 -1138
rect -1302 -1146 -1301 -1138
rect -1297 -1146 -1296 -1138
rect -1294 -1146 -1292 -1138
rect -1288 -1146 -1286 -1138
rect -1284 -1146 -1283 -1138
rect -931 -1146 -930 -1138
rect -928 -1146 -927 -1138
rect -923 -1146 -922 -1138
rect -920 -1146 -918 -1138
rect -914 -1146 -912 -1138
rect -910 -1146 -909 -1138
rect -573 -1146 -572 -1138
rect -570 -1146 -569 -1138
rect -565 -1146 -564 -1138
rect -562 -1146 -560 -1138
rect -556 -1146 -554 -1138
rect -552 -1146 -551 -1138
rect -215 -1146 -214 -1138
rect -212 -1146 -211 -1138
rect -207 -1146 -206 -1138
rect -204 -1146 -202 -1138
rect -198 -1146 -196 -1138
rect -194 -1146 -193 -1138
rect 143 -1146 144 -1138
rect 146 -1146 147 -1138
rect 151 -1146 152 -1138
rect 154 -1146 156 -1138
rect 160 -1146 162 -1138
rect 164 -1146 165 -1138
rect 499 -1146 500 -1138
rect 502 -1146 503 -1138
rect 507 -1146 508 -1138
rect 510 -1146 512 -1138
rect 516 -1146 518 -1138
rect 520 -1146 521 -1138
rect 857 -1146 858 -1138
rect 860 -1146 861 -1138
rect 865 -1146 866 -1138
rect 868 -1146 870 -1138
rect 874 -1146 876 -1138
rect 878 -1146 879 -1138
rect 1215 -1146 1216 -1138
rect 1218 -1146 1219 -1138
rect 1223 -1146 1224 -1138
rect 1226 -1146 1228 -1138
rect 1232 -1146 1234 -1138
rect 1236 -1146 1237 -1138
rect -1226 -1310 -1225 -1302
rect -1223 -1310 -1221 -1302
rect -1217 -1310 -1215 -1302
rect -1213 -1310 -1212 -1302
rect -1200 -1310 -1199 -1302
rect -1197 -1310 -1189 -1302
rect -1187 -1310 -1186 -1302
rect -1182 -1310 -1181 -1302
rect -1179 -1310 -1171 -1302
rect -1169 -1310 -1164 -1302
rect -1160 -1310 -1155 -1302
rect -1153 -1310 -1152 -1302
rect -1148 -1310 -1147 -1302
rect -1145 -1310 -1143 -1302
rect -1139 -1310 -1137 -1302
rect -1135 -1310 -1134 -1302
rect -931 -1310 -930 -1302
rect -928 -1310 -926 -1302
rect -922 -1310 -920 -1302
rect -918 -1310 -917 -1302
rect -905 -1310 -904 -1302
rect -902 -1310 -900 -1302
rect -896 -1310 -894 -1302
rect -892 -1310 -891 -1302
rect -879 -1310 -878 -1302
rect -876 -1310 -868 -1302
rect -866 -1310 -865 -1302
rect -861 -1310 -860 -1302
rect -858 -1310 -850 -1302
rect -848 -1310 -843 -1302
rect -839 -1310 -834 -1302
rect -832 -1310 -831 -1302
rect -827 -1310 -826 -1302
rect -824 -1310 -822 -1302
rect -818 -1310 -816 -1302
rect -814 -1310 -813 -1302
rect -801 -1310 -800 -1302
rect -798 -1310 -790 -1302
rect -788 -1310 -787 -1302
rect -783 -1310 -782 -1302
rect -780 -1310 -772 -1302
rect -770 -1310 -765 -1302
rect -761 -1310 -756 -1302
rect -754 -1310 -753 -1302
rect -749 -1310 -748 -1302
rect -746 -1310 -741 -1302
rect -737 -1310 -732 -1302
rect -730 -1310 -729 -1302
rect -717 -1310 -716 -1302
rect -714 -1310 -708 -1302
rect -706 -1310 -704 -1302
rect -700 -1310 -698 -1302
rect -696 -1310 -695 -1302
rect -573 -1310 -572 -1302
rect -570 -1310 -568 -1302
rect -564 -1310 -562 -1302
rect -560 -1310 -559 -1302
rect -547 -1310 -546 -1302
rect -544 -1310 -542 -1302
rect -538 -1310 -536 -1302
rect -534 -1310 -533 -1302
rect -521 -1310 -520 -1302
rect -518 -1310 -510 -1302
rect -508 -1310 -507 -1302
rect -503 -1310 -502 -1302
rect -500 -1310 -492 -1302
rect -490 -1310 -485 -1302
rect -481 -1310 -476 -1302
rect -474 -1310 -473 -1302
rect -469 -1310 -468 -1302
rect -466 -1310 -464 -1302
rect -460 -1310 -458 -1302
rect -456 -1310 -455 -1302
rect -443 -1310 -442 -1302
rect -440 -1310 -432 -1302
rect -430 -1310 -429 -1302
rect -425 -1310 -424 -1302
rect -422 -1310 -414 -1302
rect -412 -1310 -407 -1302
rect -403 -1310 -398 -1302
rect -396 -1310 -395 -1302
rect -391 -1310 -390 -1302
rect -388 -1310 -383 -1302
rect -379 -1310 -374 -1302
rect -372 -1310 -371 -1302
rect -359 -1310 -358 -1302
rect -356 -1310 -350 -1302
rect -348 -1310 -346 -1302
rect -342 -1310 -340 -1302
rect -338 -1310 -337 -1302
rect -215 -1310 -214 -1302
rect -212 -1310 -210 -1302
rect -206 -1310 -204 -1302
rect -202 -1310 -201 -1302
rect -189 -1310 -188 -1302
rect -186 -1310 -184 -1302
rect -180 -1310 -178 -1302
rect -176 -1310 -175 -1302
rect -163 -1310 -162 -1302
rect -160 -1310 -152 -1302
rect -150 -1310 -149 -1302
rect -145 -1310 -144 -1302
rect -142 -1310 -134 -1302
rect -132 -1310 -127 -1302
rect -123 -1310 -118 -1302
rect -116 -1310 -115 -1302
rect -111 -1310 -110 -1302
rect -108 -1310 -106 -1302
rect -102 -1310 -100 -1302
rect -98 -1310 -97 -1302
rect -85 -1310 -84 -1302
rect -82 -1310 -74 -1302
rect -72 -1310 -71 -1302
rect -67 -1310 -66 -1302
rect -64 -1310 -56 -1302
rect -54 -1310 -49 -1302
rect -45 -1310 -40 -1302
rect -38 -1310 -37 -1302
rect -33 -1310 -32 -1302
rect -30 -1310 -25 -1302
rect -21 -1310 -16 -1302
rect -14 -1310 -13 -1302
rect -1 -1310 0 -1302
rect 2 -1310 8 -1302
rect 10 -1310 12 -1302
rect 16 -1310 18 -1302
rect 20 -1310 21 -1302
rect 143 -1310 144 -1302
rect 146 -1310 148 -1302
rect 152 -1310 154 -1302
rect 156 -1310 157 -1302
rect 169 -1310 170 -1302
rect 172 -1310 174 -1302
rect 178 -1310 180 -1302
rect 182 -1310 183 -1302
rect 195 -1310 196 -1302
rect 198 -1310 206 -1302
rect 208 -1310 209 -1302
rect 213 -1310 214 -1302
rect 216 -1310 224 -1302
rect 226 -1310 231 -1302
rect 235 -1310 240 -1302
rect 242 -1310 243 -1302
rect 247 -1310 248 -1302
rect 250 -1310 252 -1302
rect 256 -1310 258 -1302
rect 260 -1310 261 -1302
rect 273 -1310 274 -1302
rect 276 -1310 284 -1302
rect 286 -1310 287 -1302
rect 291 -1310 292 -1302
rect 294 -1310 302 -1302
rect 304 -1310 309 -1302
rect 313 -1310 318 -1302
rect 320 -1310 321 -1302
rect 325 -1310 326 -1302
rect 328 -1310 333 -1302
rect 337 -1310 342 -1302
rect 344 -1310 345 -1302
rect 357 -1310 358 -1302
rect 360 -1310 366 -1302
rect 368 -1310 370 -1302
rect 374 -1310 376 -1302
rect 378 -1310 379 -1302
rect 499 -1310 500 -1302
rect 502 -1310 504 -1302
rect 508 -1310 510 -1302
rect 512 -1310 513 -1302
rect 525 -1310 526 -1302
rect 528 -1310 530 -1302
rect 534 -1310 536 -1302
rect 538 -1310 539 -1302
rect 551 -1310 552 -1302
rect 554 -1310 562 -1302
rect 564 -1310 565 -1302
rect 569 -1310 570 -1302
rect 572 -1310 580 -1302
rect 582 -1310 587 -1302
rect 591 -1310 596 -1302
rect 598 -1310 599 -1302
rect 603 -1310 604 -1302
rect 606 -1310 608 -1302
rect 612 -1310 614 -1302
rect 616 -1310 617 -1302
rect 629 -1310 630 -1302
rect 632 -1310 640 -1302
rect 642 -1310 643 -1302
rect 647 -1310 648 -1302
rect 650 -1310 658 -1302
rect 660 -1310 665 -1302
rect 669 -1310 674 -1302
rect 676 -1310 677 -1302
rect 681 -1310 682 -1302
rect 684 -1310 689 -1302
rect 693 -1310 698 -1302
rect 700 -1310 701 -1302
rect 713 -1310 714 -1302
rect 716 -1310 722 -1302
rect 724 -1310 726 -1302
rect 730 -1310 732 -1302
rect 734 -1310 735 -1302
rect 857 -1310 858 -1302
rect 860 -1310 862 -1302
rect 866 -1310 868 -1302
rect 870 -1310 871 -1302
rect 883 -1310 884 -1302
rect 886 -1310 888 -1302
rect 892 -1310 894 -1302
rect 896 -1310 897 -1302
rect 909 -1310 910 -1302
rect 912 -1310 920 -1302
rect 922 -1310 923 -1302
rect 927 -1310 928 -1302
rect 930 -1310 938 -1302
rect 940 -1310 945 -1302
rect 949 -1310 954 -1302
rect 956 -1310 957 -1302
rect 961 -1310 962 -1302
rect 964 -1310 966 -1302
rect 970 -1310 972 -1302
rect 974 -1310 975 -1302
rect 987 -1310 988 -1302
rect 990 -1310 998 -1302
rect 1000 -1310 1001 -1302
rect 1005 -1310 1006 -1302
rect 1008 -1310 1016 -1302
rect 1018 -1310 1023 -1302
rect 1027 -1310 1032 -1302
rect 1034 -1310 1035 -1302
rect 1039 -1310 1040 -1302
rect 1042 -1310 1047 -1302
rect 1051 -1310 1056 -1302
rect 1058 -1310 1059 -1302
rect 1071 -1310 1072 -1302
rect 1074 -1310 1080 -1302
rect 1082 -1310 1084 -1302
rect 1088 -1310 1090 -1302
rect 1092 -1310 1093 -1302
rect 1215 -1310 1216 -1302
rect 1218 -1310 1220 -1302
rect 1224 -1310 1226 -1302
rect 1228 -1310 1229 -1302
rect 1241 -1310 1242 -1302
rect 1244 -1310 1252 -1302
rect 1254 -1310 1255 -1302
rect 1259 -1310 1260 -1302
rect 1262 -1310 1270 -1302
rect 1272 -1310 1277 -1302
rect 1281 -1310 1286 -1302
rect 1288 -1310 1289 -1302
rect 1293 -1310 1294 -1302
rect 1296 -1310 1298 -1302
rect 1302 -1310 1304 -1302
rect 1306 -1310 1307 -1302
rect -1226 -1433 -1225 -1425
rect -1223 -1433 -1221 -1425
rect -1217 -1433 -1215 -1425
rect -1213 -1433 -1212 -1425
rect -1200 -1433 -1199 -1425
rect -1197 -1433 -1196 -1425
rect -1192 -1433 -1191 -1425
rect -1189 -1433 -1184 -1425
rect -1180 -1433 -1175 -1425
rect -1173 -1433 -1172 -1425
rect -1168 -1433 -1167 -1425
rect -1165 -1433 -1163 -1425
rect -1159 -1433 -1157 -1425
rect -1155 -1433 -1154 -1425
rect -1150 -1433 -1149 -1425
rect -1147 -1433 -1142 -1425
rect -1138 -1433 -1133 -1425
rect -1131 -1433 -1130 -1425
rect -1126 -1433 -1125 -1425
rect -1123 -1433 -1121 -1425
rect -1117 -1433 -1115 -1425
rect -1113 -1433 -1112 -1425
rect -1108 -1433 -1107 -1425
rect -1105 -1433 -1100 -1425
rect -1096 -1433 -1091 -1425
rect -1089 -1433 -1088 -1425
rect -1084 -1433 -1083 -1425
rect -1081 -1433 -1079 -1425
rect -1075 -1433 -1073 -1425
rect -1071 -1433 -1070 -1425
rect -1066 -1433 -1065 -1425
rect -1063 -1433 -1058 -1425
rect -1054 -1433 -1049 -1425
rect -1047 -1433 -1046 -1425
rect -1042 -1433 -1041 -1425
rect -1039 -1433 -1038 -1425
rect -931 -1433 -930 -1425
rect -928 -1433 -926 -1425
rect -922 -1433 -920 -1425
rect -918 -1433 -917 -1425
rect -905 -1433 -904 -1425
rect -902 -1433 -901 -1425
rect -897 -1433 -896 -1425
rect -894 -1433 -889 -1425
rect -885 -1433 -880 -1425
rect -878 -1433 -877 -1425
rect -873 -1433 -872 -1425
rect -870 -1433 -868 -1425
rect -864 -1433 -862 -1425
rect -860 -1433 -859 -1425
rect -855 -1433 -854 -1425
rect -852 -1433 -847 -1425
rect -843 -1433 -838 -1425
rect -836 -1433 -835 -1425
rect -831 -1433 -830 -1425
rect -828 -1433 -826 -1425
rect -822 -1433 -820 -1425
rect -818 -1433 -817 -1425
rect -813 -1433 -812 -1425
rect -810 -1433 -805 -1425
rect -801 -1433 -796 -1425
rect -794 -1433 -793 -1425
rect -789 -1433 -788 -1425
rect -786 -1433 -784 -1425
rect -780 -1433 -778 -1425
rect -776 -1433 -775 -1425
rect -771 -1433 -770 -1425
rect -768 -1433 -763 -1425
rect -759 -1433 -754 -1425
rect -752 -1433 -751 -1425
rect -747 -1433 -746 -1425
rect -744 -1433 -743 -1425
rect -573 -1433 -572 -1425
rect -570 -1433 -568 -1425
rect -564 -1433 -562 -1425
rect -560 -1433 -559 -1425
rect -547 -1433 -546 -1425
rect -544 -1433 -543 -1425
rect -539 -1433 -538 -1425
rect -536 -1433 -531 -1425
rect -527 -1433 -522 -1425
rect -520 -1433 -519 -1425
rect -515 -1433 -514 -1425
rect -512 -1433 -510 -1425
rect -506 -1433 -504 -1425
rect -502 -1433 -501 -1425
rect -497 -1433 -496 -1425
rect -494 -1433 -489 -1425
rect -485 -1433 -480 -1425
rect -478 -1433 -477 -1425
rect -473 -1433 -472 -1425
rect -470 -1433 -468 -1425
rect -464 -1433 -462 -1425
rect -460 -1433 -459 -1425
rect -455 -1433 -454 -1425
rect -452 -1433 -447 -1425
rect -443 -1433 -438 -1425
rect -436 -1433 -435 -1425
rect -431 -1433 -430 -1425
rect -428 -1433 -426 -1425
rect -422 -1433 -420 -1425
rect -418 -1433 -417 -1425
rect -413 -1433 -412 -1425
rect -410 -1433 -405 -1425
rect -401 -1433 -396 -1425
rect -394 -1433 -393 -1425
rect -389 -1433 -388 -1425
rect -386 -1433 -385 -1425
rect -215 -1433 -214 -1425
rect -212 -1433 -210 -1425
rect -206 -1433 -204 -1425
rect -202 -1433 -201 -1425
rect -189 -1433 -188 -1425
rect -186 -1433 -185 -1425
rect -181 -1433 -180 -1425
rect -178 -1433 -173 -1425
rect -169 -1433 -164 -1425
rect -162 -1433 -161 -1425
rect -157 -1433 -156 -1425
rect -154 -1433 -152 -1425
rect -148 -1433 -146 -1425
rect -144 -1433 -143 -1425
rect -139 -1433 -138 -1425
rect -136 -1433 -131 -1425
rect -127 -1433 -122 -1425
rect -120 -1433 -119 -1425
rect -115 -1433 -114 -1425
rect -112 -1433 -110 -1425
rect -106 -1433 -104 -1425
rect -102 -1433 -101 -1425
rect -97 -1433 -96 -1425
rect -94 -1433 -89 -1425
rect -85 -1433 -80 -1425
rect -78 -1433 -77 -1425
rect -73 -1433 -72 -1425
rect -70 -1433 -68 -1425
rect -64 -1433 -62 -1425
rect -60 -1433 -59 -1425
rect -55 -1433 -54 -1425
rect -52 -1433 -47 -1425
rect -43 -1433 -38 -1425
rect -36 -1433 -35 -1425
rect -31 -1433 -30 -1425
rect -28 -1433 -27 -1425
rect 143 -1433 144 -1425
rect 146 -1433 148 -1425
rect 152 -1433 154 -1425
rect 156 -1433 157 -1425
rect 169 -1433 170 -1425
rect 172 -1433 173 -1425
rect 177 -1433 178 -1425
rect 180 -1433 185 -1425
rect 189 -1433 194 -1425
rect 196 -1433 197 -1425
rect 201 -1433 202 -1425
rect 204 -1433 206 -1425
rect 210 -1433 212 -1425
rect 214 -1433 215 -1425
rect 219 -1433 220 -1425
rect 222 -1433 227 -1425
rect 231 -1433 236 -1425
rect 238 -1433 239 -1425
rect 243 -1433 244 -1425
rect 246 -1433 248 -1425
rect 252 -1433 254 -1425
rect 256 -1433 257 -1425
rect 261 -1433 262 -1425
rect 264 -1433 269 -1425
rect 273 -1433 278 -1425
rect 280 -1433 281 -1425
rect 285 -1433 286 -1425
rect 288 -1433 290 -1425
rect 294 -1433 296 -1425
rect 298 -1433 299 -1425
rect 303 -1433 304 -1425
rect 306 -1433 311 -1425
rect 315 -1433 320 -1425
rect 322 -1433 323 -1425
rect 327 -1433 328 -1425
rect 330 -1433 331 -1425
rect 499 -1433 500 -1425
rect 502 -1433 504 -1425
rect 508 -1433 510 -1425
rect 512 -1433 513 -1425
rect 525 -1433 526 -1425
rect 528 -1433 529 -1425
rect 533 -1433 534 -1425
rect 536 -1433 541 -1425
rect 545 -1433 550 -1425
rect 552 -1433 553 -1425
rect 557 -1433 558 -1425
rect 560 -1433 562 -1425
rect 566 -1433 568 -1425
rect 570 -1433 571 -1425
rect 575 -1433 576 -1425
rect 578 -1433 583 -1425
rect 587 -1433 592 -1425
rect 594 -1433 595 -1425
rect 599 -1433 600 -1425
rect 602 -1433 604 -1425
rect 608 -1433 610 -1425
rect 612 -1433 613 -1425
rect 617 -1433 618 -1425
rect 620 -1433 625 -1425
rect 629 -1433 634 -1425
rect 636 -1433 637 -1425
rect 641 -1433 642 -1425
rect 644 -1433 646 -1425
rect 650 -1433 652 -1425
rect 654 -1433 655 -1425
rect 659 -1433 660 -1425
rect 662 -1433 667 -1425
rect 671 -1433 676 -1425
rect 678 -1433 679 -1425
rect 683 -1433 684 -1425
rect 686 -1433 687 -1425
rect 857 -1433 858 -1425
rect 860 -1433 862 -1425
rect 866 -1433 868 -1425
rect 870 -1433 871 -1425
rect 883 -1433 884 -1425
rect 886 -1433 887 -1425
rect 891 -1433 892 -1425
rect 894 -1433 899 -1425
rect 903 -1433 908 -1425
rect 910 -1433 911 -1425
rect 915 -1433 916 -1425
rect 918 -1433 920 -1425
rect 924 -1433 926 -1425
rect 928 -1433 929 -1425
rect 933 -1433 934 -1425
rect 936 -1433 941 -1425
rect 945 -1433 950 -1425
rect 952 -1433 953 -1425
rect 957 -1433 958 -1425
rect 960 -1433 962 -1425
rect 966 -1433 968 -1425
rect 970 -1433 971 -1425
rect 975 -1433 976 -1425
rect 978 -1433 983 -1425
rect 987 -1433 992 -1425
rect 994 -1433 995 -1425
rect 999 -1433 1000 -1425
rect 1002 -1433 1004 -1425
rect 1008 -1433 1010 -1425
rect 1012 -1433 1013 -1425
rect 1017 -1433 1018 -1425
rect 1020 -1433 1025 -1425
rect 1029 -1433 1034 -1425
rect 1036 -1433 1037 -1425
rect 1041 -1433 1042 -1425
rect 1044 -1433 1045 -1425
rect -1226 -1604 -1225 -1596
rect -1223 -1604 -1221 -1596
rect -1217 -1604 -1215 -1596
rect -1213 -1604 -1212 -1596
rect -1200 -1604 -1199 -1596
rect -1197 -1604 -1196 -1596
rect -1192 -1604 -1191 -1596
rect -1189 -1604 -1184 -1596
rect -1180 -1604 -1175 -1596
rect -1173 -1604 -1172 -1596
rect -1168 -1604 -1167 -1596
rect -1165 -1604 -1163 -1596
rect -1159 -1604 -1157 -1596
rect -1155 -1604 -1154 -1596
rect -1150 -1604 -1149 -1596
rect -1147 -1604 -1142 -1596
rect -1138 -1604 -1133 -1596
rect -1131 -1604 -1130 -1596
rect -1126 -1604 -1125 -1596
rect -1123 -1604 -1121 -1596
rect -1117 -1604 -1115 -1596
rect -1113 -1604 -1112 -1596
rect -1108 -1604 -1107 -1596
rect -1105 -1604 -1100 -1596
rect -1096 -1604 -1091 -1596
rect -1089 -1604 -1088 -1596
rect -1084 -1604 -1083 -1596
rect -1081 -1604 -1079 -1596
rect -1075 -1604 -1073 -1596
rect -1071 -1604 -1070 -1596
rect -1066 -1604 -1065 -1596
rect -1063 -1604 -1058 -1596
rect -1054 -1604 -1049 -1596
rect -1047 -1604 -1046 -1596
rect -1042 -1604 -1041 -1596
rect -1039 -1604 -1038 -1596
rect -931 -1604 -930 -1596
rect -928 -1604 -926 -1596
rect -922 -1604 -920 -1596
rect -918 -1604 -917 -1596
rect -905 -1604 -904 -1596
rect -902 -1604 -901 -1596
rect -897 -1604 -896 -1596
rect -894 -1604 -889 -1596
rect -885 -1604 -880 -1596
rect -878 -1604 -877 -1596
rect -873 -1604 -872 -1596
rect -870 -1604 -868 -1596
rect -864 -1604 -862 -1596
rect -860 -1604 -859 -1596
rect -855 -1604 -854 -1596
rect -852 -1604 -847 -1596
rect -843 -1604 -838 -1596
rect -836 -1604 -835 -1596
rect -831 -1604 -830 -1596
rect -828 -1604 -826 -1596
rect -822 -1604 -820 -1596
rect -818 -1604 -817 -1596
rect -813 -1604 -812 -1596
rect -810 -1604 -805 -1596
rect -801 -1604 -796 -1596
rect -794 -1604 -793 -1596
rect -789 -1604 -788 -1596
rect -786 -1604 -784 -1596
rect -780 -1604 -778 -1596
rect -776 -1604 -775 -1596
rect -771 -1604 -770 -1596
rect -768 -1604 -763 -1596
rect -759 -1604 -754 -1596
rect -752 -1604 -751 -1596
rect -747 -1604 -746 -1596
rect -744 -1604 -743 -1596
rect -573 -1604 -572 -1596
rect -570 -1604 -568 -1596
rect -564 -1604 -562 -1596
rect -560 -1604 -559 -1596
rect -547 -1604 -546 -1596
rect -544 -1604 -543 -1596
rect -539 -1604 -538 -1596
rect -536 -1604 -531 -1596
rect -527 -1604 -522 -1596
rect -520 -1604 -519 -1596
rect -515 -1604 -514 -1596
rect -512 -1604 -510 -1596
rect -506 -1604 -504 -1596
rect -502 -1604 -501 -1596
rect -497 -1604 -496 -1596
rect -494 -1604 -489 -1596
rect -485 -1604 -480 -1596
rect -478 -1604 -477 -1596
rect -473 -1604 -472 -1596
rect -470 -1604 -468 -1596
rect -464 -1604 -462 -1596
rect -460 -1604 -459 -1596
rect -455 -1604 -454 -1596
rect -452 -1604 -447 -1596
rect -443 -1604 -438 -1596
rect -436 -1604 -435 -1596
rect -431 -1604 -430 -1596
rect -428 -1604 -426 -1596
rect -422 -1604 -420 -1596
rect -418 -1604 -417 -1596
rect -413 -1604 -412 -1596
rect -410 -1604 -405 -1596
rect -401 -1604 -396 -1596
rect -394 -1604 -393 -1596
rect -389 -1604 -388 -1596
rect -386 -1604 -385 -1596
rect -215 -1604 -214 -1596
rect -212 -1604 -210 -1596
rect -206 -1604 -204 -1596
rect -202 -1604 -201 -1596
rect -189 -1604 -188 -1596
rect -186 -1604 -185 -1596
rect -181 -1604 -180 -1596
rect -178 -1604 -173 -1596
rect -169 -1604 -164 -1596
rect -162 -1604 -161 -1596
rect -157 -1604 -156 -1596
rect -154 -1604 -152 -1596
rect -148 -1604 -146 -1596
rect -144 -1604 -143 -1596
rect -139 -1604 -138 -1596
rect -136 -1604 -131 -1596
rect -127 -1604 -122 -1596
rect -120 -1604 -119 -1596
rect -115 -1604 -114 -1596
rect -112 -1604 -110 -1596
rect -106 -1604 -104 -1596
rect -102 -1604 -101 -1596
rect -97 -1604 -96 -1596
rect -94 -1604 -89 -1596
rect -85 -1604 -80 -1596
rect -78 -1604 -77 -1596
rect -73 -1604 -72 -1596
rect -70 -1604 -68 -1596
rect -64 -1604 -62 -1596
rect -60 -1604 -59 -1596
rect -55 -1604 -54 -1596
rect -52 -1604 -47 -1596
rect -43 -1604 -38 -1596
rect -36 -1604 -35 -1596
rect -31 -1604 -30 -1596
rect -28 -1604 -27 -1596
rect 143 -1604 144 -1596
rect 146 -1604 148 -1596
rect 152 -1604 154 -1596
rect 156 -1604 157 -1596
rect 169 -1604 170 -1596
rect 172 -1604 173 -1596
rect 177 -1604 178 -1596
rect 180 -1604 185 -1596
rect 189 -1604 194 -1596
rect 196 -1604 197 -1596
rect 201 -1604 202 -1596
rect 204 -1604 206 -1596
rect 210 -1604 212 -1596
rect 214 -1604 215 -1596
rect 219 -1604 220 -1596
rect 222 -1604 227 -1596
rect 231 -1604 236 -1596
rect 238 -1604 239 -1596
rect 243 -1604 244 -1596
rect 246 -1604 248 -1596
rect 252 -1604 254 -1596
rect 256 -1604 257 -1596
rect 261 -1604 262 -1596
rect 264 -1604 269 -1596
rect 273 -1604 278 -1596
rect 280 -1604 281 -1596
rect 285 -1604 286 -1596
rect 288 -1604 290 -1596
rect 294 -1604 296 -1596
rect 298 -1604 299 -1596
rect 303 -1604 304 -1596
rect 306 -1604 311 -1596
rect 315 -1604 320 -1596
rect 322 -1604 323 -1596
rect 327 -1604 328 -1596
rect 330 -1604 331 -1596
rect 499 -1604 500 -1596
rect 502 -1604 504 -1596
rect 508 -1604 510 -1596
rect 512 -1604 513 -1596
rect 525 -1604 526 -1596
rect 528 -1604 529 -1596
rect 533 -1604 534 -1596
rect 536 -1604 541 -1596
rect 545 -1604 550 -1596
rect 552 -1604 553 -1596
rect 557 -1604 558 -1596
rect 560 -1604 562 -1596
rect 566 -1604 568 -1596
rect 570 -1604 571 -1596
rect 575 -1604 576 -1596
rect 578 -1604 583 -1596
rect 587 -1604 592 -1596
rect 594 -1604 595 -1596
rect 599 -1604 600 -1596
rect 602 -1604 604 -1596
rect 608 -1604 610 -1596
rect 612 -1604 613 -1596
rect 617 -1604 618 -1596
rect 620 -1604 625 -1596
rect 629 -1604 634 -1596
rect 636 -1604 637 -1596
rect 641 -1604 642 -1596
rect 644 -1604 646 -1596
rect 650 -1604 652 -1596
rect 654 -1604 655 -1596
rect 659 -1604 660 -1596
rect 662 -1604 667 -1596
rect 671 -1604 676 -1596
rect 678 -1604 679 -1596
rect 683 -1604 684 -1596
rect 686 -1604 687 -1596
rect 857 -1604 858 -1596
rect 860 -1604 862 -1596
rect 866 -1604 868 -1596
rect 870 -1604 871 -1596
rect 883 -1604 884 -1596
rect 886 -1604 887 -1596
rect 891 -1604 892 -1596
rect 894 -1604 899 -1596
rect 903 -1604 908 -1596
rect 910 -1604 911 -1596
rect 915 -1604 916 -1596
rect 918 -1604 920 -1596
rect 924 -1604 926 -1596
rect 928 -1604 929 -1596
rect 933 -1604 934 -1596
rect 936 -1604 941 -1596
rect 945 -1604 950 -1596
rect 952 -1604 953 -1596
rect 957 -1604 958 -1596
rect 960 -1604 962 -1596
rect 966 -1604 968 -1596
rect 970 -1604 971 -1596
rect 975 -1604 976 -1596
rect 978 -1604 983 -1596
rect 987 -1604 992 -1596
rect 994 -1604 995 -1596
rect 999 -1604 1000 -1596
rect 1002 -1604 1004 -1596
rect 1008 -1604 1010 -1596
rect 1012 -1604 1013 -1596
rect 1017 -1604 1018 -1596
rect 1020 -1604 1025 -1596
rect 1029 -1604 1034 -1596
rect 1036 -1604 1037 -1596
rect 1041 -1604 1042 -1596
rect 1044 -1604 1045 -1596
rect 1215 -1604 1216 -1596
rect 1218 -1604 1220 -1596
rect 1224 -1604 1226 -1596
rect 1228 -1604 1229 -1596
rect 1241 -1604 1242 -1596
rect 1244 -1604 1245 -1596
rect 1249 -1604 1250 -1596
rect 1252 -1604 1257 -1596
rect 1261 -1604 1266 -1596
rect 1268 -1604 1269 -1596
rect 1273 -1604 1274 -1596
rect 1276 -1604 1278 -1596
rect 1282 -1604 1284 -1596
rect 1286 -1604 1287 -1596
rect 1291 -1604 1292 -1596
rect 1294 -1604 1299 -1596
rect 1303 -1604 1308 -1596
rect 1310 -1604 1311 -1596
rect 1315 -1604 1316 -1596
rect 1318 -1604 1320 -1596
rect 1324 -1604 1326 -1596
rect 1328 -1604 1329 -1596
rect 1333 -1604 1334 -1596
rect 1336 -1604 1341 -1596
rect 1345 -1604 1350 -1596
rect 1352 -1604 1353 -1596
rect 1357 -1604 1358 -1596
rect 1360 -1604 1362 -1596
rect 1366 -1604 1368 -1596
rect 1370 -1604 1371 -1596
rect 1375 -1604 1376 -1596
rect 1378 -1604 1383 -1596
rect 1387 -1604 1392 -1596
rect 1394 -1604 1395 -1596
rect 1399 -1604 1400 -1596
rect 1402 -1604 1403 -1596
rect -1555 -1775 -1554 -1767
rect -1552 -1775 -1550 -1767
rect -1546 -1775 -1544 -1767
rect -1542 -1775 -1541 -1767
rect -1529 -1775 -1528 -1767
rect -1526 -1775 -1525 -1767
rect -1521 -1775 -1520 -1767
rect -1518 -1775 -1513 -1767
rect -1509 -1775 -1504 -1767
rect -1502 -1775 -1501 -1767
rect -1497 -1775 -1496 -1767
rect -1494 -1775 -1492 -1767
rect -1488 -1775 -1486 -1767
rect -1484 -1775 -1483 -1767
rect -1479 -1775 -1478 -1767
rect -1476 -1775 -1471 -1767
rect -1467 -1775 -1462 -1767
rect -1460 -1775 -1459 -1767
rect -1455 -1775 -1454 -1767
rect -1452 -1775 -1450 -1767
rect -1446 -1775 -1444 -1767
rect -1442 -1775 -1441 -1767
rect -1437 -1775 -1436 -1767
rect -1434 -1775 -1429 -1767
rect -1425 -1775 -1420 -1767
rect -1418 -1775 -1417 -1767
rect -1413 -1775 -1412 -1767
rect -1410 -1775 -1408 -1767
rect -1404 -1775 -1402 -1767
rect -1400 -1775 -1399 -1767
rect -1395 -1775 -1394 -1767
rect -1392 -1775 -1387 -1767
rect -1383 -1775 -1378 -1767
rect -1376 -1775 -1375 -1767
rect -1371 -1775 -1370 -1767
rect -1368 -1775 -1367 -1767
rect -1226 -1775 -1225 -1767
rect -1223 -1775 -1221 -1767
rect -1217 -1775 -1215 -1767
rect -1213 -1775 -1212 -1767
rect -1200 -1775 -1199 -1767
rect -1197 -1775 -1196 -1767
rect -1192 -1775 -1191 -1767
rect -1189 -1775 -1184 -1767
rect -1180 -1775 -1175 -1767
rect -1173 -1775 -1172 -1767
rect -1168 -1775 -1167 -1767
rect -1165 -1775 -1163 -1767
rect -1159 -1775 -1157 -1767
rect -1155 -1775 -1154 -1767
rect -1150 -1775 -1149 -1767
rect -1147 -1775 -1142 -1767
rect -1138 -1775 -1133 -1767
rect -1131 -1775 -1130 -1767
rect -1126 -1775 -1125 -1767
rect -1123 -1775 -1121 -1767
rect -1117 -1775 -1115 -1767
rect -1113 -1775 -1112 -1767
rect -1108 -1775 -1107 -1767
rect -1105 -1775 -1100 -1767
rect -1096 -1775 -1091 -1767
rect -1089 -1775 -1088 -1767
rect -1084 -1775 -1083 -1767
rect -1081 -1775 -1079 -1767
rect -1075 -1775 -1073 -1767
rect -1071 -1775 -1070 -1767
rect -1066 -1775 -1065 -1767
rect -1063 -1775 -1058 -1767
rect -1054 -1775 -1049 -1767
rect -1047 -1775 -1046 -1767
rect -1042 -1775 -1041 -1767
rect -1039 -1775 -1038 -1767
rect -931 -1775 -930 -1767
rect -928 -1775 -926 -1767
rect -922 -1775 -920 -1767
rect -918 -1775 -917 -1767
rect -905 -1775 -904 -1767
rect -902 -1775 -901 -1767
rect -897 -1775 -896 -1767
rect -894 -1775 -889 -1767
rect -885 -1775 -880 -1767
rect -878 -1775 -877 -1767
rect -873 -1775 -872 -1767
rect -870 -1775 -868 -1767
rect -864 -1775 -862 -1767
rect -860 -1775 -859 -1767
rect -855 -1775 -854 -1767
rect -852 -1775 -847 -1767
rect -843 -1775 -838 -1767
rect -836 -1775 -835 -1767
rect -831 -1775 -830 -1767
rect -828 -1775 -826 -1767
rect -822 -1775 -820 -1767
rect -818 -1775 -817 -1767
rect -813 -1775 -812 -1767
rect -810 -1775 -805 -1767
rect -801 -1775 -796 -1767
rect -794 -1775 -793 -1767
rect -789 -1775 -788 -1767
rect -786 -1775 -784 -1767
rect -780 -1775 -778 -1767
rect -776 -1775 -775 -1767
rect -771 -1775 -770 -1767
rect -768 -1775 -763 -1767
rect -759 -1775 -754 -1767
rect -752 -1775 -751 -1767
rect -747 -1775 -746 -1767
rect -744 -1775 -743 -1767
rect -573 -1775 -572 -1767
rect -570 -1775 -568 -1767
rect -564 -1775 -562 -1767
rect -560 -1775 -559 -1767
rect -547 -1775 -546 -1767
rect -544 -1775 -543 -1767
rect -539 -1775 -538 -1767
rect -536 -1775 -531 -1767
rect -527 -1775 -522 -1767
rect -520 -1775 -519 -1767
rect -515 -1775 -514 -1767
rect -512 -1775 -510 -1767
rect -506 -1775 -504 -1767
rect -502 -1775 -501 -1767
rect -497 -1775 -496 -1767
rect -494 -1775 -489 -1767
rect -485 -1775 -480 -1767
rect -478 -1775 -477 -1767
rect -473 -1775 -472 -1767
rect -470 -1775 -468 -1767
rect -464 -1775 -462 -1767
rect -460 -1775 -459 -1767
rect -455 -1775 -454 -1767
rect -452 -1775 -447 -1767
rect -443 -1775 -438 -1767
rect -436 -1775 -435 -1767
rect -431 -1775 -430 -1767
rect -428 -1775 -426 -1767
rect -422 -1775 -420 -1767
rect -418 -1775 -417 -1767
rect -413 -1775 -412 -1767
rect -410 -1775 -405 -1767
rect -401 -1775 -396 -1767
rect -394 -1775 -393 -1767
rect -389 -1775 -388 -1767
rect -386 -1775 -385 -1767
rect -215 -1775 -214 -1767
rect -212 -1775 -210 -1767
rect -206 -1775 -204 -1767
rect -202 -1775 -201 -1767
rect -189 -1775 -188 -1767
rect -186 -1775 -185 -1767
rect -181 -1775 -180 -1767
rect -178 -1775 -173 -1767
rect -169 -1775 -164 -1767
rect -162 -1775 -161 -1767
rect -157 -1775 -156 -1767
rect -154 -1775 -152 -1767
rect -148 -1775 -146 -1767
rect -144 -1775 -143 -1767
rect -139 -1775 -138 -1767
rect -136 -1775 -131 -1767
rect -127 -1775 -122 -1767
rect -120 -1775 -119 -1767
rect -115 -1775 -114 -1767
rect -112 -1775 -110 -1767
rect -106 -1775 -104 -1767
rect -102 -1775 -101 -1767
rect -97 -1775 -96 -1767
rect -94 -1775 -89 -1767
rect -85 -1775 -80 -1767
rect -78 -1775 -77 -1767
rect -73 -1775 -72 -1767
rect -70 -1775 -68 -1767
rect -64 -1775 -62 -1767
rect -60 -1775 -59 -1767
rect -55 -1775 -54 -1767
rect -52 -1775 -47 -1767
rect -43 -1775 -38 -1767
rect -36 -1775 -35 -1767
rect -31 -1775 -30 -1767
rect -28 -1775 -27 -1767
rect 143 -1775 144 -1767
rect 146 -1775 148 -1767
rect 152 -1775 154 -1767
rect 156 -1775 157 -1767
rect 169 -1775 170 -1767
rect 172 -1775 173 -1767
rect 177 -1775 178 -1767
rect 180 -1775 185 -1767
rect 189 -1775 194 -1767
rect 196 -1775 197 -1767
rect 201 -1775 202 -1767
rect 204 -1775 206 -1767
rect 210 -1775 212 -1767
rect 214 -1775 215 -1767
rect 219 -1775 220 -1767
rect 222 -1775 227 -1767
rect 231 -1775 236 -1767
rect 238 -1775 239 -1767
rect 243 -1775 244 -1767
rect 246 -1775 248 -1767
rect 252 -1775 254 -1767
rect 256 -1775 257 -1767
rect 261 -1775 262 -1767
rect 264 -1775 269 -1767
rect 273 -1775 278 -1767
rect 280 -1775 281 -1767
rect 285 -1775 286 -1767
rect 288 -1775 290 -1767
rect 294 -1775 296 -1767
rect 298 -1775 299 -1767
rect 303 -1775 304 -1767
rect 306 -1775 311 -1767
rect 315 -1775 320 -1767
rect 322 -1775 323 -1767
rect 327 -1775 328 -1767
rect 330 -1775 331 -1767
rect 499 -1775 500 -1767
rect 502 -1775 504 -1767
rect 508 -1775 510 -1767
rect 512 -1775 513 -1767
rect 525 -1775 526 -1767
rect 528 -1775 529 -1767
rect 533 -1775 534 -1767
rect 536 -1775 541 -1767
rect 545 -1775 550 -1767
rect 552 -1775 553 -1767
rect 557 -1775 558 -1767
rect 560 -1775 562 -1767
rect 566 -1775 568 -1767
rect 570 -1775 571 -1767
rect 575 -1775 576 -1767
rect 578 -1775 583 -1767
rect 587 -1775 592 -1767
rect 594 -1775 595 -1767
rect 599 -1775 600 -1767
rect 602 -1775 604 -1767
rect 608 -1775 610 -1767
rect 612 -1775 613 -1767
rect 617 -1775 618 -1767
rect 620 -1775 625 -1767
rect 629 -1775 634 -1767
rect 636 -1775 637 -1767
rect 641 -1775 642 -1767
rect 644 -1775 646 -1767
rect 650 -1775 652 -1767
rect 654 -1775 655 -1767
rect 659 -1775 660 -1767
rect 662 -1775 667 -1767
rect 671 -1775 676 -1767
rect 678 -1775 679 -1767
rect 683 -1775 684 -1767
rect 686 -1775 687 -1767
rect 857 -1775 858 -1767
rect 860 -1775 862 -1767
rect 866 -1775 868 -1767
rect 870 -1775 871 -1767
rect 883 -1775 884 -1767
rect 886 -1775 887 -1767
rect 891 -1775 892 -1767
rect 894 -1775 899 -1767
rect 903 -1775 908 -1767
rect 910 -1775 911 -1767
rect 915 -1775 916 -1767
rect 918 -1775 920 -1767
rect 924 -1775 926 -1767
rect 928 -1775 929 -1767
rect 933 -1775 934 -1767
rect 936 -1775 941 -1767
rect 945 -1775 950 -1767
rect 952 -1775 953 -1767
rect 957 -1775 958 -1767
rect 960 -1775 962 -1767
rect 966 -1775 968 -1767
rect 970 -1775 971 -1767
rect 975 -1775 976 -1767
rect 978 -1775 983 -1767
rect 987 -1775 992 -1767
rect 994 -1775 995 -1767
rect 999 -1775 1000 -1767
rect 1002 -1775 1004 -1767
rect 1008 -1775 1010 -1767
rect 1012 -1775 1013 -1767
rect 1017 -1775 1018 -1767
rect 1020 -1775 1025 -1767
rect 1029 -1775 1034 -1767
rect 1036 -1775 1037 -1767
rect 1041 -1775 1042 -1767
rect 1044 -1775 1045 -1767
rect 1215 -1775 1216 -1767
rect 1218 -1775 1220 -1767
rect 1224 -1775 1226 -1767
rect 1228 -1775 1229 -1767
rect 1241 -1775 1242 -1767
rect 1244 -1775 1245 -1767
rect 1249 -1775 1250 -1767
rect 1252 -1775 1257 -1767
rect 1261 -1775 1266 -1767
rect 1268 -1775 1269 -1767
rect 1273 -1775 1274 -1767
rect 1276 -1775 1278 -1767
rect 1282 -1775 1284 -1767
rect 1286 -1775 1287 -1767
rect 1291 -1775 1292 -1767
rect 1294 -1775 1299 -1767
rect 1303 -1775 1308 -1767
rect 1310 -1775 1311 -1767
rect 1315 -1775 1316 -1767
rect 1318 -1775 1320 -1767
rect 1324 -1775 1326 -1767
rect 1328 -1775 1329 -1767
rect 1333 -1775 1334 -1767
rect 1336 -1775 1341 -1767
rect 1345 -1775 1350 -1767
rect 1352 -1775 1353 -1767
rect 1357 -1775 1358 -1767
rect 1360 -1775 1362 -1767
rect 1366 -1775 1368 -1767
rect 1370 -1775 1371 -1767
rect 1375 -1775 1376 -1767
rect 1378 -1775 1383 -1767
rect 1387 -1775 1392 -1767
rect 1394 -1775 1395 -1767
rect 1399 -1775 1400 -1767
rect 1402 -1775 1403 -1767
rect -1305 -1882 -1304 -1874
rect -1302 -1882 -1301 -1874
rect -1297 -1882 -1296 -1874
rect -1294 -1882 -1292 -1874
rect -1288 -1882 -1286 -1874
rect -1284 -1882 -1283 -1874
rect -931 -1882 -930 -1874
rect -928 -1882 -927 -1874
rect -923 -1882 -922 -1874
rect -920 -1882 -918 -1874
rect -914 -1882 -912 -1874
rect -910 -1882 -909 -1874
rect -573 -1882 -572 -1874
rect -570 -1882 -569 -1874
rect -565 -1882 -564 -1874
rect -562 -1882 -560 -1874
rect -556 -1882 -554 -1874
rect -552 -1882 -551 -1874
rect -215 -1882 -214 -1874
rect -212 -1882 -211 -1874
rect -207 -1882 -206 -1874
rect -204 -1882 -202 -1874
rect -198 -1882 -196 -1874
rect -194 -1882 -193 -1874
rect 143 -1882 144 -1874
rect 146 -1882 147 -1874
rect 151 -1882 152 -1874
rect 154 -1882 156 -1874
rect 160 -1882 162 -1874
rect 164 -1882 165 -1874
rect 499 -1882 500 -1874
rect 502 -1882 503 -1874
rect 507 -1882 508 -1874
rect 510 -1882 512 -1874
rect 516 -1882 518 -1874
rect 520 -1882 521 -1874
rect 857 -1882 858 -1874
rect 860 -1882 861 -1874
rect 865 -1882 866 -1874
rect 868 -1882 870 -1874
rect 874 -1882 876 -1874
rect 878 -1882 879 -1874
rect 1215 -1882 1216 -1874
rect 1218 -1882 1219 -1874
rect 1223 -1882 1224 -1874
rect 1226 -1882 1228 -1874
rect 1232 -1882 1234 -1874
rect 1236 -1882 1237 -1874
rect -1230 -2041 -1229 -2033
rect -1227 -2041 -1225 -2033
rect -1221 -2041 -1219 -2033
rect -1217 -2041 -1216 -2033
rect -1204 -2041 -1203 -2033
rect -1201 -2041 -1193 -2033
rect -1191 -2041 -1190 -2033
rect -1186 -2041 -1185 -2033
rect -1183 -2041 -1175 -2033
rect -1173 -2041 -1168 -2033
rect -1164 -2041 -1159 -2033
rect -1157 -2041 -1156 -2033
rect -1152 -2041 -1151 -2033
rect -1149 -2041 -1147 -2033
rect -1143 -2041 -1141 -2033
rect -1139 -2041 -1138 -2033
rect -931 -2041 -930 -2033
rect -928 -2041 -926 -2033
rect -922 -2041 -920 -2033
rect -918 -2041 -917 -2033
rect -905 -2041 -904 -2033
rect -902 -2041 -900 -2033
rect -896 -2041 -894 -2033
rect -892 -2041 -891 -2033
rect -879 -2041 -878 -2033
rect -876 -2041 -868 -2033
rect -866 -2041 -865 -2033
rect -861 -2041 -860 -2033
rect -858 -2041 -850 -2033
rect -848 -2041 -843 -2033
rect -839 -2041 -834 -2033
rect -832 -2041 -831 -2033
rect -827 -2041 -826 -2033
rect -824 -2041 -822 -2033
rect -818 -2041 -816 -2033
rect -814 -2041 -813 -2033
rect -801 -2041 -800 -2033
rect -798 -2041 -790 -2033
rect -788 -2041 -787 -2033
rect -783 -2041 -782 -2033
rect -780 -2041 -772 -2033
rect -770 -2041 -765 -2033
rect -761 -2041 -756 -2033
rect -754 -2041 -753 -2033
rect -749 -2041 -748 -2033
rect -746 -2041 -741 -2033
rect -737 -2041 -732 -2033
rect -730 -2041 -729 -2033
rect -717 -2041 -716 -2033
rect -714 -2041 -708 -2033
rect -706 -2041 -704 -2033
rect -700 -2041 -698 -2033
rect -696 -2041 -695 -2033
rect -573 -2041 -572 -2033
rect -570 -2041 -568 -2033
rect -564 -2041 -562 -2033
rect -560 -2041 -559 -2033
rect -547 -2041 -546 -2033
rect -544 -2041 -542 -2033
rect -538 -2041 -536 -2033
rect -534 -2041 -533 -2033
rect -521 -2041 -520 -2033
rect -518 -2041 -510 -2033
rect -508 -2041 -507 -2033
rect -503 -2041 -502 -2033
rect -500 -2041 -492 -2033
rect -490 -2041 -485 -2033
rect -481 -2041 -476 -2033
rect -474 -2041 -473 -2033
rect -469 -2041 -468 -2033
rect -466 -2041 -464 -2033
rect -460 -2041 -458 -2033
rect -456 -2041 -455 -2033
rect -443 -2041 -442 -2033
rect -440 -2041 -432 -2033
rect -430 -2041 -429 -2033
rect -425 -2041 -424 -2033
rect -422 -2041 -414 -2033
rect -412 -2041 -407 -2033
rect -403 -2041 -398 -2033
rect -396 -2041 -395 -2033
rect -391 -2041 -390 -2033
rect -388 -2041 -383 -2033
rect -379 -2041 -374 -2033
rect -372 -2041 -371 -2033
rect -359 -2041 -358 -2033
rect -356 -2041 -350 -2033
rect -348 -2041 -346 -2033
rect -342 -2041 -340 -2033
rect -338 -2041 -337 -2033
rect -215 -2041 -214 -2033
rect -212 -2041 -210 -2033
rect -206 -2041 -204 -2033
rect -202 -2041 -201 -2033
rect -189 -2041 -188 -2033
rect -186 -2041 -184 -2033
rect -180 -2041 -178 -2033
rect -176 -2041 -175 -2033
rect -163 -2041 -162 -2033
rect -160 -2041 -152 -2033
rect -150 -2041 -149 -2033
rect -145 -2041 -144 -2033
rect -142 -2041 -134 -2033
rect -132 -2041 -127 -2033
rect -123 -2041 -118 -2033
rect -116 -2041 -115 -2033
rect -111 -2041 -110 -2033
rect -108 -2041 -106 -2033
rect -102 -2041 -100 -2033
rect -98 -2041 -97 -2033
rect -85 -2041 -84 -2033
rect -82 -2041 -74 -2033
rect -72 -2041 -71 -2033
rect -67 -2041 -66 -2033
rect -64 -2041 -56 -2033
rect -54 -2041 -49 -2033
rect -45 -2041 -40 -2033
rect -38 -2041 -37 -2033
rect -33 -2041 -32 -2033
rect -30 -2041 -25 -2033
rect -21 -2041 -16 -2033
rect -14 -2041 -13 -2033
rect -1 -2041 0 -2033
rect 2 -2041 8 -2033
rect 10 -2041 12 -2033
rect 16 -2041 18 -2033
rect 20 -2041 21 -2033
rect 143 -2041 144 -2033
rect 146 -2041 148 -2033
rect 152 -2041 154 -2033
rect 156 -2041 157 -2033
rect 169 -2041 170 -2033
rect 172 -2041 174 -2033
rect 178 -2041 180 -2033
rect 182 -2041 183 -2033
rect 195 -2041 196 -2033
rect 198 -2041 206 -2033
rect 208 -2041 209 -2033
rect 213 -2041 214 -2033
rect 216 -2041 224 -2033
rect 226 -2041 231 -2033
rect 235 -2041 240 -2033
rect 242 -2041 243 -2033
rect 247 -2041 248 -2033
rect 250 -2041 252 -2033
rect 256 -2041 258 -2033
rect 260 -2041 261 -2033
rect 273 -2041 274 -2033
rect 276 -2041 284 -2033
rect 286 -2041 287 -2033
rect 291 -2041 292 -2033
rect 294 -2041 302 -2033
rect 304 -2041 309 -2033
rect 313 -2041 318 -2033
rect 320 -2041 321 -2033
rect 325 -2041 326 -2033
rect 328 -2041 333 -2033
rect 337 -2041 342 -2033
rect 344 -2041 345 -2033
rect 357 -2041 358 -2033
rect 360 -2041 366 -2033
rect 368 -2041 370 -2033
rect 374 -2041 376 -2033
rect 378 -2041 379 -2033
rect 499 -2041 500 -2033
rect 502 -2041 504 -2033
rect 508 -2041 510 -2033
rect 512 -2041 513 -2033
rect 525 -2041 526 -2033
rect 528 -2041 530 -2033
rect 534 -2041 536 -2033
rect 538 -2041 539 -2033
rect 551 -2041 552 -2033
rect 554 -2041 562 -2033
rect 564 -2041 565 -2033
rect 569 -2041 570 -2033
rect 572 -2041 580 -2033
rect 582 -2041 587 -2033
rect 591 -2041 596 -2033
rect 598 -2041 599 -2033
rect 603 -2041 604 -2033
rect 606 -2041 608 -2033
rect 612 -2041 614 -2033
rect 616 -2041 617 -2033
rect 629 -2041 630 -2033
rect 632 -2041 640 -2033
rect 642 -2041 643 -2033
rect 647 -2041 648 -2033
rect 650 -2041 658 -2033
rect 660 -2041 665 -2033
rect 669 -2041 674 -2033
rect 676 -2041 677 -2033
rect 681 -2041 682 -2033
rect 684 -2041 689 -2033
rect 693 -2041 698 -2033
rect 700 -2041 701 -2033
rect 713 -2041 714 -2033
rect 716 -2041 722 -2033
rect 724 -2041 726 -2033
rect 730 -2041 732 -2033
rect 734 -2041 735 -2033
rect 857 -2041 858 -2033
rect 860 -2041 862 -2033
rect 866 -2041 868 -2033
rect 870 -2041 871 -2033
rect 883 -2041 884 -2033
rect 886 -2041 888 -2033
rect 892 -2041 894 -2033
rect 896 -2041 897 -2033
rect 909 -2041 910 -2033
rect 912 -2041 920 -2033
rect 922 -2041 923 -2033
rect 927 -2041 928 -2033
rect 930 -2041 938 -2033
rect 940 -2041 945 -2033
rect 949 -2041 954 -2033
rect 956 -2041 957 -2033
rect 961 -2041 962 -2033
rect 964 -2041 966 -2033
rect 970 -2041 972 -2033
rect 974 -2041 975 -2033
rect 987 -2041 988 -2033
rect 990 -2041 998 -2033
rect 1000 -2041 1001 -2033
rect 1005 -2041 1006 -2033
rect 1008 -2041 1016 -2033
rect 1018 -2041 1023 -2033
rect 1027 -2041 1032 -2033
rect 1034 -2041 1035 -2033
rect 1039 -2041 1040 -2033
rect 1042 -2041 1047 -2033
rect 1051 -2041 1056 -2033
rect 1058 -2041 1059 -2033
rect 1071 -2041 1072 -2033
rect 1074 -2041 1080 -2033
rect 1082 -2041 1084 -2033
rect 1088 -2041 1090 -2033
rect 1092 -2041 1093 -2033
rect 1215 -2041 1216 -2033
rect 1218 -2041 1220 -2033
rect 1224 -2041 1226 -2033
rect 1228 -2041 1229 -2033
rect 1241 -2041 1242 -2033
rect 1244 -2041 1246 -2033
rect 1250 -2041 1252 -2033
rect 1254 -2041 1255 -2033
rect 1267 -2041 1268 -2033
rect 1270 -2041 1278 -2033
rect 1280 -2041 1281 -2033
rect 1285 -2041 1286 -2033
rect 1288 -2041 1296 -2033
rect 1298 -2041 1303 -2033
rect 1307 -2041 1312 -2033
rect 1314 -2041 1315 -2033
rect 1319 -2041 1320 -2033
rect 1322 -2041 1324 -2033
rect 1328 -2041 1330 -2033
rect 1332 -2041 1333 -2033
rect 1345 -2041 1346 -2033
rect 1348 -2041 1356 -2033
rect 1358 -2041 1359 -2033
rect 1363 -2041 1364 -2033
rect 1366 -2041 1374 -2033
rect 1376 -2041 1381 -2033
rect 1385 -2041 1390 -2033
rect 1392 -2041 1393 -2033
rect 1397 -2041 1398 -2033
rect 1400 -2041 1405 -2033
rect 1409 -2041 1414 -2033
rect 1416 -2041 1417 -2033
rect 1429 -2041 1430 -2033
rect 1432 -2041 1438 -2033
rect 1440 -2041 1442 -2033
rect 1446 -2041 1448 -2033
rect 1450 -2041 1451 -2033
rect -1230 -2185 -1229 -2177
rect -1227 -2185 -1225 -2177
rect -1221 -2185 -1219 -2177
rect -1217 -2185 -1216 -2177
rect -1204 -2185 -1203 -2177
rect -1201 -2185 -1200 -2177
rect -1196 -2185 -1195 -2177
rect -1193 -2185 -1188 -2177
rect -1184 -2185 -1179 -2177
rect -1177 -2185 -1176 -2177
rect -1172 -2185 -1171 -2177
rect -1169 -2185 -1167 -2177
rect -1163 -2185 -1161 -2177
rect -1159 -2185 -1158 -2177
rect -1154 -2185 -1153 -2177
rect -1151 -2185 -1146 -2177
rect -1142 -2185 -1137 -2177
rect -1135 -2185 -1134 -2177
rect -1130 -2185 -1129 -2177
rect -1127 -2185 -1125 -2177
rect -1121 -2185 -1119 -2177
rect -1117 -2185 -1116 -2177
rect -1112 -2185 -1111 -2177
rect -1109 -2185 -1104 -2177
rect -1100 -2185 -1095 -2177
rect -1093 -2185 -1092 -2177
rect -1088 -2185 -1087 -2177
rect -1085 -2185 -1083 -2177
rect -1079 -2185 -1077 -2177
rect -1075 -2185 -1074 -2177
rect -1070 -2185 -1069 -2177
rect -1067 -2185 -1062 -2177
rect -1058 -2185 -1053 -2177
rect -1051 -2185 -1050 -2177
rect -1046 -2185 -1045 -2177
rect -1043 -2185 -1042 -2177
rect -931 -2185 -930 -2177
rect -928 -2185 -926 -2177
rect -922 -2185 -920 -2177
rect -918 -2185 -917 -2177
rect -905 -2185 -904 -2177
rect -902 -2185 -901 -2177
rect -897 -2185 -896 -2177
rect -894 -2185 -889 -2177
rect -885 -2185 -880 -2177
rect -878 -2185 -877 -2177
rect -873 -2185 -872 -2177
rect -870 -2185 -868 -2177
rect -864 -2185 -862 -2177
rect -860 -2185 -859 -2177
rect -855 -2185 -854 -2177
rect -852 -2185 -847 -2177
rect -843 -2185 -838 -2177
rect -836 -2185 -835 -2177
rect -831 -2185 -830 -2177
rect -828 -2185 -826 -2177
rect -822 -2185 -820 -2177
rect -818 -2185 -817 -2177
rect -813 -2185 -812 -2177
rect -810 -2185 -805 -2177
rect -801 -2185 -796 -2177
rect -794 -2185 -793 -2177
rect -789 -2185 -788 -2177
rect -786 -2185 -784 -2177
rect -780 -2185 -778 -2177
rect -776 -2185 -775 -2177
rect -771 -2185 -770 -2177
rect -768 -2185 -763 -2177
rect -759 -2185 -754 -2177
rect -752 -2185 -751 -2177
rect -747 -2185 -746 -2177
rect -744 -2185 -743 -2177
rect -573 -2185 -572 -2177
rect -570 -2185 -568 -2177
rect -564 -2185 -562 -2177
rect -560 -2185 -559 -2177
rect -547 -2185 -546 -2177
rect -544 -2185 -543 -2177
rect -539 -2185 -538 -2177
rect -536 -2185 -531 -2177
rect -527 -2185 -522 -2177
rect -520 -2185 -519 -2177
rect -515 -2185 -514 -2177
rect -512 -2185 -510 -2177
rect -506 -2185 -504 -2177
rect -502 -2185 -501 -2177
rect -497 -2185 -496 -2177
rect -494 -2185 -489 -2177
rect -485 -2185 -480 -2177
rect -478 -2185 -477 -2177
rect -473 -2185 -472 -2177
rect -470 -2185 -468 -2177
rect -464 -2185 -462 -2177
rect -460 -2185 -459 -2177
rect -455 -2185 -454 -2177
rect -452 -2185 -447 -2177
rect -443 -2185 -438 -2177
rect -436 -2185 -435 -2177
rect -431 -2185 -430 -2177
rect -428 -2185 -426 -2177
rect -422 -2185 -420 -2177
rect -418 -2185 -417 -2177
rect -413 -2185 -412 -2177
rect -410 -2185 -405 -2177
rect -401 -2185 -396 -2177
rect -394 -2185 -393 -2177
rect -389 -2185 -388 -2177
rect -386 -2185 -385 -2177
rect -215 -2185 -214 -2177
rect -212 -2185 -210 -2177
rect -206 -2185 -204 -2177
rect -202 -2185 -201 -2177
rect -189 -2185 -188 -2177
rect -186 -2185 -185 -2177
rect -181 -2185 -180 -2177
rect -178 -2185 -173 -2177
rect -169 -2185 -164 -2177
rect -162 -2185 -161 -2177
rect -157 -2185 -156 -2177
rect -154 -2185 -152 -2177
rect -148 -2185 -146 -2177
rect -144 -2185 -143 -2177
rect -139 -2185 -138 -2177
rect -136 -2185 -131 -2177
rect -127 -2185 -122 -2177
rect -120 -2185 -119 -2177
rect -115 -2185 -114 -2177
rect -112 -2185 -110 -2177
rect -106 -2185 -104 -2177
rect -102 -2185 -101 -2177
rect -97 -2185 -96 -2177
rect -94 -2185 -89 -2177
rect -85 -2185 -80 -2177
rect -78 -2185 -77 -2177
rect -73 -2185 -72 -2177
rect -70 -2185 -68 -2177
rect -64 -2185 -62 -2177
rect -60 -2185 -59 -2177
rect -55 -2185 -54 -2177
rect -52 -2185 -47 -2177
rect -43 -2185 -38 -2177
rect -36 -2185 -35 -2177
rect -31 -2185 -30 -2177
rect -28 -2185 -27 -2177
rect 143 -2185 144 -2177
rect 146 -2185 148 -2177
rect 152 -2185 154 -2177
rect 156 -2185 157 -2177
rect 169 -2185 170 -2177
rect 172 -2185 173 -2177
rect 177 -2185 178 -2177
rect 180 -2185 185 -2177
rect 189 -2185 194 -2177
rect 196 -2185 197 -2177
rect 201 -2185 202 -2177
rect 204 -2185 206 -2177
rect 210 -2185 212 -2177
rect 214 -2185 215 -2177
rect 219 -2185 220 -2177
rect 222 -2185 227 -2177
rect 231 -2185 236 -2177
rect 238 -2185 239 -2177
rect 243 -2185 244 -2177
rect 246 -2185 248 -2177
rect 252 -2185 254 -2177
rect 256 -2185 257 -2177
rect 261 -2185 262 -2177
rect 264 -2185 269 -2177
rect 273 -2185 278 -2177
rect 280 -2185 281 -2177
rect 285 -2185 286 -2177
rect 288 -2185 290 -2177
rect 294 -2185 296 -2177
rect 298 -2185 299 -2177
rect 303 -2185 304 -2177
rect 306 -2185 311 -2177
rect 315 -2185 320 -2177
rect 322 -2185 323 -2177
rect 327 -2185 328 -2177
rect 330 -2185 331 -2177
rect 499 -2185 500 -2177
rect 502 -2185 504 -2177
rect 508 -2185 510 -2177
rect 512 -2185 513 -2177
rect 525 -2185 526 -2177
rect 528 -2185 529 -2177
rect 533 -2185 534 -2177
rect 536 -2185 541 -2177
rect 545 -2185 550 -2177
rect 552 -2185 553 -2177
rect 557 -2185 558 -2177
rect 560 -2185 562 -2177
rect 566 -2185 568 -2177
rect 570 -2185 571 -2177
rect 575 -2185 576 -2177
rect 578 -2185 583 -2177
rect 587 -2185 592 -2177
rect 594 -2185 595 -2177
rect 599 -2185 600 -2177
rect 602 -2185 604 -2177
rect 608 -2185 610 -2177
rect 612 -2185 613 -2177
rect 617 -2185 618 -2177
rect 620 -2185 625 -2177
rect 629 -2185 634 -2177
rect 636 -2185 637 -2177
rect 641 -2185 642 -2177
rect 644 -2185 646 -2177
rect 650 -2185 652 -2177
rect 654 -2185 655 -2177
rect 659 -2185 660 -2177
rect 662 -2185 667 -2177
rect 671 -2185 676 -2177
rect 678 -2185 679 -2177
rect 683 -2185 684 -2177
rect 686 -2185 687 -2177
rect -1555 -2356 -1554 -2348
rect -1552 -2356 -1550 -2348
rect -1546 -2356 -1544 -2348
rect -1542 -2356 -1541 -2348
rect -1529 -2356 -1528 -2348
rect -1526 -2356 -1525 -2348
rect -1521 -2356 -1520 -2348
rect -1518 -2356 -1513 -2348
rect -1509 -2356 -1504 -2348
rect -1502 -2356 -1501 -2348
rect -1497 -2356 -1496 -2348
rect -1494 -2356 -1492 -2348
rect -1488 -2356 -1486 -2348
rect -1484 -2356 -1483 -2348
rect -1479 -2356 -1478 -2348
rect -1476 -2356 -1471 -2348
rect -1467 -2356 -1462 -2348
rect -1460 -2356 -1459 -2348
rect -1455 -2356 -1454 -2348
rect -1452 -2356 -1450 -2348
rect -1446 -2356 -1444 -2348
rect -1442 -2356 -1441 -2348
rect -1437 -2356 -1436 -2348
rect -1434 -2356 -1429 -2348
rect -1425 -2356 -1420 -2348
rect -1418 -2356 -1417 -2348
rect -1413 -2356 -1412 -2348
rect -1410 -2356 -1408 -2348
rect -1404 -2356 -1402 -2348
rect -1400 -2356 -1399 -2348
rect -1395 -2356 -1394 -2348
rect -1392 -2356 -1387 -2348
rect -1383 -2356 -1378 -2348
rect -1376 -2356 -1375 -2348
rect -1371 -2356 -1370 -2348
rect -1368 -2356 -1367 -2348
rect -1230 -2356 -1229 -2348
rect -1227 -2356 -1225 -2348
rect -1221 -2356 -1219 -2348
rect -1217 -2356 -1216 -2348
rect -1204 -2356 -1203 -2348
rect -1201 -2356 -1200 -2348
rect -1196 -2356 -1195 -2348
rect -1193 -2356 -1188 -2348
rect -1184 -2356 -1179 -2348
rect -1177 -2356 -1176 -2348
rect -1172 -2356 -1171 -2348
rect -1169 -2356 -1167 -2348
rect -1163 -2356 -1161 -2348
rect -1159 -2356 -1158 -2348
rect -1154 -2356 -1153 -2348
rect -1151 -2356 -1146 -2348
rect -1142 -2356 -1137 -2348
rect -1135 -2356 -1134 -2348
rect -1130 -2356 -1129 -2348
rect -1127 -2356 -1125 -2348
rect -1121 -2356 -1119 -2348
rect -1117 -2356 -1116 -2348
rect -1112 -2356 -1111 -2348
rect -1109 -2356 -1104 -2348
rect -1100 -2356 -1095 -2348
rect -1093 -2356 -1092 -2348
rect -1088 -2356 -1087 -2348
rect -1085 -2356 -1083 -2348
rect -1079 -2356 -1077 -2348
rect -1075 -2356 -1074 -2348
rect -1070 -2356 -1069 -2348
rect -1067 -2356 -1062 -2348
rect -1058 -2356 -1053 -2348
rect -1051 -2356 -1050 -2348
rect -1046 -2356 -1045 -2348
rect -1043 -2356 -1042 -2348
rect -931 -2356 -930 -2348
rect -928 -2356 -926 -2348
rect -922 -2356 -920 -2348
rect -918 -2356 -917 -2348
rect -905 -2356 -904 -2348
rect -902 -2356 -901 -2348
rect -897 -2356 -896 -2348
rect -894 -2356 -889 -2348
rect -885 -2356 -880 -2348
rect -878 -2356 -877 -2348
rect -873 -2356 -872 -2348
rect -870 -2356 -868 -2348
rect -864 -2356 -862 -2348
rect -860 -2356 -859 -2348
rect -855 -2356 -854 -2348
rect -852 -2356 -847 -2348
rect -843 -2356 -838 -2348
rect -836 -2356 -835 -2348
rect -831 -2356 -830 -2348
rect -828 -2356 -826 -2348
rect -822 -2356 -820 -2348
rect -818 -2356 -817 -2348
rect -813 -2356 -812 -2348
rect -810 -2356 -805 -2348
rect -801 -2356 -796 -2348
rect -794 -2356 -793 -2348
rect -789 -2356 -788 -2348
rect -786 -2356 -784 -2348
rect -780 -2356 -778 -2348
rect -776 -2356 -775 -2348
rect -771 -2356 -770 -2348
rect -768 -2356 -763 -2348
rect -759 -2356 -754 -2348
rect -752 -2356 -751 -2348
rect -747 -2356 -746 -2348
rect -744 -2356 -743 -2348
rect -573 -2356 -572 -2348
rect -570 -2356 -568 -2348
rect -564 -2356 -562 -2348
rect -560 -2356 -559 -2348
rect -547 -2356 -546 -2348
rect -544 -2356 -543 -2348
rect -539 -2356 -538 -2348
rect -536 -2356 -531 -2348
rect -527 -2356 -522 -2348
rect -520 -2356 -519 -2348
rect -515 -2356 -514 -2348
rect -512 -2356 -510 -2348
rect -506 -2356 -504 -2348
rect -502 -2356 -501 -2348
rect -497 -2356 -496 -2348
rect -494 -2356 -489 -2348
rect -485 -2356 -480 -2348
rect -478 -2356 -477 -2348
rect -473 -2356 -472 -2348
rect -470 -2356 -468 -2348
rect -464 -2356 -462 -2348
rect -460 -2356 -459 -2348
rect -455 -2356 -454 -2348
rect -452 -2356 -447 -2348
rect -443 -2356 -438 -2348
rect -436 -2356 -435 -2348
rect -431 -2356 -430 -2348
rect -428 -2356 -426 -2348
rect -422 -2356 -420 -2348
rect -418 -2356 -417 -2348
rect -413 -2356 -412 -2348
rect -410 -2356 -405 -2348
rect -401 -2356 -396 -2348
rect -394 -2356 -393 -2348
rect -389 -2356 -388 -2348
rect -386 -2356 -385 -2348
rect -215 -2356 -214 -2348
rect -212 -2356 -210 -2348
rect -206 -2356 -204 -2348
rect -202 -2356 -201 -2348
rect -189 -2356 -188 -2348
rect -186 -2356 -185 -2348
rect -181 -2356 -180 -2348
rect -178 -2356 -173 -2348
rect -169 -2356 -164 -2348
rect -162 -2356 -161 -2348
rect -157 -2356 -156 -2348
rect -154 -2356 -152 -2348
rect -148 -2356 -146 -2348
rect -144 -2356 -143 -2348
rect -139 -2356 -138 -2348
rect -136 -2356 -131 -2348
rect -127 -2356 -122 -2348
rect -120 -2356 -119 -2348
rect -115 -2356 -114 -2348
rect -112 -2356 -110 -2348
rect -106 -2356 -104 -2348
rect -102 -2356 -101 -2348
rect -97 -2356 -96 -2348
rect -94 -2356 -89 -2348
rect -85 -2356 -80 -2348
rect -78 -2356 -77 -2348
rect -73 -2356 -72 -2348
rect -70 -2356 -68 -2348
rect -64 -2356 -62 -2348
rect -60 -2356 -59 -2348
rect -55 -2356 -54 -2348
rect -52 -2356 -47 -2348
rect -43 -2356 -38 -2348
rect -36 -2356 -35 -2348
rect -31 -2356 -30 -2348
rect -28 -2356 -27 -2348
rect 143 -2356 144 -2348
rect 146 -2356 148 -2348
rect 152 -2356 154 -2348
rect 156 -2356 157 -2348
rect 169 -2356 170 -2348
rect 172 -2356 173 -2348
rect 177 -2356 178 -2348
rect 180 -2356 185 -2348
rect 189 -2356 194 -2348
rect 196 -2356 197 -2348
rect 201 -2356 202 -2348
rect 204 -2356 206 -2348
rect 210 -2356 212 -2348
rect 214 -2356 215 -2348
rect 219 -2356 220 -2348
rect 222 -2356 227 -2348
rect 231 -2356 236 -2348
rect 238 -2356 239 -2348
rect 243 -2356 244 -2348
rect 246 -2356 248 -2348
rect 252 -2356 254 -2348
rect 256 -2356 257 -2348
rect 261 -2356 262 -2348
rect 264 -2356 269 -2348
rect 273 -2356 278 -2348
rect 280 -2356 281 -2348
rect 285 -2356 286 -2348
rect 288 -2356 290 -2348
rect 294 -2356 296 -2348
rect 298 -2356 299 -2348
rect 303 -2356 304 -2348
rect 306 -2356 311 -2348
rect 315 -2356 320 -2348
rect 322 -2356 323 -2348
rect 327 -2356 328 -2348
rect 330 -2356 331 -2348
rect 499 -2356 500 -2348
rect 502 -2356 504 -2348
rect 508 -2356 510 -2348
rect 512 -2356 513 -2348
rect 525 -2356 526 -2348
rect 528 -2356 529 -2348
rect 533 -2356 534 -2348
rect 536 -2356 541 -2348
rect 545 -2356 550 -2348
rect 552 -2356 553 -2348
rect 557 -2356 558 -2348
rect 560 -2356 562 -2348
rect 566 -2356 568 -2348
rect 570 -2356 571 -2348
rect 575 -2356 576 -2348
rect 578 -2356 583 -2348
rect 587 -2356 592 -2348
rect 594 -2356 595 -2348
rect 599 -2356 600 -2348
rect 602 -2356 604 -2348
rect 608 -2356 610 -2348
rect 612 -2356 613 -2348
rect 617 -2356 618 -2348
rect 620 -2356 625 -2348
rect 629 -2356 634 -2348
rect 636 -2356 637 -2348
rect 641 -2356 642 -2348
rect 644 -2356 646 -2348
rect 650 -2356 652 -2348
rect 654 -2356 655 -2348
rect 659 -2356 660 -2348
rect 662 -2356 667 -2348
rect 671 -2356 676 -2348
rect 678 -2356 679 -2348
rect 683 -2356 684 -2348
rect 686 -2356 687 -2348
rect 857 -2356 858 -2348
rect 860 -2356 862 -2348
rect 866 -2356 868 -2348
rect 870 -2356 871 -2348
rect 883 -2356 884 -2348
rect 886 -2356 887 -2348
rect 891 -2356 892 -2348
rect 894 -2356 899 -2348
rect 903 -2356 908 -2348
rect 910 -2356 911 -2348
rect 915 -2356 916 -2348
rect 918 -2356 920 -2348
rect 924 -2356 926 -2348
rect 928 -2356 929 -2348
rect 933 -2356 934 -2348
rect 936 -2356 941 -2348
rect 945 -2356 950 -2348
rect 952 -2356 953 -2348
rect 957 -2356 958 -2348
rect 960 -2356 962 -2348
rect 966 -2356 968 -2348
rect 970 -2356 971 -2348
rect 975 -2356 976 -2348
rect 978 -2356 983 -2348
rect 987 -2356 992 -2348
rect 994 -2356 995 -2348
rect 999 -2356 1000 -2348
rect 1002 -2356 1004 -2348
rect 1008 -2356 1010 -2348
rect 1012 -2356 1013 -2348
rect 1017 -2356 1018 -2348
rect 1020 -2356 1025 -2348
rect 1029 -2356 1034 -2348
rect 1036 -2356 1037 -2348
rect 1041 -2356 1042 -2348
rect 1044 -2356 1045 -2348
rect 1215 -2356 1216 -2348
rect 1218 -2356 1220 -2348
rect 1224 -2356 1226 -2348
rect 1228 -2356 1229 -2348
rect 1241 -2356 1242 -2348
rect 1244 -2356 1245 -2348
rect 1249 -2356 1250 -2348
rect 1252 -2356 1257 -2348
rect 1261 -2356 1266 -2348
rect 1268 -2356 1269 -2348
rect 1273 -2356 1274 -2348
rect 1276 -2356 1278 -2348
rect 1282 -2356 1284 -2348
rect 1286 -2356 1287 -2348
rect 1291 -2356 1292 -2348
rect 1294 -2356 1299 -2348
rect 1303 -2356 1308 -2348
rect 1310 -2356 1311 -2348
rect 1315 -2356 1316 -2348
rect 1318 -2356 1320 -2348
rect 1324 -2356 1326 -2348
rect 1328 -2356 1329 -2348
rect 1333 -2356 1334 -2348
rect 1336 -2356 1341 -2348
rect 1345 -2356 1350 -2348
rect 1352 -2356 1353 -2348
rect 1357 -2356 1358 -2348
rect 1360 -2356 1362 -2348
rect 1366 -2356 1368 -2348
rect 1370 -2356 1371 -2348
rect 1375 -2356 1376 -2348
rect 1378 -2356 1383 -2348
rect 1387 -2356 1392 -2348
rect 1394 -2356 1395 -2348
rect 1399 -2356 1400 -2348
rect 1402 -2356 1403 -2348
rect -1555 -2527 -1554 -2519
rect -1552 -2527 -1550 -2519
rect -1546 -2527 -1544 -2519
rect -1542 -2527 -1541 -2519
rect -1529 -2527 -1528 -2519
rect -1526 -2527 -1525 -2519
rect -1521 -2527 -1520 -2519
rect -1518 -2527 -1513 -2519
rect -1509 -2527 -1504 -2519
rect -1502 -2527 -1501 -2519
rect -1497 -2527 -1496 -2519
rect -1494 -2527 -1492 -2519
rect -1488 -2527 -1486 -2519
rect -1484 -2527 -1483 -2519
rect -1479 -2527 -1478 -2519
rect -1476 -2527 -1471 -2519
rect -1467 -2527 -1462 -2519
rect -1460 -2527 -1459 -2519
rect -1455 -2527 -1454 -2519
rect -1452 -2527 -1450 -2519
rect -1446 -2527 -1444 -2519
rect -1442 -2527 -1441 -2519
rect -1437 -2527 -1436 -2519
rect -1434 -2527 -1429 -2519
rect -1425 -2527 -1420 -2519
rect -1418 -2527 -1417 -2519
rect -1413 -2527 -1412 -2519
rect -1410 -2527 -1408 -2519
rect -1404 -2527 -1402 -2519
rect -1400 -2527 -1399 -2519
rect -1395 -2527 -1394 -2519
rect -1392 -2527 -1387 -2519
rect -1383 -2527 -1378 -2519
rect -1376 -2527 -1375 -2519
rect -1371 -2527 -1370 -2519
rect -1368 -2527 -1367 -2519
rect -1230 -2527 -1229 -2519
rect -1227 -2527 -1225 -2519
rect -1221 -2527 -1219 -2519
rect -1217 -2527 -1216 -2519
rect -1204 -2527 -1203 -2519
rect -1201 -2527 -1200 -2519
rect -1196 -2527 -1195 -2519
rect -1193 -2527 -1188 -2519
rect -1184 -2527 -1179 -2519
rect -1177 -2527 -1176 -2519
rect -1172 -2527 -1171 -2519
rect -1169 -2527 -1167 -2519
rect -1163 -2527 -1161 -2519
rect -1159 -2527 -1158 -2519
rect -1154 -2527 -1153 -2519
rect -1151 -2527 -1146 -2519
rect -1142 -2527 -1137 -2519
rect -1135 -2527 -1134 -2519
rect -1130 -2527 -1129 -2519
rect -1127 -2527 -1125 -2519
rect -1121 -2527 -1119 -2519
rect -1117 -2527 -1116 -2519
rect -1112 -2527 -1111 -2519
rect -1109 -2527 -1104 -2519
rect -1100 -2527 -1095 -2519
rect -1093 -2527 -1092 -2519
rect -1088 -2527 -1087 -2519
rect -1085 -2527 -1083 -2519
rect -1079 -2527 -1077 -2519
rect -1075 -2527 -1074 -2519
rect -1070 -2527 -1069 -2519
rect -1067 -2527 -1062 -2519
rect -1058 -2527 -1053 -2519
rect -1051 -2527 -1050 -2519
rect -1046 -2527 -1045 -2519
rect -1043 -2527 -1042 -2519
rect -931 -2527 -930 -2519
rect -928 -2527 -926 -2519
rect -922 -2527 -920 -2519
rect -918 -2527 -917 -2519
rect -905 -2527 -904 -2519
rect -902 -2527 -901 -2519
rect -897 -2527 -896 -2519
rect -894 -2527 -889 -2519
rect -885 -2527 -880 -2519
rect -878 -2527 -877 -2519
rect -873 -2527 -872 -2519
rect -870 -2527 -868 -2519
rect -864 -2527 -862 -2519
rect -860 -2527 -859 -2519
rect -855 -2527 -854 -2519
rect -852 -2527 -847 -2519
rect -843 -2527 -838 -2519
rect -836 -2527 -835 -2519
rect -831 -2527 -830 -2519
rect -828 -2527 -826 -2519
rect -822 -2527 -820 -2519
rect -818 -2527 -817 -2519
rect -813 -2527 -812 -2519
rect -810 -2527 -805 -2519
rect -801 -2527 -796 -2519
rect -794 -2527 -793 -2519
rect -789 -2527 -788 -2519
rect -786 -2527 -784 -2519
rect -780 -2527 -778 -2519
rect -776 -2527 -775 -2519
rect -771 -2527 -770 -2519
rect -768 -2527 -763 -2519
rect -759 -2527 -754 -2519
rect -752 -2527 -751 -2519
rect -747 -2527 -746 -2519
rect -744 -2527 -743 -2519
rect -573 -2527 -572 -2519
rect -570 -2527 -568 -2519
rect -564 -2527 -562 -2519
rect -560 -2527 -559 -2519
rect -547 -2527 -546 -2519
rect -544 -2527 -543 -2519
rect -539 -2527 -538 -2519
rect -536 -2527 -531 -2519
rect -527 -2527 -522 -2519
rect -520 -2527 -519 -2519
rect -515 -2527 -514 -2519
rect -512 -2527 -510 -2519
rect -506 -2527 -504 -2519
rect -502 -2527 -501 -2519
rect -497 -2527 -496 -2519
rect -494 -2527 -489 -2519
rect -485 -2527 -480 -2519
rect -478 -2527 -477 -2519
rect -473 -2527 -472 -2519
rect -470 -2527 -468 -2519
rect -464 -2527 -462 -2519
rect -460 -2527 -459 -2519
rect -455 -2527 -454 -2519
rect -452 -2527 -447 -2519
rect -443 -2527 -438 -2519
rect -436 -2527 -435 -2519
rect -431 -2527 -430 -2519
rect -428 -2527 -426 -2519
rect -422 -2527 -420 -2519
rect -418 -2527 -417 -2519
rect -413 -2527 -412 -2519
rect -410 -2527 -405 -2519
rect -401 -2527 -396 -2519
rect -394 -2527 -393 -2519
rect -389 -2527 -388 -2519
rect -386 -2527 -385 -2519
rect -216 -2527 -215 -2519
rect -213 -2527 -211 -2519
rect -207 -2527 -205 -2519
rect -203 -2527 -202 -2519
rect -190 -2527 -189 -2519
rect -187 -2527 -186 -2519
rect -182 -2527 -181 -2519
rect -179 -2527 -174 -2519
rect -170 -2527 -165 -2519
rect -163 -2527 -162 -2519
rect -158 -2527 -157 -2519
rect -155 -2527 -153 -2519
rect -149 -2527 -147 -2519
rect -145 -2527 -144 -2519
rect -140 -2527 -139 -2519
rect -137 -2527 -132 -2519
rect -128 -2527 -123 -2519
rect -121 -2527 -120 -2519
rect -116 -2527 -115 -2519
rect -113 -2527 -111 -2519
rect -107 -2527 -105 -2519
rect -103 -2527 -102 -2519
rect -98 -2527 -97 -2519
rect -95 -2527 -90 -2519
rect -86 -2527 -81 -2519
rect -79 -2527 -78 -2519
rect -74 -2527 -73 -2519
rect -71 -2527 -69 -2519
rect -65 -2527 -63 -2519
rect -61 -2527 -60 -2519
rect -56 -2527 -55 -2519
rect -53 -2527 -48 -2519
rect -44 -2527 -39 -2519
rect -37 -2527 -36 -2519
rect -32 -2527 -31 -2519
rect -29 -2527 -28 -2519
rect 143 -2527 144 -2519
rect 146 -2527 148 -2519
rect 152 -2527 154 -2519
rect 156 -2527 157 -2519
rect 169 -2527 170 -2519
rect 172 -2527 173 -2519
rect 177 -2527 178 -2519
rect 180 -2527 185 -2519
rect 189 -2527 194 -2519
rect 196 -2527 197 -2519
rect 201 -2527 202 -2519
rect 204 -2527 206 -2519
rect 210 -2527 212 -2519
rect 214 -2527 215 -2519
rect 219 -2527 220 -2519
rect 222 -2527 227 -2519
rect 231 -2527 236 -2519
rect 238 -2527 239 -2519
rect 243 -2527 244 -2519
rect 246 -2527 248 -2519
rect 252 -2527 254 -2519
rect 256 -2527 257 -2519
rect 261 -2527 262 -2519
rect 264 -2527 269 -2519
rect 273 -2527 278 -2519
rect 280 -2527 281 -2519
rect 285 -2527 286 -2519
rect 288 -2527 290 -2519
rect 294 -2527 296 -2519
rect 298 -2527 299 -2519
rect 303 -2527 304 -2519
rect 306 -2527 311 -2519
rect 315 -2527 320 -2519
rect 322 -2527 323 -2519
rect 327 -2527 328 -2519
rect 330 -2527 331 -2519
rect 499 -2527 500 -2519
rect 502 -2527 504 -2519
rect 508 -2527 510 -2519
rect 512 -2527 513 -2519
rect 525 -2527 526 -2519
rect 528 -2527 529 -2519
rect 533 -2527 534 -2519
rect 536 -2527 541 -2519
rect 545 -2527 550 -2519
rect 552 -2527 553 -2519
rect 557 -2527 558 -2519
rect 560 -2527 562 -2519
rect 566 -2527 568 -2519
rect 570 -2527 571 -2519
rect 575 -2527 576 -2519
rect 578 -2527 583 -2519
rect 587 -2527 592 -2519
rect 594 -2527 595 -2519
rect 599 -2527 600 -2519
rect 602 -2527 604 -2519
rect 608 -2527 610 -2519
rect 612 -2527 613 -2519
rect 617 -2527 618 -2519
rect 620 -2527 625 -2519
rect 629 -2527 634 -2519
rect 636 -2527 637 -2519
rect 641 -2527 642 -2519
rect 644 -2527 646 -2519
rect 650 -2527 652 -2519
rect 654 -2527 655 -2519
rect 659 -2527 660 -2519
rect 662 -2527 667 -2519
rect 671 -2527 676 -2519
rect 678 -2527 679 -2519
rect 683 -2527 684 -2519
rect 686 -2527 687 -2519
rect 857 -2527 858 -2519
rect 860 -2527 862 -2519
rect 866 -2527 868 -2519
rect 870 -2527 871 -2519
rect 883 -2527 884 -2519
rect 886 -2527 887 -2519
rect 891 -2527 892 -2519
rect 894 -2527 899 -2519
rect 903 -2527 908 -2519
rect 910 -2527 911 -2519
rect 915 -2527 916 -2519
rect 918 -2527 920 -2519
rect 924 -2527 926 -2519
rect 928 -2527 929 -2519
rect 933 -2527 934 -2519
rect 936 -2527 941 -2519
rect 945 -2527 950 -2519
rect 952 -2527 953 -2519
rect 957 -2527 958 -2519
rect 960 -2527 962 -2519
rect 966 -2527 968 -2519
rect 970 -2527 971 -2519
rect 975 -2527 976 -2519
rect 978 -2527 983 -2519
rect 987 -2527 992 -2519
rect 994 -2527 995 -2519
rect 999 -2527 1000 -2519
rect 1002 -2527 1004 -2519
rect 1008 -2527 1010 -2519
rect 1012 -2527 1013 -2519
rect 1017 -2527 1018 -2519
rect 1020 -2527 1025 -2519
rect 1029 -2527 1034 -2519
rect 1036 -2527 1037 -2519
rect 1041 -2527 1042 -2519
rect 1044 -2527 1045 -2519
rect 1215 -2527 1216 -2519
rect 1218 -2527 1220 -2519
rect 1224 -2527 1226 -2519
rect 1228 -2527 1229 -2519
rect 1241 -2527 1242 -2519
rect 1244 -2527 1245 -2519
rect 1249 -2527 1250 -2519
rect 1252 -2527 1257 -2519
rect 1261 -2527 1266 -2519
rect 1268 -2527 1269 -2519
rect 1273 -2527 1274 -2519
rect 1276 -2527 1278 -2519
rect 1282 -2527 1284 -2519
rect 1286 -2527 1287 -2519
rect 1291 -2527 1292 -2519
rect 1294 -2527 1299 -2519
rect 1303 -2527 1308 -2519
rect 1310 -2527 1311 -2519
rect 1315 -2527 1316 -2519
rect 1318 -2527 1320 -2519
rect 1324 -2527 1326 -2519
rect 1328 -2527 1329 -2519
rect 1333 -2527 1334 -2519
rect 1336 -2527 1341 -2519
rect 1345 -2527 1350 -2519
rect 1352 -2527 1353 -2519
rect 1357 -2527 1358 -2519
rect 1360 -2527 1362 -2519
rect 1366 -2527 1368 -2519
rect 1370 -2527 1371 -2519
rect 1375 -2527 1376 -2519
rect 1378 -2527 1383 -2519
rect 1387 -2527 1392 -2519
rect 1394 -2527 1395 -2519
rect 1399 -2527 1400 -2519
rect 1402 -2527 1403 -2519
rect -1305 -2632 -1304 -2624
rect -1302 -2632 -1301 -2624
rect -1297 -2632 -1296 -2624
rect -1294 -2632 -1292 -2624
rect -1288 -2632 -1286 -2624
rect -1284 -2632 -1283 -2624
rect -931 -2632 -930 -2624
rect -928 -2632 -927 -2624
rect -923 -2632 -922 -2624
rect -920 -2632 -918 -2624
rect -914 -2632 -912 -2624
rect -910 -2632 -909 -2624
rect -573 -2632 -572 -2624
rect -570 -2632 -569 -2624
rect -565 -2632 -564 -2624
rect -562 -2632 -560 -2624
rect -556 -2632 -554 -2624
rect -552 -2632 -551 -2624
rect -215 -2632 -214 -2624
rect -212 -2632 -211 -2624
rect -207 -2632 -206 -2624
rect -204 -2632 -202 -2624
rect -198 -2632 -196 -2624
rect -194 -2632 -193 -2624
rect 143 -2632 144 -2624
rect 146 -2632 147 -2624
rect 151 -2632 152 -2624
rect 154 -2632 156 -2624
rect 160 -2632 162 -2624
rect 164 -2632 165 -2624
rect 499 -2632 500 -2624
rect 502 -2632 503 -2624
rect 507 -2632 508 -2624
rect 510 -2632 512 -2624
rect 516 -2632 518 -2624
rect 520 -2632 521 -2624
rect 857 -2632 858 -2624
rect 860 -2632 861 -2624
rect 865 -2632 866 -2624
rect 868 -2632 870 -2624
rect 874 -2632 876 -2624
rect 878 -2632 879 -2624
rect 1215 -2632 1216 -2624
rect 1218 -2632 1219 -2624
rect 1223 -2632 1224 -2624
rect 1226 -2632 1228 -2624
rect 1232 -2632 1234 -2624
rect 1236 -2632 1237 -2624
rect -1230 -2791 -1229 -2783
rect -1227 -2791 -1225 -2783
rect -1221 -2791 -1219 -2783
rect -1217 -2791 -1216 -2783
rect -1204 -2791 -1203 -2783
rect -1201 -2791 -1193 -2783
rect -1191 -2791 -1190 -2783
rect -1186 -2791 -1185 -2783
rect -1183 -2791 -1175 -2783
rect -1173 -2791 -1168 -2783
rect -1164 -2791 -1159 -2783
rect -1157 -2791 -1156 -2783
rect -1152 -2791 -1151 -2783
rect -1149 -2791 -1147 -2783
rect -1143 -2791 -1141 -2783
rect -1139 -2791 -1138 -2783
rect -931 -2791 -930 -2783
rect -928 -2791 -926 -2783
rect -922 -2791 -920 -2783
rect -918 -2791 -917 -2783
rect -905 -2791 -904 -2783
rect -902 -2791 -900 -2783
rect -896 -2791 -894 -2783
rect -892 -2791 -891 -2783
rect -879 -2791 -878 -2783
rect -876 -2791 -868 -2783
rect -866 -2791 -865 -2783
rect -861 -2791 -860 -2783
rect -858 -2791 -850 -2783
rect -848 -2791 -843 -2783
rect -839 -2791 -834 -2783
rect -832 -2791 -831 -2783
rect -827 -2791 -826 -2783
rect -824 -2791 -822 -2783
rect -818 -2791 -816 -2783
rect -814 -2791 -813 -2783
rect -801 -2791 -800 -2783
rect -798 -2791 -790 -2783
rect -788 -2791 -787 -2783
rect -783 -2791 -782 -2783
rect -780 -2791 -772 -2783
rect -770 -2791 -765 -2783
rect -761 -2791 -756 -2783
rect -754 -2791 -753 -2783
rect -749 -2791 -748 -2783
rect -746 -2791 -741 -2783
rect -737 -2791 -732 -2783
rect -730 -2791 -729 -2783
rect -717 -2791 -716 -2783
rect -714 -2791 -708 -2783
rect -706 -2791 -704 -2783
rect -700 -2791 -698 -2783
rect -696 -2791 -695 -2783
rect -573 -2791 -572 -2783
rect -570 -2791 -568 -2783
rect -564 -2791 -562 -2783
rect -560 -2791 -559 -2783
rect -547 -2791 -546 -2783
rect -544 -2791 -542 -2783
rect -538 -2791 -536 -2783
rect -534 -2791 -533 -2783
rect -521 -2791 -520 -2783
rect -518 -2791 -510 -2783
rect -508 -2791 -507 -2783
rect -503 -2791 -502 -2783
rect -500 -2791 -492 -2783
rect -490 -2791 -485 -2783
rect -481 -2791 -476 -2783
rect -474 -2791 -473 -2783
rect -469 -2791 -468 -2783
rect -466 -2791 -464 -2783
rect -460 -2791 -458 -2783
rect -456 -2791 -455 -2783
rect -443 -2791 -442 -2783
rect -440 -2791 -432 -2783
rect -430 -2791 -429 -2783
rect -425 -2791 -424 -2783
rect -422 -2791 -414 -2783
rect -412 -2791 -407 -2783
rect -403 -2791 -398 -2783
rect -396 -2791 -395 -2783
rect -391 -2791 -390 -2783
rect -388 -2791 -383 -2783
rect -379 -2791 -374 -2783
rect -372 -2791 -371 -2783
rect -359 -2791 -358 -2783
rect -356 -2791 -350 -2783
rect -348 -2791 -346 -2783
rect -342 -2791 -340 -2783
rect -338 -2791 -337 -2783
rect -215 -2791 -214 -2783
rect -212 -2791 -210 -2783
rect -206 -2791 -204 -2783
rect -202 -2791 -201 -2783
rect -189 -2791 -188 -2783
rect -186 -2791 -184 -2783
rect -180 -2791 -178 -2783
rect -176 -2791 -175 -2783
rect -163 -2791 -162 -2783
rect -160 -2791 -152 -2783
rect -150 -2791 -149 -2783
rect -145 -2791 -144 -2783
rect -142 -2791 -134 -2783
rect -132 -2791 -127 -2783
rect -123 -2791 -118 -2783
rect -116 -2791 -115 -2783
rect -111 -2791 -110 -2783
rect -108 -2791 -106 -2783
rect -102 -2791 -100 -2783
rect -98 -2791 -97 -2783
rect -85 -2791 -84 -2783
rect -82 -2791 -74 -2783
rect -72 -2791 -71 -2783
rect -67 -2791 -66 -2783
rect -64 -2791 -56 -2783
rect -54 -2791 -49 -2783
rect -45 -2791 -40 -2783
rect -38 -2791 -37 -2783
rect -33 -2791 -32 -2783
rect -30 -2791 -25 -2783
rect -21 -2791 -16 -2783
rect -14 -2791 -13 -2783
rect -1 -2791 0 -2783
rect 2 -2791 8 -2783
rect 10 -2791 12 -2783
rect 16 -2791 18 -2783
rect 20 -2791 21 -2783
rect 143 -2791 144 -2783
rect 146 -2791 148 -2783
rect 152 -2791 154 -2783
rect 156 -2791 157 -2783
rect 169 -2791 170 -2783
rect 172 -2791 174 -2783
rect 178 -2791 180 -2783
rect 182 -2791 183 -2783
rect 195 -2791 196 -2783
rect 198 -2791 206 -2783
rect 208 -2791 209 -2783
rect 213 -2791 214 -2783
rect 216 -2791 224 -2783
rect 226 -2791 231 -2783
rect 235 -2791 240 -2783
rect 242 -2791 243 -2783
rect 247 -2791 248 -2783
rect 250 -2791 252 -2783
rect 256 -2791 258 -2783
rect 260 -2791 261 -2783
rect 273 -2791 274 -2783
rect 276 -2791 284 -2783
rect 286 -2791 287 -2783
rect 291 -2791 292 -2783
rect 294 -2791 302 -2783
rect 304 -2791 309 -2783
rect 313 -2791 318 -2783
rect 320 -2791 321 -2783
rect 325 -2791 326 -2783
rect 328 -2791 333 -2783
rect 337 -2791 342 -2783
rect 344 -2791 345 -2783
rect 357 -2791 358 -2783
rect 360 -2791 366 -2783
rect 368 -2791 370 -2783
rect 374 -2791 376 -2783
rect 378 -2791 379 -2783
rect 499 -2791 500 -2783
rect 502 -2791 504 -2783
rect 508 -2791 510 -2783
rect 512 -2791 513 -2783
rect 525 -2791 526 -2783
rect 528 -2791 530 -2783
rect 534 -2791 536 -2783
rect 538 -2791 539 -2783
rect 551 -2791 552 -2783
rect 554 -2791 562 -2783
rect 564 -2791 565 -2783
rect 569 -2791 570 -2783
rect 572 -2791 580 -2783
rect 582 -2791 587 -2783
rect 591 -2791 596 -2783
rect 598 -2791 599 -2783
rect 603 -2791 604 -2783
rect 606 -2791 608 -2783
rect 612 -2791 614 -2783
rect 616 -2791 617 -2783
rect 629 -2791 630 -2783
rect 632 -2791 640 -2783
rect 642 -2791 643 -2783
rect 647 -2791 648 -2783
rect 650 -2791 658 -2783
rect 660 -2791 665 -2783
rect 669 -2791 674 -2783
rect 676 -2791 677 -2783
rect 681 -2791 682 -2783
rect 684 -2791 689 -2783
rect 693 -2791 698 -2783
rect 700 -2791 701 -2783
rect 713 -2791 714 -2783
rect 716 -2791 722 -2783
rect 724 -2791 726 -2783
rect 730 -2791 732 -2783
rect 734 -2791 735 -2783
rect 857 -2791 858 -2783
rect 860 -2791 862 -2783
rect 866 -2791 868 -2783
rect 870 -2791 871 -2783
rect 883 -2791 884 -2783
rect 886 -2791 888 -2783
rect 892 -2791 894 -2783
rect 896 -2791 897 -2783
rect 909 -2791 910 -2783
rect 912 -2791 920 -2783
rect 922 -2791 923 -2783
rect 927 -2791 928 -2783
rect 930 -2791 938 -2783
rect 940 -2791 945 -2783
rect 949 -2791 954 -2783
rect 956 -2791 957 -2783
rect 961 -2791 962 -2783
rect 964 -2791 966 -2783
rect 970 -2791 972 -2783
rect 974 -2791 975 -2783
rect 987 -2791 988 -2783
rect 990 -2791 998 -2783
rect 1000 -2791 1001 -2783
rect 1005 -2791 1006 -2783
rect 1008 -2791 1016 -2783
rect 1018 -2791 1023 -2783
rect 1027 -2791 1032 -2783
rect 1034 -2791 1035 -2783
rect 1039 -2791 1040 -2783
rect 1042 -2791 1047 -2783
rect 1051 -2791 1056 -2783
rect 1058 -2791 1059 -2783
rect 1071 -2791 1072 -2783
rect 1074 -2791 1080 -2783
rect 1082 -2791 1084 -2783
rect 1088 -2791 1090 -2783
rect 1092 -2791 1093 -2783
rect 1215 -2791 1216 -2783
rect 1218 -2791 1220 -2783
rect 1224 -2791 1226 -2783
rect 1228 -2791 1229 -2783
rect 1241 -2791 1242 -2783
rect 1244 -2791 1246 -2783
rect 1250 -2791 1252 -2783
rect 1254 -2791 1255 -2783
rect 1267 -2791 1268 -2783
rect 1270 -2791 1278 -2783
rect 1280 -2791 1281 -2783
rect 1285 -2791 1286 -2783
rect 1288 -2791 1296 -2783
rect 1298 -2791 1303 -2783
rect 1307 -2791 1312 -2783
rect 1314 -2791 1315 -2783
rect 1319 -2791 1320 -2783
rect 1322 -2791 1324 -2783
rect 1328 -2791 1330 -2783
rect 1332 -2791 1333 -2783
rect 1345 -2791 1346 -2783
rect 1348 -2791 1356 -2783
rect 1358 -2791 1359 -2783
rect 1363 -2791 1364 -2783
rect 1366 -2791 1374 -2783
rect 1376 -2791 1381 -2783
rect 1385 -2791 1390 -2783
rect 1392 -2791 1393 -2783
rect 1397 -2791 1398 -2783
rect 1400 -2791 1405 -2783
rect 1409 -2791 1414 -2783
rect 1416 -2791 1417 -2783
rect 1429 -2791 1430 -2783
rect 1432 -2791 1438 -2783
rect 1440 -2791 1442 -2783
rect 1446 -2791 1448 -2783
rect 1450 -2791 1451 -2783
rect -1555 -2910 -1554 -2902
rect -1552 -2910 -1550 -2902
rect -1546 -2910 -1544 -2902
rect -1542 -2910 -1541 -2902
rect -1529 -2910 -1528 -2902
rect -1526 -2910 -1525 -2902
rect -1521 -2910 -1520 -2902
rect -1518 -2910 -1513 -2902
rect -1509 -2910 -1504 -2902
rect -1502 -2910 -1501 -2902
rect -1497 -2910 -1496 -2902
rect -1494 -2910 -1492 -2902
rect -1488 -2910 -1486 -2902
rect -1484 -2910 -1483 -2902
rect -1479 -2910 -1478 -2902
rect -1476 -2910 -1471 -2902
rect -1467 -2910 -1462 -2902
rect -1460 -2910 -1459 -2902
rect -1455 -2910 -1454 -2902
rect -1452 -2910 -1450 -2902
rect -1446 -2910 -1444 -2902
rect -1442 -2910 -1441 -2902
rect -1437 -2910 -1436 -2902
rect -1434 -2910 -1429 -2902
rect -1425 -2910 -1420 -2902
rect -1418 -2910 -1417 -2902
rect -1413 -2910 -1412 -2902
rect -1410 -2910 -1408 -2902
rect -1404 -2910 -1402 -2902
rect -1400 -2910 -1399 -2902
rect -1395 -2910 -1394 -2902
rect -1392 -2910 -1387 -2902
rect -1383 -2910 -1378 -2902
rect -1376 -2910 -1375 -2902
rect -1371 -2910 -1370 -2902
rect -1368 -2910 -1367 -2902
rect -1230 -2910 -1229 -2902
rect -1227 -2910 -1225 -2902
rect -1221 -2910 -1219 -2902
rect -1217 -2910 -1216 -2902
rect -1204 -2910 -1203 -2902
rect -1201 -2910 -1200 -2902
rect -1196 -2910 -1195 -2902
rect -1193 -2910 -1188 -2902
rect -1184 -2910 -1179 -2902
rect -1177 -2910 -1176 -2902
rect -1172 -2910 -1171 -2902
rect -1169 -2910 -1167 -2902
rect -1163 -2910 -1161 -2902
rect -1159 -2910 -1158 -2902
rect -1154 -2910 -1153 -2902
rect -1151 -2910 -1146 -2902
rect -1142 -2910 -1137 -2902
rect -1135 -2910 -1134 -2902
rect -1130 -2910 -1129 -2902
rect -1127 -2910 -1125 -2902
rect -1121 -2910 -1119 -2902
rect -1117 -2910 -1116 -2902
rect -1112 -2910 -1111 -2902
rect -1109 -2910 -1104 -2902
rect -1100 -2910 -1095 -2902
rect -1093 -2910 -1092 -2902
rect -1088 -2910 -1087 -2902
rect -1085 -2910 -1083 -2902
rect -1079 -2910 -1077 -2902
rect -1075 -2910 -1074 -2902
rect -1070 -2910 -1069 -2902
rect -1067 -2910 -1062 -2902
rect -1058 -2910 -1053 -2902
rect -1051 -2910 -1050 -2902
rect -1046 -2910 -1045 -2902
rect -1043 -2910 -1042 -2902
rect -931 -2910 -930 -2902
rect -928 -2910 -926 -2902
rect -922 -2910 -920 -2902
rect -918 -2910 -917 -2902
rect -905 -2910 -904 -2902
rect -902 -2910 -901 -2902
rect -897 -2910 -896 -2902
rect -894 -2910 -889 -2902
rect -885 -2910 -880 -2902
rect -878 -2910 -877 -2902
rect -873 -2910 -872 -2902
rect -870 -2910 -868 -2902
rect -864 -2910 -862 -2902
rect -860 -2910 -859 -2902
rect -855 -2910 -854 -2902
rect -852 -2910 -847 -2902
rect -843 -2910 -838 -2902
rect -836 -2910 -835 -2902
rect -831 -2910 -830 -2902
rect -828 -2910 -826 -2902
rect -822 -2910 -820 -2902
rect -818 -2910 -817 -2902
rect -813 -2910 -812 -2902
rect -810 -2910 -805 -2902
rect -801 -2910 -796 -2902
rect -794 -2910 -793 -2902
rect -789 -2910 -788 -2902
rect -786 -2910 -784 -2902
rect -780 -2910 -778 -2902
rect -776 -2910 -775 -2902
rect -771 -2910 -770 -2902
rect -768 -2910 -763 -2902
rect -759 -2910 -754 -2902
rect -752 -2910 -751 -2902
rect -747 -2910 -746 -2902
rect -744 -2910 -743 -2902
rect -573 -2910 -572 -2902
rect -570 -2910 -568 -2902
rect -564 -2910 -562 -2902
rect -560 -2910 -559 -2902
rect -547 -2910 -546 -2902
rect -544 -2910 -543 -2902
rect -539 -2910 -538 -2902
rect -536 -2910 -531 -2902
rect -527 -2910 -522 -2902
rect -520 -2910 -519 -2902
rect -515 -2910 -514 -2902
rect -512 -2910 -510 -2902
rect -506 -2910 -504 -2902
rect -502 -2910 -501 -2902
rect -497 -2910 -496 -2902
rect -494 -2910 -489 -2902
rect -485 -2910 -480 -2902
rect -478 -2910 -477 -2902
rect -473 -2910 -472 -2902
rect -470 -2910 -468 -2902
rect -464 -2910 -462 -2902
rect -460 -2910 -459 -2902
rect -455 -2910 -454 -2902
rect -452 -2910 -447 -2902
rect -443 -2910 -438 -2902
rect -436 -2910 -435 -2902
rect -431 -2910 -430 -2902
rect -428 -2910 -426 -2902
rect -422 -2910 -420 -2902
rect -418 -2910 -417 -2902
rect -413 -2910 -412 -2902
rect -410 -2910 -405 -2902
rect -401 -2910 -396 -2902
rect -394 -2910 -393 -2902
rect -389 -2910 -388 -2902
rect -386 -2910 -385 -2902
rect -215 -2910 -214 -2902
rect -212 -2910 -210 -2902
rect -206 -2910 -204 -2902
rect -202 -2910 -201 -2902
rect -189 -2910 -188 -2902
rect -186 -2910 -185 -2902
rect -181 -2910 -180 -2902
rect -178 -2910 -173 -2902
rect -169 -2910 -164 -2902
rect -162 -2910 -161 -2902
rect -157 -2910 -156 -2902
rect -154 -2910 -152 -2902
rect -148 -2910 -146 -2902
rect -144 -2910 -143 -2902
rect -139 -2910 -138 -2902
rect -136 -2910 -131 -2902
rect -127 -2910 -122 -2902
rect -120 -2910 -119 -2902
rect -115 -2910 -114 -2902
rect -112 -2910 -110 -2902
rect -106 -2910 -104 -2902
rect -102 -2910 -101 -2902
rect -97 -2910 -96 -2902
rect -94 -2910 -89 -2902
rect -85 -2910 -80 -2902
rect -78 -2910 -77 -2902
rect -73 -2910 -72 -2902
rect -70 -2910 -68 -2902
rect -64 -2910 -62 -2902
rect -60 -2910 -59 -2902
rect -55 -2910 -54 -2902
rect -52 -2910 -47 -2902
rect -43 -2910 -38 -2902
rect -36 -2910 -35 -2902
rect -31 -2910 -30 -2902
rect -28 -2910 -27 -2902
rect 143 -2910 144 -2902
rect 146 -2910 148 -2902
rect 152 -2910 154 -2902
rect 156 -2910 157 -2902
rect 169 -2910 170 -2902
rect 172 -2910 173 -2902
rect 177 -2910 178 -2902
rect 180 -2910 185 -2902
rect 189 -2910 194 -2902
rect 196 -2910 197 -2902
rect 201 -2910 202 -2902
rect 204 -2910 206 -2902
rect 210 -2910 212 -2902
rect 214 -2910 215 -2902
rect 219 -2910 220 -2902
rect 222 -2910 227 -2902
rect 231 -2910 236 -2902
rect 238 -2910 239 -2902
rect 243 -2910 244 -2902
rect 246 -2910 248 -2902
rect 252 -2910 254 -2902
rect 256 -2910 257 -2902
rect 261 -2910 262 -2902
rect 264 -2910 269 -2902
rect 273 -2910 278 -2902
rect 280 -2910 281 -2902
rect 285 -2910 286 -2902
rect 288 -2910 290 -2902
rect 294 -2910 296 -2902
rect 298 -2910 299 -2902
rect 303 -2910 304 -2902
rect 306 -2910 311 -2902
rect 315 -2910 320 -2902
rect 322 -2910 323 -2902
rect 327 -2910 328 -2902
rect 330 -2910 331 -2902
rect -1555 -3081 -1554 -3073
rect -1552 -3081 -1550 -3073
rect -1546 -3081 -1544 -3073
rect -1542 -3081 -1541 -3073
rect -1529 -3081 -1528 -3073
rect -1526 -3081 -1525 -3073
rect -1521 -3081 -1520 -3073
rect -1518 -3081 -1513 -3073
rect -1509 -3081 -1504 -3073
rect -1502 -3081 -1501 -3073
rect -1497 -3081 -1496 -3073
rect -1494 -3081 -1492 -3073
rect -1488 -3081 -1486 -3073
rect -1484 -3081 -1483 -3073
rect -1479 -3081 -1478 -3073
rect -1476 -3081 -1471 -3073
rect -1467 -3081 -1462 -3073
rect -1460 -3081 -1459 -3073
rect -1455 -3081 -1454 -3073
rect -1452 -3081 -1450 -3073
rect -1446 -3081 -1444 -3073
rect -1442 -3081 -1441 -3073
rect -1437 -3081 -1436 -3073
rect -1434 -3081 -1429 -3073
rect -1425 -3081 -1420 -3073
rect -1418 -3081 -1417 -3073
rect -1413 -3081 -1412 -3073
rect -1410 -3081 -1408 -3073
rect -1404 -3081 -1402 -3073
rect -1400 -3081 -1399 -3073
rect -1395 -3081 -1394 -3073
rect -1392 -3081 -1387 -3073
rect -1383 -3081 -1378 -3073
rect -1376 -3081 -1375 -3073
rect -1371 -3081 -1370 -3073
rect -1368 -3081 -1367 -3073
rect -1230 -3081 -1229 -3073
rect -1227 -3081 -1225 -3073
rect -1221 -3081 -1219 -3073
rect -1217 -3081 -1216 -3073
rect -1204 -3081 -1203 -3073
rect -1201 -3081 -1200 -3073
rect -1196 -3081 -1195 -3073
rect -1193 -3081 -1188 -3073
rect -1184 -3081 -1179 -3073
rect -1177 -3081 -1176 -3073
rect -1172 -3081 -1171 -3073
rect -1169 -3081 -1167 -3073
rect -1163 -3081 -1161 -3073
rect -1159 -3081 -1158 -3073
rect -1154 -3081 -1153 -3073
rect -1151 -3081 -1146 -3073
rect -1142 -3081 -1137 -3073
rect -1135 -3081 -1134 -3073
rect -1130 -3081 -1129 -3073
rect -1127 -3081 -1125 -3073
rect -1121 -3081 -1119 -3073
rect -1117 -3081 -1116 -3073
rect -1112 -3081 -1111 -3073
rect -1109 -3081 -1104 -3073
rect -1100 -3081 -1095 -3073
rect -1093 -3081 -1092 -3073
rect -1088 -3081 -1087 -3073
rect -1085 -3081 -1083 -3073
rect -1079 -3081 -1077 -3073
rect -1075 -3081 -1074 -3073
rect -1070 -3081 -1069 -3073
rect -1067 -3081 -1062 -3073
rect -1058 -3081 -1053 -3073
rect -1051 -3081 -1050 -3073
rect -1046 -3081 -1045 -3073
rect -1043 -3081 -1042 -3073
rect -931 -3081 -930 -3073
rect -928 -3081 -926 -3073
rect -922 -3081 -920 -3073
rect -918 -3081 -917 -3073
rect -905 -3081 -904 -3073
rect -902 -3081 -901 -3073
rect -897 -3081 -896 -3073
rect -894 -3081 -889 -3073
rect -885 -3081 -880 -3073
rect -878 -3081 -877 -3073
rect -873 -3081 -872 -3073
rect -870 -3081 -868 -3073
rect -864 -3081 -862 -3073
rect -860 -3081 -859 -3073
rect -855 -3081 -854 -3073
rect -852 -3081 -847 -3073
rect -843 -3081 -838 -3073
rect -836 -3081 -835 -3073
rect -831 -3081 -830 -3073
rect -828 -3081 -826 -3073
rect -822 -3081 -820 -3073
rect -818 -3081 -817 -3073
rect -813 -3081 -812 -3073
rect -810 -3081 -805 -3073
rect -801 -3081 -796 -3073
rect -794 -3081 -793 -3073
rect -789 -3081 -788 -3073
rect -786 -3081 -784 -3073
rect -780 -3081 -778 -3073
rect -776 -3081 -775 -3073
rect -771 -3081 -770 -3073
rect -768 -3081 -763 -3073
rect -759 -3081 -754 -3073
rect -752 -3081 -751 -3073
rect -747 -3081 -746 -3073
rect -744 -3081 -743 -3073
rect -573 -3081 -572 -3073
rect -570 -3081 -568 -3073
rect -564 -3081 -562 -3073
rect -560 -3081 -559 -3073
rect -547 -3081 -546 -3073
rect -544 -3081 -543 -3073
rect -539 -3081 -538 -3073
rect -536 -3081 -531 -3073
rect -527 -3081 -522 -3073
rect -520 -3081 -519 -3073
rect -515 -3081 -514 -3073
rect -512 -3081 -510 -3073
rect -506 -3081 -504 -3073
rect -502 -3081 -501 -3073
rect -497 -3081 -496 -3073
rect -494 -3081 -489 -3073
rect -485 -3081 -480 -3073
rect -478 -3081 -477 -3073
rect -473 -3081 -472 -3073
rect -470 -3081 -468 -3073
rect -464 -3081 -462 -3073
rect -460 -3081 -459 -3073
rect -455 -3081 -454 -3073
rect -452 -3081 -447 -3073
rect -443 -3081 -438 -3073
rect -436 -3081 -435 -3073
rect -431 -3081 -430 -3073
rect -428 -3081 -426 -3073
rect -422 -3081 -420 -3073
rect -418 -3081 -417 -3073
rect -413 -3081 -412 -3073
rect -410 -3081 -405 -3073
rect -401 -3081 -396 -3073
rect -394 -3081 -393 -3073
rect -389 -3081 -388 -3073
rect -386 -3081 -385 -3073
rect -215 -3081 -214 -3073
rect -212 -3081 -210 -3073
rect -206 -3081 -204 -3073
rect -202 -3081 -201 -3073
rect -189 -3081 -188 -3073
rect -186 -3081 -185 -3073
rect -181 -3081 -180 -3073
rect -178 -3081 -173 -3073
rect -169 -3081 -164 -3073
rect -162 -3081 -161 -3073
rect -157 -3081 -156 -3073
rect -154 -3081 -152 -3073
rect -148 -3081 -146 -3073
rect -144 -3081 -143 -3073
rect -139 -3081 -138 -3073
rect -136 -3081 -131 -3073
rect -127 -3081 -122 -3073
rect -120 -3081 -119 -3073
rect -115 -3081 -114 -3073
rect -112 -3081 -110 -3073
rect -106 -3081 -104 -3073
rect -102 -3081 -101 -3073
rect -97 -3081 -96 -3073
rect -94 -3081 -89 -3073
rect -85 -3081 -80 -3073
rect -78 -3081 -77 -3073
rect -73 -3081 -72 -3073
rect -70 -3081 -68 -3073
rect -64 -3081 -62 -3073
rect -60 -3081 -59 -3073
rect -55 -3081 -54 -3073
rect -52 -3081 -47 -3073
rect -43 -3081 -38 -3073
rect -36 -3081 -35 -3073
rect -31 -3081 -30 -3073
rect -28 -3081 -27 -3073
rect 143 -3081 144 -3073
rect 146 -3081 148 -3073
rect 152 -3081 154 -3073
rect 156 -3081 157 -3073
rect 169 -3081 170 -3073
rect 172 -3081 173 -3073
rect 177 -3081 178 -3073
rect 180 -3081 185 -3073
rect 189 -3081 194 -3073
rect 196 -3081 197 -3073
rect 201 -3081 202 -3073
rect 204 -3081 206 -3073
rect 210 -3081 212 -3073
rect 214 -3081 215 -3073
rect 219 -3081 220 -3073
rect 222 -3081 227 -3073
rect 231 -3081 236 -3073
rect 238 -3081 239 -3073
rect 243 -3081 244 -3073
rect 246 -3081 248 -3073
rect 252 -3081 254 -3073
rect 256 -3081 257 -3073
rect 261 -3081 262 -3073
rect 264 -3081 269 -3073
rect 273 -3081 278 -3073
rect 280 -3081 281 -3073
rect 285 -3081 286 -3073
rect 288 -3081 290 -3073
rect 294 -3081 296 -3073
rect 298 -3081 299 -3073
rect 303 -3081 304 -3073
rect 306 -3081 311 -3073
rect 315 -3081 320 -3073
rect 322 -3081 323 -3073
rect 327 -3081 328 -3073
rect 330 -3081 331 -3073
rect 499 -3081 500 -3073
rect 502 -3081 504 -3073
rect 508 -3081 510 -3073
rect 512 -3081 513 -3073
rect 525 -3081 526 -3073
rect 528 -3081 529 -3073
rect 533 -3081 534 -3073
rect 536 -3081 541 -3073
rect 545 -3081 550 -3073
rect 552 -3081 553 -3073
rect 557 -3081 558 -3073
rect 560 -3081 562 -3073
rect 566 -3081 568 -3073
rect 570 -3081 571 -3073
rect 575 -3081 576 -3073
rect 578 -3081 583 -3073
rect 587 -3081 592 -3073
rect 594 -3081 595 -3073
rect 599 -3081 600 -3073
rect 602 -3081 604 -3073
rect 608 -3081 610 -3073
rect 612 -3081 613 -3073
rect 617 -3081 618 -3073
rect 620 -3081 625 -3073
rect 629 -3081 634 -3073
rect 636 -3081 637 -3073
rect 641 -3081 642 -3073
rect 644 -3081 646 -3073
rect 650 -3081 652 -3073
rect 654 -3081 655 -3073
rect 659 -3081 660 -3073
rect 662 -3081 667 -3073
rect 671 -3081 676 -3073
rect 678 -3081 679 -3073
rect 683 -3081 684 -3073
rect 686 -3081 687 -3073
rect 857 -3081 858 -3073
rect 860 -3081 862 -3073
rect 866 -3081 868 -3073
rect 870 -3081 871 -3073
rect 883 -3081 884 -3073
rect 886 -3081 887 -3073
rect 891 -3081 892 -3073
rect 894 -3081 899 -3073
rect 903 -3081 908 -3073
rect 910 -3081 911 -3073
rect 915 -3081 916 -3073
rect 918 -3081 920 -3073
rect 924 -3081 926 -3073
rect 928 -3081 929 -3073
rect 933 -3081 934 -3073
rect 936 -3081 941 -3073
rect 945 -3081 950 -3073
rect 952 -3081 953 -3073
rect 957 -3081 958 -3073
rect 960 -3081 962 -3073
rect 966 -3081 968 -3073
rect 970 -3081 971 -3073
rect 975 -3081 976 -3073
rect 978 -3081 983 -3073
rect 987 -3081 992 -3073
rect 994 -3081 995 -3073
rect 999 -3081 1000 -3073
rect 1002 -3081 1004 -3073
rect 1008 -3081 1010 -3073
rect 1012 -3081 1013 -3073
rect 1017 -3081 1018 -3073
rect 1020 -3081 1025 -3073
rect 1029 -3081 1034 -3073
rect 1036 -3081 1037 -3073
rect 1041 -3081 1042 -3073
rect 1044 -3081 1045 -3073
rect 1215 -3081 1216 -3073
rect 1218 -3081 1220 -3073
rect 1224 -3081 1226 -3073
rect 1228 -3081 1229 -3073
rect 1241 -3081 1242 -3073
rect 1244 -3081 1245 -3073
rect 1249 -3081 1250 -3073
rect 1252 -3081 1257 -3073
rect 1261 -3081 1266 -3073
rect 1268 -3081 1269 -3073
rect 1273 -3081 1274 -3073
rect 1276 -3081 1278 -3073
rect 1282 -3081 1284 -3073
rect 1286 -3081 1287 -3073
rect 1291 -3081 1292 -3073
rect 1294 -3081 1299 -3073
rect 1303 -3081 1308 -3073
rect 1310 -3081 1311 -3073
rect 1315 -3081 1316 -3073
rect 1318 -3081 1320 -3073
rect 1324 -3081 1326 -3073
rect 1328 -3081 1329 -3073
rect 1333 -3081 1334 -3073
rect 1336 -3081 1341 -3073
rect 1345 -3081 1350 -3073
rect 1352 -3081 1353 -3073
rect 1357 -3081 1358 -3073
rect 1360 -3081 1362 -3073
rect 1366 -3081 1368 -3073
rect 1370 -3081 1371 -3073
rect 1375 -3081 1376 -3073
rect 1378 -3081 1383 -3073
rect 1387 -3081 1392 -3073
rect 1394 -3081 1395 -3073
rect 1399 -3081 1400 -3073
rect 1402 -3081 1403 -3073
rect -1555 -3252 -1554 -3244
rect -1552 -3252 -1550 -3244
rect -1546 -3252 -1544 -3244
rect -1542 -3252 -1541 -3244
rect -1529 -3252 -1528 -3244
rect -1526 -3252 -1525 -3244
rect -1521 -3252 -1520 -3244
rect -1518 -3252 -1513 -3244
rect -1509 -3252 -1504 -3244
rect -1502 -3252 -1501 -3244
rect -1497 -3252 -1496 -3244
rect -1494 -3252 -1492 -3244
rect -1488 -3252 -1486 -3244
rect -1484 -3252 -1483 -3244
rect -1479 -3252 -1478 -3244
rect -1476 -3252 -1471 -3244
rect -1467 -3252 -1462 -3244
rect -1460 -3252 -1459 -3244
rect -1455 -3252 -1454 -3244
rect -1452 -3252 -1450 -3244
rect -1446 -3252 -1444 -3244
rect -1442 -3252 -1441 -3244
rect -1437 -3252 -1436 -3244
rect -1434 -3252 -1429 -3244
rect -1425 -3252 -1420 -3244
rect -1418 -3252 -1417 -3244
rect -1413 -3252 -1412 -3244
rect -1410 -3252 -1408 -3244
rect -1404 -3252 -1402 -3244
rect -1400 -3252 -1399 -3244
rect -1395 -3252 -1394 -3244
rect -1392 -3252 -1387 -3244
rect -1383 -3252 -1378 -3244
rect -1376 -3252 -1375 -3244
rect -1371 -3252 -1370 -3244
rect -1368 -3252 -1367 -3244
rect -1230 -3252 -1229 -3244
rect -1227 -3252 -1225 -3244
rect -1221 -3252 -1219 -3244
rect -1217 -3252 -1216 -3244
rect -1204 -3252 -1203 -3244
rect -1201 -3252 -1200 -3244
rect -1196 -3252 -1195 -3244
rect -1193 -3252 -1188 -3244
rect -1184 -3252 -1179 -3244
rect -1177 -3252 -1176 -3244
rect -1172 -3252 -1171 -3244
rect -1169 -3252 -1167 -3244
rect -1163 -3252 -1161 -3244
rect -1159 -3252 -1158 -3244
rect -1154 -3252 -1153 -3244
rect -1151 -3252 -1146 -3244
rect -1142 -3252 -1137 -3244
rect -1135 -3252 -1134 -3244
rect -1130 -3252 -1129 -3244
rect -1127 -3252 -1125 -3244
rect -1121 -3252 -1119 -3244
rect -1117 -3252 -1116 -3244
rect -1112 -3252 -1111 -3244
rect -1109 -3252 -1104 -3244
rect -1100 -3252 -1095 -3244
rect -1093 -3252 -1092 -3244
rect -1088 -3252 -1087 -3244
rect -1085 -3252 -1083 -3244
rect -1079 -3252 -1077 -3244
rect -1075 -3252 -1074 -3244
rect -1070 -3252 -1069 -3244
rect -1067 -3252 -1062 -3244
rect -1058 -3252 -1053 -3244
rect -1051 -3252 -1050 -3244
rect -1046 -3252 -1045 -3244
rect -1043 -3252 -1042 -3244
rect -931 -3252 -930 -3244
rect -928 -3252 -926 -3244
rect -922 -3252 -920 -3244
rect -918 -3252 -917 -3244
rect -905 -3252 -904 -3244
rect -902 -3252 -901 -3244
rect -897 -3252 -896 -3244
rect -894 -3252 -889 -3244
rect -885 -3252 -880 -3244
rect -878 -3252 -877 -3244
rect -873 -3252 -872 -3244
rect -870 -3252 -868 -3244
rect -864 -3252 -862 -3244
rect -860 -3252 -859 -3244
rect -855 -3252 -854 -3244
rect -852 -3252 -847 -3244
rect -843 -3252 -838 -3244
rect -836 -3252 -835 -3244
rect -831 -3252 -830 -3244
rect -828 -3252 -826 -3244
rect -822 -3252 -820 -3244
rect -818 -3252 -817 -3244
rect -813 -3252 -812 -3244
rect -810 -3252 -805 -3244
rect -801 -3252 -796 -3244
rect -794 -3252 -793 -3244
rect -789 -3252 -788 -3244
rect -786 -3252 -784 -3244
rect -780 -3252 -778 -3244
rect -776 -3252 -775 -3244
rect -771 -3252 -770 -3244
rect -768 -3252 -763 -3244
rect -759 -3252 -754 -3244
rect -752 -3252 -751 -3244
rect -747 -3252 -746 -3244
rect -744 -3252 -743 -3244
rect -573 -3252 -572 -3244
rect -570 -3252 -568 -3244
rect -564 -3252 -562 -3244
rect -560 -3252 -559 -3244
rect -547 -3252 -546 -3244
rect -544 -3252 -543 -3244
rect -539 -3252 -538 -3244
rect -536 -3252 -531 -3244
rect -527 -3252 -522 -3244
rect -520 -3252 -519 -3244
rect -515 -3252 -514 -3244
rect -512 -3252 -510 -3244
rect -506 -3252 -504 -3244
rect -502 -3252 -501 -3244
rect -497 -3252 -496 -3244
rect -494 -3252 -489 -3244
rect -485 -3252 -480 -3244
rect -478 -3252 -477 -3244
rect -473 -3252 -472 -3244
rect -470 -3252 -468 -3244
rect -464 -3252 -462 -3244
rect -460 -3252 -459 -3244
rect -455 -3252 -454 -3244
rect -452 -3252 -447 -3244
rect -443 -3252 -438 -3244
rect -436 -3252 -435 -3244
rect -431 -3252 -430 -3244
rect -428 -3252 -426 -3244
rect -422 -3252 -420 -3244
rect -418 -3252 -417 -3244
rect -413 -3252 -412 -3244
rect -410 -3252 -405 -3244
rect -401 -3252 -396 -3244
rect -394 -3252 -393 -3244
rect -389 -3252 -388 -3244
rect -386 -3252 -385 -3244
rect -215 -3252 -214 -3244
rect -212 -3252 -210 -3244
rect -206 -3252 -204 -3244
rect -202 -3252 -201 -3244
rect -189 -3252 -188 -3244
rect -186 -3252 -185 -3244
rect -181 -3252 -180 -3244
rect -178 -3252 -173 -3244
rect -169 -3252 -164 -3244
rect -162 -3252 -161 -3244
rect -157 -3252 -156 -3244
rect -154 -3252 -152 -3244
rect -148 -3252 -146 -3244
rect -144 -3252 -143 -3244
rect -139 -3252 -138 -3244
rect -136 -3252 -131 -3244
rect -127 -3252 -122 -3244
rect -120 -3252 -119 -3244
rect -115 -3252 -114 -3244
rect -112 -3252 -110 -3244
rect -106 -3252 -104 -3244
rect -102 -3252 -101 -3244
rect -97 -3252 -96 -3244
rect -94 -3252 -89 -3244
rect -85 -3252 -80 -3244
rect -78 -3252 -77 -3244
rect -73 -3252 -72 -3244
rect -70 -3252 -68 -3244
rect -64 -3252 -62 -3244
rect -60 -3252 -59 -3244
rect -55 -3252 -54 -3244
rect -52 -3252 -47 -3244
rect -43 -3252 -38 -3244
rect -36 -3252 -35 -3244
rect -31 -3252 -30 -3244
rect -28 -3252 -27 -3244
rect 143 -3252 144 -3244
rect 146 -3252 148 -3244
rect 152 -3252 154 -3244
rect 156 -3252 157 -3244
rect 169 -3252 170 -3244
rect 172 -3252 173 -3244
rect 177 -3252 178 -3244
rect 180 -3252 185 -3244
rect 189 -3252 194 -3244
rect 196 -3252 197 -3244
rect 201 -3252 202 -3244
rect 204 -3252 206 -3244
rect 210 -3252 212 -3244
rect 214 -3252 215 -3244
rect 219 -3252 220 -3244
rect 222 -3252 227 -3244
rect 231 -3252 236 -3244
rect 238 -3252 239 -3244
rect 243 -3252 244 -3244
rect 246 -3252 248 -3244
rect 252 -3252 254 -3244
rect 256 -3252 257 -3244
rect 261 -3252 262 -3244
rect 264 -3252 269 -3244
rect 273 -3252 278 -3244
rect 280 -3252 281 -3244
rect 285 -3252 286 -3244
rect 288 -3252 290 -3244
rect 294 -3252 296 -3244
rect 298 -3252 299 -3244
rect 303 -3252 304 -3244
rect 306 -3252 311 -3244
rect 315 -3252 320 -3244
rect 322 -3252 323 -3244
rect 327 -3252 328 -3244
rect 330 -3252 331 -3244
rect 499 -3252 500 -3244
rect 502 -3252 504 -3244
rect 508 -3252 510 -3244
rect 512 -3252 513 -3244
rect 525 -3252 526 -3244
rect 528 -3252 529 -3244
rect 533 -3252 534 -3244
rect 536 -3252 541 -3244
rect 545 -3252 550 -3244
rect 552 -3252 553 -3244
rect 557 -3252 558 -3244
rect 560 -3252 562 -3244
rect 566 -3252 568 -3244
rect 570 -3252 571 -3244
rect 575 -3252 576 -3244
rect 578 -3252 583 -3244
rect 587 -3252 592 -3244
rect 594 -3252 595 -3244
rect 599 -3252 600 -3244
rect 602 -3252 604 -3244
rect 608 -3252 610 -3244
rect 612 -3252 613 -3244
rect 617 -3252 618 -3244
rect 620 -3252 625 -3244
rect 629 -3252 634 -3244
rect 636 -3252 637 -3244
rect 641 -3252 642 -3244
rect 644 -3252 646 -3244
rect 650 -3252 652 -3244
rect 654 -3252 655 -3244
rect 659 -3252 660 -3244
rect 662 -3252 667 -3244
rect 671 -3252 676 -3244
rect 678 -3252 679 -3244
rect 683 -3252 684 -3244
rect 686 -3252 687 -3244
rect 857 -3252 858 -3244
rect 860 -3252 862 -3244
rect 866 -3252 868 -3244
rect 870 -3252 871 -3244
rect 883 -3252 884 -3244
rect 886 -3252 887 -3244
rect 891 -3252 892 -3244
rect 894 -3252 899 -3244
rect 903 -3252 908 -3244
rect 910 -3252 911 -3244
rect 915 -3252 916 -3244
rect 918 -3252 920 -3244
rect 924 -3252 926 -3244
rect 928 -3252 929 -3244
rect 933 -3252 934 -3244
rect 936 -3252 941 -3244
rect 945 -3252 950 -3244
rect 952 -3252 953 -3244
rect 957 -3252 958 -3244
rect 960 -3252 962 -3244
rect 966 -3252 968 -3244
rect 970 -3252 971 -3244
rect 975 -3252 976 -3244
rect 978 -3252 983 -3244
rect 987 -3252 992 -3244
rect 994 -3252 995 -3244
rect 999 -3252 1000 -3244
rect 1002 -3252 1004 -3244
rect 1008 -3252 1010 -3244
rect 1012 -3252 1013 -3244
rect 1017 -3252 1018 -3244
rect 1020 -3252 1025 -3244
rect 1029 -3252 1034 -3244
rect 1036 -3252 1037 -3244
rect 1041 -3252 1042 -3244
rect 1044 -3252 1045 -3244
rect 1215 -3252 1216 -3244
rect 1218 -3252 1220 -3244
rect 1224 -3252 1226 -3244
rect 1228 -3252 1229 -3244
rect 1241 -3252 1242 -3244
rect 1244 -3252 1245 -3244
rect 1249 -3252 1250 -3244
rect 1252 -3252 1257 -3244
rect 1261 -3252 1266 -3244
rect 1268 -3252 1269 -3244
rect 1273 -3252 1274 -3244
rect 1276 -3252 1278 -3244
rect 1282 -3252 1284 -3244
rect 1286 -3252 1287 -3244
rect 1291 -3252 1292 -3244
rect 1294 -3252 1299 -3244
rect 1303 -3252 1308 -3244
rect 1310 -3252 1311 -3244
rect 1315 -3252 1316 -3244
rect 1318 -3252 1320 -3244
rect 1324 -3252 1326 -3244
rect 1328 -3252 1329 -3244
rect 1333 -3252 1334 -3244
rect 1336 -3252 1341 -3244
rect 1345 -3252 1350 -3244
rect 1352 -3252 1353 -3244
rect 1357 -3252 1358 -3244
rect 1360 -3252 1362 -3244
rect 1366 -3252 1368 -3244
rect 1370 -3252 1371 -3244
rect 1375 -3252 1376 -3244
rect 1378 -3252 1383 -3244
rect 1387 -3252 1392 -3244
rect 1394 -3252 1395 -3244
rect 1399 -3252 1400 -3244
rect 1402 -3252 1403 -3244
rect -1305 -3363 -1304 -3355
rect -1302 -3363 -1301 -3355
rect -1297 -3363 -1296 -3355
rect -1294 -3363 -1292 -3355
rect -1288 -3363 -1286 -3355
rect -1284 -3363 -1283 -3355
rect -931 -3363 -930 -3355
rect -928 -3363 -927 -3355
rect -923 -3363 -922 -3355
rect -920 -3363 -918 -3355
rect -914 -3363 -912 -3355
rect -910 -3363 -909 -3355
rect -573 -3363 -572 -3355
rect -570 -3363 -569 -3355
rect -565 -3363 -564 -3355
rect -562 -3363 -560 -3355
rect -556 -3363 -554 -3355
rect -552 -3363 -551 -3355
rect -215 -3363 -214 -3355
rect -212 -3363 -211 -3355
rect -207 -3363 -206 -3355
rect -204 -3363 -202 -3355
rect -198 -3363 -196 -3355
rect -194 -3363 -193 -3355
rect 143 -3363 144 -3355
rect 146 -3363 147 -3355
rect 151 -3363 152 -3355
rect 154 -3363 156 -3355
rect 160 -3363 162 -3355
rect 164 -3363 165 -3355
rect 499 -3363 500 -3355
rect 502 -3363 503 -3355
rect 507 -3363 508 -3355
rect 510 -3363 512 -3355
rect 516 -3363 518 -3355
rect 520 -3363 521 -3355
rect 857 -3363 858 -3355
rect 860 -3363 861 -3355
rect 865 -3363 866 -3355
rect 868 -3363 870 -3355
rect 874 -3363 876 -3355
rect 878 -3363 879 -3355
rect 1215 -3363 1216 -3355
rect 1218 -3363 1219 -3355
rect 1223 -3363 1224 -3355
rect 1226 -3363 1228 -3355
rect 1232 -3363 1234 -3355
rect 1236 -3363 1237 -3355
rect -1230 -3522 -1229 -3514
rect -1227 -3522 -1225 -3514
rect -1221 -3522 -1219 -3514
rect -1217 -3522 -1216 -3514
rect -1204 -3522 -1203 -3514
rect -1201 -3522 -1193 -3514
rect -1191 -3522 -1190 -3514
rect -1186 -3522 -1185 -3514
rect -1183 -3522 -1175 -3514
rect -1173 -3522 -1168 -3514
rect -1164 -3522 -1159 -3514
rect -1157 -3522 -1156 -3514
rect -1152 -3522 -1151 -3514
rect -1149 -3522 -1147 -3514
rect -1143 -3522 -1141 -3514
rect -1139 -3522 -1138 -3514
rect -931 -3522 -930 -3514
rect -928 -3522 -926 -3514
rect -922 -3522 -920 -3514
rect -918 -3522 -917 -3514
rect -905 -3522 -904 -3514
rect -902 -3522 -900 -3514
rect -896 -3522 -894 -3514
rect -892 -3522 -891 -3514
rect -879 -3522 -878 -3514
rect -876 -3522 -868 -3514
rect -866 -3522 -865 -3514
rect -861 -3522 -860 -3514
rect -858 -3522 -850 -3514
rect -848 -3522 -843 -3514
rect -839 -3522 -834 -3514
rect -832 -3522 -831 -3514
rect -827 -3522 -826 -3514
rect -824 -3522 -822 -3514
rect -818 -3522 -816 -3514
rect -814 -3522 -813 -3514
rect -801 -3522 -800 -3514
rect -798 -3522 -790 -3514
rect -788 -3522 -787 -3514
rect -783 -3522 -782 -3514
rect -780 -3522 -772 -3514
rect -770 -3522 -765 -3514
rect -761 -3522 -756 -3514
rect -754 -3522 -753 -3514
rect -749 -3522 -748 -3514
rect -746 -3522 -741 -3514
rect -737 -3522 -732 -3514
rect -730 -3522 -729 -3514
rect -717 -3522 -716 -3514
rect -714 -3522 -708 -3514
rect -706 -3522 -704 -3514
rect -700 -3522 -698 -3514
rect -696 -3522 -695 -3514
rect -573 -3522 -572 -3514
rect -570 -3522 -568 -3514
rect -564 -3522 -562 -3514
rect -560 -3522 -559 -3514
rect -547 -3522 -546 -3514
rect -544 -3522 -542 -3514
rect -538 -3522 -536 -3514
rect -534 -3522 -533 -3514
rect -521 -3522 -520 -3514
rect -518 -3522 -510 -3514
rect -508 -3522 -507 -3514
rect -503 -3522 -502 -3514
rect -500 -3522 -492 -3514
rect -490 -3522 -485 -3514
rect -481 -3522 -476 -3514
rect -474 -3522 -473 -3514
rect -469 -3522 -468 -3514
rect -466 -3522 -464 -3514
rect -460 -3522 -458 -3514
rect -456 -3522 -455 -3514
rect -443 -3522 -442 -3514
rect -440 -3522 -432 -3514
rect -430 -3522 -429 -3514
rect -425 -3522 -424 -3514
rect -422 -3522 -414 -3514
rect -412 -3522 -407 -3514
rect -403 -3522 -398 -3514
rect -396 -3522 -395 -3514
rect -391 -3522 -390 -3514
rect -388 -3522 -383 -3514
rect -379 -3522 -374 -3514
rect -372 -3522 -371 -3514
rect -359 -3522 -358 -3514
rect -356 -3522 -350 -3514
rect -348 -3522 -346 -3514
rect -342 -3522 -340 -3514
rect -338 -3522 -337 -3514
rect -215 -3522 -214 -3514
rect -212 -3522 -210 -3514
rect -206 -3522 -204 -3514
rect -202 -3522 -201 -3514
rect -189 -3522 -188 -3514
rect -186 -3522 -184 -3514
rect -180 -3522 -178 -3514
rect -176 -3522 -175 -3514
rect -163 -3522 -162 -3514
rect -160 -3522 -152 -3514
rect -150 -3522 -149 -3514
rect -145 -3522 -144 -3514
rect -142 -3522 -134 -3514
rect -132 -3522 -127 -3514
rect -123 -3522 -118 -3514
rect -116 -3522 -115 -3514
rect -111 -3522 -110 -3514
rect -108 -3522 -106 -3514
rect -102 -3522 -100 -3514
rect -98 -3522 -97 -3514
rect -85 -3522 -84 -3514
rect -82 -3522 -74 -3514
rect -72 -3522 -71 -3514
rect -67 -3522 -66 -3514
rect -64 -3522 -56 -3514
rect -54 -3522 -49 -3514
rect -45 -3522 -40 -3514
rect -38 -3522 -37 -3514
rect -33 -3522 -32 -3514
rect -30 -3522 -25 -3514
rect -21 -3522 -16 -3514
rect -14 -3522 -13 -3514
rect -1 -3522 0 -3514
rect 2 -3522 8 -3514
rect 10 -3522 12 -3514
rect 16 -3522 18 -3514
rect 20 -3522 21 -3514
rect 143 -3522 144 -3514
rect 146 -3522 148 -3514
rect 152 -3522 154 -3514
rect 156 -3522 157 -3514
rect 169 -3522 170 -3514
rect 172 -3522 174 -3514
rect 178 -3522 180 -3514
rect 182 -3522 183 -3514
rect 195 -3522 196 -3514
rect 198 -3522 206 -3514
rect 208 -3522 209 -3514
rect 213 -3522 214 -3514
rect 216 -3522 224 -3514
rect 226 -3522 231 -3514
rect 235 -3522 240 -3514
rect 242 -3522 243 -3514
rect 247 -3522 248 -3514
rect 250 -3522 252 -3514
rect 256 -3522 258 -3514
rect 260 -3522 261 -3514
rect 273 -3522 274 -3514
rect 276 -3522 284 -3514
rect 286 -3522 287 -3514
rect 291 -3522 292 -3514
rect 294 -3522 302 -3514
rect 304 -3522 309 -3514
rect 313 -3522 318 -3514
rect 320 -3522 321 -3514
rect 325 -3522 326 -3514
rect 328 -3522 333 -3514
rect 337 -3522 342 -3514
rect 344 -3522 345 -3514
rect 357 -3522 358 -3514
rect 360 -3522 366 -3514
rect 368 -3522 370 -3514
rect 374 -3522 376 -3514
rect 378 -3522 379 -3514
rect 499 -3522 500 -3514
rect 502 -3522 504 -3514
rect 508 -3522 510 -3514
rect 512 -3522 513 -3514
rect 525 -3522 526 -3514
rect 528 -3522 530 -3514
rect 534 -3522 536 -3514
rect 538 -3522 539 -3514
rect 551 -3522 552 -3514
rect 554 -3522 562 -3514
rect 564 -3522 565 -3514
rect 569 -3522 570 -3514
rect 572 -3522 580 -3514
rect 582 -3522 587 -3514
rect 591 -3522 596 -3514
rect 598 -3522 599 -3514
rect 603 -3522 604 -3514
rect 606 -3522 608 -3514
rect 612 -3522 614 -3514
rect 616 -3522 617 -3514
rect 629 -3522 630 -3514
rect 632 -3522 640 -3514
rect 642 -3522 643 -3514
rect 647 -3522 648 -3514
rect 650 -3522 658 -3514
rect 660 -3522 665 -3514
rect 669 -3522 674 -3514
rect 676 -3522 677 -3514
rect 681 -3522 682 -3514
rect 684 -3522 689 -3514
rect 693 -3522 698 -3514
rect 700 -3522 701 -3514
rect 713 -3522 714 -3514
rect 716 -3522 722 -3514
rect 724 -3522 726 -3514
rect 730 -3522 732 -3514
rect 734 -3522 735 -3514
rect 857 -3522 858 -3514
rect 860 -3522 862 -3514
rect 866 -3522 868 -3514
rect 870 -3522 871 -3514
rect 883 -3522 884 -3514
rect 886 -3522 888 -3514
rect 892 -3522 894 -3514
rect 896 -3522 897 -3514
rect 909 -3522 910 -3514
rect 912 -3522 920 -3514
rect 922 -3522 923 -3514
rect 927 -3522 928 -3514
rect 930 -3522 938 -3514
rect 940 -3522 945 -3514
rect 949 -3522 954 -3514
rect 956 -3522 957 -3514
rect 961 -3522 962 -3514
rect 964 -3522 966 -3514
rect 970 -3522 972 -3514
rect 974 -3522 975 -3514
rect 987 -3522 988 -3514
rect 990 -3522 998 -3514
rect 1000 -3522 1001 -3514
rect 1005 -3522 1006 -3514
rect 1008 -3522 1016 -3514
rect 1018 -3522 1023 -3514
rect 1027 -3522 1032 -3514
rect 1034 -3522 1035 -3514
rect 1039 -3522 1040 -3514
rect 1042 -3522 1047 -3514
rect 1051 -3522 1056 -3514
rect 1058 -3522 1059 -3514
rect 1071 -3522 1072 -3514
rect 1074 -3522 1080 -3514
rect 1082 -3522 1084 -3514
rect 1088 -3522 1090 -3514
rect 1092 -3522 1093 -3514
rect 1215 -3522 1216 -3514
rect 1218 -3522 1220 -3514
rect 1224 -3522 1226 -3514
rect 1228 -3522 1229 -3514
rect 1241 -3522 1242 -3514
rect 1244 -3522 1246 -3514
rect 1250 -3522 1252 -3514
rect 1254 -3522 1255 -3514
rect 1267 -3522 1268 -3514
rect 1270 -3522 1278 -3514
rect 1280 -3522 1281 -3514
rect 1285 -3522 1286 -3514
rect 1288 -3522 1296 -3514
rect 1298 -3522 1303 -3514
rect 1307 -3522 1312 -3514
rect 1314 -3522 1315 -3514
rect 1319 -3522 1320 -3514
rect 1322 -3522 1324 -3514
rect 1328 -3522 1330 -3514
rect 1332 -3522 1333 -3514
rect 1345 -3522 1346 -3514
rect 1348 -3522 1356 -3514
rect 1358 -3522 1359 -3514
rect 1363 -3522 1364 -3514
rect 1366 -3522 1374 -3514
rect 1376 -3522 1381 -3514
rect 1385 -3522 1390 -3514
rect 1392 -3522 1393 -3514
rect 1397 -3522 1398 -3514
rect 1400 -3522 1405 -3514
rect 1409 -3522 1414 -3514
rect 1416 -3522 1417 -3514
rect 1429 -3522 1430 -3514
rect 1432 -3522 1438 -3514
rect 1440 -3522 1442 -3514
rect 1446 -3522 1448 -3514
rect 1450 -3522 1451 -3514
rect -1818 -3652 -1817 -3644
rect -1815 -3652 -1813 -3644
rect -1809 -3652 -1807 -3644
rect -1805 -3652 -1804 -3644
rect -1792 -3652 -1791 -3644
rect -1789 -3652 -1788 -3644
rect -1784 -3652 -1783 -3644
rect -1781 -3652 -1776 -3644
rect -1772 -3652 -1767 -3644
rect -1765 -3652 -1764 -3644
rect -1760 -3652 -1759 -3644
rect -1757 -3652 -1755 -3644
rect -1751 -3652 -1749 -3644
rect -1747 -3652 -1746 -3644
rect -1742 -3652 -1741 -3644
rect -1739 -3652 -1734 -3644
rect -1730 -3652 -1725 -3644
rect -1723 -3652 -1722 -3644
rect -1718 -3652 -1717 -3644
rect -1715 -3652 -1713 -3644
rect -1709 -3652 -1707 -3644
rect -1705 -3652 -1704 -3644
rect -1700 -3652 -1699 -3644
rect -1697 -3652 -1692 -3644
rect -1688 -3652 -1683 -3644
rect -1681 -3652 -1680 -3644
rect -1676 -3652 -1675 -3644
rect -1673 -3652 -1671 -3644
rect -1667 -3652 -1665 -3644
rect -1663 -3652 -1662 -3644
rect -1658 -3652 -1657 -3644
rect -1655 -3652 -1650 -3644
rect -1646 -3652 -1641 -3644
rect -1639 -3652 -1638 -3644
rect -1634 -3652 -1633 -3644
rect -1631 -3652 -1630 -3644
rect -1555 -3652 -1554 -3644
rect -1552 -3652 -1550 -3644
rect -1546 -3652 -1544 -3644
rect -1542 -3652 -1541 -3644
rect -1529 -3652 -1528 -3644
rect -1526 -3652 -1525 -3644
rect -1521 -3652 -1520 -3644
rect -1518 -3652 -1513 -3644
rect -1509 -3652 -1504 -3644
rect -1502 -3652 -1501 -3644
rect -1497 -3652 -1496 -3644
rect -1494 -3652 -1492 -3644
rect -1488 -3652 -1486 -3644
rect -1484 -3652 -1483 -3644
rect -1479 -3652 -1478 -3644
rect -1476 -3652 -1471 -3644
rect -1467 -3652 -1462 -3644
rect -1460 -3652 -1459 -3644
rect -1455 -3652 -1454 -3644
rect -1452 -3652 -1450 -3644
rect -1446 -3652 -1444 -3644
rect -1442 -3652 -1441 -3644
rect -1437 -3652 -1436 -3644
rect -1434 -3652 -1429 -3644
rect -1425 -3652 -1420 -3644
rect -1418 -3652 -1417 -3644
rect -1413 -3652 -1412 -3644
rect -1410 -3652 -1408 -3644
rect -1404 -3652 -1402 -3644
rect -1400 -3652 -1399 -3644
rect -1395 -3652 -1394 -3644
rect -1392 -3652 -1387 -3644
rect -1383 -3652 -1378 -3644
rect -1376 -3652 -1375 -3644
rect -1371 -3652 -1370 -3644
rect -1368 -3652 -1367 -3644
rect -1230 -3652 -1229 -3644
rect -1227 -3652 -1225 -3644
rect -1221 -3652 -1219 -3644
rect -1217 -3652 -1216 -3644
rect -1204 -3652 -1203 -3644
rect -1201 -3652 -1200 -3644
rect -1196 -3652 -1195 -3644
rect -1193 -3652 -1188 -3644
rect -1184 -3652 -1179 -3644
rect -1177 -3652 -1176 -3644
rect -1172 -3652 -1171 -3644
rect -1169 -3652 -1167 -3644
rect -1163 -3652 -1161 -3644
rect -1159 -3652 -1158 -3644
rect -1154 -3652 -1153 -3644
rect -1151 -3652 -1146 -3644
rect -1142 -3652 -1137 -3644
rect -1135 -3652 -1134 -3644
rect -1130 -3652 -1129 -3644
rect -1127 -3652 -1125 -3644
rect -1121 -3652 -1119 -3644
rect -1117 -3652 -1116 -3644
rect -1112 -3652 -1111 -3644
rect -1109 -3652 -1104 -3644
rect -1100 -3652 -1095 -3644
rect -1093 -3652 -1092 -3644
rect -1088 -3652 -1087 -3644
rect -1085 -3652 -1083 -3644
rect -1079 -3652 -1077 -3644
rect -1075 -3652 -1074 -3644
rect -1070 -3652 -1069 -3644
rect -1067 -3652 -1062 -3644
rect -1058 -3652 -1053 -3644
rect -1051 -3652 -1050 -3644
rect -1046 -3652 -1045 -3644
rect -1043 -3652 -1042 -3644
rect -930 -3652 -929 -3644
rect -927 -3652 -925 -3644
rect -921 -3652 -919 -3644
rect -917 -3652 -916 -3644
rect -904 -3652 -903 -3644
rect -901 -3652 -900 -3644
rect -896 -3652 -895 -3644
rect -893 -3652 -888 -3644
rect -884 -3652 -879 -3644
rect -877 -3652 -876 -3644
rect -872 -3652 -871 -3644
rect -869 -3652 -867 -3644
rect -863 -3652 -861 -3644
rect -859 -3652 -858 -3644
rect -854 -3652 -853 -3644
rect -851 -3652 -846 -3644
rect -842 -3652 -837 -3644
rect -835 -3652 -834 -3644
rect -830 -3652 -829 -3644
rect -827 -3652 -825 -3644
rect -821 -3652 -819 -3644
rect -817 -3652 -816 -3644
rect -812 -3652 -811 -3644
rect -809 -3652 -804 -3644
rect -800 -3652 -795 -3644
rect -793 -3652 -792 -3644
rect -788 -3652 -787 -3644
rect -785 -3652 -783 -3644
rect -779 -3652 -777 -3644
rect -775 -3652 -774 -3644
rect -770 -3652 -769 -3644
rect -767 -3652 -762 -3644
rect -758 -3652 -753 -3644
rect -751 -3652 -750 -3644
rect -746 -3652 -745 -3644
rect -743 -3652 -742 -3644
rect -573 -3652 -572 -3644
rect -570 -3652 -568 -3644
rect -564 -3652 -562 -3644
rect -560 -3652 -559 -3644
rect -547 -3652 -546 -3644
rect -544 -3652 -543 -3644
rect -539 -3652 -538 -3644
rect -536 -3652 -531 -3644
rect -527 -3652 -522 -3644
rect -520 -3652 -519 -3644
rect -515 -3652 -514 -3644
rect -512 -3652 -510 -3644
rect -506 -3652 -504 -3644
rect -502 -3652 -501 -3644
rect -497 -3652 -496 -3644
rect -494 -3652 -489 -3644
rect -485 -3652 -480 -3644
rect -478 -3652 -477 -3644
rect -473 -3652 -472 -3644
rect -470 -3652 -468 -3644
rect -464 -3652 -462 -3644
rect -460 -3652 -459 -3644
rect -455 -3652 -454 -3644
rect -452 -3652 -447 -3644
rect -443 -3652 -438 -3644
rect -436 -3652 -435 -3644
rect -431 -3652 -430 -3644
rect -428 -3652 -426 -3644
rect -422 -3652 -420 -3644
rect -418 -3652 -417 -3644
rect -413 -3652 -412 -3644
rect -410 -3652 -405 -3644
rect -401 -3652 -396 -3644
rect -394 -3652 -393 -3644
rect -389 -3652 -388 -3644
rect -386 -3652 -385 -3644
rect -215 -3652 -214 -3644
rect -212 -3652 -210 -3644
rect -206 -3652 -204 -3644
rect -202 -3652 -201 -3644
rect -189 -3652 -188 -3644
rect -186 -3652 -185 -3644
rect -181 -3652 -180 -3644
rect -178 -3652 -173 -3644
rect -169 -3652 -164 -3644
rect -162 -3652 -161 -3644
rect -157 -3652 -156 -3644
rect -154 -3652 -152 -3644
rect -148 -3652 -146 -3644
rect -144 -3652 -143 -3644
rect -139 -3652 -138 -3644
rect -136 -3652 -131 -3644
rect -127 -3652 -122 -3644
rect -120 -3652 -119 -3644
rect -115 -3652 -114 -3644
rect -112 -3652 -110 -3644
rect -106 -3652 -104 -3644
rect -102 -3652 -101 -3644
rect -97 -3652 -96 -3644
rect -94 -3652 -89 -3644
rect -85 -3652 -80 -3644
rect -78 -3652 -77 -3644
rect -73 -3652 -72 -3644
rect -70 -3652 -68 -3644
rect -64 -3652 -62 -3644
rect -60 -3652 -59 -3644
rect -55 -3652 -54 -3644
rect -52 -3652 -47 -3644
rect -43 -3652 -38 -3644
rect -36 -3652 -35 -3644
rect -31 -3652 -30 -3644
rect -28 -3652 -27 -3644
rect -1555 -3823 -1554 -3815
rect -1552 -3823 -1550 -3815
rect -1546 -3823 -1544 -3815
rect -1542 -3823 -1541 -3815
rect -1529 -3823 -1528 -3815
rect -1526 -3823 -1525 -3815
rect -1521 -3823 -1520 -3815
rect -1518 -3823 -1513 -3815
rect -1509 -3823 -1504 -3815
rect -1502 -3823 -1501 -3815
rect -1497 -3823 -1496 -3815
rect -1494 -3823 -1492 -3815
rect -1488 -3823 -1486 -3815
rect -1484 -3823 -1483 -3815
rect -1479 -3823 -1478 -3815
rect -1476 -3823 -1471 -3815
rect -1467 -3823 -1462 -3815
rect -1460 -3823 -1459 -3815
rect -1455 -3823 -1454 -3815
rect -1452 -3823 -1450 -3815
rect -1446 -3823 -1444 -3815
rect -1442 -3823 -1441 -3815
rect -1437 -3823 -1436 -3815
rect -1434 -3823 -1429 -3815
rect -1425 -3823 -1420 -3815
rect -1418 -3823 -1417 -3815
rect -1413 -3823 -1412 -3815
rect -1410 -3823 -1408 -3815
rect -1404 -3823 -1402 -3815
rect -1400 -3823 -1399 -3815
rect -1395 -3823 -1394 -3815
rect -1392 -3823 -1387 -3815
rect -1383 -3823 -1378 -3815
rect -1376 -3823 -1375 -3815
rect -1371 -3823 -1370 -3815
rect -1368 -3823 -1367 -3815
rect -1230 -3823 -1229 -3815
rect -1227 -3823 -1225 -3815
rect -1221 -3823 -1219 -3815
rect -1217 -3823 -1216 -3815
rect -1204 -3823 -1203 -3815
rect -1201 -3823 -1200 -3815
rect -1196 -3823 -1195 -3815
rect -1193 -3823 -1188 -3815
rect -1184 -3823 -1179 -3815
rect -1177 -3823 -1176 -3815
rect -1172 -3823 -1171 -3815
rect -1169 -3823 -1167 -3815
rect -1163 -3823 -1161 -3815
rect -1159 -3823 -1158 -3815
rect -1154 -3823 -1153 -3815
rect -1151 -3823 -1146 -3815
rect -1142 -3823 -1137 -3815
rect -1135 -3823 -1134 -3815
rect -1130 -3823 -1129 -3815
rect -1127 -3823 -1125 -3815
rect -1121 -3823 -1119 -3815
rect -1117 -3823 -1116 -3815
rect -1112 -3823 -1111 -3815
rect -1109 -3823 -1104 -3815
rect -1100 -3823 -1095 -3815
rect -1093 -3823 -1092 -3815
rect -1088 -3823 -1087 -3815
rect -1085 -3823 -1083 -3815
rect -1079 -3823 -1077 -3815
rect -1075 -3823 -1074 -3815
rect -1070 -3823 -1069 -3815
rect -1067 -3823 -1062 -3815
rect -1058 -3823 -1053 -3815
rect -1051 -3823 -1050 -3815
rect -1046 -3823 -1045 -3815
rect -1043 -3823 -1042 -3815
rect -930 -3823 -929 -3815
rect -927 -3823 -925 -3815
rect -921 -3823 -919 -3815
rect -917 -3823 -916 -3815
rect -904 -3823 -903 -3815
rect -901 -3823 -900 -3815
rect -896 -3823 -895 -3815
rect -893 -3823 -888 -3815
rect -884 -3823 -879 -3815
rect -877 -3823 -876 -3815
rect -872 -3823 -871 -3815
rect -869 -3823 -867 -3815
rect -863 -3823 -861 -3815
rect -859 -3823 -858 -3815
rect -854 -3823 -853 -3815
rect -851 -3823 -846 -3815
rect -842 -3823 -837 -3815
rect -835 -3823 -834 -3815
rect -830 -3823 -829 -3815
rect -827 -3823 -825 -3815
rect -821 -3823 -819 -3815
rect -817 -3823 -816 -3815
rect -812 -3823 -811 -3815
rect -809 -3823 -804 -3815
rect -800 -3823 -795 -3815
rect -793 -3823 -792 -3815
rect -788 -3823 -787 -3815
rect -785 -3823 -783 -3815
rect -779 -3823 -777 -3815
rect -775 -3823 -774 -3815
rect -770 -3823 -769 -3815
rect -767 -3823 -762 -3815
rect -758 -3823 -753 -3815
rect -751 -3823 -750 -3815
rect -746 -3823 -745 -3815
rect -743 -3823 -742 -3815
rect -573 -3823 -572 -3815
rect -570 -3823 -568 -3815
rect -564 -3823 -562 -3815
rect -560 -3823 -559 -3815
rect -547 -3823 -546 -3815
rect -544 -3823 -543 -3815
rect -539 -3823 -538 -3815
rect -536 -3823 -531 -3815
rect -527 -3823 -522 -3815
rect -520 -3823 -519 -3815
rect -515 -3823 -514 -3815
rect -512 -3823 -510 -3815
rect -506 -3823 -504 -3815
rect -502 -3823 -501 -3815
rect -497 -3823 -496 -3815
rect -494 -3823 -489 -3815
rect -485 -3823 -480 -3815
rect -478 -3823 -477 -3815
rect -473 -3823 -472 -3815
rect -470 -3823 -468 -3815
rect -464 -3823 -462 -3815
rect -460 -3823 -459 -3815
rect -455 -3823 -454 -3815
rect -452 -3823 -447 -3815
rect -443 -3823 -438 -3815
rect -436 -3823 -435 -3815
rect -431 -3823 -430 -3815
rect -428 -3823 -426 -3815
rect -422 -3823 -420 -3815
rect -418 -3823 -417 -3815
rect -413 -3823 -412 -3815
rect -410 -3823 -405 -3815
rect -401 -3823 -396 -3815
rect -394 -3823 -393 -3815
rect -389 -3823 -388 -3815
rect -386 -3823 -385 -3815
rect -215 -3823 -214 -3815
rect -212 -3823 -210 -3815
rect -206 -3823 -204 -3815
rect -202 -3823 -201 -3815
rect -189 -3823 -188 -3815
rect -186 -3823 -185 -3815
rect -181 -3823 -180 -3815
rect -178 -3823 -173 -3815
rect -169 -3823 -164 -3815
rect -162 -3823 -161 -3815
rect -157 -3823 -156 -3815
rect -154 -3823 -152 -3815
rect -148 -3823 -146 -3815
rect -144 -3823 -143 -3815
rect -139 -3823 -138 -3815
rect -136 -3823 -131 -3815
rect -127 -3823 -122 -3815
rect -120 -3823 -119 -3815
rect -115 -3823 -114 -3815
rect -112 -3823 -110 -3815
rect -106 -3823 -104 -3815
rect -102 -3823 -101 -3815
rect -97 -3823 -96 -3815
rect -94 -3823 -89 -3815
rect -85 -3823 -80 -3815
rect -78 -3823 -77 -3815
rect -73 -3823 -72 -3815
rect -70 -3823 -68 -3815
rect -64 -3823 -62 -3815
rect -60 -3823 -59 -3815
rect -55 -3823 -54 -3815
rect -52 -3823 -47 -3815
rect -43 -3823 -38 -3815
rect -36 -3823 -35 -3815
rect -31 -3823 -30 -3815
rect -28 -3823 -27 -3815
rect 143 -3823 144 -3815
rect 146 -3823 148 -3815
rect 152 -3823 154 -3815
rect 156 -3823 157 -3815
rect 169 -3823 170 -3815
rect 172 -3823 173 -3815
rect 177 -3823 178 -3815
rect 180 -3823 185 -3815
rect 189 -3823 194 -3815
rect 196 -3823 197 -3815
rect 201 -3823 202 -3815
rect 204 -3823 206 -3815
rect 210 -3823 212 -3815
rect 214 -3823 215 -3815
rect 219 -3823 220 -3815
rect 222 -3823 227 -3815
rect 231 -3823 236 -3815
rect 238 -3823 239 -3815
rect 243 -3823 244 -3815
rect 246 -3823 248 -3815
rect 252 -3823 254 -3815
rect 256 -3823 257 -3815
rect 261 -3823 262 -3815
rect 264 -3823 269 -3815
rect 273 -3823 278 -3815
rect 280 -3823 281 -3815
rect 285 -3823 286 -3815
rect 288 -3823 290 -3815
rect 294 -3823 296 -3815
rect 298 -3823 299 -3815
rect 303 -3823 304 -3815
rect 306 -3823 311 -3815
rect 315 -3823 320 -3815
rect 322 -3823 323 -3815
rect 327 -3823 328 -3815
rect 330 -3823 331 -3815
rect 499 -3823 500 -3815
rect 502 -3823 504 -3815
rect 508 -3823 510 -3815
rect 512 -3823 513 -3815
rect 525 -3823 526 -3815
rect 528 -3823 529 -3815
rect 533 -3823 534 -3815
rect 536 -3823 541 -3815
rect 545 -3823 550 -3815
rect 552 -3823 553 -3815
rect 557 -3823 558 -3815
rect 560 -3823 562 -3815
rect 566 -3823 568 -3815
rect 570 -3823 571 -3815
rect 575 -3823 576 -3815
rect 578 -3823 583 -3815
rect 587 -3823 592 -3815
rect 594 -3823 595 -3815
rect 599 -3823 600 -3815
rect 602 -3823 604 -3815
rect 608 -3823 610 -3815
rect 612 -3823 613 -3815
rect 617 -3823 618 -3815
rect 620 -3823 625 -3815
rect 629 -3823 634 -3815
rect 636 -3823 637 -3815
rect 641 -3823 642 -3815
rect 644 -3823 646 -3815
rect 650 -3823 652 -3815
rect 654 -3823 655 -3815
rect 659 -3823 660 -3815
rect 662 -3823 667 -3815
rect 671 -3823 676 -3815
rect 678 -3823 679 -3815
rect 683 -3823 684 -3815
rect 686 -3823 687 -3815
rect 857 -3823 858 -3815
rect 860 -3823 862 -3815
rect 866 -3823 868 -3815
rect 870 -3823 871 -3815
rect 883 -3823 884 -3815
rect 886 -3823 887 -3815
rect 891 -3823 892 -3815
rect 894 -3823 899 -3815
rect 903 -3823 908 -3815
rect 910 -3823 911 -3815
rect 915 -3823 916 -3815
rect 918 -3823 920 -3815
rect 924 -3823 926 -3815
rect 928 -3823 929 -3815
rect 933 -3823 934 -3815
rect 936 -3823 941 -3815
rect 945 -3823 950 -3815
rect 952 -3823 953 -3815
rect 957 -3823 958 -3815
rect 960 -3823 962 -3815
rect 966 -3823 968 -3815
rect 970 -3823 971 -3815
rect 975 -3823 976 -3815
rect 978 -3823 983 -3815
rect 987 -3823 992 -3815
rect 994 -3823 995 -3815
rect 999 -3823 1000 -3815
rect 1002 -3823 1004 -3815
rect 1008 -3823 1010 -3815
rect 1012 -3823 1013 -3815
rect 1017 -3823 1018 -3815
rect 1020 -3823 1025 -3815
rect 1029 -3823 1034 -3815
rect 1036 -3823 1037 -3815
rect 1041 -3823 1042 -3815
rect 1044 -3823 1045 -3815
rect 1215 -3823 1216 -3815
rect 1218 -3823 1220 -3815
rect 1224 -3823 1226 -3815
rect 1228 -3823 1229 -3815
rect 1241 -3823 1242 -3815
rect 1244 -3823 1245 -3815
rect 1249 -3823 1250 -3815
rect 1252 -3823 1257 -3815
rect 1261 -3823 1266 -3815
rect 1268 -3823 1269 -3815
rect 1273 -3823 1274 -3815
rect 1276 -3823 1278 -3815
rect 1282 -3823 1284 -3815
rect 1286 -3823 1287 -3815
rect 1291 -3823 1292 -3815
rect 1294 -3823 1299 -3815
rect 1303 -3823 1308 -3815
rect 1310 -3823 1311 -3815
rect 1315 -3823 1316 -3815
rect 1318 -3823 1320 -3815
rect 1324 -3823 1326 -3815
rect 1328 -3823 1329 -3815
rect 1333 -3823 1334 -3815
rect 1336 -3823 1341 -3815
rect 1345 -3823 1350 -3815
rect 1352 -3823 1353 -3815
rect 1357 -3823 1358 -3815
rect 1360 -3823 1362 -3815
rect 1366 -3823 1368 -3815
rect 1370 -3823 1371 -3815
rect 1375 -3823 1376 -3815
rect 1378 -3823 1383 -3815
rect 1387 -3823 1392 -3815
rect 1394 -3823 1395 -3815
rect 1399 -3823 1400 -3815
rect 1402 -3823 1403 -3815
rect -1555 -3998 -1554 -3990
rect -1552 -3998 -1550 -3990
rect -1546 -3998 -1544 -3990
rect -1542 -3998 -1541 -3990
rect -1529 -3998 -1528 -3990
rect -1526 -3998 -1525 -3990
rect -1521 -3998 -1520 -3990
rect -1518 -3998 -1513 -3990
rect -1509 -3998 -1504 -3990
rect -1502 -3998 -1501 -3990
rect -1497 -3998 -1496 -3990
rect -1494 -3998 -1492 -3990
rect -1488 -3998 -1486 -3990
rect -1484 -3998 -1483 -3990
rect -1479 -3998 -1478 -3990
rect -1476 -3998 -1471 -3990
rect -1467 -3998 -1462 -3990
rect -1460 -3998 -1459 -3990
rect -1455 -3998 -1454 -3990
rect -1452 -3998 -1450 -3990
rect -1446 -3998 -1444 -3990
rect -1442 -3998 -1441 -3990
rect -1437 -3998 -1436 -3990
rect -1434 -3998 -1429 -3990
rect -1425 -3998 -1420 -3990
rect -1418 -3998 -1417 -3990
rect -1413 -3998 -1412 -3990
rect -1410 -3998 -1408 -3990
rect -1404 -3998 -1402 -3990
rect -1400 -3998 -1399 -3990
rect -1395 -3998 -1394 -3990
rect -1392 -3998 -1387 -3990
rect -1383 -3998 -1378 -3990
rect -1376 -3998 -1375 -3990
rect -1371 -3998 -1370 -3990
rect -1368 -3998 -1367 -3990
rect -1230 -3998 -1229 -3990
rect -1227 -3998 -1225 -3990
rect -1221 -3998 -1219 -3990
rect -1217 -3998 -1216 -3990
rect -1204 -3998 -1203 -3990
rect -1201 -3998 -1200 -3990
rect -1196 -3998 -1195 -3990
rect -1193 -3998 -1188 -3990
rect -1184 -3998 -1179 -3990
rect -1177 -3998 -1176 -3990
rect -1172 -3998 -1171 -3990
rect -1169 -3998 -1167 -3990
rect -1163 -3998 -1161 -3990
rect -1159 -3998 -1158 -3990
rect -1154 -3998 -1153 -3990
rect -1151 -3998 -1146 -3990
rect -1142 -3998 -1137 -3990
rect -1135 -3998 -1134 -3990
rect -1130 -3998 -1129 -3990
rect -1127 -3998 -1125 -3990
rect -1121 -3998 -1119 -3990
rect -1117 -3998 -1116 -3990
rect -1112 -3998 -1111 -3990
rect -1109 -3998 -1104 -3990
rect -1100 -3998 -1095 -3990
rect -1093 -3998 -1092 -3990
rect -1088 -3998 -1087 -3990
rect -1085 -3998 -1083 -3990
rect -1079 -3998 -1077 -3990
rect -1075 -3998 -1074 -3990
rect -1070 -3998 -1069 -3990
rect -1067 -3998 -1062 -3990
rect -1058 -3998 -1053 -3990
rect -1051 -3998 -1050 -3990
rect -1046 -3998 -1045 -3990
rect -1043 -3998 -1042 -3990
rect -931 -3998 -930 -3990
rect -928 -3998 -926 -3990
rect -922 -3998 -920 -3990
rect -918 -3998 -917 -3990
rect -905 -3998 -904 -3990
rect -902 -3998 -901 -3990
rect -897 -3998 -896 -3990
rect -894 -3998 -889 -3990
rect -885 -3998 -880 -3990
rect -878 -3998 -877 -3990
rect -873 -3998 -872 -3990
rect -870 -3998 -868 -3990
rect -864 -3998 -862 -3990
rect -860 -3998 -859 -3990
rect -855 -3998 -854 -3990
rect -852 -3998 -847 -3990
rect -843 -3998 -838 -3990
rect -836 -3998 -835 -3990
rect -831 -3998 -830 -3990
rect -828 -3998 -826 -3990
rect -822 -3998 -820 -3990
rect -818 -3998 -817 -3990
rect -813 -3998 -812 -3990
rect -810 -3998 -805 -3990
rect -801 -3998 -796 -3990
rect -794 -3998 -793 -3990
rect -789 -3998 -788 -3990
rect -786 -3998 -784 -3990
rect -780 -3998 -778 -3990
rect -776 -3998 -775 -3990
rect -771 -3998 -770 -3990
rect -768 -3998 -763 -3990
rect -759 -3998 -754 -3990
rect -752 -3998 -751 -3990
rect -747 -3998 -746 -3990
rect -744 -3998 -743 -3990
rect -573 -3998 -572 -3990
rect -570 -3998 -568 -3990
rect -564 -3998 -562 -3990
rect -560 -3998 -559 -3990
rect -547 -3998 -546 -3990
rect -544 -3998 -543 -3990
rect -539 -3998 -538 -3990
rect -536 -3998 -531 -3990
rect -527 -3998 -522 -3990
rect -520 -3998 -519 -3990
rect -515 -3998 -514 -3990
rect -512 -3998 -510 -3990
rect -506 -3998 -504 -3990
rect -502 -3998 -501 -3990
rect -497 -3998 -496 -3990
rect -494 -3998 -489 -3990
rect -485 -3998 -480 -3990
rect -478 -3998 -477 -3990
rect -473 -3998 -472 -3990
rect -470 -3998 -468 -3990
rect -464 -3998 -462 -3990
rect -460 -3998 -459 -3990
rect -455 -3998 -454 -3990
rect -452 -3998 -447 -3990
rect -443 -3998 -438 -3990
rect -436 -3998 -435 -3990
rect -431 -3998 -430 -3990
rect -428 -3998 -426 -3990
rect -422 -3998 -420 -3990
rect -418 -3998 -417 -3990
rect -413 -3998 -412 -3990
rect -410 -3998 -405 -3990
rect -401 -3998 -396 -3990
rect -394 -3998 -393 -3990
rect -389 -3998 -388 -3990
rect -386 -3998 -385 -3990
rect -215 -3998 -214 -3990
rect -212 -3998 -210 -3990
rect -206 -3998 -204 -3990
rect -202 -3998 -201 -3990
rect -189 -3998 -188 -3990
rect -186 -3998 -185 -3990
rect -181 -3998 -180 -3990
rect -178 -3998 -173 -3990
rect -169 -3998 -164 -3990
rect -162 -3998 -161 -3990
rect -157 -3998 -156 -3990
rect -154 -3998 -152 -3990
rect -148 -3998 -146 -3990
rect -144 -3998 -143 -3990
rect -139 -3998 -138 -3990
rect -136 -3998 -131 -3990
rect -127 -3998 -122 -3990
rect -120 -3998 -119 -3990
rect -115 -3998 -114 -3990
rect -112 -3998 -110 -3990
rect -106 -3998 -104 -3990
rect -102 -3998 -101 -3990
rect -97 -3998 -96 -3990
rect -94 -3998 -89 -3990
rect -85 -3998 -80 -3990
rect -78 -3998 -77 -3990
rect -73 -3998 -72 -3990
rect -70 -3998 -68 -3990
rect -64 -3998 -62 -3990
rect -60 -3998 -59 -3990
rect -55 -3998 -54 -3990
rect -52 -3998 -47 -3990
rect -43 -3998 -38 -3990
rect -36 -3998 -35 -3990
rect -31 -3998 -30 -3990
rect -28 -3998 -27 -3990
rect 143 -3998 144 -3990
rect 146 -3998 148 -3990
rect 152 -3998 154 -3990
rect 156 -3998 157 -3990
rect 169 -3998 170 -3990
rect 172 -3998 173 -3990
rect 177 -3998 178 -3990
rect 180 -3998 185 -3990
rect 189 -3998 194 -3990
rect 196 -3998 197 -3990
rect 201 -3998 202 -3990
rect 204 -3998 206 -3990
rect 210 -3998 212 -3990
rect 214 -3998 215 -3990
rect 219 -3998 220 -3990
rect 222 -3998 227 -3990
rect 231 -3998 236 -3990
rect 238 -3998 239 -3990
rect 243 -3998 244 -3990
rect 246 -3998 248 -3990
rect 252 -3998 254 -3990
rect 256 -3998 257 -3990
rect 261 -3998 262 -3990
rect 264 -3998 269 -3990
rect 273 -3998 278 -3990
rect 280 -3998 281 -3990
rect 285 -3998 286 -3990
rect 288 -3998 290 -3990
rect 294 -3998 296 -3990
rect 298 -3998 299 -3990
rect 303 -3998 304 -3990
rect 306 -3998 311 -3990
rect 315 -3998 320 -3990
rect 322 -3998 323 -3990
rect 327 -3998 328 -3990
rect 330 -3998 331 -3990
rect 499 -3998 500 -3990
rect 502 -3998 504 -3990
rect 508 -3998 510 -3990
rect 512 -3998 513 -3990
rect 525 -3998 526 -3990
rect 528 -3998 529 -3990
rect 533 -3998 534 -3990
rect 536 -3998 541 -3990
rect 545 -3998 550 -3990
rect 552 -3998 553 -3990
rect 557 -3998 558 -3990
rect 560 -3998 562 -3990
rect 566 -3998 568 -3990
rect 570 -3998 571 -3990
rect 575 -3998 576 -3990
rect 578 -3998 583 -3990
rect 587 -3998 592 -3990
rect 594 -3998 595 -3990
rect 599 -3998 600 -3990
rect 602 -3998 604 -3990
rect 608 -3998 610 -3990
rect 612 -3998 613 -3990
rect 617 -3998 618 -3990
rect 620 -3998 625 -3990
rect 629 -3998 634 -3990
rect 636 -3998 637 -3990
rect 641 -3998 642 -3990
rect 644 -3998 646 -3990
rect 650 -3998 652 -3990
rect 654 -3998 655 -3990
rect 659 -3998 660 -3990
rect 662 -3998 667 -3990
rect 671 -3998 676 -3990
rect 678 -3998 679 -3990
rect 683 -3998 684 -3990
rect 686 -3998 687 -3990
rect 857 -3998 858 -3990
rect 860 -3998 862 -3990
rect 866 -3998 868 -3990
rect 870 -3998 871 -3990
rect 883 -3998 884 -3990
rect 886 -3998 887 -3990
rect 891 -3998 892 -3990
rect 894 -3998 899 -3990
rect 903 -3998 908 -3990
rect 910 -3998 911 -3990
rect 915 -3998 916 -3990
rect 918 -3998 920 -3990
rect 924 -3998 926 -3990
rect 928 -3998 929 -3990
rect 933 -3998 934 -3990
rect 936 -3998 941 -3990
rect 945 -3998 950 -3990
rect 952 -3998 953 -3990
rect 957 -3998 958 -3990
rect 960 -3998 962 -3990
rect 966 -3998 968 -3990
rect 970 -3998 971 -3990
rect 975 -3998 976 -3990
rect 978 -3998 983 -3990
rect 987 -3998 992 -3990
rect 994 -3998 995 -3990
rect 999 -3998 1000 -3990
rect 1002 -3998 1004 -3990
rect 1008 -3998 1010 -3990
rect 1012 -3998 1013 -3990
rect 1017 -3998 1018 -3990
rect 1020 -3998 1025 -3990
rect 1029 -3998 1034 -3990
rect 1036 -3998 1037 -3990
rect 1041 -3998 1042 -3990
rect 1044 -3998 1045 -3990
rect 1215 -3998 1216 -3990
rect 1218 -3998 1220 -3990
rect 1224 -3998 1226 -3990
rect 1228 -3998 1229 -3990
rect 1241 -3998 1242 -3990
rect 1244 -3998 1245 -3990
rect 1249 -3998 1250 -3990
rect 1252 -3998 1257 -3990
rect 1261 -3998 1266 -3990
rect 1268 -3998 1269 -3990
rect 1273 -3998 1274 -3990
rect 1276 -3998 1278 -3990
rect 1282 -3998 1284 -3990
rect 1286 -3998 1287 -3990
rect 1291 -3998 1292 -3990
rect 1294 -3998 1299 -3990
rect 1303 -3998 1308 -3990
rect 1310 -3998 1311 -3990
rect 1315 -3998 1316 -3990
rect 1318 -3998 1320 -3990
rect 1324 -3998 1326 -3990
rect 1328 -3998 1329 -3990
rect 1333 -3998 1334 -3990
rect 1336 -3998 1341 -3990
rect 1345 -3998 1350 -3990
rect 1352 -3998 1353 -3990
rect 1357 -3998 1358 -3990
rect 1360 -3998 1362 -3990
rect 1366 -3998 1368 -3990
rect 1370 -3998 1371 -3990
rect 1375 -3998 1376 -3990
rect 1378 -3998 1383 -3990
rect 1387 -3998 1392 -3990
rect 1394 -3998 1395 -3990
rect 1399 -3998 1400 -3990
rect 1402 -3998 1403 -3990
rect -1305 -4113 -1304 -4105
rect -1302 -4113 -1301 -4105
rect -1297 -4113 -1296 -4105
rect -1294 -4113 -1292 -4105
rect -1288 -4113 -1286 -4105
rect -1284 -4113 -1283 -4105
rect -931 -4113 -930 -4105
rect -928 -4113 -927 -4105
rect -923 -4113 -922 -4105
rect -920 -4113 -918 -4105
rect -914 -4113 -912 -4105
rect -910 -4113 -909 -4105
rect -573 -4113 -572 -4105
rect -570 -4113 -569 -4105
rect -565 -4113 -564 -4105
rect -562 -4113 -560 -4105
rect -556 -4113 -554 -4105
rect -552 -4113 -551 -4105
rect -215 -4113 -214 -4105
rect -212 -4113 -211 -4105
rect -207 -4113 -206 -4105
rect -204 -4113 -202 -4105
rect -198 -4113 -196 -4105
rect -194 -4113 -193 -4105
rect 143 -4113 144 -4105
rect 146 -4113 147 -4105
rect 151 -4113 152 -4105
rect 154 -4113 156 -4105
rect 160 -4113 162 -4105
rect 164 -4113 165 -4105
rect 499 -4113 500 -4105
rect 502 -4113 503 -4105
rect 507 -4113 508 -4105
rect 510 -4113 512 -4105
rect 516 -4113 518 -4105
rect 520 -4113 521 -4105
rect 857 -4113 858 -4105
rect 860 -4113 861 -4105
rect 865 -4113 866 -4105
rect 868 -4113 870 -4105
rect 874 -4113 876 -4105
rect 878 -4113 879 -4105
rect 1215 -4113 1216 -4105
rect 1218 -4113 1219 -4105
rect 1223 -4113 1224 -4105
rect 1226 -4113 1228 -4105
rect 1232 -4113 1234 -4105
rect 1236 -4113 1237 -4105
rect -1230 -4272 -1229 -4264
rect -1227 -4272 -1225 -4264
rect -1221 -4272 -1219 -4264
rect -1217 -4272 -1216 -4264
rect -1204 -4272 -1203 -4264
rect -1201 -4272 -1193 -4264
rect -1191 -4272 -1190 -4264
rect -1186 -4272 -1185 -4264
rect -1183 -4272 -1175 -4264
rect -1173 -4272 -1168 -4264
rect -1164 -4272 -1159 -4264
rect -1157 -4272 -1156 -4264
rect -1152 -4272 -1151 -4264
rect -1149 -4272 -1147 -4264
rect -1143 -4272 -1141 -4264
rect -1139 -4272 -1138 -4264
rect -931 -4272 -930 -4264
rect -928 -4272 -926 -4264
rect -922 -4272 -920 -4264
rect -918 -4272 -917 -4264
rect -905 -4272 -904 -4264
rect -902 -4272 -900 -4264
rect -896 -4272 -894 -4264
rect -892 -4272 -891 -4264
rect -879 -4272 -878 -4264
rect -876 -4272 -868 -4264
rect -866 -4272 -865 -4264
rect -861 -4272 -860 -4264
rect -858 -4272 -850 -4264
rect -848 -4272 -843 -4264
rect -839 -4272 -834 -4264
rect -832 -4272 -831 -4264
rect -827 -4272 -826 -4264
rect -824 -4272 -822 -4264
rect -818 -4272 -816 -4264
rect -814 -4272 -813 -4264
rect -801 -4272 -800 -4264
rect -798 -4272 -790 -4264
rect -788 -4272 -787 -4264
rect -783 -4272 -782 -4264
rect -780 -4272 -772 -4264
rect -770 -4272 -765 -4264
rect -761 -4272 -756 -4264
rect -754 -4272 -753 -4264
rect -749 -4272 -748 -4264
rect -746 -4272 -741 -4264
rect -737 -4272 -732 -4264
rect -730 -4272 -729 -4264
rect -717 -4272 -716 -4264
rect -714 -4272 -708 -4264
rect -706 -4272 -704 -4264
rect -700 -4272 -698 -4264
rect -696 -4272 -695 -4264
rect -573 -4272 -572 -4264
rect -570 -4272 -568 -4264
rect -564 -4272 -562 -4264
rect -560 -4272 -559 -4264
rect -547 -4272 -546 -4264
rect -544 -4272 -542 -4264
rect -538 -4272 -536 -4264
rect -534 -4272 -533 -4264
rect -521 -4272 -520 -4264
rect -518 -4272 -510 -4264
rect -508 -4272 -507 -4264
rect -503 -4272 -502 -4264
rect -500 -4272 -492 -4264
rect -490 -4272 -485 -4264
rect -481 -4272 -476 -4264
rect -474 -4272 -473 -4264
rect -469 -4272 -468 -4264
rect -466 -4272 -464 -4264
rect -460 -4272 -458 -4264
rect -456 -4272 -455 -4264
rect -443 -4272 -442 -4264
rect -440 -4272 -432 -4264
rect -430 -4272 -429 -4264
rect -425 -4272 -424 -4264
rect -422 -4272 -414 -4264
rect -412 -4272 -407 -4264
rect -403 -4272 -398 -4264
rect -396 -4272 -395 -4264
rect -391 -4272 -390 -4264
rect -388 -4272 -383 -4264
rect -379 -4272 -374 -4264
rect -372 -4272 -371 -4264
rect -359 -4272 -358 -4264
rect -356 -4272 -350 -4264
rect -348 -4272 -346 -4264
rect -342 -4272 -340 -4264
rect -338 -4272 -337 -4264
rect -215 -4272 -214 -4264
rect -212 -4272 -210 -4264
rect -206 -4272 -204 -4264
rect -202 -4272 -201 -4264
rect -189 -4272 -188 -4264
rect -186 -4272 -184 -4264
rect -180 -4272 -178 -4264
rect -176 -4272 -175 -4264
rect -163 -4272 -162 -4264
rect -160 -4272 -152 -4264
rect -150 -4272 -149 -4264
rect -145 -4272 -144 -4264
rect -142 -4272 -134 -4264
rect -132 -4272 -127 -4264
rect -123 -4272 -118 -4264
rect -116 -4272 -115 -4264
rect -111 -4272 -110 -4264
rect -108 -4272 -106 -4264
rect -102 -4272 -100 -4264
rect -98 -4272 -97 -4264
rect -85 -4272 -84 -4264
rect -82 -4272 -74 -4264
rect -72 -4272 -71 -4264
rect -67 -4272 -66 -4264
rect -64 -4272 -56 -4264
rect -54 -4272 -49 -4264
rect -45 -4272 -40 -4264
rect -38 -4272 -37 -4264
rect -33 -4272 -32 -4264
rect -30 -4272 -25 -4264
rect -21 -4272 -16 -4264
rect -14 -4272 -13 -4264
rect -1 -4272 0 -4264
rect 2 -4272 8 -4264
rect 10 -4272 12 -4264
rect 16 -4272 18 -4264
rect 20 -4272 21 -4264
rect 143 -4272 144 -4264
rect 146 -4272 148 -4264
rect 152 -4272 154 -4264
rect 156 -4272 157 -4264
rect 169 -4272 170 -4264
rect 172 -4272 174 -4264
rect 178 -4272 180 -4264
rect 182 -4272 183 -4264
rect 195 -4272 196 -4264
rect 198 -4272 206 -4264
rect 208 -4272 209 -4264
rect 213 -4272 214 -4264
rect 216 -4272 224 -4264
rect 226 -4272 231 -4264
rect 235 -4272 240 -4264
rect 242 -4272 243 -4264
rect 247 -4272 248 -4264
rect 250 -4272 252 -4264
rect 256 -4272 258 -4264
rect 260 -4272 261 -4264
rect 273 -4272 274 -4264
rect 276 -4272 284 -4264
rect 286 -4272 287 -4264
rect 291 -4272 292 -4264
rect 294 -4272 302 -4264
rect 304 -4272 309 -4264
rect 313 -4272 318 -4264
rect 320 -4272 321 -4264
rect 325 -4272 326 -4264
rect 328 -4272 333 -4264
rect 337 -4272 342 -4264
rect 344 -4272 345 -4264
rect 357 -4272 358 -4264
rect 360 -4272 366 -4264
rect 368 -4272 370 -4264
rect 374 -4272 376 -4264
rect 378 -4272 379 -4264
rect 499 -4272 500 -4264
rect 502 -4272 504 -4264
rect 508 -4272 510 -4264
rect 512 -4272 513 -4264
rect 525 -4272 526 -4264
rect 528 -4272 530 -4264
rect 534 -4272 536 -4264
rect 538 -4272 539 -4264
rect 551 -4272 552 -4264
rect 554 -4272 562 -4264
rect 564 -4272 565 -4264
rect 569 -4272 570 -4264
rect 572 -4272 580 -4264
rect 582 -4272 587 -4264
rect 591 -4272 596 -4264
rect 598 -4272 599 -4264
rect 603 -4272 604 -4264
rect 606 -4272 608 -4264
rect 612 -4272 614 -4264
rect 616 -4272 617 -4264
rect 629 -4272 630 -4264
rect 632 -4272 640 -4264
rect 642 -4272 643 -4264
rect 647 -4272 648 -4264
rect 650 -4272 658 -4264
rect 660 -4272 665 -4264
rect 669 -4272 674 -4264
rect 676 -4272 677 -4264
rect 681 -4272 682 -4264
rect 684 -4272 689 -4264
rect 693 -4272 698 -4264
rect 700 -4272 701 -4264
rect 713 -4272 714 -4264
rect 716 -4272 722 -4264
rect 724 -4272 726 -4264
rect 730 -4272 732 -4264
rect 734 -4272 735 -4264
rect 857 -4272 858 -4264
rect 860 -4272 862 -4264
rect 866 -4272 868 -4264
rect 870 -4272 871 -4264
rect 883 -4272 884 -4264
rect 886 -4272 888 -4264
rect 892 -4272 894 -4264
rect 896 -4272 897 -4264
rect 909 -4272 910 -4264
rect 912 -4272 920 -4264
rect 922 -4272 923 -4264
rect 927 -4272 928 -4264
rect 930 -4272 938 -4264
rect 940 -4272 945 -4264
rect 949 -4272 954 -4264
rect 956 -4272 957 -4264
rect 961 -4272 962 -4264
rect 964 -4272 966 -4264
rect 970 -4272 972 -4264
rect 974 -4272 975 -4264
rect 987 -4272 988 -4264
rect 990 -4272 998 -4264
rect 1000 -4272 1001 -4264
rect 1005 -4272 1006 -4264
rect 1008 -4272 1016 -4264
rect 1018 -4272 1023 -4264
rect 1027 -4272 1032 -4264
rect 1034 -4272 1035 -4264
rect 1039 -4272 1040 -4264
rect 1042 -4272 1047 -4264
rect 1051 -4272 1056 -4264
rect 1058 -4272 1059 -4264
rect 1071 -4272 1072 -4264
rect 1074 -4272 1080 -4264
rect 1082 -4272 1084 -4264
rect 1088 -4272 1090 -4264
rect 1092 -4272 1093 -4264
rect 1215 -4272 1216 -4264
rect 1218 -4272 1220 -4264
rect 1224 -4272 1226 -4264
rect 1228 -4272 1229 -4264
rect 1241 -4272 1242 -4264
rect 1244 -4272 1246 -4264
rect 1250 -4272 1252 -4264
rect 1254 -4272 1255 -4264
rect 1267 -4272 1268 -4264
rect 1270 -4272 1278 -4264
rect 1280 -4272 1281 -4264
rect 1285 -4272 1286 -4264
rect 1288 -4272 1296 -4264
rect 1298 -4272 1303 -4264
rect 1307 -4272 1312 -4264
rect 1314 -4272 1315 -4264
rect 1319 -4272 1320 -4264
rect 1322 -4272 1324 -4264
rect 1328 -4272 1330 -4264
rect 1332 -4272 1333 -4264
rect 1345 -4272 1346 -4264
rect 1348 -4272 1356 -4264
rect 1358 -4272 1359 -4264
rect 1363 -4272 1364 -4264
rect 1366 -4272 1374 -4264
rect 1376 -4272 1381 -4264
rect 1385 -4272 1390 -4264
rect 1392 -4272 1393 -4264
rect 1397 -4272 1398 -4264
rect 1400 -4272 1405 -4264
rect 1409 -4272 1414 -4264
rect 1416 -4272 1417 -4264
rect 1429 -4272 1430 -4264
rect 1432 -4272 1438 -4264
rect 1440 -4272 1442 -4264
rect 1446 -4272 1448 -4264
rect 1450 -4272 1451 -4264
rect -1810 -4395 -1809 -4387
rect -1807 -4395 -1805 -4387
rect -1801 -4395 -1799 -4387
rect -1797 -4395 -1796 -4387
rect -1784 -4395 -1783 -4387
rect -1781 -4395 -1780 -4387
rect -1776 -4395 -1775 -4387
rect -1773 -4395 -1768 -4387
rect -1764 -4395 -1759 -4387
rect -1757 -4395 -1756 -4387
rect -1752 -4395 -1751 -4387
rect -1749 -4395 -1747 -4387
rect -1743 -4395 -1741 -4387
rect -1739 -4395 -1738 -4387
rect -1734 -4395 -1733 -4387
rect -1731 -4395 -1726 -4387
rect -1722 -4395 -1717 -4387
rect -1715 -4395 -1714 -4387
rect -1710 -4395 -1709 -4387
rect -1707 -4395 -1705 -4387
rect -1701 -4395 -1699 -4387
rect -1697 -4395 -1696 -4387
rect -1692 -4395 -1691 -4387
rect -1689 -4395 -1684 -4387
rect -1680 -4395 -1675 -4387
rect -1673 -4395 -1672 -4387
rect -1668 -4395 -1667 -4387
rect -1665 -4395 -1663 -4387
rect -1659 -4395 -1657 -4387
rect -1655 -4395 -1654 -4387
rect -1650 -4395 -1649 -4387
rect -1647 -4395 -1642 -4387
rect -1638 -4395 -1633 -4387
rect -1631 -4395 -1630 -4387
rect -1626 -4395 -1625 -4387
rect -1623 -4395 -1622 -4387
rect -1547 -4395 -1546 -4387
rect -1544 -4395 -1542 -4387
rect -1538 -4395 -1536 -4387
rect -1534 -4395 -1533 -4387
rect -1521 -4395 -1520 -4387
rect -1518 -4395 -1517 -4387
rect -1513 -4395 -1512 -4387
rect -1510 -4395 -1505 -4387
rect -1501 -4395 -1496 -4387
rect -1494 -4395 -1493 -4387
rect -1489 -4395 -1488 -4387
rect -1486 -4395 -1484 -4387
rect -1480 -4395 -1478 -4387
rect -1476 -4395 -1475 -4387
rect -1471 -4395 -1470 -4387
rect -1468 -4395 -1463 -4387
rect -1459 -4395 -1454 -4387
rect -1452 -4395 -1451 -4387
rect -1447 -4395 -1446 -4387
rect -1444 -4395 -1442 -4387
rect -1438 -4395 -1436 -4387
rect -1434 -4395 -1433 -4387
rect -1429 -4395 -1428 -4387
rect -1426 -4395 -1421 -4387
rect -1417 -4395 -1412 -4387
rect -1410 -4395 -1409 -4387
rect -1405 -4395 -1404 -4387
rect -1402 -4395 -1400 -4387
rect -1396 -4395 -1394 -4387
rect -1392 -4395 -1391 -4387
rect -1387 -4395 -1386 -4387
rect -1384 -4395 -1379 -4387
rect -1375 -4395 -1370 -4387
rect -1368 -4395 -1367 -4387
rect -1363 -4395 -1362 -4387
rect -1360 -4395 -1359 -4387
rect -1230 -4395 -1229 -4387
rect -1227 -4395 -1225 -4387
rect -1221 -4395 -1219 -4387
rect -1217 -4395 -1216 -4387
rect -1204 -4395 -1203 -4387
rect -1201 -4395 -1200 -4387
rect -1196 -4395 -1195 -4387
rect -1193 -4395 -1188 -4387
rect -1184 -4395 -1179 -4387
rect -1177 -4395 -1176 -4387
rect -1172 -4395 -1171 -4387
rect -1169 -4395 -1167 -4387
rect -1163 -4395 -1161 -4387
rect -1159 -4395 -1158 -4387
rect -1154 -4395 -1153 -4387
rect -1151 -4395 -1146 -4387
rect -1142 -4395 -1137 -4387
rect -1135 -4395 -1134 -4387
rect -1130 -4395 -1129 -4387
rect -1127 -4395 -1125 -4387
rect -1121 -4395 -1119 -4387
rect -1117 -4395 -1116 -4387
rect -1112 -4395 -1111 -4387
rect -1109 -4395 -1104 -4387
rect -1100 -4395 -1095 -4387
rect -1093 -4395 -1092 -4387
rect -1088 -4395 -1087 -4387
rect -1085 -4395 -1083 -4387
rect -1079 -4395 -1077 -4387
rect -1075 -4395 -1074 -4387
rect -1070 -4395 -1069 -4387
rect -1067 -4395 -1062 -4387
rect -1058 -4395 -1053 -4387
rect -1051 -4395 -1050 -4387
rect -1046 -4395 -1045 -4387
rect -1043 -4395 -1042 -4387
rect -931 -4395 -930 -4387
rect -928 -4395 -926 -4387
rect -922 -4395 -920 -4387
rect -918 -4395 -917 -4387
rect -905 -4395 -904 -4387
rect -902 -4395 -901 -4387
rect -897 -4395 -896 -4387
rect -894 -4395 -889 -4387
rect -885 -4395 -880 -4387
rect -878 -4395 -877 -4387
rect -873 -4395 -872 -4387
rect -870 -4395 -868 -4387
rect -864 -4395 -862 -4387
rect -860 -4395 -859 -4387
rect -855 -4395 -854 -4387
rect -852 -4395 -847 -4387
rect -843 -4395 -838 -4387
rect -836 -4395 -835 -4387
rect -831 -4395 -830 -4387
rect -828 -4395 -826 -4387
rect -822 -4395 -820 -4387
rect -818 -4395 -817 -4387
rect -813 -4395 -812 -4387
rect -810 -4395 -805 -4387
rect -801 -4395 -796 -4387
rect -794 -4395 -793 -4387
rect -789 -4395 -788 -4387
rect -786 -4395 -784 -4387
rect -780 -4395 -778 -4387
rect -776 -4395 -775 -4387
rect -771 -4395 -770 -4387
rect -768 -4395 -763 -4387
rect -759 -4395 -754 -4387
rect -752 -4395 -751 -4387
rect -747 -4395 -746 -4387
rect -744 -4395 -743 -4387
rect -573 -4395 -572 -4387
rect -570 -4395 -568 -4387
rect -564 -4395 -562 -4387
rect -560 -4395 -559 -4387
rect -547 -4395 -546 -4387
rect -544 -4395 -543 -4387
rect -539 -4395 -538 -4387
rect -536 -4395 -531 -4387
rect -527 -4395 -522 -4387
rect -520 -4395 -519 -4387
rect -515 -4395 -514 -4387
rect -512 -4395 -510 -4387
rect -506 -4395 -504 -4387
rect -502 -4395 -501 -4387
rect -497 -4395 -496 -4387
rect -494 -4395 -489 -4387
rect -485 -4395 -480 -4387
rect -478 -4395 -477 -4387
rect -473 -4395 -472 -4387
rect -470 -4395 -468 -4387
rect -464 -4395 -462 -4387
rect -460 -4395 -459 -4387
rect -455 -4395 -454 -4387
rect -452 -4395 -447 -4387
rect -443 -4395 -438 -4387
rect -436 -4395 -435 -4387
rect -431 -4395 -430 -4387
rect -428 -4395 -426 -4387
rect -422 -4395 -420 -4387
rect -418 -4395 -417 -4387
rect -413 -4395 -412 -4387
rect -410 -4395 -405 -4387
rect -401 -4395 -396 -4387
rect -394 -4395 -393 -4387
rect -389 -4395 -388 -4387
rect -386 -4395 -385 -4387
rect -1810 -4566 -1809 -4558
rect -1807 -4566 -1805 -4558
rect -1801 -4566 -1799 -4558
rect -1797 -4566 -1796 -4558
rect -1784 -4566 -1783 -4558
rect -1781 -4566 -1780 -4558
rect -1776 -4566 -1775 -4558
rect -1773 -4566 -1768 -4558
rect -1764 -4566 -1759 -4558
rect -1757 -4566 -1756 -4558
rect -1752 -4566 -1751 -4558
rect -1749 -4566 -1747 -4558
rect -1743 -4566 -1741 -4558
rect -1739 -4566 -1738 -4558
rect -1734 -4566 -1733 -4558
rect -1731 -4566 -1726 -4558
rect -1722 -4566 -1717 -4558
rect -1715 -4566 -1714 -4558
rect -1710 -4566 -1709 -4558
rect -1707 -4566 -1705 -4558
rect -1701 -4566 -1699 -4558
rect -1697 -4566 -1696 -4558
rect -1692 -4566 -1691 -4558
rect -1689 -4566 -1684 -4558
rect -1680 -4566 -1675 -4558
rect -1673 -4566 -1672 -4558
rect -1668 -4566 -1667 -4558
rect -1665 -4566 -1663 -4558
rect -1659 -4566 -1657 -4558
rect -1655 -4566 -1654 -4558
rect -1650 -4566 -1649 -4558
rect -1647 -4566 -1642 -4558
rect -1638 -4566 -1633 -4558
rect -1631 -4566 -1630 -4558
rect -1626 -4566 -1625 -4558
rect -1623 -4566 -1622 -4558
rect -1547 -4566 -1546 -4558
rect -1544 -4566 -1542 -4558
rect -1538 -4566 -1536 -4558
rect -1534 -4566 -1533 -4558
rect -1521 -4566 -1520 -4558
rect -1518 -4566 -1517 -4558
rect -1513 -4566 -1512 -4558
rect -1510 -4566 -1505 -4558
rect -1501 -4566 -1496 -4558
rect -1494 -4566 -1493 -4558
rect -1489 -4566 -1488 -4558
rect -1486 -4566 -1484 -4558
rect -1480 -4566 -1478 -4558
rect -1476 -4566 -1475 -4558
rect -1471 -4566 -1470 -4558
rect -1468 -4566 -1463 -4558
rect -1459 -4566 -1454 -4558
rect -1452 -4566 -1451 -4558
rect -1447 -4566 -1446 -4558
rect -1444 -4566 -1442 -4558
rect -1438 -4566 -1436 -4558
rect -1434 -4566 -1433 -4558
rect -1429 -4566 -1428 -4558
rect -1426 -4566 -1421 -4558
rect -1417 -4566 -1412 -4558
rect -1410 -4566 -1409 -4558
rect -1405 -4566 -1404 -4558
rect -1402 -4566 -1400 -4558
rect -1396 -4566 -1394 -4558
rect -1392 -4566 -1391 -4558
rect -1387 -4566 -1386 -4558
rect -1384 -4566 -1379 -4558
rect -1375 -4566 -1370 -4558
rect -1368 -4566 -1367 -4558
rect -1363 -4566 -1362 -4558
rect -1360 -4566 -1359 -4558
rect -1230 -4566 -1229 -4558
rect -1227 -4566 -1225 -4558
rect -1221 -4566 -1219 -4558
rect -1217 -4566 -1216 -4558
rect -1204 -4566 -1203 -4558
rect -1201 -4566 -1200 -4558
rect -1196 -4566 -1195 -4558
rect -1193 -4566 -1188 -4558
rect -1184 -4566 -1179 -4558
rect -1177 -4566 -1176 -4558
rect -1172 -4566 -1171 -4558
rect -1169 -4566 -1167 -4558
rect -1163 -4566 -1161 -4558
rect -1159 -4566 -1158 -4558
rect -1154 -4566 -1153 -4558
rect -1151 -4566 -1146 -4558
rect -1142 -4566 -1137 -4558
rect -1135 -4566 -1134 -4558
rect -1130 -4566 -1129 -4558
rect -1127 -4566 -1125 -4558
rect -1121 -4566 -1119 -4558
rect -1117 -4566 -1116 -4558
rect -1112 -4566 -1111 -4558
rect -1109 -4566 -1104 -4558
rect -1100 -4566 -1095 -4558
rect -1093 -4566 -1092 -4558
rect -1088 -4566 -1087 -4558
rect -1085 -4566 -1083 -4558
rect -1079 -4566 -1077 -4558
rect -1075 -4566 -1074 -4558
rect -1070 -4566 -1069 -4558
rect -1067 -4566 -1062 -4558
rect -1058 -4566 -1053 -4558
rect -1051 -4566 -1050 -4558
rect -1046 -4566 -1045 -4558
rect -1043 -4566 -1042 -4558
rect -931 -4566 -930 -4558
rect -928 -4566 -926 -4558
rect -922 -4566 -920 -4558
rect -918 -4566 -917 -4558
rect -905 -4566 -904 -4558
rect -902 -4566 -901 -4558
rect -897 -4566 -896 -4558
rect -894 -4566 -889 -4558
rect -885 -4566 -880 -4558
rect -878 -4566 -877 -4558
rect -873 -4566 -872 -4558
rect -870 -4566 -868 -4558
rect -864 -4566 -862 -4558
rect -860 -4566 -859 -4558
rect -855 -4566 -854 -4558
rect -852 -4566 -847 -4558
rect -843 -4566 -838 -4558
rect -836 -4566 -835 -4558
rect -831 -4566 -830 -4558
rect -828 -4566 -826 -4558
rect -822 -4566 -820 -4558
rect -818 -4566 -817 -4558
rect -813 -4566 -812 -4558
rect -810 -4566 -805 -4558
rect -801 -4566 -796 -4558
rect -794 -4566 -793 -4558
rect -789 -4566 -788 -4558
rect -786 -4566 -784 -4558
rect -780 -4566 -778 -4558
rect -776 -4566 -775 -4558
rect -771 -4566 -770 -4558
rect -768 -4566 -763 -4558
rect -759 -4566 -754 -4558
rect -752 -4566 -751 -4558
rect -747 -4566 -746 -4558
rect -744 -4566 -743 -4558
rect -573 -4566 -572 -4558
rect -570 -4566 -568 -4558
rect -564 -4566 -562 -4558
rect -560 -4566 -559 -4558
rect -547 -4566 -546 -4558
rect -544 -4566 -543 -4558
rect -539 -4566 -538 -4558
rect -536 -4566 -531 -4558
rect -527 -4566 -522 -4558
rect -520 -4566 -519 -4558
rect -515 -4566 -514 -4558
rect -512 -4566 -510 -4558
rect -506 -4566 -504 -4558
rect -502 -4566 -501 -4558
rect -497 -4566 -496 -4558
rect -494 -4566 -489 -4558
rect -485 -4566 -480 -4558
rect -478 -4566 -477 -4558
rect -473 -4566 -472 -4558
rect -470 -4566 -468 -4558
rect -464 -4566 -462 -4558
rect -460 -4566 -459 -4558
rect -455 -4566 -454 -4558
rect -452 -4566 -447 -4558
rect -443 -4566 -438 -4558
rect -436 -4566 -435 -4558
rect -431 -4566 -430 -4558
rect -428 -4566 -426 -4558
rect -422 -4566 -420 -4558
rect -418 -4566 -417 -4558
rect -413 -4566 -412 -4558
rect -410 -4566 -405 -4558
rect -401 -4566 -396 -4558
rect -394 -4566 -393 -4558
rect -389 -4566 -388 -4558
rect -386 -4566 -385 -4558
rect -215 -4566 -214 -4558
rect -212 -4566 -210 -4558
rect -206 -4566 -204 -4558
rect -202 -4566 -201 -4558
rect -189 -4566 -188 -4558
rect -186 -4566 -185 -4558
rect -181 -4566 -180 -4558
rect -178 -4566 -173 -4558
rect -169 -4566 -164 -4558
rect -162 -4566 -161 -4558
rect -157 -4566 -156 -4558
rect -154 -4566 -152 -4558
rect -148 -4566 -146 -4558
rect -144 -4566 -143 -4558
rect -139 -4566 -138 -4558
rect -136 -4566 -131 -4558
rect -127 -4566 -122 -4558
rect -120 -4566 -119 -4558
rect -115 -4566 -114 -4558
rect -112 -4566 -110 -4558
rect -106 -4566 -104 -4558
rect -102 -4566 -101 -4558
rect -97 -4566 -96 -4558
rect -94 -4566 -89 -4558
rect -85 -4566 -80 -4558
rect -78 -4566 -77 -4558
rect -73 -4566 -72 -4558
rect -70 -4566 -68 -4558
rect -64 -4566 -62 -4558
rect -60 -4566 -59 -4558
rect -55 -4566 -54 -4558
rect -52 -4566 -47 -4558
rect -43 -4566 -38 -4558
rect -36 -4566 -35 -4558
rect -31 -4566 -30 -4558
rect -28 -4566 -27 -4558
rect 143 -4566 144 -4558
rect 146 -4566 148 -4558
rect 152 -4566 154 -4558
rect 156 -4566 157 -4558
rect 169 -4566 170 -4558
rect 172 -4566 173 -4558
rect 177 -4566 178 -4558
rect 180 -4566 185 -4558
rect 189 -4566 194 -4558
rect 196 -4566 197 -4558
rect 201 -4566 202 -4558
rect 204 -4566 206 -4558
rect 210 -4566 212 -4558
rect 214 -4566 215 -4558
rect 219 -4566 220 -4558
rect 222 -4566 227 -4558
rect 231 -4566 236 -4558
rect 238 -4566 239 -4558
rect 243 -4566 244 -4558
rect 246 -4566 248 -4558
rect 252 -4566 254 -4558
rect 256 -4566 257 -4558
rect 261 -4566 262 -4558
rect 264 -4566 269 -4558
rect 273 -4566 278 -4558
rect 280 -4566 281 -4558
rect 285 -4566 286 -4558
rect 288 -4566 290 -4558
rect 294 -4566 296 -4558
rect 298 -4566 299 -4558
rect 303 -4566 304 -4558
rect 306 -4566 311 -4558
rect 315 -4566 320 -4558
rect 322 -4566 323 -4558
rect 327 -4566 328 -4558
rect 330 -4566 331 -4558
rect 499 -4566 500 -4558
rect 502 -4566 504 -4558
rect 508 -4566 510 -4558
rect 512 -4566 513 -4558
rect 525 -4566 526 -4558
rect 528 -4566 529 -4558
rect 533 -4566 534 -4558
rect 536 -4566 541 -4558
rect 545 -4566 550 -4558
rect 552 -4566 553 -4558
rect 557 -4566 558 -4558
rect 560 -4566 562 -4558
rect 566 -4566 568 -4558
rect 570 -4566 571 -4558
rect 575 -4566 576 -4558
rect 578 -4566 583 -4558
rect 587 -4566 592 -4558
rect 594 -4566 595 -4558
rect 599 -4566 600 -4558
rect 602 -4566 604 -4558
rect 608 -4566 610 -4558
rect 612 -4566 613 -4558
rect 617 -4566 618 -4558
rect 620 -4566 625 -4558
rect 629 -4566 634 -4558
rect 636 -4566 637 -4558
rect 641 -4566 642 -4558
rect 644 -4566 646 -4558
rect 650 -4566 652 -4558
rect 654 -4566 655 -4558
rect 659 -4566 660 -4558
rect 662 -4566 667 -4558
rect 671 -4566 676 -4558
rect 678 -4566 679 -4558
rect 683 -4566 684 -4558
rect 686 -4566 687 -4558
rect 857 -4566 858 -4558
rect 860 -4566 862 -4558
rect 866 -4566 868 -4558
rect 870 -4566 871 -4558
rect 883 -4566 884 -4558
rect 886 -4566 887 -4558
rect 891 -4566 892 -4558
rect 894 -4566 899 -4558
rect 903 -4566 908 -4558
rect 910 -4566 911 -4558
rect 915 -4566 916 -4558
rect 918 -4566 920 -4558
rect 924 -4566 926 -4558
rect 928 -4566 929 -4558
rect 933 -4566 934 -4558
rect 936 -4566 941 -4558
rect 945 -4566 950 -4558
rect 952 -4566 953 -4558
rect 957 -4566 958 -4558
rect 960 -4566 962 -4558
rect 966 -4566 968 -4558
rect 970 -4566 971 -4558
rect 975 -4566 976 -4558
rect 978 -4566 983 -4558
rect 987 -4566 992 -4558
rect 994 -4566 995 -4558
rect 999 -4566 1000 -4558
rect 1002 -4566 1004 -4558
rect 1008 -4566 1010 -4558
rect 1012 -4566 1013 -4558
rect 1017 -4566 1018 -4558
rect 1020 -4566 1025 -4558
rect 1029 -4566 1034 -4558
rect 1036 -4566 1037 -4558
rect 1041 -4566 1042 -4558
rect 1044 -4566 1045 -4558
rect 1215 -4566 1216 -4558
rect 1218 -4566 1220 -4558
rect 1224 -4566 1226 -4558
rect 1228 -4566 1229 -4558
rect 1241 -4566 1242 -4558
rect 1244 -4566 1245 -4558
rect 1249 -4566 1250 -4558
rect 1252 -4566 1257 -4558
rect 1261 -4566 1266 -4558
rect 1268 -4566 1269 -4558
rect 1273 -4566 1274 -4558
rect 1276 -4566 1278 -4558
rect 1282 -4566 1284 -4558
rect 1286 -4566 1287 -4558
rect 1291 -4566 1292 -4558
rect 1294 -4566 1299 -4558
rect 1303 -4566 1308 -4558
rect 1310 -4566 1311 -4558
rect 1315 -4566 1316 -4558
rect 1318 -4566 1320 -4558
rect 1324 -4566 1326 -4558
rect 1328 -4566 1329 -4558
rect 1333 -4566 1334 -4558
rect 1336 -4566 1341 -4558
rect 1345 -4566 1350 -4558
rect 1352 -4566 1353 -4558
rect 1357 -4566 1358 -4558
rect 1360 -4566 1362 -4558
rect 1366 -4566 1368 -4558
rect 1370 -4566 1371 -4558
rect 1375 -4566 1376 -4558
rect 1378 -4566 1383 -4558
rect 1387 -4566 1392 -4558
rect 1394 -4566 1395 -4558
rect 1399 -4566 1400 -4558
rect 1402 -4566 1403 -4558
rect -1547 -4737 -1546 -4729
rect -1544 -4737 -1542 -4729
rect -1538 -4737 -1536 -4729
rect -1534 -4737 -1533 -4729
rect -1521 -4737 -1520 -4729
rect -1518 -4737 -1517 -4729
rect -1513 -4737 -1512 -4729
rect -1510 -4737 -1505 -4729
rect -1501 -4737 -1496 -4729
rect -1494 -4737 -1493 -4729
rect -1489 -4737 -1488 -4729
rect -1486 -4737 -1484 -4729
rect -1480 -4737 -1478 -4729
rect -1476 -4737 -1475 -4729
rect -1471 -4737 -1470 -4729
rect -1468 -4737 -1463 -4729
rect -1459 -4737 -1454 -4729
rect -1452 -4737 -1451 -4729
rect -1447 -4737 -1446 -4729
rect -1444 -4737 -1442 -4729
rect -1438 -4737 -1436 -4729
rect -1434 -4737 -1433 -4729
rect -1429 -4737 -1428 -4729
rect -1426 -4737 -1421 -4729
rect -1417 -4737 -1412 -4729
rect -1410 -4737 -1409 -4729
rect -1405 -4737 -1404 -4729
rect -1402 -4737 -1400 -4729
rect -1396 -4737 -1394 -4729
rect -1392 -4737 -1391 -4729
rect -1387 -4737 -1386 -4729
rect -1384 -4737 -1379 -4729
rect -1375 -4737 -1370 -4729
rect -1368 -4737 -1367 -4729
rect -1363 -4737 -1362 -4729
rect -1360 -4737 -1359 -4729
rect -1230 -4737 -1229 -4729
rect -1227 -4737 -1225 -4729
rect -1221 -4737 -1219 -4729
rect -1217 -4737 -1216 -4729
rect -1204 -4737 -1203 -4729
rect -1201 -4737 -1200 -4729
rect -1196 -4737 -1195 -4729
rect -1193 -4737 -1188 -4729
rect -1184 -4737 -1179 -4729
rect -1177 -4737 -1176 -4729
rect -1172 -4737 -1171 -4729
rect -1169 -4737 -1167 -4729
rect -1163 -4737 -1161 -4729
rect -1159 -4737 -1158 -4729
rect -1154 -4737 -1153 -4729
rect -1151 -4737 -1146 -4729
rect -1142 -4737 -1137 -4729
rect -1135 -4737 -1134 -4729
rect -1130 -4737 -1129 -4729
rect -1127 -4737 -1125 -4729
rect -1121 -4737 -1119 -4729
rect -1117 -4737 -1116 -4729
rect -1112 -4737 -1111 -4729
rect -1109 -4737 -1104 -4729
rect -1100 -4737 -1095 -4729
rect -1093 -4737 -1092 -4729
rect -1088 -4737 -1087 -4729
rect -1085 -4737 -1083 -4729
rect -1079 -4737 -1077 -4729
rect -1075 -4737 -1074 -4729
rect -1070 -4737 -1069 -4729
rect -1067 -4737 -1062 -4729
rect -1058 -4737 -1053 -4729
rect -1051 -4737 -1050 -4729
rect -1046 -4737 -1045 -4729
rect -1043 -4737 -1042 -4729
rect -931 -4737 -930 -4729
rect -928 -4737 -926 -4729
rect -922 -4737 -920 -4729
rect -918 -4737 -917 -4729
rect -905 -4737 -904 -4729
rect -902 -4737 -901 -4729
rect -897 -4737 -896 -4729
rect -894 -4737 -889 -4729
rect -885 -4737 -880 -4729
rect -878 -4737 -877 -4729
rect -873 -4737 -872 -4729
rect -870 -4737 -868 -4729
rect -864 -4737 -862 -4729
rect -860 -4737 -859 -4729
rect -855 -4737 -854 -4729
rect -852 -4737 -847 -4729
rect -843 -4737 -838 -4729
rect -836 -4737 -835 -4729
rect -831 -4737 -830 -4729
rect -828 -4737 -826 -4729
rect -822 -4737 -820 -4729
rect -818 -4737 -817 -4729
rect -813 -4737 -812 -4729
rect -810 -4737 -805 -4729
rect -801 -4737 -796 -4729
rect -794 -4737 -793 -4729
rect -789 -4737 -788 -4729
rect -786 -4737 -784 -4729
rect -780 -4737 -778 -4729
rect -776 -4737 -775 -4729
rect -771 -4737 -770 -4729
rect -768 -4737 -763 -4729
rect -759 -4737 -754 -4729
rect -752 -4737 -751 -4729
rect -747 -4737 -746 -4729
rect -744 -4737 -743 -4729
rect -573 -4737 -572 -4729
rect -570 -4737 -568 -4729
rect -564 -4737 -562 -4729
rect -560 -4737 -559 -4729
rect -547 -4737 -546 -4729
rect -544 -4737 -543 -4729
rect -539 -4737 -538 -4729
rect -536 -4737 -531 -4729
rect -527 -4737 -522 -4729
rect -520 -4737 -519 -4729
rect -515 -4737 -514 -4729
rect -512 -4737 -510 -4729
rect -506 -4737 -504 -4729
rect -502 -4737 -501 -4729
rect -497 -4737 -496 -4729
rect -494 -4737 -489 -4729
rect -485 -4737 -480 -4729
rect -478 -4737 -477 -4729
rect -473 -4737 -472 -4729
rect -470 -4737 -468 -4729
rect -464 -4737 -462 -4729
rect -460 -4737 -459 -4729
rect -455 -4737 -454 -4729
rect -452 -4737 -447 -4729
rect -443 -4737 -438 -4729
rect -436 -4737 -435 -4729
rect -431 -4737 -430 -4729
rect -428 -4737 -426 -4729
rect -422 -4737 -420 -4729
rect -418 -4737 -417 -4729
rect -413 -4737 -412 -4729
rect -410 -4737 -405 -4729
rect -401 -4737 -396 -4729
rect -394 -4737 -393 -4729
rect -389 -4737 -388 -4729
rect -386 -4737 -385 -4729
rect -215 -4737 -214 -4729
rect -212 -4737 -210 -4729
rect -206 -4737 -204 -4729
rect -202 -4737 -201 -4729
rect -189 -4737 -188 -4729
rect -186 -4737 -185 -4729
rect -181 -4737 -180 -4729
rect -178 -4737 -173 -4729
rect -169 -4737 -164 -4729
rect -162 -4737 -161 -4729
rect -157 -4737 -156 -4729
rect -154 -4737 -152 -4729
rect -148 -4737 -146 -4729
rect -144 -4737 -143 -4729
rect -139 -4737 -138 -4729
rect -136 -4737 -131 -4729
rect -127 -4737 -122 -4729
rect -120 -4737 -119 -4729
rect -115 -4737 -114 -4729
rect -112 -4737 -110 -4729
rect -106 -4737 -104 -4729
rect -102 -4737 -101 -4729
rect -97 -4737 -96 -4729
rect -94 -4737 -89 -4729
rect -85 -4737 -80 -4729
rect -78 -4737 -77 -4729
rect -73 -4737 -72 -4729
rect -70 -4737 -68 -4729
rect -64 -4737 -62 -4729
rect -60 -4737 -59 -4729
rect -55 -4737 -54 -4729
rect -52 -4737 -47 -4729
rect -43 -4737 -38 -4729
rect -36 -4737 -35 -4729
rect -31 -4737 -30 -4729
rect -28 -4737 -27 -4729
rect 143 -4737 144 -4729
rect 146 -4737 148 -4729
rect 152 -4737 154 -4729
rect 156 -4737 157 -4729
rect 169 -4737 170 -4729
rect 172 -4737 173 -4729
rect 177 -4737 178 -4729
rect 180 -4737 185 -4729
rect 189 -4737 194 -4729
rect 196 -4737 197 -4729
rect 201 -4737 202 -4729
rect 204 -4737 206 -4729
rect 210 -4737 212 -4729
rect 214 -4737 215 -4729
rect 219 -4737 220 -4729
rect 222 -4737 227 -4729
rect 231 -4737 236 -4729
rect 238 -4737 239 -4729
rect 243 -4737 244 -4729
rect 246 -4737 248 -4729
rect 252 -4737 254 -4729
rect 256 -4737 257 -4729
rect 261 -4737 262 -4729
rect 264 -4737 269 -4729
rect 273 -4737 278 -4729
rect 280 -4737 281 -4729
rect 285 -4737 286 -4729
rect 288 -4737 290 -4729
rect 294 -4737 296 -4729
rect 298 -4737 299 -4729
rect 303 -4737 304 -4729
rect 306 -4737 311 -4729
rect 315 -4737 320 -4729
rect 322 -4737 323 -4729
rect 327 -4737 328 -4729
rect 330 -4737 331 -4729
rect 499 -4737 500 -4729
rect 502 -4737 504 -4729
rect 508 -4737 510 -4729
rect 512 -4737 513 -4729
rect 525 -4737 526 -4729
rect 528 -4737 529 -4729
rect 533 -4737 534 -4729
rect 536 -4737 541 -4729
rect 545 -4737 550 -4729
rect 552 -4737 553 -4729
rect 557 -4737 558 -4729
rect 560 -4737 562 -4729
rect 566 -4737 568 -4729
rect 570 -4737 571 -4729
rect 575 -4737 576 -4729
rect 578 -4737 583 -4729
rect 587 -4737 592 -4729
rect 594 -4737 595 -4729
rect 599 -4737 600 -4729
rect 602 -4737 604 -4729
rect 608 -4737 610 -4729
rect 612 -4737 613 -4729
rect 617 -4737 618 -4729
rect 620 -4737 625 -4729
rect 629 -4737 634 -4729
rect 636 -4737 637 -4729
rect 641 -4737 642 -4729
rect 644 -4737 646 -4729
rect 650 -4737 652 -4729
rect 654 -4737 655 -4729
rect 659 -4737 660 -4729
rect 662 -4737 667 -4729
rect 671 -4737 676 -4729
rect 678 -4737 679 -4729
rect 683 -4737 684 -4729
rect 686 -4737 687 -4729
rect 857 -4737 858 -4729
rect 860 -4737 862 -4729
rect 866 -4737 868 -4729
rect 870 -4737 871 -4729
rect 883 -4737 884 -4729
rect 886 -4737 887 -4729
rect 891 -4737 892 -4729
rect 894 -4737 899 -4729
rect 903 -4737 908 -4729
rect 910 -4737 911 -4729
rect 915 -4737 916 -4729
rect 918 -4737 920 -4729
rect 924 -4737 926 -4729
rect 928 -4737 929 -4729
rect 933 -4737 934 -4729
rect 936 -4737 941 -4729
rect 945 -4737 950 -4729
rect 952 -4737 953 -4729
rect 957 -4737 958 -4729
rect 960 -4737 962 -4729
rect 966 -4737 968 -4729
rect 970 -4737 971 -4729
rect 975 -4737 976 -4729
rect 978 -4737 983 -4729
rect 987 -4737 992 -4729
rect 994 -4737 995 -4729
rect 999 -4737 1000 -4729
rect 1002 -4737 1004 -4729
rect 1008 -4737 1010 -4729
rect 1012 -4737 1013 -4729
rect 1017 -4737 1018 -4729
rect 1020 -4737 1025 -4729
rect 1029 -4737 1034 -4729
rect 1036 -4737 1037 -4729
rect 1041 -4737 1042 -4729
rect 1044 -4737 1045 -4729
rect 1215 -4737 1216 -4729
rect 1218 -4737 1220 -4729
rect 1224 -4737 1226 -4729
rect 1228 -4737 1229 -4729
rect 1241 -4737 1242 -4729
rect 1244 -4737 1245 -4729
rect 1249 -4737 1250 -4729
rect 1252 -4737 1257 -4729
rect 1261 -4737 1266 -4729
rect 1268 -4737 1269 -4729
rect 1273 -4737 1274 -4729
rect 1276 -4737 1278 -4729
rect 1282 -4737 1284 -4729
rect 1286 -4737 1287 -4729
rect 1291 -4737 1292 -4729
rect 1294 -4737 1299 -4729
rect 1303 -4737 1308 -4729
rect 1310 -4737 1311 -4729
rect 1315 -4737 1316 -4729
rect 1318 -4737 1320 -4729
rect 1324 -4737 1326 -4729
rect 1328 -4737 1329 -4729
rect 1333 -4737 1334 -4729
rect 1336 -4737 1341 -4729
rect 1345 -4737 1350 -4729
rect 1352 -4737 1353 -4729
rect 1357 -4737 1358 -4729
rect 1360 -4737 1362 -4729
rect 1366 -4737 1368 -4729
rect 1370 -4737 1371 -4729
rect 1375 -4737 1376 -4729
rect 1378 -4737 1383 -4729
rect 1387 -4737 1392 -4729
rect 1394 -4737 1395 -4729
rect 1399 -4737 1400 -4729
rect 1402 -4737 1403 -4729
rect -1305 -4852 -1304 -4844
rect -1302 -4852 -1301 -4844
rect -1297 -4852 -1296 -4844
rect -1294 -4852 -1292 -4844
rect -1288 -4852 -1286 -4844
rect -1284 -4852 -1283 -4844
rect -931 -4852 -930 -4844
rect -928 -4852 -927 -4844
rect -923 -4852 -922 -4844
rect -920 -4852 -918 -4844
rect -914 -4852 -912 -4844
rect -910 -4852 -909 -4844
rect -573 -4852 -572 -4844
rect -570 -4852 -569 -4844
rect -565 -4852 -564 -4844
rect -562 -4852 -560 -4844
rect -556 -4852 -554 -4844
rect -552 -4852 -551 -4844
rect -215 -4852 -214 -4844
rect -212 -4852 -211 -4844
rect -207 -4852 -206 -4844
rect -204 -4852 -202 -4844
rect -198 -4852 -196 -4844
rect -194 -4852 -193 -4844
rect 143 -4852 144 -4844
rect 146 -4852 147 -4844
rect 151 -4852 152 -4844
rect 154 -4852 156 -4844
rect 160 -4852 162 -4844
rect 164 -4852 165 -4844
rect 499 -4852 500 -4844
rect 502 -4852 503 -4844
rect 507 -4852 508 -4844
rect 510 -4852 512 -4844
rect 516 -4852 518 -4844
rect 520 -4852 521 -4844
rect 857 -4852 858 -4844
rect 860 -4852 861 -4844
rect 865 -4852 866 -4844
rect 868 -4852 870 -4844
rect 874 -4852 876 -4844
rect 878 -4852 879 -4844
rect 1215 -4852 1216 -4844
rect 1218 -4852 1219 -4844
rect 1223 -4852 1224 -4844
rect 1226 -4852 1228 -4844
rect 1232 -4852 1234 -4844
rect 1236 -4852 1237 -4844
rect -1230 -5011 -1229 -5003
rect -1227 -5011 -1225 -5003
rect -1221 -5011 -1219 -5003
rect -1217 -5011 -1216 -5003
rect -1204 -5011 -1203 -5003
rect -1201 -5011 -1193 -5003
rect -1191 -5011 -1190 -5003
rect -1186 -5011 -1185 -5003
rect -1183 -5011 -1175 -5003
rect -1173 -5011 -1168 -5003
rect -1164 -5011 -1159 -5003
rect -1157 -5011 -1156 -5003
rect -1152 -5011 -1151 -5003
rect -1149 -5011 -1147 -5003
rect -1143 -5011 -1141 -5003
rect -1139 -5011 -1138 -5003
rect -931 -5011 -930 -5003
rect -928 -5011 -926 -5003
rect -922 -5011 -920 -5003
rect -918 -5011 -917 -5003
rect -905 -5011 -904 -5003
rect -902 -5011 -900 -5003
rect -896 -5011 -894 -5003
rect -892 -5011 -891 -5003
rect -879 -5011 -878 -5003
rect -876 -5011 -868 -5003
rect -866 -5011 -865 -5003
rect -861 -5011 -860 -5003
rect -858 -5011 -850 -5003
rect -848 -5011 -843 -5003
rect -839 -5011 -834 -5003
rect -832 -5011 -831 -5003
rect -827 -5011 -826 -5003
rect -824 -5011 -822 -5003
rect -818 -5011 -816 -5003
rect -814 -5011 -813 -5003
rect -801 -5011 -800 -5003
rect -798 -5011 -790 -5003
rect -788 -5011 -787 -5003
rect -783 -5011 -782 -5003
rect -780 -5011 -772 -5003
rect -770 -5011 -765 -5003
rect -761 -5011 -756 -5003
rect -754 -5011 -753 -5003
rect -749 -5011 -748 -5003
rect -746 -5011 -741 -5003
rect -737 -5011 -732 -5003
rect -730 -5011 -729 -5003
rect -717 -5011 -716 -5003
rect -714 -5011 -708 -5003
rect -706 -5011 -704 -5003
rect -700 -5011 -698 -5003
rect -696 -5011 -695 -5003
rect -573 -5011 -572 -5003
rect -570 -5011 -568 -5003
rect -564 -5011 -562 -5003
rect -560 -5011 -559 -5003
rect -547 -5011 -546 -5003
rect -544 -5011 -542 -5003
rect -538 -5011 -536 -5003
rect -534 -5011 -533 -5003
rect -521 -5011 -520 -5003
rect -518 -5011 -510 -5003
rect -508 -5011 -507 -5003
rect -503 -5011 -502 -5003
rect -500 -5011 -492 -5003
rect -490 -5011 -485 -5003
rect -481 -5011 -476 -5003
rect -474 -5011 -473 -5003
rect -469 -5011 -468 -5003
rect -466 -5011 -464 -5003
rect -460 -5011 -458 -5003
rect -456 -5011 -455 -5003
rect -443 -5011 -442 -5003
rect -440 -5011 -432 -5003
rect -430 -5011 -429 -5003
rect -425 -5011 -424 -5003
rect -422 -5011 -414 -5003
rect -412 -5011 -407 -5003
rect -403 -5011 -398 -5003
rect -396 -5011 -395 -5003
rect -391 -5011 -390 -5003
rect -388 -5011 -383 -5003
rect -379 -5011 -374 -5003
rect -372 -5011 -371 -5003
rect -359 -5011 -358 -5003
rect -356 -5011 -350 -5003
rect -348 -5011 -346 -5003
rect -342 -5011 -340 -5003
rect -338 -5011 -337 -5003
rect -215 -5011 -214 -5003
rect -212 -5011 -210 -5003
rect -206 -5011 -204 -5003
rect -202 -5011 -201 -5003
rect -189 -5011 -188 -5003
rect -186 -5011 -184 -5003
rect -180 -5011 -178 -5003
rect -176 -5011 -175 -5003
rect -163 -5011 -162 -5003
rect -160 -5011 -152 -5003
rect -150 -5011 -149 -5003
rect -145 -5011 -144 -5003
rect -142 -5011 -134 -5003
rect -132 -5011 -127 -5003
rect -123 -5011 -118 -5003
rect -116 -5011 -115 -5003
rect -111 -5011 -110 -5003
rect -108 -5011 -106 -5003
rect -102 -5011 -100 -5003
rect -98 -5011 -97 -5003
rect -85 -5011 -84 -5003
rect -82 -5011 -74 -5003
rect -72 -5011 -71 -5003
rect -67 -5011 -66 -5003
rect -64 -5011 -56 -5003
rect -54 -5011 -49 -5003
rect -45 -5011 -40 -5003
rect -38 -5011 -37 -5003
rect -33 -5011 -32 -5003
rect -30 -5011 -25 -5003
rect -21 -5011 -16 -5003
rect -14 -5011 -13 -5003
rect -1 -5011 0 -5003
rect 2 -5011 8 -5003
rect 10 -5011 12 -5003
rect 16 -5011 18 -5003
rect 20 -5011 21 -5003
rect 143 -5011 144 -5003
rect 146 -5011 148 -5003
rect 152 -5011 154 -5003
rect 156 -5011 157 -5003
rect 169 -5011 170 -5003
rect 172 -5011 174 -5003
rect 178 -5011 180 -5003
rect 182 -5011 183 -5003
rect 195 -5011 196 -5003
rect 198 -5011 206 -5003
rect 208 -5011 209 -5003
rect 213 -5011 214 -5003
rect 216 -5011 224 -5003
rect 226 -5011 231 -5003
rect 235 -5011 240 -5003
rect 242 -5011 243 -5003
rect 247 -5011 248 -5003
rect 250 -5011 252 -5003
rect 256 -5011 258 -5003
rect 260 -5011 261 -5003
rect 273 -5011 274 -5003
rect 276 -5011 284 -5003
rect 286 -5011 287 -5003
rect 291 -5011 292 -5003
rect 294 -5011 302 -5003
rect 304 -5011 309 -5003
rect 313 -5011 318 -5003
rect 320 -5011 321 -5003
rect 325 -5011 326 -5003
rect 328 -5011 333 -5003
rect 337 -5011 342 -5003
rect 344 -5011 345 -5003
rect 357 -5011 358 -5003
rect 360 -5011 366 -5003
rect 368 -5011 370 -5003
rect 374 -5011 376 -5003
rect 378 -5011 379 -5003
rect 499 -5011 500 -5003
rect 502 -5011 504 -5003
rect 508 -5011 510 -5003
rect 512 -5011 513 -5003
rect 525 -5011 526 -5003
rect 528 -5011 530 -5003
rect 534 -5011 536 -5003
rect 538 -5011 539 -5003
rect 551 -5011 552 -5003
rect 554 -5011 562 -5003
rect 564 -5011 565 -5003
rect 569 -5011 570 -5003
rect 572 -5011 580 -5003
rect 582 -5011 587 -5003
rect 591 -5011 596 -5003
rect 598 -5011 599 -5003
rect 603 -5011 604 -5003
rect 606 -5011 608 -5003
rect 612 -5011 614 -5003
rect 616 -5011 617 -5003
rect 629 -5011 630 -5003
rect 632 -5011 640 -5003
rect 642 -5011 643 -5003
rect 647 -5011 648 -5003
rect 650 -5011 658 -5003
rect 660 -5011 665 -5003
rect 669 -5011 674 -5003
rect 676 -5011 677 -5003
rect 681 -5011 682 -5003
rect 684 -5011 689 -5003
rect 693 -5011 698 -5003
rect 700 -5011 701 -5003
rect 713 -5011 714 -5003
rect 716 -5011 722 -5003
rect 724 -5011 726 -5003
rect 730 -5011 732 -5003
rect 734 -5011 735 -5003
rect 857 -5011 858 -5003
rect 860 -5011 862 -5003
rect 866 -5011 868 -5003
rect 870 -5011 871 -5003
rect 883 -5011 884 -5003
rect 886 -5011 888 -5003
rect 892 -5011 894 -5003
rect 896 -5011 897 -5003
rect 909 -5011 910 -5003
rect 912 -5011 920 -5003
rect 922 -5011 923 -5003
rect 927 -5011 928 -5003
rect 930 -5011 938 -5003
rect 940 -5011 945 -5003
rect 949 -5011 954 -5003
rect 956 -5011 957 -5003
rect 961 -5011 962 -5003
rect 964 -5011 966 -5003
rect 970 -5011 972 -5003
rect 974 -5011 975 -5003
rect 987 -5011 988 -5003
rect 990 -5011 998 -5003
rect 1000 -5011 1001 -5003
rect 1005 -5011 1006 -5003
rect 1008 -5011 1016 -5003
rect 1018 -5011 1023 -5003
rect 1027 -5011 1032 -5003
rect 1034 -5011 1035 -5003
rect 1039 -5011 1040 -5003
rect 1042 -5011 1047 -5003
rect 1051 -5011 1056 -5003
rect 1058 -5011 1059 -5003
rect 1071 -5011 1072 -5003
rect 1074 -5011 1080 -5003
rect 1082 -5011 1084 -5003
rect 1088 -5011 1090 -5003
rect 1092 -5011 1093 -5003
rect 1215 -5011 1216 -5003
rect 1218 -5011 1220 -5003
rect 1224 -5011 1226 -5003
rect 1228 -5011 1229 -5003
rect 1241 -5011 1242 -5003
rect 1244 -5011 1246 -5003
rect 1250 -5011 1252 -5003
rect 1254 -5011 1255 -5003
rect 1267 -5011 1268 -5003
rect 1270 -5011 1278 -5003
rect 1280 -5011 1281 -5003
rect 1285 -5011 1286 -5003
rect 1288 -5011 1296 -5003
rect 1298 -5011 1303 -5003
rect 1307 -5011 1312 -5003
rect 1314 -5011 1315 -5003
rect 1319 -5011 1320 -5003
rect 1322 -5011 1324 -5003
rect 1328 -5011 1330 -5003
rect 1332 -5011 1333 -5003
rect 1345 -5011 1346 -5003
rect 1348 -5011 1356 -5003
rect 1358 -5011 1359 -5003
rect 1363 -5011 1364 -5003
rect 1366 -5011 1374 -5003
rect 1376 -5011 1381 -5003
rect 1385 -5011 1390 -5003
rect 1392 -5011 1393 -5003
rect 1397 -5011 1398 -5003
rect 1400 -5011 1405 -5003
rect 1409 -5011 1414 -5003
rect 1416 -5011 1417 -5003
rect 1429 -5011 1430 -5003
rect 1432 -5011 1438 -5003
rect 1440 -5011 1442 -5003
rect 1446 -5011 1448 -5003
rect 1450 -5011 1451 -5003
rect -1806 -5130 -1805 -5122
rect -1803 -5130 -1801 -5122
rect -1797 -5130 -1795 -5122
rect -1793 -5130 -1792 -5122
rect -1780 -5130 -1779 -5122
rect -1777 -5130 -1776 -5122
rect -1772 -5130 -1771 -5122
rect -1769 -5130 -1764 -5122
rect -1760 -5130 -1755 -5122
rect -1753 -5130 -1752 -5122
rect -1748 -5130 -1747 -5122
rect -1745 -5130 -1743 -5122
rect -1739 -5130 -1737 -5122
rect -1735 -5130 -1734 -5122
rect -1730 -5130 -1729 -5122
rect -1727 -5130 -1722 -5122
rect -1718 -5130 -1713 -5122
rect -1711 -5130 -1710 -5122
rect -1706 -5130 -1705 -5122
rect -1703 -5130 -1701 -5122
rect -1697 -5130 -1695 -5122
rect -1693 -5130 -1692 -5122
rect -1688 -5130 -1687 -5122
rect -1685 -5130 -1680 -5122
rect -1676 -5130 -1671 -5122
rect -1669 -5130 -1668 -5122
rect -1664 -5130 -1663 -5122
rect -1661 -5130 -1659 -5122
rect -1655 -5130 -1653 -5122
rect -1651 -5130 -1650 -5122
rect -1646 -5130 -1645 -5122
rect -1643 -5130 -1638 -5122
rect -1634 -5130 -1629 -5122
rect -1627 -5130 -1626 -5122
rect -1622 -5130 -1621 -5122
rect -1619 -5130 -1618 -5122
rect -1543 -5130 -1542 -5122
rect -1540 -5130 -1538 -5122
rect -1534 -5130 -1532 -5122
rect -1530 -5130 -1529 -5122
rect -1517 -5130 -1516 -5122
rect -1514 -5130 -1513 -5122
rect -1509 -5130 -1508 -5122
rect -1506 -5130 -1501 -5122
rect -1497 -5130 -1492 -5122
rect -1490 -5130 -1489 -5122
rect -1485 -5130 -1484 -5122
rect -1482 -5130 -1480 -5122
rect -1476 -5130 -1474 -5122
rect -1472 -5130 -1471 -5122
rect -1467 -5130 -1466 -5122
rect -1464 -5130 -1459 -5122
rect -1455 -5130 -1450 -5122
rect -1448 -5130 -1447 -5122
rect -1443 -5130 -1442 -5122
rect -1440 -5130 -1438 -5122
rect -1434 -5130 -1432 -5122
rect -1430 -5130 -1429 -5122
rect -1425 -5130 -1424 -5122
rect -1422 -5130 -1417 -5122
rect -1413 -5130 -1408 -5122
rect -1406 -5130 -1405 -5122
rect -1401 -5130 -1400 -5122
rect -1398 -5130 -1396 -5122
rect -1392 -5130 -1390 -5122
rect -1388 -5130 -1387 -5122
rect -1383 -5130 -1382 -5122
rect -1380 -5130 -1375 -5122
rect -1371 -5130 -1366 -5122
rect -1364 -5130 -1363 -5122
rect -1359 -5130 -1358 -5122
rect -1356 -5130 -1355 -5122
rect -1230 -5130 -1229 -5122
rect -1227 -5130 -1225 -5122
rect -1221 -5130 -1219 -5122
rect -1217 -5130 -1216 -5122
rect -1204 -5130 -1203 -5122
rect -1201 -5130 -1200 -5122
rect -1196 -5130 -1195 -5122
rect -1193 -5130 -1188 -5122
rect -1184 -5130 -1179 -5122
rect -1177 -5130 -1176 -5122
rect -1172 -5130 -1171 -5122
rect -1169 -5130 -1167 -5122
rect -1163 -5130 -1161 -5122
rect -1159 -5130 -1158 -5122
rect -1154 -5130 -1153 -5122
rect -1151 -5130 -1146 -5122
rect -1142 -5130 -1137 -5122
rect -1135 -5130 -1134 -5122
rect -1130 -5130 -1129 -5122
rect -1127 -5130 -1125 -5122
rect -1121 -5130 -1119 -5122
rect -1117 -5130 -1116 -5122
rect -1112 -5130 -1111 -5122
rect -1109 -5130 -1104 -5122
rect -1100 -5130 -1095 -5122
rect -1093 -5130 -1092 -5122
rect -1088 -5130 -1087 -5122
rect -1085 -5130 -1083 -5122
rect -1079 -5130 -1077 -5122
rect -1075 -5130 -1074 -5122
rect -1070 -5130 -1069 -5122
rect -1067 -5130 -1062 -5122
rect -1058 -5130 -1053 -5122
rect -1051 -5130 -1050 -5122
rect -1046 -5130 -1045 -5122
rect -1043 -5130 -1042 -5122
rect -931 -5130 -930 -5122
rect -928 -5130 -926 -5122
rect -922 -5130 -920 -5122
rect -918 -5130 -917 -5122
rect -905 -5130 -904 -5122
rect -902 -5130 -901 -5122
rect -897 -5130 -896 -5122
rect -894 -5130 -889 -5122
rect -885 -5130 -880 -5122
rect -878 -5130 -877 -5122
rect -873 -5130 -872 -5122
rect -870 -5130 -868 -5122
rect -864 -5130 -862 -5122
rect -860 -5130 -859 -5122
rect -855 -5130 -854 -5122
rect -852 -5130 -847 -5122
rect -843 -5130 -838 -5122
rect -836 -5130 -835 -5122
rect -831 -5130 -830 -5122
rect -828 -5130 -826 -5122
rect -822 -5130 -820 -5122
rect -818 -5130 -817 -5122
rect -813 -5130 -812 -5122
rect -810 -5130 -805 -5122
rect -801 -5130 -796 -5122
rect -794 -5130 -793 -5122
rect -789 -5130 -788 -5122
rect -786 -5130 -784 -5122
rect -780 -5130 -778 -5122
rect -776 -5130 -775 -5122
rect -771 -5130 -770 -5122
rect -768 -5130 -763 -5122
rect -759 -5130 -754 -5122
rect -752 -5130 -751 -5122
rect -747 -5130 -746 -5122
rect -744 -5130 -743 -5122
rect -1806 -5301 -1805 -5293
rect -1803 -5301 -1801 -5293
rect -1797 -5301 -1795 -5293
rect -1793 -5301 -1792 -5293
rect -1780 -5301 -1779 -5293
rect -1777 -5301 -1776 -5293
rect -1772 -5301 -1771 -5293
rect -1769 -5301 -1764 -5293
rect -1760 -5301 -1755 -5293
rect -1753 -5301 -1752 -5293
rect -1748 -5301 -1747 -5293
rect -1745 -5301 -1743 -5293
rect -1739 -5301 -1737 -5293
rect -1735 -5301 -1734 -5293
rect -1730 -5301 -1729 -5293
rect -1727 -5301 -1722 -5293
rect -1718 -5301 -1713 -5293
rect -1711 -5301 -1710 -5293
rect -1706 -5301 -1705 -5293
rect -1703 -5301 -1701 -5293
rect -1697 -5301 -1695 -5293
rect -1693 -5301 -1692 -5293
rect -1688 -5301 -1687 -5293
rect -1685 -5301 -1680 -5293
rect -1676 -5301 -1671 -5293
rect -1669 -5301 -1668 -5293
rect -1664 -5301 -1663 -5293
rect -1661 -5301 -1659 -5293
rect -1655 -5301 -1653 -5293
rect -1651 -5301 -1650 -5293
rect -1646 -5301 -1645 -5293
rect -1643 -5301 -1638 -5293
rect -1634 -5301 -1629 -5293
rect -1627 -5301 -1626 -5293
rect -1622 -5301 -1621 -5293
rect -1619 -5301 -1618 -5293
rect -1543 -5301 -1542 -5293
rect -1540 -5301 -1538 -5293
rect -1534 -5301 -1532 -5293
rect -1530 -5301 -1529 -5293
rect -1517 -5301 -1516 -5293
rect -1514 -5301 -1513 -5293
rect -1509 -5301 -1508 -5293
rect -1506 -5301 -1501 -5293
rect -1497 -5301 -1492 -5293
rect -1490 -5301 -1489 -5293
rect -1485 -5301 -1484 -5293
rect -1482 -5301 -1480 -5293
rect -1476 -5301 -1474 -5293
rect -1472 -5301 -1471 -5293
rect -1467 -5301 -1466 -5293
rect -1464 -5301 -1459 -5293
rect -1455 -5301 -1450 -5293
rect -1448 -5301 -1447 -5293
rect -1443 -5301 -1442 -5293
rect -1440 -5301 -1438 -5293
rect -1434 -5301 -1432 -5293
rect -1430 -5301 -1429 -5293
rect -1425 -5301 -1424 -5293
rect -1422 -5301 -1417 -5293
rect -1413 -5301 -1408 -5293
rect -1406 -5301 -1405 -5293
rect -1401 -5301 -1400 -5293
rect -1398 -5301 -1396 -5293
rect -1392 -5301 -1390 -5293
rect -1388 -5301 -1387 -5293
rect -1383 -5301 -1382 -5293
rect -1380 -5301 -1375 -5293
rect -1371 -5301 -1366 -5293
rect -1364 -5301 -1363 -5293
rect -1359 -5301 -1358 -5293
rect -1356 -5301 -1355 -5293
rect -1230 -5301 -1229 -5293
rect -1227 -5301 -1225 -5293
rect -1221 -5301 -1219 -5293
rect -1217 -5301 -1216 -5293
rect -1204 -5301 -1203 -5293
rect -1201 -5301 -1200 -5293
rect -1196 -5301 -1195 -5293
rect -1193 -5301 -1188 -5293
rect -1184 -5301 -1179 -5293
rect -1177 -5301 -1176 -5293
rect -1172 -5301 -1171 -5293
rect -1169 -5301 -1167 -5293
rect -1163 -5301 -1161 -5293
rect -1159 -5301 -1158 -5293
rect -1154 -5301 -1153 -5293
rect -1151 -5301 -1146 -5293
rect -1142 -5301 -1137 -5293
rect -1135 -5301 -1134 -5293
rect -1130 -5301 -1129 -5293
rect -1127 -5301 -1125 -5293
rect -1121 -5301 -1119 -5293
rect -1117 -5301 -1116 -5293
rect -1112 -5301 -1111 -5293
rect -1109 -5301 -1104 -5293
rect -1100 -5301 -1095 -5293
rect -1093 -5301 -1092 -5293
rect -1088 -5301 -1087 -5293
rect -1085 -5301 -1083 -5293
rect -1079 -5301 -1077 -5293
rect -1075 -5301 -1074 -5293
rect -1070 -5301 -1069 -5293
rect -1067 -5301 -1062 -5293
rect -1058 -5301 -1053 -5293
rect -1051 -5301 -1050 -5293
rect -1046 -5301 -1045 -5293
rect -1043 -5301 -1042 -5293
rect -931 -5301 -930 -5293
rect -928 -5301 -926 -5293
rect -922 -5301 -920 -5293
rect -918 -5301 -917 -5293
rect -905 -5301 -904 -5293
rect -902 -5301 -901 -5293
rect -897 -5301 -896 -5293
rect -894 -5301 -889 -5293
rect -885 -5301 -880 -5293
rect -878 -5301 -877 -5293
rect -873 -5301 -872 -5293
rect -870 -5301 -868 -5293
rect -864 -5301 -862 -5293
rect -860 -5301 -859 -5293
rect -855 -5301 -854 -5293
rect -852 -5301 -847 -5293
rect -843 -5301 -838 -5293
rect -836 -5301 -835 -5293
rect -831 -5301 -830 -5293
rect -828 -5301 -826 -5293
rect -822 -5301 -820 -5293
rect -818 -5301 -817 -5293
rect -813 -5301 -812 -5293
rect -810 -5301 -805 -5293
rect -801 -5301 -796 -5293
rect -794 -5301 -793 -5293
rect -789 -5301 -788 -5293
rect -786 -5301 -784 -5293
rect -780 -5301 -778 -5293
rect -776 -5301 -775 -5293
rect -771 -5301 -770 -5293
rect -768 -5301 -763 -5293
rect -759 -5301 -754 -5293
rect -752 -5301 -751 -5293
rect -747 -5301 -746 -5293
rect -744 -5301 -743 -5293
rect -573 -5301 -572 -5293
rect -570 -5301 -568 -5293
rect -564 -5301 -562 -5293
rect -560 -5301 -559 -5293
rect -547 -5301 -546 -5293
rect -544 -5301 -543 -5293
rect -539 -5301 -538 -5293
rect -536 -5301 -531 -5293
rect -527 -5301 -522 -5293
rect -520 -5301 -519 -5293
rect -515 -5301 -514 -5293
rect -512 -5301 -510 -5293
rect -506 -5301 -504 -5293
rect -502 -5301 -501 -5293
rect -497 -5301 -496 -5293
rect -494 -5301 -489 -5293
rect -485 -5301 -480 -5293
rect -478 -5301 -477 -5293
rect -473 -5301 -472 -5293
rect -470 -5301 -468 -5293
rect -464 -5301 -462 -5293
rect -460 -5301 -459 -5293
rect -455 -5301 -454 -5293
rect -452 -5301 -447 -5293
rect -443 -5301 -438 -5293
rect -436 -5301 -435 -5293
rect -431 -5301 -430 -5293
rect -428 -5301 -426 -5293
rect -422 -5301 -420 -5293
rect -418 -5301 -417 -5293
rect -413 -5301 -412 -5293
rect -410 -5301 -405 -5293
rect -401 -5301 -396 -5293
rect -394 -5301 -393 -5293
rect -389 -5301 -388 -5293
rect -386 -5301 -385 -5293
rect -215 -5301 -214 -5293
rect -212 -5301 -210 -5293
rect -206 -5301 -204 -5293
rect -202 -5301 -201 -5293
rect -189 -5301 -188 -5293
rect -186 -5301 -185 -5293
rect -181 -5301 -180 -5293
rect -178 -5301 -173 -5293
rect -169 -5301 -164 -5293
rect -162 -5301 -161 -5293
rect -157 -5301 -156 -5293
rect -154 -5301 -152 -5293
rect -148 -5301 -146 -5293
rect -144 -5301 -143 -5293
rect -139 -5301 -138 -5293
rect -136 -5301 -131 -5293
rect -127 -5301 -122 -5293
rect -120 -5301 -119 -5293
rect -115 -5301 -114 -5293
rect -112 -5301 -110 -5293
rect -106 -5301 -104 -5293
rect -102 -5301 -101 -5293
rect -97 -5301 -96 -5293
rect -94 -5301 -89 -5293
rect -85 -5301 -80 -5293
rect -78 -5301 -77 -5293
rect -73 -5301 -72 -5293
rect -70 -5301 -68 -5293
rect -64 -5301 -62 -5293
rect -60 -5301 -59 -5293
rect -55 -5301 -54 -5293
rect -52 -5301 -47 -5293
rect -43 -5301 -38 -5293
rect -36 -5301 -35 -5293
rect -31 -5301 -30 -5293
rect -28 -5301 -27 -5293
rect 143 -5301 144 -5293
rect 146 -5301 148 -5293
rect 152 -5301 154 -5293
rect 156 -5301 157 -5293
rect 169 -5301 170 -5293
rect 172 -5301 173 -5293
rect 177 -5301 178 -5293
rect 180 -5301 185 -5293
rect 189 -5301 194 -5293
rect 196 -5301 197 -5293
rect 201 -5301 202 -5293
rect 204 -5301 206 -5293
rect 210 -5301 212 -5293
rect 214 -5301 215 -5293
rect 219 -5301 220 -5293
rect 222 -5301 227 -5293
rect 231 -5301 236 -5293
rect 238 -5301 239 -5293
rect 243 -5301 244 -5293
rect 246 -5301 248 -5293
rect 252 -5301 254 -5293
rect 256 -5301 257 -5293
rect 261 -5301 262 -5293
rect 264 -5301 269 -5293
rect 273 -5301 278 -5293
rect 280 -5301 281 -5293
rect 285 -5301 286 -5293
rect 288 -5301 290 -5293
rect 294 -5301 296 -5293
rect 298 -5301 299 -5293
rect 303 -5301 304 -5293
rect 306 -5301 311 -5293
rect 315 -5301 320 -5293
rect 322 -5301 323 -5293
rect 327 -5301 328 -5293
rect 330 -5301 331 -5293
rect 499 -5301 500 -5293
rect 502 -5301 504 -5293
rect 508 -5301 510 -5293
rect 512 -5301 513 -5293
rect 525 -5301 526 -5293
rect 528 -5301 529 -5293
rect 533 -5301 534 -5293
rect 536 -5301 541 -5293
rect 545 -5301 550 -5293
rect 552 -5301 553 -5293
rect 557 -5301 558 -5293
rect 560 -5301 562 -5293
rect 566 -5301 568 -5293
rect 570 -5301 571 -5293
rect 575 -5301 576 -5293
rect 578 -5301 583 -5293
rect 587 -5301 592 -5293
rect 594 -5301 595 -5293
rect 599 -5301 600 -5293
rect 602 -5301 604 -5293
rect 608 -5301 610 -5293
rect 612 -5301 613 -5293
rect 617 -5301 618 -5293
rect 620 -5301 625 -5293
rect 629 -5301 634 -5293
rect 636 -5301 637 -5293
rect 641 -5301 642 -5293
rect 644 -5301 646 -5293
rect 650 -5301 652 -5293
rect 654 -5301 655 -5293
rect 659 -5301 660 -5293
rect 662 -5301 667 -5293
rect 671 -5301 676 -5293
rect 678 -5301 679 -5293
rect 683 -5301 684 -5293
rect 686 -5301 687 -5293
rect 857 -5301 858 -5293
rect 860 -5301 862 -5293
rect 866 -5301 868 -5293
rect 870 -5301 871 -5293
rect 883 -5301 884 -5293
rect 886 -5301 887 -5293
rect 891 -5301 892 -5293
rect 894 -5301 899 -5293
rect 903 -5301 908 -5293
rect 910 -5301 911 -5293
rect 915 -5301 916 -5293
rect 918 -5301 920 -5293
rect 924 -5301 926 -5293
rect 928 -5301 929 -5293
rect 933 -5301 934 -5293
rect 936 -5301 941 -5293
rect 945 -5301 950 -5293
rect 952 -5301 953 -5293
rect 957 -5301 958 -5293
rect 960 -5301 962 -5293
rect 966 -5301 968 -5293
rect 970 -5301 971 -5293
rect 975 -5301 976 -5293
rect 978 -5301 983 -5293
rect 987 -5301 992 -5293
rect 994 -5301 995 -5293
rect 999 -5301 1000 -5293
rect 1002 -5301 1004 -5293
rect 1008 -5301 1010 -5293
rect 1012 -5301 1013 -5293
rect 1017 -5301 1018 -5293
rect 1020 -5301 1025 -5293
rect 1029 -5301 1034 -5293
rect 1036 -5301 1037 -5293
rect 1041 -5301 1042 -5293
rect 1044 -5301 1045 -5293
rect 1215 -5301 1216 -5293
rect 1218 -5301 1220 -5293
rect 1224 -5301 1226 -5293
rect 1228 -5301 1229 -5293
rect 1241 -5301 1242 -5293
rect 1244 -5301 1245 -5293
rect 1249 -5301 1250 -5293
rect 1252 -5301 1257 -5293
rect 1261 -5301 1266 -5293
rect 1268 -5301 1269 -5293
rect 1273 -5301 1274 -5293
rect 1276 -5301 1278 -5293
rect 1282 -5301 1284 -5293
rect 1286 -5301 1287 -5293
rect 1291 -5301 1292 -5293
rect 1294 -5301 1299 -5293
rect 1303 -5301 1308 -5293
rect 1310 -5301 1311 -5293
rect 1315 -5301 1316 -5293
rect 1318 -5301 1320 -5293
rect 1324 -5301 1326 -5293
rect 1328 -5301 1329 -5293
rect 1333 -5301 1334 -5293
rect 1336 -5301 1341 -5293
rect 1345 -5301 1350 -5293
rect 1352 -5301 1353 -5293
rect 1357 -5301 1358 -5293
rect 1360 -5301 1362 -5293
rect 1366 -5301 1368 -5293
rect 1370 -5301 1371 -5293
rect 1375 -5301 1376 -5293
rect 1378 -5301 1383 -5293
rect 1387 -5301 1392 -5293
rect 1394 -5301 1395 -5293
rect 1399 -5301 1400 -5293
rect 1402 -5301 1403 -5293
rect -1806 -5461 -1805 -5453
rect -1803 -5461 -1801 -5453
rect -1797 -5461 -1795 -5453
rect -1793 -5461 -1792 -5453
rect -1780 -5461 -1779 -5453
rect -1777 -5461 -1776 -5453
rect -1772 -5461 -1771 -5453
rect -1769 -5461 -1764 -5453
rect -1760 -5461 -1755 -5453
rect -1753 -5461 -1752 -5453
rect -1748 -5461 -1747 -5453
rect -1745 -5461 -1743 -5453
rect -1739 -5461 -1737 -5453
rect -1735 -5461 -1734 -5453
rect -1730 -5461 -1729 -5453
rect -1727 -5461 -1722 -5453
rect -1718 -5461 -1713 -5453
rect -1711 -5461 -1710 -5453
rect -1706 -5461 -1705 -5453
rect -1703 -5461 -1701 -5453
rect -1697 -5461 -1695 -5453
rect -1693 -5461 -1692 -5453
rect -1688 -5461 -1687 -5453
rect -1685 -5461 -1680 -5453
rect -1676 -5461 -1671 -5453
rect -1669 -5461 -1668 -5453
rect -1664 -5461 -1663 -5453
rect -1661 -5461 -1659 -5453
rect -1655 -5461 -1653 -5453
rect -1651 -5461 -1650 -5453
rect -1646 -5461 -1645 -5453
rect -1643 -5461 -1638 -5453
rect -1634 -5461 -1629 -5453
rect -1627 -5461 -1626 -5453
rect -1622 -5461 -1621 -5453
rect -1619 -5461 -1618 -5453
rect -1543 -5461 -1542 -5453
rect -1540 -5461 -1538 -5453
rect -1534 -5461 -1532 -5453
rect -1530 -5461 -1529 -5453
rect -1517 -5461 -1516 -5453
rect -1514 -5461 -1513 -5453
rect -1509 -5461 -1508 -5453
rect -1506 -5461 -1501 -5453
rect -1497 -5461 -1492 -5453
rect -1490 -5461 -1489 -5453
rect -1485 -5461 -1484 -5453
rect -1482 -5461 -1480 -5453
rect -1476 -5461 -1474 -5453
rect -1472 -5461 -1471 -5453
rect -1467 -5461 -1466 -5453
rect -1464 -5461 -1459 -5453
rect -1455 -5461 -1450 -5453
rect -1448 -5461 -1447 -5453
rect -1443 -5461 -1442 -5453
rect -1440 -5461 -1438 -5453
rect -1434 -5461 -1432 -5453
rect -1430 -5461 -1429 -5453
rect -1425 -5461 -1424 -5453
rect -1422 -5461 -1417 -5453
rect -1413 -5461 -1408 -5453
rect -1406 -5461 -1405 -5453
rect -1401 -5461 -1400 -5453
rect -1398 -5461 -1396 -5453
rect -1392 -5461 -1390 -5453
rect -1388 -5461 -1387 -5453
rect -1383 -5461 -1382 -5453
rect -1380 -5461 -1375 -5453
rect -1371 -5461 -1366 -5453
rect -1364 -5461 -1363 -5453
rect -1359 -5461 -1358 -5453
rect -1356 -5461 -1355 -5453
rect -1230 -5461 -1229 -5453
rect -1227 -5461 -1225 -5453
rect -1221 -5461 -1219 -5453
rect -1217 -5461 -1216 -5453
rect -1204 -5461 -1203 -5453
rect -1201 -5461 -1200 -5453
rect -1196 -5461 -1195 -5453
rect -1193 -5461 -1188 -5453
rect -1184 -5461 -1179 -5453
rect -1177 -5461 -1176 -5453
rect -1172 -5461 -1171 -5453
rect -1169 -5461 -1167 -5453
rect -1163 -5461 -1161 -5453
rect -1159 -5461 -1158 -5453
rect -1154 -5461 -1153 -5453
rect -1151 -5461 -1146 -5453
rect -1142 -5461 -1137 -5453
rect -1135 -5461 -1134 -5453
rect -1130 -5461 -1129 -5453
rect -1127 -5461 -1125 -5453
rect -1121 -5461 -1119 -5453
rect -1117 -5461 -1116 -5453
rect -1112 -5461 -1111 -5453
rect -1109 -5461 -1104 -5453
rect -1100 -5461 -1095 -5453
rect -1093 -5461 -1092 -5453
rect -1088 -5461 -1087 -5453
rect -1085 -5461 -1083 -5453
rect -1079 -5461 -1077 -5453
rect -1075 -5461 -1074 -5453
rect -1070 -5461 -1069 -5453
rect -1067 -5461 -1062 -5453
rect -1058 -5461 -1053 -5453
rect -1051 -5461 -1050 -5453
rect -1046 -5461 -1045 -5453
rect -1043 -5461 -1042 -5453
rect -931 -5461 -930 -5453
rect -928 -5461 -926 -5453
rect -922 -5461 -920 -5453
rect -918 -5461 -917 -5453
rect -905 -5461 -904 -5453
rect -902 -5461 -901 -5453
rect -897 -5461 -896 -5453
rect -894 -5461 -889 -5453
rect -885 -5461 -880 -5453
rect -878 -5461 -877 -5453
rect -873 -5461 -872 -5453
rect -870 -5461 -868 -5453
rect -864 -5461 -862 -5453
rect -860 -5461 -859 -5453
rect -855 -5461 -854 -5453
rect -852 -5461 -847 -5453
rect -843 -5461 -838 -5453
rect -836 -5461 -835 -5453
rect -831 -5461 -830 -5453
rect -828 -5461 -826 -5453
rect -822 -5461 -820 -5453
rect -818 -5461 -817 -5453
rect -813 -5461 -812 -5453
rect -810 -5461 -805 -5453
rect -801 -5461 -796 -5453
rect -794 -5461 -793 -5453
rect -789 -5461 -788 -5453
rect -786 -5461 -784 -5453
rect -780 -5461 -778 -5453
rect -776 -5461 -775 -5453
rect -771 -5461 -770 -5453
rect -768 -5461 -763 -5453
rect -759 -5461 -754 -5453
rect -752 -5461 -751 -5453
rect -747 -5461 -746 -5453
rect -744 -5461 -743 -5453
rect -573 -5461 -572 -5453
rect -570 -5461 -568 -5453
rect -564 -5461 -562 -5453
rect -560 -5461 -559 -5453
rect -547 -5461 -546 -5453
rect -544 -5461 -543 -5453
rect -539 -5461 -538 -5453
rect -536 -5461 -531 -5453
rect -527 -5461 -522 -5453
rect -520 -5461 -519 -5453
rect -515 -5461 -514 -5453
rect -512 -5461 -510 -5453
rect -506 -5461 -504 -5453
rect -502 -5461 -501 -5453
rect -497 -5461 -496 -5453
rect -494 -5461 -489 -5453
rect -485 -5461 -480 -5453
rect -478 -5461 -477 -5453
rect -473 -5461 -472 -5453
rect -470 -5461 -468 -5453
rect -464 -5461 -462 -5453
rect -460 -5461 -459 -5453
rect -455 -5461 -454 -5453
rect -452 -5461 -447 -5453
rect -443 -5461 -438 -5453
rect -436 -5461 -435 -5453
rect -431 -5461 -430 -5453
rect -428 -5461 -426 -5453
rect -422 -5461 -420 -5453
rect -418 -5461 -417 -5453
rect -413 -5461 -412 -5453
rect -410 -5461 -405 -5453
rect -401 -5461 -396 -5453
rect -394 -5461 -393 -5453
rect -389 -5461 -388 -5453
rect -386 -5461 -385 -5453
rect -215 -5461 -214 -5453
rect -212 -5461 -210 -5453
rect -206 -5461 -204 -5453
rect -202 -5461 -201 -5453
rect -189 -5461 -188 -5453
rect -186 -5461 -185 -5453
rect -181 -5461 -180 -5453
rect -178 -5461 -173 -5453
rect -169 -5461 -164 -5453
rect -162 -5461 -161 -5453
rect -157 -5461 -156 -5453
rect -154 -5461 -152 -5453
rect -148 -5461 -146 -5453
rect -144 -5461 -143 -5453
rect -139 -5461 -138 -5453
rect -136 -5461 -131 -5453
rect -127 -5461 -122 -5453
rect -120 -5461 -119 -5453
rect -115 -5461 -114 -5453
rect -112 -5461 -110 -5453
rect -106 -5461 -104 -5453
rect -102 -5461 -101 -5453
rect -97 -5461 -96 -5453
rect -94 -5461 -89 -5453
rect -85 -5461 -80 -5453
rect -78 -5461 -77 -5453
rect -73 -5461 -72 -5453
rect -70 -5461 -68 -5453
rect -64 -5461 -62 -5453
rect -60 -5461 -59 -5453
rect -55 -5461 -54 -5453
rect -52 -5461 -47 -5453
rect -43 -5461 -38 -5453
rect -36 -5461 -35 -5453
rect -31 -5461 -30 -5453
rect -28 -5461 -27 -5453
rect 143 -5461 144 -5453
rect 146 -5461 148 -5453
rect 152 -5461 154 -5453
rect 156 -5461 157 -5453
rect 169 -5461 170 -5453
rect 172 -5461 173 -5453
rect 177 -5461 178 -5453
rect 180 -5461 185 -5453
rect 189 -5461 194 -5453
rect 196 -5461 197 -5453
rect 201 -5461 202 -5453
rect 204 -5461 206 -5453
rect 210 -5461 212 -5453
rect 214 -5461 215 -5453
rect 219 -5461 220 -5453
rect 222 -5461 227 -5453
rect 231 -5461 236 -5453
rect 238 -5461 239 -5453
rect 243 -5461 244 -5453
rect 246 -5461 248 -5453
rect 252 -5461 254 -5453
rect 256 -5461 257 -5453
rect 261 -5461 262 -5453
rect 264 -5461 269 -5453
rect 273 -5461 278 -5453
rect 280 -5461 281 -5453
rect 285 -5461 286 -5453
rect 288 -5461 290 -5453
rect 294 -5461 296 -5453
rect 298 -5461 299 -5453
rect 303 -5461 304 -5453
rect 306 -5461 311 -5453
rect 315 -5461 320 -5453
rect 322 -5461 323 -5453
rect 327 -5461 328 -5453
rect 330 -5461 331 -5453
rect 499 -5461 500 -5453
rect 502 -5461 504 -5453
rect 508 -5461 510 -5453
rect 512 -5461 513 -5453
rect 525 -5461 526 -5453
rect 528 -5461 529 -5453
rect 533 -5461 534 -5453
rect 536 -5461 541 -5453
rect 545 -5461 550 -5453
rect 552 -5461 553 -5453
rect 557 -5461 558 -5453
rect 560 -5461 562 -5453
rect 566 -5461 568 -5453
rect 570 -5461 571 -5453
rect 575 -5461 576 -5453
rect 578 -5461 583 -5453
rect 587 -5461 592 -5453
rect 594 -5461 595 -5453
rect 599 -5461 600 -5453
rect 602 -5461 604 -5453
rect 608 -5461 610 -5453
rect 612 -5461 613 -5453
rect 617 -5461 618 -5453
rect 620 -5461 625 -5453
rect 629 -5461 634 -5453
rect 636 -5461 637 -5453
rect 641 -5461 642 -5453
rect 644 -5461 646 -5453
rect 650 -5461 652 -5453
rect 654 -5461 655 -5453
rect 659 -5461 660 -5453
rect 662 -5461 667 -5453
rect 671 -5461 676 -5453
rect 678 -5461 679 -5453
rect 683 -5461 684 -5453
rect 686 -5461 687 -5453
rect 857 -5461 858 -5453
rect 860 -5461 862 -5453
rect 866 -5461 868 -5453
rect 870 -5461 871 -5453
rect 883 -5461 884 -5453
rect 886 -5461 887 -5453
rect 891 -5461 892 -5453
rect 894 -5461 899 -5453
rect 903 -5461 908 -5453
rect 910 -5461 911 -5453
rect 915 -5461 916 -5453
rect 918 -5461 920 -5453
rect 924 -5461 926 -5453
rect 928 -5461 929 -5453
rect 933 -5461 934 -5453
rect 936 -5461 941 -5453
rect 945 -5461 950 -5453
rect 952 -5461 953 -5453
rect 957 -5461 958 -5453
rect 960 -5461 962 -5453
rect 966 -5461 968 -5453
rect 970 -5461 971 -5453
rect 975 -5461 976 -5453
rect 978 -5461 983 -5453
rect 987 -5461 992 -5453
rect 994 -5461 995 -5453
rect 999 -5461 1000 -5453
rect 1002 -5461 1004 -5453
rect 1008 -5461 1010 -5453
rect 1012 -5461 1013 -5453
rect 1017 -5461 1018 -5453
rect 1020 -5461 1025 -5453
rect 1029 -5461 1034 -5453
rect 1036 -5461 1037 -5453
rect 1041 -5461 1042 -5453
rect 1044 -5461 1045 -5453
rect 1215 -5461 1216 -5453
rect 1218 -5461 1220 -5453
rect 1224 -5461 1226 -5453
rect 1228 -5461 1229 -5453
rect 1241 -5461 1242 -5453
rect 1244 -5461 1245 -5453
rect 1249 -5461 1250 -5453
rect 1252 -5461 1257 -5453
rect 1261 -5461 1266 -5453
rect 1268 -5461 1269 -5453
rect 1273 -5461 1274 -5453
rect 1276 -5461 1278 -5453
rect 1282 -5461 1284 -5453
rect 1286 -5461 1287 -5453
rect 1291 -5461 1292 -5453
rect 1294 -5461 1299 -5453
rect 1303 -5461 1308 -5453
rect 1310 -5461 1311 -5453
rect 1315 -5461 1316 -5453
rect 1318 -5461 1320 -5453
rect 1324 -5461 1326 -5453
rect 1328 -5461 1329 -5453
rect 1333 -5461 1334 -5453
rect 1336 -5461 1341 -5453
rect 1345 -5461 1350 -5453
rect 1352 -5461 1353 -5453
rect 1357 -5461 1358 -5453
rect 1360 -5461 1362 -5453
rect 1366 -5461 1368 -5453
rect 1370 -5461 1371 -5453
rect 1375 -5461 1376 -5453
rect 1378 -5461 1383 -5453
rect 1387 -5461 1392 -5453
rect 1394 -5461 1395 -5453
rect 1399 -5461 1400 -5453
rect 1402 -5461 1403 -5453
rect -1305 -5575 -1304 -5567
rect -1302 -5575 -1301 -5567
rect -1297 -5575 -1296 -5567
rect -1294 -5575 -1292 -5567
rect -1288 -5575 -1286 -5567
rect -1284 -5575 -1283 -5567
rect -931 -5575 -930 -5567
rect -928 -5575 -927 -5567
rect -923 -5575 -922 -5567
rect -920 -5575 -918 -5567
rect -914 -5575 -912 -5567
rect -910 -5575 -909 -5567
rect -573 -5575 -572 -5567
rect -570 -5575 -569 -5567
rect -565 -5575 -564 -5567
rect -562 -5575 -560 -5567
rect -556 -5575 -554 -5567
rect -552 -5575 -551 -5567
rect -215 -5575 -214 -5567
rect -212 -5575 -211 -5567
rect -207 -5575 -206 -5567
rect -204 -5575 -202 -5567
rect -198 -5575 -196 -5567
rect -194 -5575 -193 -5567
rect 143 -5575 144 -5567
rect 146 -5575 147 -5567
rect 151 -5575 152 -5567
rect 154 -5575 156 -5567
rect 160 -5575 162 -5567
rect 164 -5575 165 -5567
rect 499 -5575 500 -5567
rect 502 -5575 503 -5567
rect 507 -5575 508 -5567
rect 510 -5575 512 -5567
rect 516 -5575 518 -5567
rect 520 -5575 521 -5567
rect 857 -5575 858 -5567
rect 860 -5575 861 -5567
rect 865 -5575 866 -5567
rect 868 -5575 870 -5567
rect 874 -5575 876 -5567
rect 878 -5575 879 -5567
rect 1215 -5575 1216 -5567
rect 1218 -5575 1219 -5567
rect 1223 -5575 1224 -5567
rect 1226 -5575 1228 -5567
rect 1232 -5575 1234 -5567
rect 1236 -5575 1237 -5567
rect -1230 -5734 -1229 -5726
rect -1227 -5734 -1225 -5726
rect -1221 -5734 -1219 -5726
rect -1217 -5734 -1216 -5726
rect -1204 -5734 -1203 -5726
rect -1201 -5734 -1193 -5726
rect -1191 -5734 -1190 -5726
rect -1186 -5734 -1185 -5726
rect -1183 -5734 -1175 -5726
rect -1173 -5734 -1168 -5726
rect -1164 -5734 -1159 -5726
rect -1157 -5734 -1156 -5726
rect -1152 -5734 -1151 -5726
rect -1149 -5734 -1147 -5726
rect -1143 -5734 -1141 -5726
rect -1139 -5734 -1138 -5726
rect -931 -5734 -930 -5726
rect -928 -5734 -926 -5726
rect -922 -5734 -920 -5726
rect -918 -5734 -917 -5726
rect -905 -5734 -904 -5726
rect -902 -5734 -900 -5726
rect -896 -5734 -894 -5726
rect -892 -5734 -891 -5726
rect -879 -5734 -878 -5726
rect -876 -5734 -868 -5726
rect -866 -5734 -865 -5726
rect -861 -5734 -860 -5726
rect -858 -5734 -850 -5726
rect -848 -5734 -843 -5726
rect -839 -5734 -834 -5726
rect -832 -5734 -831 -5726
rect -827 -5734 -826 -5726
rect -824 -5734 -822 -5726
rect -818 -5734 -816 -5726
rect -814 -5734 -813 -5726
rect -801 -5734 -800 -5726
rect -798 -5734 -790 -5726
rect -788 -5734 -787 -5726
rect -783 -5734 -782 -5726
rect -780 -5734 -772 -5726
rect -770 -5734 -765 -5726
rect -761 -5734 -756 -5726
rect -754 -5734 -753 -5726
rect -749 -5734 -748 -5726
rect -746 -5734 -741 -5726
rect -737 -5734 -732 -5726
rect -730 -5734 -729 -5726
rect -717 -5734 -716 -5726
rect -714 -5734 -708 -5726
rect -706 -5734 -704 -5726
rect -700 -5734 -698 -5726
rect -696 -5734 -695 -5726
rect -573 -5734 -572 -5726
rect -570 -5734 -568 -5726
rect -564 -5734 -562 -5726
rect -560 -5734 -559 -5726
rect -547 -5734 -546 -5726
rect -544 -5734 -542 -5726
rect -538 -5734 -536 -5726
rect -534 -5734 -533 -5726
rect -521 -5734 -520 -5726
rect -518 -5734 -510 -5726
rect -508 -5734 -507 -5726
rect -503 -5734 -502 -5726
rect -500 -5734 -492 -5726
rect -490 -5734 -485 -5726
rect -481 -5734 -476 -5726
rect -474 -5734 -473 -5726
rect -469 -5734 -468 -5726
rect -466 -5734 -464 -5726
rect -460 -5734 -458 -5726
rect -456 -5734 -455 -5726
rect -443 -5734 -442 -5726
rect -440 -5734 -432 -5726
rect -430 -5734 -429 -5726
rect -425 -5734 -424 -5726
rect -422 -5734 -414 -5726
rect -412 -5734 -407 -5726
rect -403 -5734 -398 -5726
rect -396 -5734 -395 -5726
rect -391 -5734 -390 -5726
rect -388 -5734 -383 -5726
rect -379 -5734 -374 -5726
rect -372 -5734 -371 -5726
rect -359 -5734 -358 -5726
rect -356 -5734 -350 -5726
rect -348 -5734 -346 -5726
rect -342 -5734 -340 -5726
rect -338 -5734 -337 -5726
rect -215 -5734 -214 -5726
rect -212 -5734 -210 -5726
rect -206 -5734 -204 -5726
rect -202 -5734 -201 -5726
rect -189 -5734 -188 -5726
rect -186 -5734 -184 -5726
rect -180 -5734 -178 -5726
rect -176 -5734 -175 -5726
rect -163 -5734 -162 -5726
rect -160 -5734 -152 -5726
rect -150 -5734 -149 -5726
rect -145 -5734 -144 -5726
rect -142 -5734 -134 -5726
rect -132 -5734 -127 -5726
rect -123 -5734 -118 -5726
rect -116 -5734 -115 -5726
rect -111 -5734 -110 -5726
rect -108 -5734 -106 -5726
rect -102 -5734 -100 -5726
rect -98 -5734 -97 -5726
rect -85 -5734 -84 -5726
rect -82 -5734 -74 -5726
rect -72 -5734 -71 -5726
rect -67 -5734 -66 -5726
rect -64 -5734 -56 -5726
rect -54 -5734 -49 -5726
rect -45 -5734 -40 -5726
rect -38 -5734 -37 -5726
rect -33 -5734 -32 -5726
rect -30 -5734 -25 -5726
rect -21 -5734 -16 -5726
rect -14 -5734 -13 -5726
rect -1 -5734 0 -5726
rect 2 -5734 8 -5726
rect 10 -5734 12 -5726
rect 16 -5734 18 -5726
rect 20 -5734 21 -5726
rect 143 -5734 144 -5726
rect 146 -5734 148 -5726
rect 152 -5734 154 -5726
rect 156 -5734 157 -5726
rect 169 -5734 170 -5726
rect 172 -5734 174 -5726
rect 178 -5734 180 -5726
rect 182 -5734 183 -5726
rect 195 -5734 196 -5726
rect 198 -5734 206 -5726
rect 208 -5734 209 -5726
rect 213 -5734 214 -5726
rect 216 -5734 224 -5726
rect 226 -5734 231 -5726
rect 235 -5734 240 -5726
rect 242 -5734 243 -5726
rect 247 -5734 248 -5726
rect 250 -5734 252 -5726
rect 256 -5734 258 -5726
rect 260 -5734 261 -5726
rect 273 -5734 274 -5726
rect 276 -5734 284 -5726
rect 286 -5734 287 -5726
rect 291 -5734 292 -5726
rect 294 -5734 302 -5726
rect 304 -5734 309 -5726
rect 313 -5734 318 -5726
rect 320 -5734 321 -5726
rect 325 -5734 326 -5726
rect 328 -5734 333 -5726
rect 337 -5734 342 -5726
rect 344 -5734 345 -5726
rect 357 -5734 358 -5726
rect 360 -5734 366 -5726
rect 368 -5734 370 -5726
rect 374 -5734 376 -5726
rect 378 -5734 379 -5726
rect 499 -5734 500 -5726
rect 502 -5734 504 -5726
rect 508 -5734 510 -5726
rect 512 -5734 513 -5726
rect 525 -5734 526 -5726
rect 528 -5734 530 -5726
rect 534 -5734 536 -5726
rect 538 -5734 539 -5726
rect 551 -5734 552 -5726
rect 554 -5734 562 -5726
rect 564 -5734 565 -5726
rect 569 -5734 570 -5726
rect 572 -5734 580 -5726
rect 582 -5734 587 -5726
rect 591 -5734 596 -5726
rect 598 -5734 599 -5726
rect 603 -5734 604 -5726
rect 606 -5734 608 -5726
rect 612 -5734 614 -5726
rect 616 -5734 617 -5726
rect 629 -5734 630 -5726
rect 632 -5734 640 -5726
rect 642 -5734 643 -5726
rect 647 -5734 648 -5726
rect 650 -5734 658 -5726
rect 660 -5734 665 -5726
rect 669 -5734 674 -5726
rect 676 -5734 677 -5726
rect 681 -5734 682 -5726
rect 684 -5734 689 -5726
rect 693 -5734 698 -5726
rect 700 -5734 701 -5726
rect 713 -5734 714 -5726
rect 716 -5734 722 -5726
rect 724 -5734 726 -5726
rect 730 -5734 732 -5726
rect 734 -5734 735 -5726
rect 857 -5734 858 -5726
rect 860 -5734 862 -5726
rect 866 -5734 868 -5726
rect 870 -5734 871 -5726
rect 883 -5734 884 -5726
rect 886 -5734 888 -5726
rect 892 -5734 894 -5726
rect 896 -5734 897 -5726
rect 909 -5734 910 -5726
rect 912 -5734 920 -5726
rect 922 -5734 923 -5726
rect 927 -5734 928 -5726
rect 930 -5734 938 -5726
rect 940 -5734 945 -5726
rect 949 -5734 954 -5726
rect 956 -5734 957 -5726
rect 961 -5734 962 -5726
rect 964 -5734 966 -5726
rect 970 -5734 972 -5726
rect 974 -5734 975 -5726
rect 987 -5734 988 -5726
rect 990 -5734 998 -5726
rect 1000 -5734 1001 -5726
rect 1005 -5734 1006 -5726
rect 1008 -5734 1016 -5726
rect 1018 -5734 1023 -5726
rect 1027 -5734 1032 -5726
rect 1034 -5734 1035 -5726
rect 1039 -5734 1040 -5726
rect 1042 -5734 1047 -5726
rect 1051 -5734 1056 -5726
rect 1058 -5734 1059 -5726
rect 1071 -5734 1072 -5726
rect 1074 -5734 1080 -5726
rect 1082 -5734 1084 -5726
rect 1088 -5734 1090 -5726
rect 1092 -5734 1093 -5726
rect 1215 -5734 1216 -5726
rect 1218 -5734 1220 -5726
rect 1224 -5734 1226 -5726
rect 1228 -5734 1229 -5726
rect 1241 -5734 1242 -5726
rect 1244 -5734 1246 -5726
rect 1250 -5734 1252 -5726
rect 1254 -5734 1255 -5726
rect 1267 -5734 1268 -5726
rect 1270 -5734 1278 -5726
rect 1280 -5734 1281 -5726
rect 1285 -5734 1286 -5726
rect 1288 -5734 1296 -5726
rect 1298 -5734 1303 -5726
rect 1307 -5734 1312 -5726
rect 1314 -5734 1315 -5726
rect 1319 -5734 1320 -5726
rect 1322 -5734 1324 -5726
rect 1328 -5734 1330 -5726
rect 1332 -5734 1333 -5726
rect 1345 -5734 1346 -5726
rect 1348 -5734 1356 -5726
rect 1358 -5734 1359 -5726
rect 1363 -5734 1364 -5726
rect 1366 -5734 1374 -5726
rect 1376 -5734 1381 -5726
rect 1385 -5734 1390 -5726
rect 1392 -5734 1393 -5726
rect 1397 -5734 1398 -5726
rect 1400 -5734 1405 -5726
rect 1409 -5734 1414 -5726
rect 1416 -5734 1417 -5726
rect 1429 -5734 1430 -5726
rect 1432 -5734 1438 -5726
rect 1440 -5734 1442 -5726
rect 1446 -5734 1448 -5726
rect 1450 -5734 1451 -5726
rect -1230 -5857 -1229 -5849
rect -1227 -5857 -1225 -5849
rect -1221 -5857 -1219 -5849
rect -1217 -5857 -1216 -5849
rect -1204 -5857 -1203 -5849
rect -1201 -5857 -1200 -5849
rect -1196 -5857 -1195 -5849
rect -1193 -5857 -1188 -5849
rect -1184 -5857 -1179 -5849
rect -1177 -5857 -1176 -5849
rect -1172 -5857 -1171 -5849
rect -1169 -5857 -1167 -5849
rect -1163 -5857 -1161 -5849
rect -1159 -5857 -1158 -5849
rect -1154 -5857 -1153 -5849
rect -1151 -5857 -1146 -5849
rect -1142 -5857 -1137 -5849
rect -1135 -5857 -1134 -5849
rect -1130 -5857 -1129 -5849
rect -1127 -5857 -1125 -5849
rect -1121 -5857 -1119 -5849
rect -1117 -5857 -1116 -5849
rect -1112 -5857 -1111 -5849
rect -1109 -5857 -1104 -5849
rect -1100 -5857 -1095 -5849
rect -1093 -5857 -1092 -5849
rect -1088 -5857 -1087 -5849
rect -1085 -5857 -1083 -5849
rect -1079 -5857 -1077 -5849
rect -1075 -5857 -1074 -5849
rect -1070 -5857 -1069 -5849
rect -1067 -5857 -1062 -5849
rect -1058 -5857 -1053 -5849
rect -1051 -5857 -1050 -5849
rect -1046 -5857 -1045 -5849
rect -1043 -5857 -1042 -5849
rect -931 -5857 -930 -5849
rect -928 -5857 -926 -5849
rect -922 -5857 -920 -5849
rect -918 -5857 -917 -5849
rect -905 -5857 -904 -5849
rect -902 -5857 -901 -5849
rect -897 -5857 -896 -5849
rect -894 -5857 -889 -5849
rect -885 -5857 -880 -5849
rect -878 -5857 -877 -5849
rect -873 -5857 -872 -5849
rect -870 -5857 -868 -5849
rect -864 -5857 -862 -5849
rect -860 -5857 -859 -5849
rect -855 -5857 -854 -5849
rect -852 -5857 -847 -5849
rect -843 -5857 -838 -5849
rect -836 -5857 -835 -5849
rect -831 -5857 -830 -5849
rect -828 -5857 -826 -5849
rect -822 -5857 -820 -5849
rect -818 -5857 -817 -5849
rect -813 -5857 -812 -5849
rect -810 -5857 -805 -5849
rect -801 -5857 -796 -5849
rect -794 -5857 -793 -5849
rect -789 -5857 -788 -5849
rect -786 -5857 -784 -5849
rect -780 -5857 -778 -5849
rect -776 -5857 -775 -5849
rect -771 -5857 -770 -5849
rect -768 -5857 -763 -5849
rect -759 -5857 -754 -5849
rect -752 -5857 -751 -5849
rect -747 -5857 -746 -5849
rect -744 -5857 -743 -5849
rect -573 -5857 -572 -5849
rect -570 -5857 -568 -5849
rect -564 -5857 -562 -5849
rect -560 -5857 -559 -5849
rect -547 -5857 -546 -5849
rect -544 -5857 -543 -5849
rect -539 -5857 -538 -5849
rect -536 -5857 -531 -5849
rect -527 -5857 -522 -5849
rect -520 -5857 -519 -5849
rect -515 -5857 -514 -5849
rect -512 -5857 -510 -5849
rect -506 -5857 -504 -5849
rect -502 -5857 -501 -5849
rect -497 -5857 -496 -5849
rect -494 -5857 -489 -5849
rect -485 -5857 -480 -5849
rect -478 -5857 -477 -5849
rect -473 -5857 -472 -5849
rect -470 -5857 -468 -5849
rect -464 -5857 -462 -5849
rect -460 -5857 -459 -5849
rect -455 -5857 -454 -5849
rect -452 -5857 -447 -5849
rect -443 -5857 -438 -5849
rect -436 -5857 -435 -5849
rect -431 -5857 -430 -5849
rect -428 -5857 -426 -5849
rect -422 -5857 -420 -5849
rect -418 -5857 -417 -5849
rect -413 -5857 -412 -5849
rect -410 -5857 -405 -5849
rect -401 -5857 -396 -5849
rect -394 -5857 -393 -5849
rect -389 -5857 -388 -5849
rect -386 -5857 -385 -5849
rect -215 -5857 -214 -5849
rect -212 -5857 -210 -5849
rect -206 -5857 -204 -5849
rect -202 -5857 -201 -5849
rect -189 -5857 -188 -5849
rect -186 -5857 -185 -5849
rect -181 -5857 -180 -5849
rect -178 -5857 -173 -5849
rect -169 -5857 -164 -5849
rect -162 -5857 -161 -5849
rect -157 -5857 -156 -5849
rect -154 -5857 -152 -5849
rect -148 -5857 -146 -5849
rect -144 -5857 -143 -5849
rect -139 -5857 -138 -5849
rect -136 -5857 -131 -5849
rect -127 -5857 -122 -5849
rect -120 -5857 -119 -5849
rect -115 -5857 -114 -5849
rect -112 -5857 -110 -5849
rect -106 -5857 -104 -5849
rect -102 -5857 -101 -5849
rect -97 -5857 -96 -5849
rect -94 -5857 -89 -5849
rect -85 -5857 -80 -5849
rect -78 -5857 -77 -5849
rect -73 -5857 -72 -5849
rect -70 -5857 -68 -5849
rect -64 -5857 -62 -5849
rect -60 -5857 -59 -5849
rect -55 -5857 -54 -5849
rect -52 -5857 -47 -5849
rect -43 -5857 -38 -5849
rect -36 -5857 -35 -5849
rect -31 -5857 -30 -5849
rect -28 -5857 -27 -5849
rect 143 -5857 144 -5849
rect 146 -5857 148 -5849
rect 152 -5857 154 -5849
rect 156 -5857 157 -5849
rect 169 -5857 170 -5849
rect 172 -5857 173 -5849
rect 177 -5857 178 -5849
rect 180 -5857 185 -5849
rect 189 -5857 194 -5849
rect 196 -5857 197 -5849
rect 201 -5857 202 -5849
rect 204 -5857 206 -5849
rect 210 -5857 212 -5849
rect 214 -5857 215 -5849
rect 219 -5857 220 -5849
rect 222 -5857 227 -5849
rect 231 -5857 236 -5849
rect 238 -5857 239 -5849
rect 243 -5857 244 -5849
rect 246 -5857 248 -5849
rect 252 -5857 254 -5849
rect 256 -5857 257 -5849
rect 261 -5857 262 -5849
rect 264 -5857 269 -5849
rect 273 -5857 278 -5849
rect 280 -5857 281 -5849
rect 285 -5857 286 -5849
rect 288 -5857 290 -5849
rect 294 -5857 296 -5849
rect 298 -5857 299 -5849
rect 303 -5857 304 -5849
rect 306 -5857 311 -5849
rect 315 -5857 320 -5849
rect 322 -5857 323 -5849
rect 327 -5857 328 -5849
rect 330 -5857 331 -5849
rect 499 -5857 500 -5849
rect 502 -5857 504 -5849
rect 508 -5857 510 -5849
rect 512 -5857 513 -5849
rect 525 -5857 526 -5849
rect 528 -5857 529 -5849
rect 533 -5857 534 -5849
rect 536 -5857 541 -5849
rect 545 -5857 550 -5849
rect 552 -5857 553 -5849
rect 557 -5857 558 -5849
rect 560 -5857 562 -5849
rect 566 -5857 568 -5849
rect 570 -5857 571 -5849
rect 575 -5857 576 -5849
rect 578 -5857 583 -5849
rect 587 -5857 592 -5849
rect 594 -5857 595 -5849
rect 599 -5857 600 -5849
rect 602 -5857 604 -5849
rect 608 -5857 610 -5849
rect 612 -5857 613 -5849
rect 617 -5857 618 -5849
rect 620 -5857 625 -5849
rect 629 -5857 634 -5849
rect 636 -5857 637 -5849
rect 641 -5857 642 -5849
rect 644 -5857 646 -5849
rect 650 -5857 652 -5849
rect 654 -5857 655 -5849
rect 659 -5857 660 -5849
rect 662 -5857 667 -5849
rect 671 -5857 676 -5849
rect 678 -5857 679 -5849
rect 683 -5857 684 -5849
rect 686 -5857 687 -5849
rect 857 -5857 858 -5849
rect 860 -5857 862 -5849
rect 866 -5857 868 -5849
rect 870 -5857 871 -5849
rect 883 -5857 884 -5849
rect 886 -5857 887 -5849
rect 891 -5857 892 -5849
rect 894 -5857 899 -5849
rect 903 -5857 908 -5849
rect 910 -5857 911 -5849
rect 915 -5857 916 -5849
rect 918 -5857 920 -5849
rect 924 -5857 926 -5849
rect 928 -5857 929 -5849
rect 933 -5857 934 -5849
rect 936 -5857 941 -5849
rect 945 -5857 950 -5849
rect 952 -5857 953 -5849
rect 957 -5857 958 -5849
rect 960 -5857 962 -5849
rect 966 -5857 968 -5849
rect 970 -5857 971 -5849
rect 975 -5857 976 -5849
rect 978 -5857 983 -5849
rect 987 -5857 992 -5849
rect 994 -5857 995 -5849
rect 999 -5857 1000 -5849
rect 1002 -5857 1004 -5849
rect 1008 -5857 1010 -5849
rect 1012 -5857 1013 -5849
rect 1017 -5857 1018 -5849
rect 1020 -5857 1025 -5849
rect 1029 -5857 1034 -5849
rect 1036 -5857 1037 -5849
rect 1041 -5857 1042 -5849
rect 1044 -5857 1045 -5849
rect 1215 -5857 1216 -5849
rect 1218 -5857 1220 -5849
rect 1224 -5857 1226 -5849
rect 1228 -5857 1229 -5849
rect 1241 -5857 1242 -5849
rect 1244 -5857 1245 -5849
rect 1249 -5857 1250 -5849
rect 1252 -5857 1257 -5849
rect 1261 -5857 1266 -5849
rect 1268 -5857 1269 -5849
rect 1273 -5857 1274 -5849
rect 1276 -5857 1278 -5849
rect 1282 -5857 1284 -5849
rect 1286 -5857 1287 -5849
rect 1291 -5857 1292 -5849
rect 1294 -5857 1299 -5849
rect 1303 -5857 1308 -5849
rect 1310 -5857 1311 -5849
rect 1315 -5857 1316 -5849
rect 1318 -5857 1320 -5849
rect 1324 -5857 1326 -5849
rect 1328 -5857 1329 -5849
rect 1333 -5857 1334 -5849
rect 1336 -5857 1341 -5849
rect 1345 -5857 1350 -5849
rect 1352 -5857 1353 -5849
rect 1357 -5857 1358 -5849
rect 1360 -5857 1362 -5849
rect 1366 -5857 1368 -5849
rect 1370 -5857 1371 -5849
rect 1375 -5857 1376 -5849
rect 1378 -5857 1383 -5849
rect 1387 -5857 1392 -5849
rect 1394 -5857 1395 -5849
rect 1399 -5857 1400 -5849
rect 1402 -5857 1403 -5849
rect 1559 -5857 1560 -5849
rect 1562 -5857 1564 -5849
rect 1568 -5857 1570 -5849
rect 1572 -5857 1573 -5849
rect 1585 -5857 1586 -5849
rect 1588 -5857 1589 -5849
rect 1593 -5857 1594 -5849
rect 1596 -5857 1601 -5849
rect 1605 -5857 1610 -5849
rect 1612 -5857 1613 -5849
rect 1617 -5857 1618 -5849
rect 1620 -5857 1622 -5849
rect 1626 -5857 1628 -5849
rect 1630 -5857 1631 -5849
rect 1635 -5857 1636 -5849
rect 1638 -5857 1643 -5849
rect 1647 -5857 1652 -5849
rect 1654 -5857 1655 -5849
rect 1659 -5857 1660 -5849
rect 1662 -5857 1664 -5849
rect 1668 -5857 1670 -5849
rect 1672 -5857 1673 -5849
rect 1677 -5857 1678 -5849
rect 1680 -5857 1685 -5849
rect 1689 -5857 1694 -5849
rect 1696 -5857 1697 -5849
rect 1701 -5857 1702 -5849
rect 1704 -5857 1706 -5849
rect 1710 -5857 1712 -5849
rect 1714 -5857 1715 -5849
rect 1719 -5857 1720 -5849
rect 1722 -5857 1727 -5849
rect 1731 -5857 1736 -5849
rect 1738 -5857 1739 -5849
rect 1743 -5857 1744 -5849
rect 1746 -5857 1747 -5849
<< metal1 >>
rect -1319 -812 -1315 -748
rect -1307 -788 -1303 -784
rect -1290 -788 -1286 -784
rect -1299 -799 -1295 -796
rect -1299 -803 -1284 -799
rect -1319 -816 -1306 -812
rect -1319 -1162 -1315 -816
rect -1288 -842 -1284 -803
rect -1288 -857 -1284 -846
rect -1307 -861 -1284 -857
rect -1307 -864 -1303 -861
rect -1281 -864 -1277 -796
rect -949 -812 -945 -748
rect -936 -788 -932 -784
rect -919 -788 -915 -784
rect -928 -799 -924 -796
rect -928 -803 -913 -799
rect -949 -816 -935 -812
rect -1290 -872 -1286 -868
rect -1281 -1070 -1277 -868
rect -1309 -1138 -1305 -1134
rect -1292 -1138 -1288 -1134
rect -1301 -1149 -1297 -1146
rect -1301 -1153 -1286 -1149
rect -1319 -1166 -1308 -1162
rect -1550 -1767 -1546 -1763
rect -1533 -1767 -1529 -1763
rect -1513 -1767 -1509 -1763
rect -1492 -1767 -1488 -1763
rect -1471 -1767 -1467 -1763
rect -1450 -1767 -1446 -1763
rect -1429 -1767 -1425 -1763
rect -1408 -1767 -1404 -1763
rect -1387 -1767 -1383 -1763
rect -1367 -1767 -1363 -1763
rect -1559 -1822 -1555 -1775
rect -1559 -1843 -1555 -1826
rect -1541 -1836 -1537 -1775
rect -1525 -1836 -1521 -1775
rect -1501 -1815 -1497 -1775
rect -1501 -1836 -1497 -1819
rect -1483 -1836 -1479 -1775
rect -1459 -1822 -1455 -1775
rect -1459 -1836 -1455 -1826
rect -1441 -1815 -1437 -1775
rect -1441 -1836 -1437 -1819
rect -1417 -1829 -1413 -1775
rect -1399 -1799 -1395 -1775
rect -1399 -1815 -1395 -1803
rect -1417 -1836 -1413 -1833
rect -1541 -1840 -1532 -1836
rect -1525 -1840 -1517 -1836
rect -1541 -1843 -1537 -1840
rect -1517 -1843 -1513 -1840
rect -1509 -1840 -1497 -1836
rect -1483 -1840 -1475 -1836
rect -1509 -1843 -1505 -1840
rect -1475 -1843 -1471 -1840
rect -1467 -1840 -1455 -1836
rect -1441 -1840 -1429 -1836
rect -1467 -1843 -1463 -1840
rect -1433 -1843 -1429 -1840
rect -1425 -1840 -1413 -1836
rect -1399 -1836 -1395 -1819
rect -1375 -1822 -1371 -1775
rect -1375 -1836 -1371 -1826
rect -1399 -1840 -1387 -1836
rect -1425 -1843 -1421 -1840
rect -1391 -1843 -1387 -1840
rect -1383 -1840 -1371 -1836
rect -1383 -1843 -1379 -1840
rect -1550 -1851 -1546 -1847
rect -1533 -1851 -1529 -1847
rect -1492 -1851 -1488 -1847
rect -1450 -1851 -1446 -1847
rect -1408 -1851 -1404 -1847
rect -1367 -1851 -1363 -1847
rect -1351 -1906 -1347 -1803
rect -1319 -1815 -1315 -1166
rect -1290 -1192 -1286 -1153
rect -1290 -1207 -1286 -1196
rect -1309 -1211 -1286 -1207
rect -1309 -1214 -1305 -1211
rect -1283 -1214 -1279 -1146
rect -1292 -1222 -1288 -1218
rect -1283 -1357 -1279 -1218
rect -1251 -1350 -1247 -840
rect -1221 -1022 -1217 -1018
rect -1204 -1022 -1200 -1018
rect -1184 -1022 -1180 -1018
rect -1163 -1022 -1159 -1018
rect -1142 -1022 -1138 -1018
rect -1121 -1022 -1117 -1018
rect -1100 -1022 -1096 -1018
rect -1079 -1022 -1075 -1018
rect -1058 -1022 -1054 -1018
rect -1038 -1022 -1034 -1018
rect -1230 -1077 -1226 -1030
rect -1230 -1098 -1226 -1081
rect -1212 -1091 -1208 -1030
rect -1196 -1091 -1192 -1030
rect -1172 -1070 -1168 -1030
rect -1172 -1091 -1168 -1074
rect -1154 -1091 -1150 -1030
rect -1130 -1077 -1126 -1030
rect -1130 -1091 -1126 -1081
rect -1112 -1070 -1108 -1030
rect -1112 -1091 -1108 -1074
rect -1088 -1084 -1084 -1030
rect -1070 -1062 -1066 -1030
rect -1070 -1070 -1066 -1066
rect -1088 -1091 -1084 -1088
rect -1212 -1095 -1203 -1091
rect -1196 -1095 -1188 -1091
rect -1212 -1098 -1208 -1095
rect -1188 -1098 -1184 -1095
rect -1180 -1095 -1168 -1091
rect -1154 -1095 -1146 -1091
rect -1180 -1098 -1176 -1095
rect -1146 -1098 -1142 -1095
rect -1138 -1095 -1126 -1091
rect -1112 -1095 -1100 -1091
rect -1138 -1098 -1134 -1095
rect -1104 -1098 -1100 -1095
rect -1096 -1095 -1084 -1091
rect -1070 -1091 -1066 -1074
rect -1046 -1077 -1042 -1030
rect -1046 -1091 -1042 -1081
rect -1070 -1095 -1058 -1091
rect -1096 -1098 -1092 -1095
rect -1062 -1098 -1058 -1095
rect -1054 -1095 -1042 -1091
rect -1054 -1098 -1050 -1095
rect -1221 -1106 -1217 -1102
rect -1204 -1106 -1200 -1102
rect -1163 -1106 -1159 -1102
rect -1121 -1106 -1117 -1102
rect -1079 -1106 -1075 -1102
rect -1038 -1106 -1034 -1102
rect -1221 -1302 -1217 -1298
rect -1204 -1302 -1200 -1298
rect -1164 -1302 -1160 -1298
rect -1143 -1302 -1139 -1298
rect -1230 -1343 -1226 -1310
rect -1230 -1378 -1226 -1347
rect -1212 -1337 -1208 -1310
rect -1212 -1341 -1203 -1337
rect -1212 -1378 -1208 -1341
rect -1186 -1364 -1182 -1310
rect -1186 -1371 -1182 -1368
rect -1152 -1371 -1148 -1310
rect -1134 -1342 -1130 -1310
rect -1204 -1378 -1200 -1375
rect -1195 -1375 -1182 -1371
rect -1195 -1378 -1191 -1375
rect -1168 -1378 -1164 -1375
rect -1160 -1375 -1141 -1371
rect -1160 -1378 -1156 -1375
rect -1134 -1378 -1130 -1346
rect -976 -1349 -972 -1187
rect -964 -1334 -960 -832
rect -949 -1162 -945 -816
rect -917 -844 -913 -803
rect -917 -857 -913 -848
rect -936 -861 -913 -857
rect -910 -836 -906 -796
rect -591 -812 -587 -749
rect -577 -788 -573 -784
rect -560 -788 -556 -784
rect -569 -799 -565 -796
rect -569 -803 -554 -799
rect -591 -816 -576 -812
rect -936 -864 -932 -861
rect -910 -864 -906 -840
rect -919 -872 -915 -868
rect -926 -1022 -922 -1018
rect -909 -1022 -905 -1018
rect -889 -1022 -885 -1018
rect -868 -1022 -864 -1018
rect -847 -1022 -843 -1018
rect -826 -1022 -822 -1018
rect -805 -1022 -801 -1018
rect -784 -1022 -780 -1018
rect -763 -1022 -759 -1018
rect -743 -1022 -739 -1018
rect -935 -1077 -931 -1030
rect -935 -1098 -931 -1081
rect -917 -1091 -913 -1030
rect -901 -1091 -897 -1030
rect -877 -1070 -873 -1030
rect -877 -1091 -873 -1074
rect -859 -1091 -855 -1030
rect -835 -1077 -831 -1030
rect -835 -1091 -831 -1081
rect -817 -1070 -813 -1030
rect -817 -1091 -813 -1074
rect -793 -1084 -789 -1030
rect -775 -1062 -771 -1030
rect -775 -1070 -771 -1066
rect -793 -1091 -789 -1088
rect -917 -1095 -908 -1091
rect -901 -1095 -893 -1091
rect -917 -1098 -913 -1095
rect -893 -1098 -889 -1095
rect -885 -1095 -873 -1091
rect -859 -1095 -851 -1091
rect -885 -1098 -881 -1095
rect -851 -1098 -847 -1095
rect -843 -1095 -831 -1091
rect -817 -1095 -805 -1091
rect -843 -1098 -839 -1095
rect -809 -1098 -805 -1095
rect -801 -1095 -789 -1091
rect -775 -1091 -771 -1074
rect -751 -1077 -747 -1030
rect -751 -1091 -747 -1081
rect -775 -1095 -763 -1091
rect -801 -1098 -797 -1095
rect -767 -1098 -763 -1095
rect -759 -1095 -747 -1091
rect -759 -1098 -755 -1095
rect -926 -1106 -922 -1102
rect -909 -1106 -905 -1102
rect -868 -1106 -864 -1102
rect -826 -1106 -822 -1102
rect -784 -1106 -780 -1102
rect -743 -1106 -739 -1102
rect -935 -1138 -931 -1134
rect -918 -1138 -914 -1134
rect -927 -1149 -923 -1146
rect -927 -1153 -912 -1149
rect -949 -1166 -934 -1162
rect -1221 -1386 -1217 -1382
rect -1177 -1386 -1173 -1382
rect -1143 -1386 -1139 -1382
rect -1257 -1644 -1253 -1397
rect -1124 -1400 -1120 -1368
rect -1244 -1473 -1240 -1404
rect -1221 -1425 -1217 -1421
rect -1204 -1425 -1200 -1421
rect -1184 -1425 -1180 -1421
rect -1163 -1425 -1159 -1421
rect -1142 -1425 -1138 -1421
rect -1121 -1425 -1117 -1421
rect -1100 -1425 -1096 -1421
rect -1079 -1425 -1075 -1421
rect -1058 -1425 -1054 -1421
rect -1038 -1425 -1034 -1421
rect -1230 -1480 -1226 -1433
rect -1230 -1501 -1226 -1484
rect -1212 -1494 -1208 -1433
rect -1196 -1494 -1192 -1433
rect -1172 -1473 -1168 -1433
rect -1172 -1494 -1168 -1477
rect -1154 -1494 -1150 -1433
rect -1130 -1480 -1126 -1433
rect -1130 -1494 -1126 -1484
rect -1112 -1473 -1108 -1433
rect -1112 -1494 -1108 -1477
rect -1088 -1487 -1084 -1433
rect -1070 -1465 -1066 -1433
rect -1070 -1473 -1066 -1469
rect -1088 -1494 -1084 -1491
rect -1212 -1498 -1203 -1494
rect -1196 -1498 -1188 -1494
rect -1212 -1501 -1208 -1498
rect -1188 -1501 -1184 -1498
rect -1180 -1498 -1168 -1494
rect -1154 -1498 -1146 -1494
rect -1180 -1501 -1176 -1498
rect -1146 -1501 -1142 -1498
rect -1138 -1498 -1126 -1494
rect -1112 -1498 -1100 -1494
rect -1138 -1501 -1134 -1498
rect -1104 -1501 -1100 -1498
rect -1096 -1498 -1084 -1494
rect -1070 -1494 -1066 -1477
rect -1046 -1480 -1042 -1433
rect -1046 -1494 -1042 -1484
rect -1070 -1498 -1058 -1494
rect -1096 -1501 -1092 -1498
rect -1062 -1501 -1058 -1498
rect -1054 -1498 -1042 -1494
rect -1054 -1501 -1050 -1498
rect -1221 -1509 -1217 -1505
rect -1204 -1509 -1200 -1505
rect -1163 -1509 -1159 -1505
rect -1121 -1509 -1117 -1505
rect -1079 -1509 -1075 -1505
rect -1038 -1509 -1034 -1505
rect -1221 -1596 -1217 -1592
rect -1204 -1596 -1200 -1592
rect -1184 -1596 -1180 -1592
rect -1163 -1596 -1159 -1592
rect -1142 -1596 -1138 -1592
rect -1121 -1596 -1117 -1592
rect -1100 -1596 -1096 -1592
rect -1079 -1596 -1075 -1592
rect -1058 -1596 -1054 -1592
rect -1038 -1596 -1034 -1592
rect -1230 -1651 -1226 -1604
rect -1230 -1672 -1226 -1655
rect -1212 -1665 -1208 -1604
rect -1196 -1665 -1192 -1604
rect -1172 -1644 -1168 -1604
rect -1172 -1665 -1168 -1648
rect -1154 -1665 -1150 -1604
rect -1130 -1651 -1126 -1604
rect -1130 -1665 -1126 -1655
rect -1112 -1644 -1108 -1604
rect -1112 -1665 -1108 -1648
rect -1088 -1658 -1084 -1604
rect -1070 -1636 -1066 -1604
rect -1070 -1644 -1066 -1640
rect -1088 -1665 -1084 -1662
rect -1212 -1669 -1203 -1665
rect -1196 -1669 -1188 -1665
rect -1212 -1672 -1208 -1669
rect -1188 -1672 -1184 -1669
rect -1180 -1669 -1168 -1665
rect -1154 -1669 -1146 -1665
rect -1180 -1672 -1176 -1669
rect -1146 -1672 -1142 -1669
rect -1138 -1669 -1126 -1665
rect -1112 -1669 -1100 -1665
rect -1138 -1672 -1134 -1669
rect -1104 -1672 -1100 -1669
rect -1096 -1669 -1084 -1665
rect -1070 -1665 -1066 -1648
rect -1046 -1651 -1042 -1604
rect -1046 -1665 -1042 -1655
rect -1070 -1669 -1058 -1665
rect -1096 -1672 -1092 -1669
rect -1062 -1672 -1058 -1669
rect -1054 -1669 -1042 -1665
rect -1054 -1672 -1050 -1669
rect -1221 -1680 -1217 -1676
rect -1204 -1680 -1200 -1676
rect -1163 -1680 -1159 -1676
rect -1121 -1680 -1117 -1676
rect -1079 -1680 -1075 -1676
rect -1038 -1680 -1034 -1676
rect -1023 -1687 -1019 -1640
rect -976 -1644 -972 -1404
rect -1309 -1874 -1305 -1870
rect -1292 -1874 -1288 -1870
rect -1301 -1885 -1297 -1882
rect -1301 -1889 -1286 -1885
rect -1319 -1902 -1308 -1898
rect -1550 -2348 -1546 -2344
rect -1533 -2348 -1529 -2344
rect -1513 -2348 -1509 -2344
rect -1492 -2348 -1488 -2344
rect -1471 -2348 -1467 -2344
rect -1450 -2348 -1446 -2344
rect -1429 -2348 -1425 -2344
rect -1408 -2348 -1404 -2344
rect -1387 -2348 -1383 -2344
rect -1367 -2348 -1363 -2344
rect -1559 -2403 -1555 -2356
rect -1559 -2424 -1555 -2407
rect -1541 -2417 -1537 -2356
rect -1525 -2417 -1521 -2356
rect -1501 -2396 -1497 -2356
rect -1501 -2417 -1497 -2400
rect -1483 -2417 -1479 -2356
rect -1459 -2403 -1455 -2356
rect -1459 -2417 -1455 -2407
rect -1441 -2396 -1437 -2356
rect -1441 -2417 -1437 -2400
rect -1417 -2410 -1413 -2356
rect -1399 -2388 -1395 -2356
rect -1399 -2396 -1395 -2392
rect -1417 -2417 -1413 -2414
rect -1541 -2421 -1532 -2417
rect -1525 -2421 -1517 -2417
rect -1541 -2424 -1537 -2421
rect -1517 -2424 -1513 -2421
rect -1509 -2421 -1497 -2417
rect -1483 -2421 -1475 -2417
rect -1509 -2424 -1505 -2421
rect -1475 -2424 -1471 -2421
rect -1467 -2421 -1455 -2417
rect -1441 -2421 -1429 -2417
rect -1467 -2424 -1463 -2421
rect -1433 -2424 -1429 -2421
rect -1425 -2421 -1413 -2417
rect -1399 -2417 -1395 -2400
rect -1375 -2403 -1371 -2356
rect -1375 -2417 -1371 -2407
rect -1399 -2421 -1387 -2417
rect -1425 -2424 -1421 -2421
rect -1391 -2424 -1387 -2421
rect -1383 -2421 -1371 -2417
rect -1383 -2424 -1379 -2421
rect -1550 -2432 -1546 -2428
rect -1533 -2432 -1529 -2428
rect -1492 -2432 -1488 -2428
rect -1450 -2432 -1446 -2428
rect -1408 -2432 -1404 -2428
rect -1367 -2432 -1363 -2428
rect -1350 -2440 -1346 -2392
rect -1581 -2567 -1577 -2444
rect -1550 -2519 -1546 -2515
rect -1533 -2519 -1529 -2515
rect -1513 -2519 -1509 -2515
rect -1492 -2519 -1488 -2515
rect -1471 -2519 -1467 -2515
rect -1450 -2519 -1446 -2515
rect -1429 -2519 -1425 -2515
rect -1408 -2519 -1404 -2515
rect -1387 -2519 -1383 -2515
rect -1367 -2519 -1363 -2515
rect -1559 -2574 -1555 -2527
rect -1559 -2595 -1555 -2578
rect -1541 -2588 -1537 -2527
rect -1525 -2588 -1521 -2527
rect -1501 -2567 -1497 -2527
rect -1501 -2588 -1497 -2571
rect -1483 -2588 -1479 -2527
rect -1459 -2574 -1455 -2527
rect -1459 -2588 -1455 -2578
rect -1441 -2567 -1437 -2527
rect -1441 -2588 -1437 -2571
rect -1417 -2581 -1413 -2527
rect -1399 -2559 -1395 -2527
rect -1399 -2567 -1395 -2563
rect -1417 -2588 -1413 -2585
rect -1541 -2592 -1532 -2588
rect -1525 -2592 -1517 -2588
rect -1541 -2595 -1537 -2592
rect -1517 -2595 -1513 -2592
rect -1509 -2592 -1497 -2588
rect -1483 -2592 -1475 -2588
rect -1509 -2595 -1505 -2592
rect -1475 -2595 -1471 -2592
rect -1467 -2592 -1455 -2588
rect -1441 -2592 -1429 -2588
rect -1467 -2595 -1463 -2592
rect -1433 -2595 -1429 -2592
rect -1425 -2592 -1413 -2588
rect -1399 -2588 -1395 -2571
rect -1375 -2574 -1371 -2527
rect -1375 -2588 -1371 -2578
rect -1399 -2592 -1387 -2588
rect -1425 -2595 -1421 -2592
rect -1391 -2595 -1387 -2592
rect -1383 -2592 -1371 -2588
rect -1383 -2595 -1379 -2592
rect -1550 -2603 -1546 -2599
rect -1533 -2603 -1529 -2599
rect -1492 -2603 -1488 -2599
rect -1450 -2603 -1446 -2599
rect -1408 -2603 -1404 -2599
rect -1367 -2603 -1363 -2599
rect -1355 -2656 -1351 -2563
rect -1319 -2567 -1315 -1902
rect -1290 -1928 -1286 -1889
rect -1290 -1943 -1286 -1932
rect -1309 -1947 -1286 -1943
rect -1309 -1950 -1305 -1947
rect -1283 -1950 -1279 -1882
rect -1292 -1958 -1288 -1954
rect -1283 -2088 -1279 -1954
rect -1257 -2081 -1253 -1691
rect -1221 -1767 -1217 -1763
rect -1204 -1767 -1200 -1763
rect -1184 -1767 -1180 -1763
rect -1163 -1767 -1159 -1763
rect -1142 -1767 -1138 -1763
rect -1121 -1767 -1117 -1763
rect -1100 -1767 -1096 -1763
rect -1079 -1767 -1075 -1763
rect -1058 -1767 -1054 -1763
rect -1038 -1767 -1034 -1763
rect -1230 -1822 -1226 -1775
rect -1230 -1843 -1226 -1826
rect -1212 -1836 -1208 -1775
rect -1196 -1836 -1192 -1775
rect -1172 -1815 -1168 -1775
rect -1172 -1836 -1168 -1819
rect -1154 -1836 -1150 -1775
rect -1130 -1822 -1126 -1775
rect -1130 -1836 -1126 -1826
rect -1112 -1815 -1108 -1775
rect -1112 -1836 -1108 -1819
rect -1088 -1829 -1084 -1775
rect -1070 -1807 -1066 -1775
rect -1070 -1815 -1066 -1811
rect -1088 -1836 -1084 -1833
rect -1212 -1840 -1203 -1836
rect -1196 -1840 -1188 -1836
rect -1212 -1843 -1208 -1840
rect -1188 -1843 -1184 -1840
rect -1180 -1840 -1168 -1836
rect -1154 -1840 -1146 -1836
rect -1180 -1843 -1176 -1840
rect -1146 -1843 -1142 -1840
rect -1138 -1840 -1126 -1836
rect -1112 -1840 -1100 -1836
rect -1138 -1843 -1134 -1840
rect -1104 -1843 -1100 -1840
rect -1096 -1840 -1084 -1836
rect -1070 -1836 -1066 -1819
rect -1046 -1822 -1042 -1775
rect -1046 -1836 -1042 -1826
rect -1070 -1840 -1058 -1836
rect -1096 -1843 -1092 -1840
rect -1062 -1843 -1058 -1840
rect -1054 -1840 -1042 -1836
rect -1054 -1843 -1050 -1840
rect -1221 -1851 -1217 -1847
rect -1204 -1851 -1200 -1847
rect -1163 -1851 -1159 -1847
rect -1121 -1851 -1117 -1847
rect -1079 -1851 -1075 -1847
rect -1038 -1851 -1034 -1847
rect -1016 -1898 -1012 -1811
rect -1225 -2033 -1221 -2029
rect -1208 -2033 -1204 -2029
rect -1168 -2033 -1164 -2029
rect -1147 -2033 -1143 -2029
rect -1234 -2074 -1230 -2041
rect -1234 -2109 -1230 -2078
rect -1216 -2068 -1212 -2041
rect -1216 -2072 -1207 -2068
rect -1216 -2109 -1212 -2072
rect -1190 -2095 -1186 -2041
rect -1190 -2102 -1186 -2099
rect -1156 -2102 -1152 -2041
rect -1138 -2073 -1134 -2041
rect -976 -2065 -972 -1692
rect -949 -1815 -945 -1166
rect -916 -1192 -912 -1153
rect -916 -1207 -912 -1196
rect -935 -1211 -912 -1207
rect -909 -1183 -905 -1146
rect -935 -1214 -931 -1211
rect -909 -1214 -905 -1187
rect -918 -1222 -914 -1218
rect -926 -1302 -922 -1298
rect -900 -1302 -896 -1298
rect -883 -1302 -879 -1298
rect -843 -1302 -839 -1298
rect -822 -1302 -818 -1298
rect -805 -1302 -801 -1298
rect -765 -1302 -761 -1298
rect -741 -1302 -737 -1298
rect -704 -1302 -700 -1298
rect -935 -1327 -931 -1310
rect -935 -1378 -931 -1331
rect -917 -1320 -913 -1310
rect -917 -1378 -913 -1324
rect -909 -1349 -905 -1310
rect -891 -1342 -887 -1310
rect -909 -1378 -905 -1353
rect -891 -1378 -887 -1346
rect -865 -1334 -861 -1310
rect -865 -1371 -861 -1338
rect -831 -1371 -827 -1310
rect -813 -1327 -809 -1310
rect -883 -1378 -879 -1375
rect -875 -1375 -861 -1371
rect -875 -1378 -871 -1375
rect -847 -1378 -843 -1375
rect -839 -1375 -820 -1371
rect -839 -1378 -835 -1375
rect -813 -1378 -809 -1331
rect -787 -1342 -783 -1310
rect -787 -1371 -783 -1346
rect -753 -1364 -749 -1310
rect -753 -1368 -736 -1364
rect -805 -1378 -801 -1375
rect -796 -1375 -783 -1371
rect -796 -1378 -792 -1375
rect -769 -1378 -765 -1375
rect -745 -1378 -741 -1368
rect -729 -1371 -725 -1310
rect -721 -1364 -717 -1310
rect -695 -1334 -691 -1310
rect -721 -1368 -702 -1364
rect -737 -1375 -720 -1371
rect -737 -1378 -733 -1375
rect -713 -1378 -709 -1368
rect -695 -1378 -691 -1338
rect -926 -1386 -922 -1382
rect -900 -1386 -896 -1382
rect -857 -1386 -853 -1382
rect -822 -1386 -818 -1382
rect -778 -1386 -774 -1382
rect -761 -1386 -757 -1382
rect -725 -1386 -721 -1382
rect -704 -1386 -700 -1382
rect -688 -1393 -684 -1346
rect -618 -1349 -614 -1187
rect -605 -1334 -601 -840
rect -591 -1162 -587 -816
rect -558 -844 -554 -803
rect -558 -857 -554 -848
rect -577 -861 -554 -857
rect -551 -828 -547 -796
rect -233 -812 -229 -748
rect -219 -788 -215 -784
rect -202 -788 -198 -784
rect -211 -799 -207 -796
rect -211 -803 -196 -799
rect -233 -816 -218 -812
rect -577 -864 -573 -861
rect -551 -864 -547 -832
rect -560 -872 -556 -868
rect -568 -1022 -564 -1018
rect -551 -1022 -547 -1018
rect -531 -1022 -527 -1018
rect -510 -1022 -506 -1018
rect -489 -1022 -485 -1018
rect -468 -1022 -464 -1018
rect -447 -1022 -443 -1018
rect -426 -1022 -422 -1018
rect -405 -1022 -401 -1018
rect -385 -1022 -381 -1018
rect -577 -1077 -573 -1030
rect -577 -1098 -573 -1081
rect -559 -1091 -555 -1030
rect -543 -1091 -539 -1030
rect -519 -1070 -515 -1030
rect -519 -1091 -515 -1074
rect -501 -1091 -497 -1030
rect -477 -1077 -473 -1030
rect -477 -1091 -473 -1081
rect -459 -1070 -455 -1030
rect -459 -1091 -455 -1074
rect -435 -1084 -431 -1030
rect -417 -1062 -413 -1030
rect -417 -1070 -413 -1066
rect -435 -1091 -431 -1088
rect -559 -1095 -550 -1091
rect -543 -1095 -535 -1091
rect -559 -1098 -555 -1095
rect -535 -1098 -531 -1095
rect -527 -1095 -515 -1091
rect -501 -1095 -493 -1091
rect -527 -1098 -523 -1095
rect -493 -1098 -489 -1095
rect -485 -1095 -473 -1091
rect -459 -1095 -447 -1091
rect -485 -1098 -481 -1095
rect -451 -1098 -447 -1095
rect -443 -1095 -431 -1091
rect -417 -1091 -413 -1074
rect -393 -1077 -389 -1030
rect -393 -1091 -389 -1081
rect -417 -1095 -405 -1091
rect -443 -1098 -439 -1095
rect -409 -1098 -405 -1095
rect -401 -1095 -389 -1091
rect -401 -1098 -397 -1095
rect -568 -1106 -564 -1102
rect -551 -1106 -547 -1102
rect -510 -1106 -506 -1102
rect -468 -1106 -464 -1102
rect -426 -1106 -422 -1102
rect -385 -1106 -381 -1102
rect -577 -1138 -573 -1134
rect -560 -1138 -556 -1134
rect -569 -1149 -565 -1146
rect -569 -1153 -554 -1149
rect -591 -1166 -576 -1162
rect -926 -1425 -922 -1421
rect -909 -1425 -905 -1421
rect -889 -1425 -885 -1421
rect -868 -1425 -864 -1421
rect -847 -1425 -843 -1421
rect -826 -1425 -822 -1421
rect -805 -1425 -801 -1421
rect -784 -1425 -780 -1421
rect -763 -1425 -759 -1421
rect -743 -1425 -739 -1421
rect -935 -1480 -931 -1433
rect -935 -1501 -931 -1484
rect -917 -1494 -913 -1433
rect -901 -1494 -897 -1433
rect -877 -1473 -873 -1433
rect -877 -1494 -873 -1477
rect -859 -1494 -855 -1433
rect -835 -1480 -831 -1433
rect -835 -1494 -831 -1484
rect -817 -1473 -813 -1433
rect -817 -1494 -813 -1477
rect -793 -1487 -789 -1433
rect -775 -1465 -771 -1433
rect -775 -1473 -771 -1469
rect -793 -1494 -789 -1491
rect -917 -1498 -908 -1494
rect -901 -1498 -893 -1494
rect -917 -1501 -913 -1498
rect -893 -1501 -889 -1498
rect -885 -1498 -873 -1494
rect -859 -1498 -851 -1494
rect -885 -1501 -881 -1498
rect -851 -1501 -847 -1498
rect -843 -1498 -831 -1494
rect -817 -1498 -805 -1494
rect -843 -1501 -839 -1498
rect -809 -1501 -805 -1498
rect -801 -1498 -789 -1494
rect -775 -1494 -771 -1477
rect -751 -1480 -747 -1433
rect -751 -1494 -747 -1484
rect -775 -1498 -763 -1494
rect -801 -1501 -797 -1498
rect -767 -1501 -763 -1498
rect -759 -1498 -747 -1494
rect -759 -1501 -755 -1498
rect -926 -1509 -922 -1505
rect -909 -1509 -905 -1505
rect -868 -1509 -864 -1505
rect -826 -1509 -822 -1505
rect -784 -1509 -780 -1505
rect -743 -1509 -739 -1505
rect -926 -1596 -922 -1592
rect -909 -1596 -905 -1592
rect -889 -1596 -885 -1592
rect -868 -1596 -864 -1592
rect -847 -1596 -843 -1592
rect -826 -1596 -822 -1592
rect -805 -1596 -801 -1592
rect -784 -1596 -780 -1592
rect -763 -1596 -759 -1592
rect -743 -1596 -739 -1592
rect -935 -1651 -931 -1604
rect -935 -1672 -931 -1655
rect -917 -1665 -913 -1604
rect -901 -1665 -897 -1604
rect -877 -1644 -873 -1604
rect -877 -1665 -873 -1648
rect -859 -1665 -855 -1604
rect -835 -1651 -831 -1604
rect -835 -1665 -831 -1655
rect -817 -1644 -813 -1604
rect -817 -1665 -813 -1648
rect -793 -1658 -789 -1604
rect -775 -1636 -771 -1604
rect -775 -1644 -771 -1640
rect -793 -1665 -789 -1662
rect -917 -1669 -908 -1665
rect -901 -1669 -893 -1665
rect -917 -1672 -913 -1669
rect -893 -1672 -889 -1669
rect -885 -1669 -873 -1665
rect -859 -1669 -851 -1665
rect -885 -1672 -881 -1669
rect -851 -1672 -847 -1669
rect -843 -1669 -831 -1665
rect -817 -1669 -805 -1665
rect -843 -1672 -839 -1669
rect -809 -1672 -805 -1669
rect -801 -1669 -789 -1665
rect -775 -1665 -771 -1648
rect -751 -1651 -747 -1604
rect -751 -1665 -747 -1655
rect -775 -1669 -763 -1665
rect -801 -1672 -797 -1669
rect -767 -1672 -763 -1669
rect -759 -1669 -747 -1665
rect -759 -1672 -755 -1669
rect -926 -1680 -922 -1676
rect -909 -1680 -905 -1676
rect -868 -1680 -864 -1676
rect -826 -1680 -822 -1676
rect -784 -1680 -780 -1676
rect -743 -1680 -739 -1676
rect -730 -1688 -726 -1640
rect -605 -1644 -601 -1411
rect -926 -1767 -922 -1763
rect -909 -1767 -905 -1763
rect -889 -1767 -885 -1763
rect -868 -1767 -864 -1763
rect -847 -1767 -843 -1763
rect -826 -1767 -822 -1763
rect -805 -1767 -801 -1763
rect -784 -1767 -780 -1763
rect -763 -1767 -759 -1763
rect -743 -1767 -739 -1763
rect -935 -1822 -931 -1775
rect -935 -1843 -931 -1826
rect -917 -1836 -913 -1775
rect -901 -1836 -897 -1775
rect -877 -1815 -873 -1775
rect -877 -1836 -873 -1819
rect -859 -1836 -855 -1775
rect -835 -1822 -831 -1775
rect -835 -1836 -831 -1826
rect -817 -1815 -813 -1775
rect -817 -1836 -813 -1819
rect -793 -1829 -789 -1775
rect -775 -1807 -771 -1775
rect -775 -1815 -771 -1811
rect -793 -1836 -789 -1833
rect -917 -1840 -908 -1836
rect -901 -1840 -893 -1836
rect -917 -1843 -913 -1840
rect -893 -1843 -889 -1840
rect -885 -1840 -873 -1836
rect -859 -1840 -851 -1836
rect -885 -1843 -881 -1840
rect -851 -1843 -847 -1840
rect -843 -1840 -831 -1836
rect -817 -1840 -805 -1836
rect -843 -1843 -839 -1840
rect -809 -1843 -805 -1840
rect -801 -1840 -789 -1836
rect -775 -1836 -771 -1819
rect -751 -1822 -747 -1775
rect -751 -1836 -747 -1826
rect -775 -1840 -763 -1836
rect -801 -1843 -797 -1840
rect -767 -1843 -763 -1840
rect -759 -1840 -747 -1836
rect -759 -1843 -755 -1840
rect -926 -1851 -922 -1847
rect -909 -1851 -905 -1847
rect -868 -1851 -864 -1847
rect -826 -1851 -822 -1847
rect -784 -1851 -780 -1847
rect -743 -1851 -739 -1847
rect -935 -1874 -931 -1870
rect -918 -1874 -914 -1870
rect -927 -1885 -923 -1882
rect -927 -1889 -912 -1885
rect -949 -1902 -934 -1898
rect -1208 -2109 -1204 -2106
rect -1199 -2106 -1186 -2102
rect -1199 -2109 -1195 -2106
rect -1172 -2109 -1168 -2106
rect -1164 -2106 -1145 -2102
rect -1164 -2109 -1160 -2106
rect -1138 -2109 -1134 -2077
rect -968 -2080 -964 -1923
rect -1225 -2117 -1221 -2113
rect -1181 -2117 -1177 -2113
rect -1147 -2117 -1143 -2113
rect -1257 -2396 -1253 -2128
rect -1115 -2131 -1111 -2099
rect -1245 -2225 -1241 -2135
rect -1225 -2177 -1221 -2173
rect -1208 -2177 -1204 -2173
rect -1188 -2177 -1184 -2173
rect -1167 -2177 -1163 -2173
rect -1146 -2177 -1142 -2173
rect -1125 -2177 -1121 -2173
rect -1104 -2177 -1100 -2173
rect -1083 -2177 -1079 -2173
rect -1062 -2177 -1058 -2173
rect -1042 -2177 -1038 -2173
rect -1234 -2232 -1230 -2185
rect -1234 -2253 -1230 -2236
rect -1216 -2246 -1212 -2185
rect -1200 -2246 -1196 -2185
rect -1176 -2225 -1172 -2185
rect -1176 -2246 -1172 -2229
rect -1158 -2246 -1154 -2185
rect -1134 -2232 -1130 -2185
rect -1134 -2246 -1130 -2236
rect -1116 -2225 -1112 -2185
rect -1116 -2246 -1112 -2229
rect -1092 -2239 -1088 -2185
rect -1074 -2217 -1070 -2185
rect -1074 -2225 -1070 -2221
rect -1092 -2246 -1088 -2243
rect -1216 -2250 -1207 -2246
rect -1200 -2250 -1192 -2246
rect -1216 -2253 -1212 -2250
rect -1192 -2253 -1188 -2250
rect -1184 -2250 -1172 -2246
rect -1158 -2250 -1150 -2246
rect -1184 -2253 -1180 -2250
rect -1150 -2253 -1146 -2250
rect -1142 -2250 -1130 -2246
rect -1116 -2250 -1104 -2246
rect -1142 -2253 -1138 -2250
rect -1108 -2253 -1104 -2250
rect -1100 -2250 -1088 -2246
rect -1074 -2246 -1070 -2229
rect -1050 -2232 -1046 -2185
rect -1050 -2246 -1046 -2236
rect -1074 -2250 -1062 -2246
rect -1100 -2253 -1096 -2250
rect -1066 -2253 -1062 -2250
rect -1058 -2250 -1046 -2246
rect -1058 -2253 -1054 -2250
rect -1225 -2261 -1221 -2257
rect -1208 -2261 -1204 -2257
rect -1167 -2261 -1163 -2257
rect -1125 -2261 -1121 -2257
rect -1083 -2261 -1079 -2257
rect -1042 -2261 -1038 -2257
rect -1225 -2348 -1221 -2344
rect -1208 -2348 -1204 -2344
rect -1188 -2348 -1184 -2344
rect -1167 -2348 -1163 -2344
rect -1146 -2348 -1142 -2344
rect -1125 -2348 -1121 -2344
rect -1104 -2348 -1100 -2344
rect -1083 -2348 -1079 -2344
rect -1062 -2348 -1058 -2344
rect -1042 -2348 -1038 -2344
rect -1234 -2403 -1230 -2356
rect -1234 -2424 -1230 -2407
rect -1216 -2417 -1212 -2356
rect -1200 -2417 -1196 -2356
rect -1176 -2396 -1172 -2356
rect -1176 -2417 -1172 -2400
rect -1158 -2417 -1154 -2356
rect -1134 -2403 -1130 -2356
rect -1134 -2417 -1130 -2407
rect -1116 -2396 -1112 -2356
rect -1116 -2417 -1112 -2400
rect -1092 -2410 -1088 -2356
rect -1074 -2388 -1070 -2356
rect -1074 -2396 -1070 -2392
rect -1092 -2417 -1088 -2414
rect -1216 -2421 -1207 -2417
rect -1200 -2421 -1192 -2417
rect -1216 -2424 -1212 -2421
rect -1192 -2424 -1188 -2421
rect -1184 -2421 -1172 -2417
rect -1158 -2421 -1150 -2417
rect -1184 -2424 -1180 -2421
rect -1150 -2424 -1146 -2421
rect -1142 -2421 -1130 -2417
rect -1116 -2421 -1104 -2417
rect -1142 -2424 -1138 -2421
rect -1108 -2424 -1104 -2421
rect -1100 -2421 -1088 -2417
rect -1074 -2417 -1070 -2400
rect -1050 -2403 -1046 -2356
rect -1050 -2417 -1046 -2407
rect -1074 -2421 -1062 -2417
rect -1100 -2424 -1096 -2421
rect -1066 -2424 -1062 -2421
rect -1058 -2421 -1046 -2417
rect -1058 -2424 -1054 -2421
rect -1225 -2432 -1221 -2428
rect -1208 -2432 -1204 -2428
rect -1167 -2432 -1163 -2428
rect -1125 -2432 -1121 -2428
rect -1083 -2432 -1079 -2428
rect -1042 -2432 -1038 -2428
rect -1024 -2440 -1020 -2392
rect -963 -2396 -959 -2135
rect -1309 -2624 -1305 -2620
rect -1292 -2624 -1288 -2620
rect -1301 -2635 -1297 -2632
rect -1301 -2639 -1286 -2635
rect -1319 -2652 -1308 -2648
rect -1550 -2902 -1546 -2898
rect -1533 -2902 -1529 -2898
rect -1513 -2902 -1509 -2898
rect -1492 -2902 -1488 -2898
rect -1471 -2902 -1467 -2898
rect -1450 -2902 -1446 -2898
rect -1429 -2902 -1425 -2898
rect -1408 -2902 -1404 -2898
rect -1387 -2902 -1383 -2898
rect -1367 -2902 -1363 -2898
rect -1559 -2957 -1555 -2910
rect -1559 -2978 -1555 -2961
rect -1541 -2971 -1537 -2910
rect -1525 -2971 -1521 -2910
rect -1501 -2950 -1497 -2910
rect -1501 -2971 -1497 -2954
rect -1483 -2971 -1479 -2910
rect -1459 -2957 -1455 -2910
rect -1459 -2971 -1455 -2961
rect -1441 -2950 -1437 -2910
rect -1441 -2971 -1437 -2954
rect -1417 -2964 -1413 -2910
rect -1399 -2942 -1395 -2910
rect -1399 -2950 -1395 -2946
rect -1417 -2971 -1413 -2968
rect -1541 -2975 -1532 -2971
rect -1525 -2975 -1517 -2971
rect -1541 -2978 -1537 -2975
rect -1517 -2978 -1513 -2975
rect -1509 -2975 -1497 -2971
rect -1483 -2975 -1475 -2971
rect -1509 -2978 -1505 -2975
rect -1475 -2978 -1471 -2975
rect -1467 -2975 -1455 -2971
rect -1441 -2975 -1429 -2971
rect -1467 -2978 -1463 -2975
rect -1433 -2978 -1429 -2975
rect -1425 -2975 -1413 -2971
rect -1399 -2971 -1395 -2954
rect -1375 -2957 -1371 -2910
rect -1375 -2971 -1371 -2961
rect -1399 -2975 -1387 -2971
rect -1425 -2978 -1421 -2975
rect -1391 -2978 -1387 -2975
rect -1383 -2975 -1371 -2971
rect -1383 -2978 -1379 -2975
rect -1550 -2986 -1546 -2982
rect -1533 -2986 -1529 -2982
rect -1492 -2986 -1488 -2982
rect -1450 -2986 -1446 -2982
rect -1408 -2986 -1404 -2982
rect -1367 -2986 -1363 -2982
rect -1352 -2993 -1348 -2946
rect -1581 -3121 -1577 -2997
rect -1550 -3073 -1546 -3069
rect -1533 -3073 -1529 -3069
rect -1513 -3073 -1509 -3069
rect -1492 -3073 -1488 -3069
rect -1471 -3073 -1467 -3069
rect -1450 -3073 -1446 -3069
rect -1429 -3073 -1425 -3069
rect -1408 -3073 -1404 -3069
rect -1387 -3073 -1383 -3069
rect -1367 -3073 -1363 -3069
rect -1559 -3128 -1555 -3081
rect -1559 -3149 -1555 -3132
rect -1541 -3142 -1537 -3081
rect -1525 -3142 -1521 -3081
rect -1501 -3121 -1497 -3081
rect -1501 -3142 -1497 -3125
rect -1483 -3142 -1479 -3081
rect -1459 -3128 -1455 -3081
rect -1459 -3142 -1455 -3132
rect -1441 -3121 -1437 -3081
rect -1441 -3142 -1437 -3125
rect -1417 -3135 -1413 -3081
rect -1399 -3113 -1395 -3081
rect -1399 -3121 -1395 -3117
rect -1417 -3142 -1413 -3139
rect -1541 -3146 -1532 -3142
rect -1525 -3146 -1517 -3142
rect -1541 -3149 -1537 -3146
rect -1517 -3149 -1513 -3146
rect -1509 -3146 -1497 -3142
rect -1483 -3146 -1475 -3142
rect -1509 -3149 -1505 -3146
rect -1475 -3149 -1471 -3146
rect -1467 -3146 -1455 -3142
rect -1441 -3146 -1429 -3142
rect -1467 -3149 -1463 -3146
rect -1433 -3149 -1429 -3146
rect -1425 -3146 -1413 -3142
rect -1399 -3142 -1395 -3125
rect -1375 -3128 -1371 -3081
rect -1375 -3142 -1371 -3132
rect -1399 -3146 -1387 -3142
rect -1425 -3149 -1421 -3146
rect -1391 -3149 -1387 -3146
rect -1383 -3146 -1371 -3142
rect -1383 -3149 -1379 -3146
rect -1550 -3157 -1546 -3153
rect -1533 -3157 -1529 -3153
rect -1492 -3157 -1488 -3153
rect -1450 -3157 -1446 -3153
rect -1408 -3157 -1404 -3153
rect -1367 -3157 -1363 -3153
rect -1355 -3164 -1351 -3117
rect -1582 -3292 -1578 -3168
rect -1550 -3244 -1546 -3240
rect -1533 -3244 -1529 -3240
rect -1513 -3244 -1509 -3240
rect -1492 -3244 -1488 -3240
rect -1471 -3244 -1467 -3240
rect -1450 -3244 -1446 -3240
rect -1429 -3244 -1425 -3240
rect -1408 -3244 -1404 -3240
rect -1387 -3244 -1383 -3240
rect -1367 -3244 -1363 -3240
rect -1559 -3299 -1555 -3252
rect -1559 -3320 -1555 -3303
rect -1541 -3313 -1537 -3252
rect -1525 -3313 -1521 -3252
rect -1501 -3292 -1497 -3252
rect -1501 -3313 -1497 -3296
rect -1483 -3313 -1479 -3252
rect -1459 -3299 -1455 -3252
rect -1459 -3313 -1455 -3303
rect -1441 -3292 -1437 -3252
rect -1441 -3313 -1437 -3296
rect -1417 -3306 -1413 -3252
rect -1399 -3284 -1395 -3252
rect -1399 -3292 -1395 -3288
rect -1417 -3313 -1413 -3310
rect -1541 -3317 -1532 -3313
rect -1525 -3317 -1517 -3313
rect -1541 -3320 -1537 -3317
rect -1517 -3320 -1513 -3317
rect -1509 -3317 -1497 -3313
rect -1483 -3317 -1475 -3313
rect -1509 -3320 -1505 -3317
rect -1475 -3320 -1471 -3317
rect -1467 -3317 -1455 -3313
rect -1441 -3317 -1429 -3313
rect -1467 -3320 -1463 -3317
rect -1433 -3320 -1429 -3317
rect -1425 -3317 -1413 -3313
rect -1399 -3313 -1395 -3296
rect -1375 -3299 -1371 -3252
rect -1375 -3313 -1371 -3303
rect -1399 -3317 -1387 -3313
rect -1425 -3320 -1421 -3317
rect -1391 -3320 -1387 -3317
rect -1383 -3317 -1371 -3313
rect -1383 -3320 -1379 -3317
rect -1550 -3328 -1546 -3324
rect -1533 -3328 -1529 -3324
rect -1492 -3328 -1488 -3324
rect -1450 -3328 -1446 -3324
rect -1408 -3328 -1404 -3324
rect -1367 -3328 -1363 -3324
rect -1355 -3387 -1351 -3288
rect -1319 -3292 -1315 -2652
rect -1290 -2678 -1286 -2639
rect -1290 -2693 -1286 -2682
rect -1309 -2697 -1286 -2693
rect -1309 -2700 -1305 -2697
rect -1283 -2700 -1279 -2632
rect -1292 -2708 -1288 -2704
rect -1283 -2838 -1279 -2704
rect -1257 -2831 -1253 -2444
rect -1225 -2519 -1221 -2515
rect -1208 -2519 -1204 -2515
rect -1188 -2519 -1184 -2515
rect -1167 -2519 -1163 -2515
rect -1146 -2519 -1142 -2515
rect -1125 -2519 -1121 -2515
rect -1104 -2519 -1100 -2515
rect -1083 -2519 -1079 -2515
rect -1062 -2519 -1058 -2515
rect -1042 -2519 -1038 -2515
rect -1234 -2574 -1230 -2527
rect -1234 -2595 -1230 -2578
rect -1216 -2588 -1212 -2527
rect -1200 -2588 -1196 -2527
rect -1176 -2567 -1172 -2527
rect -1176 -2588 -1172 -2571
rect -1158 -2588 -1154 -2527
rect -1134 -2574 -1130 -2527
rect -1134 -2588 -1130 -2578
rect -1116 -2567 -1112 -2527
rect -1116 -2588 -1112 -2571
rect -1092 -2581 -1088 -2527
rect -1074 -2559 -1070 -2527
rect -1074 -2567 -1070 -2563
rect -1092 -2588 -1088 -2585
rect -1216 -2592 -1207 -2588
rect -1200 -2592 -1192 -2588
rect -1216 -2595 -1212 -2592
rect -1192 -2595 -1188 -2592
rect -1184 -2592 -1172 -2588
rect -1158 -2592 -1150 -2588
rect -1184 -2595 -1180 -2592
rect -1150 -2595 -1146 -2592
rect -1142 -2592 -1130 -2588
rect -1116 -2592 -1104 -2588
rect -1142 -2595 -1138 -2592
rect -1108 -2595 -1104 -2592
rect -1100 -2592 -1088 -2588
rect -1074 -2588 -1070 -2571
rect -1050 -2574 -1046 -2527
rect -1050 -2588 -1046 -2578
rect -1074 -2592 -1062 -2588
rect -1100 -2595 -1096 -2592
rect -1066 -2595 -1062 -2592
rect -1058 -2592 -1046 -2588
rect -1058 -2595 -1054 -2592
rect -1225 -2603 -1221 -2599
rect -1208 -2603 -1204 -2599
rect -1167 -2603 -1163 -2599
rect -1125 -2603 -1121 -2599
rect -1083 -2603 -1079 -2599
rect -1042 -2603 -1038 -2599
rect -1026 -2648 -1022 -2563
rect -1225 -2783 -1221 -2779
rect -1208 -2783 -1204 -2779
rect -1168 -2783 -1164 -2779
rect -1147 -2783 -1143 -2779
rect -1234 -2824 -1230 -2791
rect -1234 -2859 -1230 -2828
rect -1216 -2818 -1212 -2791
rect -1216 -2822 -1207 -2818
rect -1216 -2859 -1212 -2822
rect -1190 -2845 -1186 -2791
rect -1190 -2852 -1186 -2849
rect -1156 -2852 -1152 -2791
rect -1138 -2823 -1134 -2791
rect -979 -2815 -975 -2673
rect -1208 -2859 -1204 -2856
rect -1199 -2856 -1186 -2852
rect -1199 -2859 -1195 -2856
rect -1172 -2859 -1168 -2856
rect -1164 -2856 -1145 -2852
rect -1164 -2859 -1160 -2856
rect -1138 -2859 -1134 -2827
rect -963 -2830 -959 -2443
rect -949 -2567 -945 -1902
rect -916 -1928 -912 -1889
rect -916 -1943 -912 -1932
rect -935 -1947 -912 -1943
rect -909 -1919 -905 -1882
rect -723 -1898 -719 -1811
rect -935 -1950 -931 -1947
rect -909 -1950 -905 -1923
rect -918 -1958 -914 -1954
rect -926 -2033 -922 -2029
rect -900 -2033 -896 -2029
rect -883 -2033 -879 -2029
rect -843 -2033 -839 -2029
rect -822 -2033 -818 -2029
rect -805 -2033 -801 -2029
rect -765 -2033 -761 -2029
rect -741 -2033 -737 -2029
rect -704 -2033 -700 -2029
rect -935 -2058 -931 -2041
rect -935 -2109 -931 -2062
rect -917 -2051 -913 -2041
rect -917 -2109 -913 -2055
rect -909 -2080 -905 -2041
rect -891 -2073 -887 -2041
rect -909 -2109 -905 -2084
rect -891 -2109 -887 -2077
rect -865 -2065 -861 -2041
rect -865 -2102 -861 -2069
rect -831 -2102 -827 -2041
rect -813 -2058 -809 -2041
rect -883 -2109 -879 -2106
rect -875 -2106 -861 -2102
rect -875 -2109 -871 -2106
rect -847 -2109 -843 -2106
rect -839 -2106 -820 -2102
rect -839 -2109 -835 -2106
rect -813 -2109 -809 -2062
rect -787 -2073 -783 -2041
rect -787 -2102 -783 -2077
rect -753 -2095 -749 -2041
rect -753 -2099 -736 -2095
rect -805 -2109 -801 -2106
rect -796 -2106 -783 -2102
rect -796 -2109 -792 -2106
rect -769 -2109 -765 -2106
rect -745 -2109 -741 -2099
rect -729 -2102 -725 -2041
rect -721 -2095 -717 -2041
rect -695 -2065 -691 -2041
rect -721 -2099 -702 -2095
rect -737 -2106 -720 -2102
rect -737 -2109 -733 -2106
rect -713 -2109 -709 -2099
rect -695 -2109 -691 -2069
rect -926 -2117 -922 -2113
rect -900 -2117 -896 -2113
rect -857 -2117 -853 -2113
rect -822 -2117 -818 -2113
rect -778 -2117 -774 -2113
rect -761 -2117 -757 -2113
rect -725 -2117 -721 -2113
rect -704 -2117 -700 -2113
rect -687 -2124 -683 -2077
rect -618 -2080 -614 -1923
rect -605 -2065 -601 -1692
rect -591 -1815 -587 -1166
rect -558 -1192 -554 -1153
rect -558 -1207 -554 -1196
rect -577 -1211 -554 -1207
rect -551 -1183 -547 -1146
rect -577 -1214 -573 -1211
rect -551 -1214 -547 -1187
rect -560 -1222 -556 -1218
rect -568 -1302 -564 -1298
rect -542 -1302 -538 -1298
rect -525 -1302 -521 -1298
rect -485 -1302 -481 -1298
rect -464 -1302 -460 -1298
rect -447 -1302 -443 -1298
rect -407 -1302 -403 -1298
rect -383 -1302 -379 -1298
rect -346 -1302 -342 -1298
rect -577 -1327 -573 -1310
rect -577 -1378 -573 -1331
rect -559 -1320 -555 -1310
rect -559 -1378 -555 -1324
rect -551 -1349 -547 -1310
rect -533 -1342 -529 -1310
rect -551 -1378 -547 -1353
rect -533 -1378 -529 -1346
rect -507 -1334 -503 -1310
rect -507 -1371 -503 -1338
rect -473 -1371 -469 -1310
rect -455 -1327 -451 -1310
rect -525 -1378 -521 -1375
rect -517 -1375 -503 -1371
rect -517 -1378 -513 -1375
rect -489 -1378 -485 -1375
rect -481 -1375 -462 -1371
rect -481 -1378 -477 -1375
rect -455 -1378 -451 -1331
rect -429 -1342 -425 -1310
rect -429 -1371 -425 -1346
rect -395 -1364 -391 -1310
rect -395 -1368 -378 -1364
rect -447 -1378 -443 -1375
rect -438 -1375 -425 -1371
rect -438 -1378 -434 -1375
rect -411 -1378 -407 -1375
rect -387 -1378 -383 -1368
rect -371 -1371 -367 -1310
rect -363 -1364 -359 -1310
rect -337 -1334 -333 -1310
rect -363 -1368 -344 -1364
rect -379 -1375 -362 -1371
rect -379 -1378 -375 -1375
rect -355 -1378 -351 -1368
rect -337 -1378 -333 -1338
rect -568 -1386 -564 -1382
rect -542 -1386 -538 -1382
rect -499 -1386 -495 -1382
rect -464 -1386 -460 -1382
rect -420 -1386 -416 -1382
rect -403 -1386 -399 -1382
rect -367 -1386 -363 -1382
rect -346 -1386 -342 -1382
rect -328 -1400 -324 -1346
rect -267 -1349 -263 -1187
rect -244 -1334 -240 -832
rect -233 -1162 -229 -816
rect -200 -844 -196 -803
rect -200 -857 -196 -848
rect -219 -861 -196 -857
rect -193 -836 -189 -796
rect 125 -812 129 -748
rect 138 -788 142 -784
rect 155 -788 159 -784
rect 146 -799 150 -796
rect 146 -803 161 -799
rect 125 -816 139 -812
rect -219 -864 -215 -861
rect -193 -864 -189 -840
rect -202 -872 -198 -868
rect -210 -1022 -206 -1018
rect -193 -1022 -189 -1018
rect -173 -1022 -169 -1018
rect -152 -1022 -148 -1018
rect -131 -1022 -127 -1018
rect -110 -1022 -106 -1018
rect -89 -1022 -85 -1018
rect -68 -1022 -64 -1018
rect -47 -1022 -43 -1018
rect -27 -1022 -23 -1018
rect -219 -1077 -215 -1030
rect -219 -1098 -215 -1081
rect -201 -1091 -197 -1030
rect -185 -1091 -181 -1030
rect -161 -1070 -157 -1030
rect -161 -1091 -157 -1074
rect -143 -1091 -139 -1030
rect -119 -1077 -115 -1030
rect -119 -1091 -115 -1081
rect -101 -1070 -97 -1030
rect -101 -1091 -97 -1074
rect -77 -1084 -73 -1030
rect -59 -1062 -55 -1030
rect -59 -1070 -55 -1066
rect -77 -1091 -73 -1088
rect -201 -1095 -192 -1091
rect -185 -1095 -177 -1091
rect -201 -1098 -197 -1095
rect -177 -1098 -173 -1095
rect -169 -1095 -157 -1091
rect -143 -1095 -135 -1091
rect -169 -1098 -165 -1095
rect -135 -1098 -131 -1095
rect -127 -1095 -115 -1091
rect -101 -1095 -89 -1091
rect -127 -1098 -123 -1095
rect -93 -1098 -89 -1095
rect -85 -1095 -73 -1091
rect -59 -1091 -55 -1074
rect -35 -1077 -31 -1030
rect -35 -1091 -31 -1081
rect -59 -1095 -47 -1091
rect -85 -1098 -81 -1095
rect -51 -1098 -47 -1095
rect -43 -1095 -31 -1091
rect -43 -1098 -39 -1095
rect -210 -1106 -206 -1102
rect -193 -1106 -189 -1102
rect -152 -1106 -148 -1102
rect -110 -1106 -106 -1102
rect -68 -1106 -64 -1102
rect -27 -1106 -23 -1102
rect -219 -1138 -215 -1134
rect -202 -1138 -198 -1134
rect -211 -1149 -207 -1146
rect -211 -1153 -196 -1149
rect -233 -1166 -218 -1162
rect -568 -1425 -564 -1421
rect -551 -1425 -547 -1421
rect -531 -1425 -527 -1421
rect -510 -1425 -506 -1421
rect -489 -1425 -485 -1421
rect -468 -1425 -464 -1421
rect -447 -1425 -443 -1421
rect -426 -1425 -422 -1421
rect -405 -1425 -401 -1421
rect -385 -1425 -381 -1421
rect -577 -1480 -573 -1433
rect -577 -1501 -573 -1484
rect -559 -1494 -555 -1433
rect -543 -1494 -539 -1433
rect -519 -1473 -515 -1433
rect -519 -1494 -515 -1477
rect -501 -1494 -497 -1433
rect -477 -1480 -473 -1433
rect -477 -1494 -473 -1484
rect -459 -1473 -455 -1433
rect -459 -1494 -455 -1477
rect -435 -1487 -431 -1433
rect -417 -1465 -413 -1433
rect -417 -1473 -413 -1469
rect -435 -1494 -431 -1491
rect -559 -1498 -550 -1494
rect -543 -1498 -535 -1494
rect -559 -1501 -555 -1498
rect -535 -1501 -531 -1498
rect -527 -1498 -515 -1494
rect -501 -1498 -493 -1494
rect -527 -1501 -523 -1498
rect -493 -1501 -489 -1498
rect -485 -1498 -473 -1494
rect -459 -1498 -447 -1494
rect -485 -1501 -481 -1498
rect -451 -1501 -447 -1498
rect -443 -1498 -431 -1494
rect -417 -1494 -413 -1477
rect -393 -1480 -389 -1433
rect -393 -1494 -389 -1484
rect -417 -1498 -405 -1494
rect -443 -1501 -439 -1498
rect -409 -1501 -405 -1498
rect -401 -1498 -389 -1494
rect -401 -1501 -397 -1498
rect -568 -1509 -564 -1505
rect -551 -1509 -547 -1505
rect -510 -1509 -506 -1505
rect -468 -1509 -464 -1505
rect -426 -1509 -422 -1505
rect -385 -1509 -381 -1505
rect -568 -1596 -564 -1592
rect -551 -1596 -547 -1592
rect -531 -1596 -527 -1592
rect -510 -1596 -506 -1592
rect -489 -1596 -485 -1592
rect -468 -1596 -464 -1592
rect -447 -1596 -443 -1592
rect -426 -1596 -422 -1592
rect -405 -1596 -401 -1592
rect -385 -1596 -381 -1592
rect -577 -1651 -573 -1604
rect -577 -1672 -573 -1655
rect -559 -1665 -555 -1604
rect -543 -1665 -539 -1604
rect -519 -1644 -515 -1604
rect -519 -1665 -515 -1648
rect -501 -1665 -497 -1604
rect -477 -1651 -473 -1604
rect -477 -1665 -473 -1655
rect -459 -1644 -455 -1604
rect -459 -1665 -455 -1648
rect -435 -1658 -431 -1604
rect -417 -1636 -413 -1604
rect -417 -1644 -413 -1640
rect -435 -1665 -431 -1662
rect -559 -1669 -550 -1665
rect -543 -1669 -535 -1665
rect -559 -1672 -555 -1669
rect -535 -1672 -531 -1669
rect -527 -1669 -515 -1665
rect -501 -1669 -493 -1665
rect -527 -1672 -523 -1669
rect -493 -1672 -489 -1669
rect -485 -1669 -473 -1665
rect -459 -1669 -447 -1665
rect -485 -1672 -481 -1669
rect -451 -1672 -447 -1669
rect -443 -1669 -431 -1665
rect -417 -1665 -413 -1648
rect -393 -1651 -389 -1604
rect -393 -1665 -389 -1655
rect -417 -1669 -405 -1665
rect -443 -1672 -439 -1669
rect -409 -1672 -405 -1669
rect -401 -1669 -389 -1665
rect -401 -1672 -397 -1669
rect -568 -1680 -564 -1676
rect -551 -1680 -547 -1676
rect -510 -1680 -506 -1676
rect -468 -1680 -464 -1676
rect -426 -1680 -422 -1676
rect -385 -1680 -381 -1676
rect -368 -1688 -364 -1640
rect -244 -1644 -240 -1404
rect -568 -1767 -564 -1763
rect -551 -1767 -547 -1763
rect -531 -1767 -527 -1763
rect -510 -1767 -506 -1763
rect -489 -1767 -485 -1763
rect -468 -1767 -464 -1763
rect -447 -1767 -443 -1763
rect -426 -1767 -422 -1763
rect -405 -1767 -401 -1763
rect -385 -1767 -381 -1763
rect -577 -1822 -573 -1775
rect -577 -1843 -573 -1826
rect -559 -1836 -555 -1775
rect -543 -1836 -539 -1775
rect -519 -1815 -515 -1775
rect -519 -1836 -515 -1819
rect -501 -1836 -497 -1775
rect -477 -1822 -473 -1775
rect -477 -1836 -473 -1826
rect -459 -1815 -455 -1775
rect -459 -1836 -455 -1819
rect -435 -1829 -431 -1775
rect -417 -1807 -413 -1775
rect -417 -1815 -413 -1811
rect -435 -1836 -431 -1833
rect -559 -1840 -550 -1836
rect -543 -1840 -535 -1836
rect -559 -1843 -555 -1840
rect -535 -1843 -531 -1840
rect -527 -1840 -515 -1836
rect -501 -1840 -493 -1836
rect -527 -1843 -523 -1840
rect -493 -1843 -489 -1840
rect -485 -1840 -473 -1836
rect -459 -1840 -447 -1836
rect -485 -1843 -481 -1840
rect -451 -1843 -447 -1840
rect -443 -1840 -431 -1836
rect -417 -1836 -413 -1819
rect -393 -1822 -389 -1775
rect -393 -1836 -389 -1826
rect -417 -1840 -405 -1836
rect -443 -1843 -439 -1840
rect -409 -1843 -405 -1840
rect -401 -1840 -389 -1836
rect -401 -1843 -397 -1840
rect -568 -1851 -564 -1847
rect -551 -1851 -547 -1847
rect -510 -1851 -506 -1847
rect -468 -1851 -464 -1847
rect -426 -1851 -422 -1847
rect -385 -1851 -381 -1847
rect -577 -1874 -573 -1870
rect -560 -1874 -556 -1870
rect -569 -1885 -565 -1882
rect -569 -1889 -554 -1885
rect -591 -1902 -576 -1898
rect -926 -2177 -922 -2173
rect -909 -2177 -905 -2173
rect -889 -2177 -885 -2173
rect -868 -2177 -864 -2173
rect -847 -2177 -843 -2173
rect -826 -2177 -822 -2173
rect -805 -2177 -801 -2173
rect -784 -2177 -780 -2173
rect -763 -2177 -759 -2173
rect -743 -2177 -739 -2173
rect -935 -2232 -931 -2185
rect -935 -2253 -931 -2236
rect -917 -2246 -913 -2185
rect -901 -2246 -897 -2185
rect -877 -2225 -873 -2185
rect -877 -2246 -873 -2229
rect -859 -2246 -855 -2185
rect -835 -2232 -831 -2185
rect -835 -2246 -831 -2236
rect -817 -2225 -813 -2185
rect -817 -2246 -813 -2229
rect -793 -2239 -789 -2185
rect -775 -2217 -771 -2185
rect -775 -2225 -771 -2221
rect -793 -2246 -789 -2243
rect -917 -2250 -908 -2246
rect -901 -2250 -893 -2246
rect -917 -2253 -913 -2250
rect -893 -2253 -889 -2250
rect -885 -2250 -873 -2246
rect -859 -2250 -851 -2246
rect -885 -2253 -881 -2250
rect -851 -2253 -847 -2250
rect -843 -2250 -831 -2246
rect -817 -2250 -805 -2246
rect -843 -2253 -839 -2250
rect -809 -2253 -805 -2250
rect -801 -2250 -789 -2246
rect -775 -2246 -771 -2229
rect -751 -2232 -747 -2185
rect -751 -2246 -747 -2236
rect -775 -2250 -763 -2246
rect -801 -2253 -797 -2250
rect -767 -2253 -763 -2250
rect -759 -2250 -747 -2246
rect -759 -2253 -755 -2250
rect -926 -2261 -922 -2257
rect -909 -2261 -905 -2257
rect -868 -2261 -864 -2257
rect -826 -2261 -822 -2257
rect -784 -2261 -780 -2257
rect -743 -2261 -739 -2257
rect -926 -2348 -922 -2344
rect -909 -2348 -905 -2344
rect -889 -2348 -885 -2344
rect -868 -2348 -864 -2344
rect -847 -2348 -843 -2344
rect -826 -2348 -822 -2344
rect -805 -2348 -801 -2344
rect -784 -2348 -780 -2344
rect -763 -2348 -759 -2344
rect -743 -2348 -739 -2344
rect -935 -2403 -931 -2356
rect -935 -2424 -931 -2407
rect -917 -2417 -913 -2356
rect -901 -2417 -897 -2356
rect -877 -2396 -873 -2356
rect -877 -2417 -873 -2400
rect -859 -2417 -855 -2356
rect -835 -2403 -831 -2356
rect -835 -2417 -831 -2407
rect -817 -2396 -813 -2356
rect -817 -2417 -813 -2400
rect -793 -2410 -789 -2356
rect -775 -2388 -771 -2356
rect -775 -2396 -771 -2392
rect -793 -2417 -789 -2414
rect -917 -2421 -908 -2417
rect -901 -2421 -893 -2417
rect -917 -2424 -913 -2421
rect -893 -2424 -889 -2421
rect -885 -2421 -873 -2417
rect -859 -2421 -851 -2417
rect -885 -2424 -881 -2421
rect -851 -2424 -847 -2421
rect -843 -2421 -831 -2417
rect -817 -2421 -805 -2417
rect -843 -2424 -839 -2421
rect -809 -2424 -805 -2421
rect -801 -2421 -789 -2417
rect -775 -2417 -771 -2400
rect -751 -2403 -747 -2356
rect -751 -2417 -747 -2407
rect -775 -2421 -763 -2417
rect -801 -2424 -797 -2421
rect -767 -2424 -763 -2421
rect -759 -2421 -747 -2417
rect -759 -2424 -755 -2421
rect -926 -2432 -922 -2428
rect -909 -2432 -905 -2428
rect -868 -2432 -864 -2428
rect -826 -2432 -822 -2428
rect -784 -2432 -780 -2428
rect -743 -2432 -739 -2428
rect -723 -2439 -719 -2392
rect -603 -2396 -599 -2128
rect -926 -2519 -922 -2515
rect -909 -2519 -905 -2515
rect -889 -2519 -885 -2515
rect -868 -2519 -864 -2515
rect -847 -2519 -843 -2515
rect -826 -2519 -822 -2515
rect -805 -2519 -801 -2515
rect -784 -2519 -780 -2515
rect -763 -2519 -759 -2515
rect -743 -2519 -739 -2515
rect -935 -2574 -931 -2527
rect -935 -2595 -931 -2578
rect -917 -2588 -913 -2527
rect -901 -2588 -897 -2527
rect -877 -2567 -873 -2527
rect -877 -2588 -873 -2571
rect -859 -2588 -855 -2527
rect -835 -2574 -831 -2527
rect -835 -2588 -831 -2578
rect -817 -2567 -813 -2527
rect -817 -2588 -813 -2571
rect -793 -2581 -789 -2527
rect -775 -2559 -771 -2527
rect -775 -2567 -771 -2563
rect -793 -2588 -789 -2585
rect -917 -2592 -908 -2588
rect -901 -2592 -893 -2588
rect -917 -2595 -913 -2592
rect -893 -2595 -889 -2592
rect -885 -2592 -873 -2588
rect -859 -2592 -851 -2588
rect -885 -2595 -881 -2592
rect -851 -2595 -847 -2592
rect -843 -2592 -831 -2588
rect -817 -2592 -805 -2588
rect -843 -2595 -839 -2592
rect -809 -2595 -805 -2592
rect -801 -2592 -789 -2588
rect -775 -2588 -771 -2571
rect -751 -2574 -747 -2527
rect -751 -2588 -747 -2578
rect -775 -2592 -763 -2588
rect -801 -2595 -797 -2592
rect -767 -2595 -763 -2592
rect -759 -2592 -747 -2588
rect -759 -2595 -755 -2592
rect -926 -2603 -922 -2599
rect -909 -2603 -905 -2599
rect -868 -2603 -864 -2599
rect -826 -2603 -822 -2599
rect -784 -2603 -780 -2599
rect -743 -2603 -739 -2599
rect -935 -2624 -931 -2620
rect -918 -2624 -914 -2620
rect -927 -2635 -923 -2632
rect -927 -2639 -912 -2635
rect -949 -2652 -934 -2648
rect -1225 -2867 -1221 -2863
rect -1181 -2867 -1177 -2863
rect -1147 -2867 -1143 -2863
rect -1257 -3121 -1253 -2878
rect -1117 -2882 -1113 -2849
rect -1246 -2950 -1242 -2886
rect -1225 -2902 -1221 -2898
rect -1208 -2902 -1204 -2898
rect -1188 -2902 -1184 -2898
rect -1167 -2902 -1163 -2898
rect -1146 -2902 -1142 -2898
rect -1125 -2902 -1121 -2898
rect -1104 -2902 -1100 -2898
rect -1083 -2902 -1079 -2898
rect -1062 -2902 -1058 -2898
rect -1042 -2902 -1038 -2898
rect -1234 -2957 -1230 -2910
rect -1234 -2978 -1230 -2961
rect -1216 -2971 -1212 -2910
rect -1200 -2971 -1196 -2910
rect -1176 -2950 -1172 -2910
rect -1176 -2971 -1172 -2954
rect -1158 -2971 -1154 -2910
rect -1134 -2957 -1130 -2910
rect -1134 -2971 -1130 -2961
rect -1116 -2950 -1112 -2910
rect -1116 -2971 -1112 -2954
rect -1092 -2964 -1088 -2910
rect -1074 -2942 -1070 -2910
rect -1074 -2950 -1070 -2946
rect -1092 -2971 -1088 -2968
rect -1216 -2975 -1207 -2971
rect -1200 -2975 -1192 -2971
rect -1216 -2978 -1212 -2975
rect -1192 -2978 -1188 -2975
rect -1184 -2975 -1172 -2971
rect -1158 -2975 -1150 -2971
rect -1184 -2978 -1180 -2975
rect -1150 -2978 -1146 -2975
rect -1142 -2975 -1130 -2971
rect -1116 -2975 -1104 -2971
rect -1142 -2978 -1138 -2975
rect -1108 -2978 -1104 -2975
rect -1100 -2975 -1088 -2971
rect -1074 -2971 -1070 -2954
rect -1050 -2957 -1046 -2910
rect -1050 -2971 -1046 -2961
rect -1074 -2975 -1062 -2971
rect -1100 -2978 -1096 -2975
rect -1066 -2978 -1062 -2975
rect -1058 -2975 -1046 -2971
rect -1058 -2978 -1054 -2975
rect -1225 -2986 -1221 -2982
rect -1208 -2986 -1204 -2982
rect -1167 -2986 -1163 -2982
rect -1125 -2986 -1121 -2982
rect -1083 -2986 -1079 -2982
rect -1042 -2986 -1038 -2982
rect -1225 -3073 -1221 -3069
rect -1208 -3073 -1204 -3069
rect -1188 -3073 -1184 -3069
rect -1167 -3073 -1163 -3069
rect -1146 -3073 -1142 -3069
rect -1125 -3073 -1121 -3069
rect -1104 -3073 -1100 -3069
rect -1083 -3073 -1079 -3069
rect -1062 -3073 -1058 -3069
rect -1042 -3073 -1038 -3069
rect -1234 -3128 -1230 -3081
rect -1234 -3149 -1230 -3132
rect -1216 -3142 -1212 -3081
rect -1200 -3142 -1196 -3081
rect -1176 -3121 -1172 -3081
rect -1176 -3142 -1172 -3125
rect -1158 -3142 -1154 -3081
rect -1134 -3128 -1130 -3081
rect -1134 -3142 -1130 -3132
rect -1116 -3121 -1112 -3081
rect -1116 -3142 -1112 -3125
rect -1092 -3135 -1088 -3081
rect -1074 -3113 -1070 -3081
rect -1074 -3121 -1070 -3117
rect -1092 -3142 -1088 -3139
rect -1216 -3146 -1207 -3142
rect -1200 -3146 -1192 -3142
rect -1216 -3149 -1212 -3146
rect -1192 -3149 -1188 -3146
rect -1184 -3146 -1172 -3142
rect -1158 -3146 -1150 -3142
rect -1184 -3149 -1180 -3146
rect -1150 -3149 -1146 -3146
rect -1142 -3146 -1130 -3142
rect -1116 -3146 -1104 -3142
rect -1142 -3149 -1138 -3146
rect -1108 -3149 -1104 -3146
rect -1100 -3146 -1088 -3142
rect -1074 -3142 -1070 -3125
rect -1050 -3128 -1046 -3081
rect -1050 -3142 -1046 -3132
rect -1074 -3146 -1062 -3142
rect -1100 -3149 -1096 -3146
rect -1066 -3149 -1062 -3146
rect -1058 -3146 -1046 -3142
rect -1058 -3149 -1054 -3146
rect -1225 -3157 -1221 -3153
rect -1208 -3157 -1204 -3153
rect -1167 -3157 -1163 -3153
rect -1125 -3157 -1121 -3153
rect -1083 -3157 -1079 -3153
rect -1042 -3157 -1038 -3153
rect -1026 -3165 -1022 -3117
rect -963 -3121 -959 -2885
rect -1309 -3355 -1305 -3351
rect -1292 -3355 -1288 -3351
rect -1301 -3366 -1297 -3363
rect -1301 -3370 -1286 -3366
rect -1319 -3383 -1308 -3379
rect -1813 -3644 -1809 -3640
rect -1796 -3644 -1792 -3640
rect -1776 -3644 -1772 -3640
rect -1755 -3644 -1751 -3640
rect -1734 -3644 -1730 -3640
rect -1713 -3644 -1709 -3640
rect -1692 -3644 -1688 -3640
rect -1671 -3644 -1667 -3640
rect -1650 -3644 -1646 -3640
rect -1630 -3644 -1626 -3640
rect -1550 -3644 -1546 -3640
rect -1533 -3644 -1529 -3640
rect -1513 -3644 -1509 -3640
rect -1492 -3644 -1488 -3640
rect -1471 -3644 -1467 -3640
rect -1450 -3644 -1446 -3640
rect -1429 -3644 -1425 -3640
rect -1408 -3644 -1404 -3640
rect -1387 -3644 -1383 -3640
rect -1367 -3644 -1363 -3640
rect -1822 -3699 -1818 -3652
rect -1822 -3720 -1818 -3703
rect -1804 -3713 -1800 -3652
rect -1788 -3713 -1784 -3652
rect -1764 -3692 -1760 -3652
rect -1764 -3713 -1760 -3696
rect -1746 -3713 -1742 -3652
rect -1722 -3699 -1718 -3652
rect -1722 -3713 -1718 -3703
rect -1704 -3692 -1700 -3652
rect -1704 -3713 -1700 -3696
rect -1680 -3706 -1676 -3652
rect -1662 -3684 -1658 -3652
rect -1662 -3692 -1658 -3688
rect -1680 -3713 -1676 -3710
rect -1804 -3717 -1795 -3713
rect -1788 -3717 -1780 -3713
rect -1804 -3720 -1800 -3717
rect -1780 -3720 -1776 -3717
rect -1772 -3717 -1760 -3713
rect -1746 -3717 -1738 -3713
rect -1772 -3720 -1768 -3717
rect -1738 -3720 -1734 -3717
rect -1730 -3717 -1718 -3713
rect -1704 -3717 -1692 -3713
rect -1730 -3720 -1726 -3717
rect -1696 -3720 -1692 -3717
rect -1688 -3717 -1676 -3713
rect -1662 -3713 -1658 -3696
rect -1638 -3699 -1634 -3652
rect -1638 -3713 -1634 -3703
rect -1662 -3717 -1650 -3713
rect -1688 -3720 -1684 -3717
rect -1654 -3720 -1650 -3717
rect -1646 -3717 -1634 -3713
rect -1559 -3699 -1555 -3652
rect -1646 -3720 -1642 -3717
rect -1559 -3720 -1555 -3703
rect -1541 -3713 -1537 -3652
rect -1525 -3713 -1521 -3652
rect -1501 -3692 -1497 -3652
rect -1501 -3713 -1497 -3696
rect -1483 -3713 -1479 -3652
rect -1459 -3699 -1455 -3652
rect -1459 -3713 -1455 -3703
rect -1441 -3692 -1437 -3652
rect -1441 -3713 -1437 -3696
rect -1417 -3706 -1413 -3652
rect -1399 -3684 -1395 -3652
rect -1399 -3692 -1395 -3688
rect -1417 -3713 -1413 -3710
rect -1541 -3717 -1532 -3713
rect -1525 -3717 -1517 -3713
rect -1541 -3720 -1537 -3717
rect -1517 -3720 -1513 -3717
rect -1509 -3717 -1497 -3713
rect -1483 -3717 -1475 -3713
rect -1509 -3720 -1505 -3717
rect -1475 -3720 -1471 -3717
rect -1467 -3717 -1455 -3713
rect -1441 -3717 -1429 -3713
rect -1467 -3720 -1463 -3717
rect -1433 -3720 -1429 -3717
rect -1425 -3717 -1413 -3713
rect -1399 -3713 -1395 -3696
rect -1375 -3699 -1371 -3652
rect -1375 -3713 -1371 -3703
rect -1399 -3717 -1387 -3713
rect -1425 -3720 -1421 -3717
rect -1391 -3720 -1387 -3717
rect -1383 -3717 -1371 -3713
rect -1383 -3720 -1379 -3717
rect -1813 -3728 -1809 -3724
rect -1796 -3728 -1792 -3724
rect -1755 -3728 -1751 -3724
rect -1713 -3728 -1709 -3724
rect -1671 -3728 -1667 -3724
rect -1630 -3728 -1626 -3724
rect -1550 -3728 -1546 -3724
rect -1533 -3728 -1529 -3724
rect -1492 -3728 -1488 -3724
rect -1450 -3728 -1446 -3724
rect -1408 -3728 -1404 -3724
rect -1367 -3728 -1363 -3724
rect -1353 -3736 -1349 -3688
rect -1572 -3863 -1568 -3740
rect -1550 -3815 -1546 -3811
rect -1533 -3815 -1529 -3811
rect -1513 -3815 -1509 -3811
rect -1492 -3815 -1488 -3811
rect -1471 -3815 -1467 -3811
rect -1450 -3815 -1446 -3811
rect -1429 -3815 -1425 -3811
rect -1408 -3815 -1404 -3811
rect -1387 -3815 -1383 -3811
rect -1367 -3815 -1363 -3811
rect -1559 -3870 -1555 -3823
rect -1559 -3891 -1555 -3874
rect -1541 -3884 -1537 -3823
rect -1525 -3884 -1521 -3823
rect -1501 -3863 -1497 -3823
rect -1501 -3884 -1497 -3867
rect -1483 -3884 -1479 -3823
rect -1459 -3870 -1455 -3823
rect -1459 -3884 -1455 -3874
rect -1441 -3863 -1437 -3823
rect -1441 -3884 -1437 -3867
rect -1417 -3877 -1413 -3823
rect -1399 -3855 -1395 -3823
rect -1399 -3863 -1395 -3859
rect -1417 -3884 -1413 -3881
rect -1541 -3888 -1532 -3884
rect -1525 -3888 -1517 -3884
rect -1541 -3891 -1537 -3888
rect -1517 -3891 -1513 -3888
rect -1509 -3888 -1497 -3884
rect -1483 -3888 -1475 -3884
rect -1509 -3891 -1505 -3888
rect -1475 -3891 -1471 -3888
rect -1467 -3888 -1455 -3884
rect -1441 -3888 -1429 -3884
rect -1467 -3891 -1463 -3888
rect -1433 -3891 -1429 -3888
rect -1425 -3888 -1413 -3884
rect -1399 -3884 -1395 -3867
rect -1375 -3870 -1371 -3823
rect -1375 -3884 -1371 -3874
rect -1399 -3888 -1387 -3884
rect -1425 -3891 -1421 -3888
rect -1391 -3891 -1387 -3888
rect -1383 -3888 -1371 -3884
rect -1383 -3891 -1379 -3888
rect -1550 -3899 -1546 -3895
rect -1533 -3899 -1529 -3895
rect -1492 -3899 -1488 -3895
rect -1450 -3899 -1446 -3895
rect -1408 -3899 -1404 -3895
rect -1367 -3899 -1363 -3895
rect -1355 -3907 -1351 -3859
rect -1575 -4038 -1571 -3911
rect -1550 -3990 -1546 -3986
rect -1533 -3990 -1529 -3986
rect -1513 -3990 -1509 -3986
rect -1492 -3990 -1488 -3986
rect -1471 -3990 -1467 -3986
rect -1450 -3990 -1446 -3986
rect -1429 -3990 -1425 -3986
rect -1408 -3990 -1404 -3986
rect -1387 -3990 -1383 -3986
rect -1367 -3990 -1363 -3986
rect -1559 -4045 -1555 -3998
rect -1559 -4066 -1555 -4049
rect -1541 -4059 -1537 -3998
rect -1525 -4059 -1521 -3998
rect -1501 -4038 -1497 -3998
rect -1501 -4059 -1497 -4042
rect -1483 -4059 -1479 -3998
rect -1459 -4045 -1455 -3998
rect -1459 -4059 -1455 -4049
rect -1441 -4038 -1437 -3998
rect -1441 -4059 -1437 -4042
rect -1417 -4052 -1413 -3998
rect -1399 -4030 -1395 -3998
rect -1399 -4038 -1395 -4034
rect -1417 -4059 -1413 -4056
rect -1541 -4063 -1532 -4059
rect -1525 -4063 -1517 -4059
rect -1541 -4066 -1537 -4063
rect -1517 -4066 -1513 -4063
rect -1509 -4063 -1497 -4059
rect -1483 -4063 -1475 -4059
rect -1509 -4066 -1505 -4063
rect -1475 -4066 -1471 -4063
rect -1467 -4063 -1455 -4059
rect -1441 -4063 -1429 -4059
rect -1467 -4066 -1463 -4063
rect -1433 -4066 -1429 -4063
rect -1425 -4063 -1413 -4059
rect -1399 -4059 -1395 -4042
rect -1375 -4045 -1371 -3998
rect -1375 -4059 -1371 -4049
rect -1399 -4063 -1387 -4059
rect -1425 -4066 -1421 -4063
rect -1391 -4066 -1387 -4063
rect -1383 -4063 -1371 -4059
rect -1383 -4066 -1379 -4063
rect -1550 -4074 -1546 -4070
rect -1533 -4074 -1529 -4070
rect -1492 -4074 -1488 -4070
rect -1450 -4074 -1446 -4070
rect -1408 -4074 -1404 -4070
rect -1367 -4074 -1363 -4070
rect -1357 -4137 -1353 -4034
rect -1319 -4038 -1315 -3383
rect -1290 -3409 -1286 -3370
rect -1290 -3424 -1286 -3413
rect -1309 -3428 -1286 -3424
rect -1309 -3431 -1305 -3428
rect -1283 -3431 -1279 -3363
rect -1292 -3439 -1288 -3435
rect -1283 -3569 -1279 -3435
rect -1257 -3562 -1253 -3169
rect -1225 -3244 -1221 -3240
rect -1208 -3244 -1204 -3240
rect -1188 -3244 -1184 -3240
rect -1167 -3244 -1163 -3240
rect -1146 -3244 -1142 -3240
rect -1125 -3244 -1121 -3240
rect -1104 -3244 -1100 -3240
rect -1083 -3244 -1079 -3240
rect -1062 -3244 -1058 -3240
rect -1042 -3244 -1038 -3240
rect -1234 -3299 -1230 -3252
rect -1234 -3320 -1230 -3303
rect -1216 -3313 -1212 -3252
rect -1200 -3313 -1196 -3252
rect -1176 -3292 -1172 -3252
rect -1176 -3313 -1172 -3296
rect -1158 -3313 -1154 -3252
rect -1134 -3299 -1130 -3252
rect -1134 -3313 -1130 -3303
rect -1116 -3292 -1112 -3252
rect -1116 -3313 -1112 -3296
rect -1092 -3306 -1088 -3252
rect -1074 -3284 -1070 -3252
rect -1074 -3292 -1070 -3288
rect -1092 -3313 -1088 -3310
rect -1216 -3317 -1207 -3313
rect -1200 -3317 -1192 -3313
rect -1216 -3320 -1212 -3317
rect -1192 -3320 -1188 -3317
rect -1184 -3317 -1172 -3313
rect -1158 -3317 -1150 -3313
rect -1184 -3320 -1180 -3317
rect -1150 -3320 -1146 -3317
rect -1142 -3317 -1130 -3313
rect -1116 -3317 -1104 -3313
rect -1142 -3320 -1138 -3317
rect -1108 -3320 -1104 -3317
rect -1100 -3317 -1088 -3313
rect -1074 -3313 -1070 -3296
rect -1050 -3299 -1046 -3252
rect -1050 -3313 -1046 -3303
rect -1074 -3317 -1062 -3313
rect -1100 -3320 -1096 -3317
rect -1066 -3320 -1062 -3317
rect -1058 -3317 -1046 -3313
rect -1058 -3320 -1054 -3317
rect -1225 -3328 -1221 -3324
rect -1208 -3328 -1204 -3324
rect -1167 -3328 -1163 -3324
rect -1125 -3328 -1121 -3324
rect -1083 -3328 -1079 -3324
rect -1042 -3328 -1038 -3324
rect -1026 -3379 -1022 -3288
rect -1225 -3514 -1221 -3510
rect -1208 -3514 -1204 -3510
rect -1168 -3514 -1164 -3510
rect -1147 -3514 -1143 -3510
rect -1234 -3555 -1230 -3522
rect -1234 -3590 -1230 -3559
rect -1216 -3549 -1212 -3522
rect -1216 -3553 -1207 -3549
rect -1216 -3590 -1212 -3553
rect -1190 -3576 -1186 -3522
rect -1190 -3583 -1186 -3580
rect -1156 -3583 -1152 -3522
rect -1138 -3554 -1134 -3522
rect -979 -3546 -975 -3404
rect -1208 -3590 -1204 -3587
rect -1199 -3587 -1186 -3583
rect -1199 -3590 -1195 -3587
rect -1172 -3590 -1168 -3587
rect -1164 -3587 -1145 -3583
rect -1164 -3590 -1160 -3587
rect -1138 -3590 -1134 -3558
rect -963 -3561 -959 -3169
rect -949 -3292 -945 -2652
rect -916 -2678 -912 -2639
rect -916 -2693 -912 -2682
rect -935 -2697 -912 -2693
rect -909 -2669 -905 -2632
rect -720 -2648 -716 -2563
rect -935 -2700 -931 -2697
rect -909 -2700 -905 -2673
rect -918 -2708 -914 -2704
rect -926 -2783 -922 -2779
rect -900 -2783 -896 -2779
rect -883 -2783 -879 -2779
rect -843 -2783 -839 -2779
rect -822 -2783 -818 -2779
rect -805 -2783 -801 -2779
rect -765 -2783 -761 -2779
rect -741 -2783 -737 -2779
rect -704 -2783 -700 -2779
rect -935 -2808 -931 -2791
rect -935 -2859 -931 -2812
rect -917 -2801 -913 -2791
rect -917 -2859 -913 -2805
rect -909 -2830 -905 -2791
rect -891 -2823 -887 -2791
rect -909 -2859 -905 -2834
rect -891 -2859 -887 -2827
rect -865 -2815 -861 -2791
rect -865 -2852 -861 -2819
rect -831 -2852 -827 -2791
rect -813 -2808 -809 -2791
rect -883 -2859 -879 -2856
rect -875 -2856 -861 -2852
rect -875 -2859 -871 -2856
rect -847 -2859 -843 -2856
rect -839 -2856 -820 -2852
rect -839 -2859 -835 -2856
rect -813 -2859 -809 -2812
rect -787 -2823 -783 -2791
rect -787 -2852 -783 -2827
rect -753 -2845 -749 -2791
rect -753 -2849 -736 -2845
rect -805 -2859 -801 -2856
rect -796 -2856 -783 -2852
rect -796 -2859 -792 -2856
rect -769 -2859 -765 -2856
rect -745 -2859 -741 -2849
rect -729 -2852 -725 -2791
rect -721 -2845 -717 -2791
rect -695 -2815 -691 -2791
rect -721 -2849 -702 -2845
rect -737 -2856 -720 -2852
rect -737 -2859 -733 -2856
rect -713 -2859 -709 -2849
rect -695 -2859 -691 -2819
rect -926 -2867 -922 -2863
rect -900 -2867 -896 -2863
rect -857 -2867 -853 -2863
rect -822 -2867 -818 -2863
rect -778 -2867 -774 -2863
rect -761 -2867 -757 -2863
rect -725 -2867 -721 -2863
rect -704 -2867 -700 -2863
rect -688 -2874 -684 -2827
rect -616 -2830 -612 -2673
rect -603 -2815 -599 -2444
rect -591 -2567 -587 -1902
rect -558 -1928 -554 -1889
rect -558 -1943 -554 -1932
rect -577 -1947 -554 -1943
rect -551 -1919 -547 -1882
rect -366 -1898 -362 -1811
rect -577 -1950 -573 -1947
rect -551 -1950 -547 -1923
rect -560 -1958 -556 -1954
rect -568 -2033 -564 -2029
rect -542 -2033 -538 -2029
rect -525 -2033 -521 -2029
rect -485 -2033 -481 -2029
rect -464 -2033 -460 -2029
rect -447 -2033 -443 -2029
rect -407 -2033 -403 -2029
rect -383 -2033 -379 -2029
rect -346 -2033 -342 -2029
rect -577 -2058 -573 -2041
rect -577 -2109 -573 -2062
rect -559 -2051 -555 -2041
rect -559 -2109 -555 -2055
rect -551 -2080 -547 -2041
rect -533 -2073 -529 -2041
rect -551 -2109 -547 -2084
rect -533 -2109 -529 -2077
rect -507 -2065 -503 -2041
rect -507 -2102 -503 -2069
rect -473 -2102 -469 -2041
rect -455 -2058 -451 -2041
rect -525 -2109 -521 -2106
rect -517 -2106 -503 -2102
rect -517 -2109 -513 -2106
rect -489 -2109 -485 -2106
rect -481 -2106 -462 -2102
rect -481 -2109 -477 -2106
rect -455 -2109 -451 -2062
rect -429 -2073 -425 -2041
rect -429 -2102 -425 -2077
rect -395 -2095 -391 -2041
rect -395 -2099 -378 -2095
rect -447 -2109 -443 -2106
rect -438 -2106 -425 -2102
rect -438 -2109 -434 -2106
rect -411 -2109 -407 -2106
rect -387 -2109 -383 -2099
rect -371 -2102 -367 -2041
rect -363 -2095 -359 -2041
rect -337 -2062 -333 -2041
rect -363 -2099 -344 -2095
rect -379 -2106 -362 -2102
rect -379 -2109 -375 -2106
rect -355 -2109 -351 -2099
rect -337 -2109 -333 -2066
rect -568 -2117 -564 -2113
rect -542 -2117 -538 -2113
rect -499 -2117 -495 -2113
rect -464 -2117 -460 -2113
rect -420 -2117 -416 -2113
rect -403 -2117 -399 -2113
rect -367 -2117 -363 -2113
rect -346 -2117 -342 -2113
rect -328 -2131 -324 -2077
rect -262 -2080 -258 -1923
rect -244 -2065 -240 -1691
rect -233 -1815 -229 -1166
rect -200 -1192 -196 -1153
rect -200 -1207 -196 -1196
rect -219 -1211 -196 -1207
rect -193 -1183 -189 -1146
rect -219 -1214 -215 -1211
rect -193 -1214 -189 -1187
rect -202 -1222 -198 -1218
rect -210 -1302 -206 -1298
rect -184 -1302 -180 -1298
rect -167 -1302 -163 -1298
rect -127 -1302 -123 -1298
rect -106 -1302 -102 -1298
rect -89 -1302 -85 -1298
rect -49 -1302 -45 -1298
rect -25 -1302 -21 -1298
rect 12 -1302 16 -1298
rect -219 -1327 -215 -1310
rect -219 -1378 -215 -1331
rect -201 -1320 -197 -1310
rect -201 -1378 -197 -1324
rect -193 -1349 -189 -1310
rect -175 -1342 -171 -1310
rect -193 -1378 -189 -1353
rect -175 -1378 -171 -1346
rect -149 -1334 -145 -1310
rect -149 -1371 -145 -1338
rect -115 -1371 -111 -1310
rect -97 -1327 -93 -1310
rect -167 -1378 -163 -1375
rect -159 -1375 -145 -1371
rect -159 -1378 -155 -1375
rect -131 -1378 -127 -1375
rect -123 -1375 -104 -1371
rect -123 -1378 -119 -1375
rect -97 -1378 -93 -1331
rect -71 -1342 -67 -1310
rect -71 -1371 -67 -1346
rect -37 -1364 -33 -1310
rect -37 -1368 -20 -1364
rect -89 -1378 -85 -1375
rect -80 -1375 -67 -1371
rect -80 -1378 -76 -1375
rect -53 -1378 -49 -1375
rect -29 -1378 -25 -1368
rect -13 -1371 -9 -1310
rect -5 -1364 -1 -1310
rect 21 -1334 25 -1310
rect -5 -1368 14 -1364
rect -21 -1375 -4 -1371
rect -21 -1378 -17 -1375
rect 3 -1378 7 -1368
rect 21 -1378 25 -1338
rect -210 -1386 -206 -1382
rect -184 -1386 -180 -1382
rect -141 -1386 -137 -1382
rect -106 -1386 -102 -1382
rect -62 -1386 -58 -1382
rect -45 -1386 -41 -1382
rect -9 -1386 -5 -1382
rect 12 -1386 16 -1382
rect 29 -1407 33 -1346
rect 91 -1349 95 -1187
rect 107 -1334 111 -840
rect 125 -1162 129 -816
rect 157 -857 161 -803
rect 138 -861 157 -857
rect 164 -828 168 -796
rect 481 -812 485 -748
rect 495 -788 499 -784
rect 512 -788 516 -784
rect 503 -799 507 -796
rect 503 -803 518 -799
rect 481 -816 496 -812
rect 138 -864 142 -861
rect 164 -864 168 -832
rect 155 -872 159 -868
rect 148 -1022 152 -1018
rect 165 -1022 169 -1018
rect 185 -1022 189 -1018
rect 206 -1022 210 -1018
rect 227 -1022 231 -1018
rect 248 -1022 252 -1018
rect 269 -1022 273 -1018
rect 290 -1022 294 -1018
rect 311 -1022 315 -1018
rect 331 -1022 335 -1018
rect 139 -1077 143 -1030
rect 139 -1098 143 -1081
rect 157 -1091 161 -1030
rect 173 -1091 177 -1030
rect 197 -1070 201 -1030
rect 197 -1091 201 -1074
rect 215 -1091 219 -1030
rect 239 -1077 243 -1030
rect 239 -1091 243 -1081
rect 257 -1070 261 -1030
rect 257 -1091 261 -1074
rect 281 -1084 285 -1030
rect 299 -1062 303 -1030
rect 299 -1070 303 -1066
rect 281 -1091 285 -1088
rect 157 -1095 166 -1091
rect 173 -1095 181 -1091
rect 157 -1098 161 -1095
rect 181 -1098 185 -1095
rect 189 -1095 201 -1091
rect 215 -1095 223 -1091
rect 189 -1098 193 -1095
rect 223 -1098 227 -1095
rect 231 -1095 243 -1091
rect 257 -1095 269 -1091
rect 231 -1098 235 -1095
rect 265 -1098 269 -1095
rect 273 -1095 285 -1091
rect 299 -1091 303 -1074
rect 323 -1077 327 -1030
rect 323 -1091 327 -1081
rect 299 -1095 311 -1091
rect 273 -1098 277 -1095
rect 307 -1098 311 -1095
rect 315 -1095 327 -1091
rect 315 -1098 319 -1095
rect 148 -1106 152 -1102
rect 165 -1106 169 -1102
rect 206 -1106 210 -1102
rect 248 -1106 252 -1102
rect 290 -1106 294 -1102
rect 331 -1106 335 -1102
rect 139 -1138 143 -1134
rect 156 -1138 160 -1134
rect 147 -1149 151 -1146
rect 147 -1153 162 -1149
rect 125 -1166 140 -1162
rect -210 -1425 -206 -1421
rect -193 -1425 -189 -1421
rect -173 -1425 -169 -1421
rect -152 -1425 -148 -1421
rect -131 -1425 -127 -1421
rect -110 -1425 -106 -1421
rect -89 -1425 -85 -1421
rect -68 -1425 -64 -1421
rect -47 -1425 -43 -1421
rect -27 -1425 -23 -1421
rect -219 -1480 -215 -1433
rect -219 -1501 -215 -1484
rect -201 -1494 -197 -1433
rect -185 -1494 -181 -1433
rect -161 -1473 -157 -1433
rect -161 -1494 -157 -1477
rect -143 -1494 -139 -1433
rect -119 -1480 -115 -1433
rect -119 -1494 -115 -1484
rect -101 -1473 -97 -1433
rect -101 -1494 -97 -1477
rect -77 -1487 -73 -1433
rect -59 -1465 -55 -1433
rect -59 -1473 -55 -1469
rect -77 -1494 -73 -1491
rect -201 -1498 -192 -1494
rect -185 -1498 -177 -1494
rect -201 -1501 -197 -1498
rect -177 -1501 -173 -1498
rect -169 -1498 -157 -1494
rect -143 -1498 -135 -1494
rect -169 -1501 -165 -1498
rect -135 -1501 -131 -1498
rect -127 -1498 -115 -1494
rect -101 -1498 -89 -1494
rect -127 -1501 -123 -1498
rect -93 -1501 -89 -1498
rect -85 -1498 -73 -1494
rect -59 -1494 -55 -1477
rect -35 -1480 -31 -1433
rect -35 -1494 -31 -1484
rect -59 -1498 -47 -1494
rect -85 -1501 -81 -1498
rect -51 -1501 -47 -1498
rect -43 -1498 -31 -1494
rect -43 -1501 -39 -1498
rect -210 -1509 -206 -1505
rect -193 -1509 -189 -1505
rect -152 -1509 -148 -1505
rect -110 -1509 -106 -1505
rect -68 -1509 -64 -1505
rect -27 -1509 -23 -1505
rect -210 -1596 -206 -1592
rect -193 -1596 -189 -1592
rect -173 -1596 -169 -1592
rect -152 -1596 -148 -1592
rect -131 -1596 -127 -1592
rect -110 -1596 -106 -1592
rect -89 -1596 -85 -1592
rect -68 -1596 -64 -1592
rect -47 -1596 -43 -1592
rect -27 -1596 -23 -1592
rect -219 -1651 -215 -1604
rect -219 -1672 -215 -1655
rect -201 -1665 -197 -1604
rect -185 -1665 -181 -1604
rect -161 -1644 -157 -1604
rect -161 -1665 -157 -1648
rect -143 -1665 -139 -1604
rect -119 -1651 -115 -1604
rect -119 -1665 -115 -1655
rect -101 -1644 -97 -1604
rect -101 -1665 -97 -1648
rect -77 -1658 -73 -1604
rect -59 -1636 -55 -1604
rect -59 -1644 -55 -1640
rect -77 -1665 -73 -1662
rect -201 -1669 -192 -1665
rect -185 -1669 -177 -1665
rect -201 -1672 -197 -1669
rect -177 -1672 -173 -1669
rect -169 -1669 -157 -1665
rect -143 -1669 -135 -1665
rect -169 -1672 -165 -1669
rect -135 -1672 -131 -1669
rect -127 -1669 -115 -1665
rect -101 -1669 -89 -1665
rect -127 -1672 -123 -1669
rect -93 -1672 -89 -1669
rect -85 -1669 -73 -1665
rect -59 -1665 -55 -1648
rect -35 -1651 -31 -1604
rect -35 -1665 -31 -1655
rect -59 -1669 -47 -1665
rect -85 -1672 -81 -1669
rect -51 -1672 -47 -1669
rect -43 -1669 -31 -1665
rect -43 -1672 -39 -1669
rect -210 -1680 -206 -1676
rect -193 -1680 -189 -1676
rect -152 -1680 -148 -1676
rect -110 -1680 -106 -1676
rect -68 -1680 -64 -1676
rect -27 -1680 -23 -1676
rect -12 -1687 -8 -1640
rect 107 -1644 111 -1411
rect -210 -1767 -206 -1763
rect -193 -1767 -189 -1763
rect -173 -1767 -169 -1763
rect -152 -1767 -148 -1763
rect -131 -1767 -127 -1763
rect -110 -1767 -106 -1763
rect -89 -1767 -85 -1763
rect -68 -1767 -64 -1763
rect -47 -1767 -43 -1763
rect -27 -1767 -23 -1763
rect -219 -1822 -215 -1775
rect -219 -1843 -215 -1826
rect -201 -1836 -197 -1775
rect -185 -1836 -181 -1775
rect -161 -1815 -157 -1775
rect -161 -1836 -157 -1819
rect -143 -1836 -139 -1775
rect -119 -1822 -115 -1775
rect -119 -1836 -115 -1826
rect -101 -1815 -97 -1775
rect -101 -1836 -97 -1819
rect -77 -1829 -73 -1775
rect -59 -1807 -55 -1775
rect -59 -1815 -55 -1811
rect -77 -1836 -73 -1833
rect -201 -1840 -192 -1836
rect -185 -1840 -177 -1836
rect -201 -1843 -197 -1840
rect -177 -1843 -173 -1840
rect -169 -1840 -157 -1836
rect -143 -1840 -135 -1836
rect -169 -1843 -165 -1840
rect -135 -1843 -131 -1840
rect -127 -1840 -115 -1836
rect -101 -1840 -89 -1836
rect -127 -1843 -123 -1840
rect -93 -1843 -89 -1840
rect -85 -1840 -73 -1836
rect -59 -1836 -55 -1819
rect -35 -1822 -31 -1775
rect -35 -1836 -31 -1826
rect -59 -1840 -47 -1836
rect -85 -1843 -81 -1840
rect -51 -1843 -47 -1840
rect -43 -1840 -31 -1836
rect -43 -1843 -39 -1840
rect -210 -1851 -206 -1847
rect -193 -1851 -189 -1847
rect -152 -1851 -148 -1847
rect -110 -1851 -106 -1847
rect -68 -1851 -64 -1847
rect -27 -1851 -23 -1847
rect -219 -1874 -215 -1870
rect -202 -1874 -198 -1870
rect -211 -1885 -207 -1882
rect -211 -1889 -196 -1885
rect -233 -1902 -218 -1898
rect -568 -2177 -564 -2173
rect -551 -2177 -547 -2173
rect -531 -2177 -527 -2173
rect -510 -2177 -506 -2173
rect -489 -2177 -485 -2173
rect -468 -2177 -464 -2173
rect -447 -2177 -443 -2173
rect -426 -2177 -422 -2173
rect -405 -2177 -401 -2173
rect -385 -2177 -381 -2173
rect -577 -2232 -573 -2185
rect -577 -2253 -573 -2236
rect -559 -2246 -555 -2185
rect -543 -2246 -539 -2185
rect -519 -2225 -515 -2185
rect -519 -2246 -515 -2229
rect -501 -2246 -497 -2185
rect -477 -2232 -473 -2185
rect -477 -2246 -473 -2236
rect -459 -2225 -455 -2185
rect -459 -2246 -455 -2229
rect -435 -2239 -431 -2185
rect -417 -2217 -413 -2185
rect -417 -2225 -413 -2221
rect -435 -2246 -431 -2243
rect -559 -2250 -550 -2246
rect -543 -2250 -535 -2246
rect -559 -2253 -555 -2250
rect -535 -2253 -531 -2250
rect -527 -2250 -515 -2246
rect -501 -2250 -493 -2246
rect -527 -2253 -523 -2250
rect -493 -2253 -489 -2250
rect -485 -2250 -473 -2246
rect -459 -2250 -447 -2246
rect -485 -2253 -481 -2250
rect -451 -2253 -447 -2250
rect -443 -2250 -431 -2246
rect -417 -2246 -413 -2229
rect -393 -2232 -389 -2185
rect -393 -2246 -389 -2236
rect -417 -2250 -405 -2246
rect -443 -2253 -439 -2250
rect -409 -2253 -405 -2250
rect -401 -2250 -389 -2246
rect -401 -2253 -397 -2250
rect -568 -2261 -564 -2257
rect -551 -2261 -547 -2257
rect -510 -2261 -506 -2257
rect -468 -2261 -464 -2257
rect -426 -2261 -422 -2257
rect -385 -2261 -381 -2257
rect -568 -2348 -564 -2344
rect -551 -2348 -547 -2344
rect -531 -2348 -527 -2344
rect -510 -2348 -506 -2344
rect -489 -2348 -485 -2344
rect -468 -2348 -464 -2344
rect -447 -2348 -443 -2344
rect -426 -2348 -422 -2344
rect -405 -2348 -401 -2344
rect -385 -2348 -381 -2344
rect -577 -2403 -573 -2356
rect -577 -2424 -573 -2407
rect -559 -2417 -555 -2356
rect -543 -2417 -539 -2356
rect -519 -2396 -515 -2356
rect -519 -2417 -515 -2400
rect -501 -2417 -497 -2356
rect -477 -2403 -473 -2356
rect -477 -2417 -473 -2407
rect -459 -2396 -455 -2356
rect -459 -2417 -455 -2400
rect -435 -2410 -431 -2356
rect -417 -2388 -413 -2356
rect -417 -2396 -413 -2392
rect -435 -2417 -431 -2414
rect -559 -2421 -550 -2417
rect -543 -2421 -535 -2417
rect -559 -2424 -555 -2421
rect -535 -2424 -531 -2421
rect -527 -2421 -515 -2417
rect -501 -2421 -493 -2417
rect -527 -2424 -523 -2421
rect -493 -2424 -489 -2421
rect -485 -2421 -473 -2417
rect -459 -2421 -447 -2417
rect -485 -2424 -481 -2421
rect -451 -2424 -447 -2421
rect -443 -2421 -431 -2417
rect -417 -2417 -413 -2400
rect -393 -2403 -389 -2356
rect -393 -2417 -389 -2407
rect -417 -2421 -405 -2417
rect -443 -2424 -439 -2421
rect -409 -2424 -405 -2421
rect -401 -2421 -389 -2417
rect -401 -2424 -397 -2421
rect -568 -2432 -564 -2428
rect -551 -2432 -547 -2428
rect -510 -2432 -506 -2428
rect -468 -2432 -464 -2428
rect -426 -2432 -422 -2428
rect -385 -2432 -381 -2428
rect -366 -2440 -362 -2392
rect -249 -2396 -245 -2135
rect -568 -2519 -564 -2515
rect -551 -2519 -547 -2515
rect -531 -2519 -527 -2515
rect -510 -2519 -506 -2515
rect -489 -2519 -485 -2515
rect -468 -2519 -464 -2515
rect -447 -2519 -443 -2515
rect -426 -2519 -422 -2515
rect -405 -2519 -401 -2515
rect -385 -2519 -381 -2515
rect -577 -2574 -573 -2527
rect -577 -2595 -573 -2578
rect -559 -2588 -555 -2527
rect -543 -2588 -539 -2527
rect -519 -2567 -515 -2527
rect -519 -2588 -515 -2571
rect -501 -2588 -497 -2527
rect -477 -2574 -473 -2527
rect -477 -2588 -473 -2578
rect -459 -2567 -455 -2527
rect -459 -2588 -455 -2571
rect -435 -2581 -431 -2527
rect -417 -2559 -413 -2527
rect -417 -2567 -413 -2563
rect -435 -2588 -431 -2585
rect -559 -2592 -550 -2588
rect -543 -2592 -535 -2588
rect -559 -2595 -555 -2592
rect -535 -2595 -531 -2592
rect -527 -2592 -515 -2588
rect -501 -2592 -493 -2588
rect -527 -2595 -523 -2592
rect -493 -2595 -489 -2592
rect -485 -2592 -473 -2588
rect -459 -2592 -447 -2588
rect -485 -2595 -481 -2592
rect -451 -2595 -447 -2592
rect -443 -2592 -431 -2588
rect -417 -2588 -413 -2571
rect -393 -2574 -389 -2527
rect -393 -2588 -389 -2578
rect -417 -2592 -405 -2588
rect -443 -2595 -439 -2592
rect -409 -2595 -405 -2592
rect -401 -2592 -389 -2588
rect -401 -2595 -397 -2592
rect -568 -2603 -564 -2599
rect -551 -2603 -547 -2599
rect -510 -2603 -506 -2599
rect -468 -2603 -464 -2599
rect -426 -2603 -422 -2599
rect -385 -2603 -381 -2599
rect -577 -2624 -573 -2620
rect -560 -2624 -556 -2620
rect -569 -2635 -565 -2632
rect -569 -2639 -554 -2635
rect -591 -2652 -576 -2648
rect -926 -2902 -922 -2898
rect -909 -2902 -905 -2898
rect -889 -2902 -885 -2898
rect -868 -2902 -864 -2898
rect -847 -2902 -843 -2898
rect -826 -2902 -822 -2898
rect -805 -2902 -801 -2898
rect -784 -2902 -780 -2898
rect -763 -2902 -759 -2898
rect -743 -2902 -739 -2898
rect -935 -2957 -931 -2910
rect -935 -2978 -931 -2961
rect -917 -2971 -913 -2910
rect -901 -2971 -897 -2910
rect -877 -2950 -873 -2910
rect -877 -2971 -873 -2954
rect -859 -2971 -855 -2910
rect -835 -2957 -831 -2910
rect -835 -2971 -831 -2961
rect -817 -2950 -813 -2910
rect -817 -2971 -813 -2954
rect -793 -2964 -789 -2910
rect -775 -2942 -771 -2910
rect -775 -2950 -771 -2946
rect -793 -2971 -789 -2968
rect -917 -2975 -908 -2971
rect -901 -2975 -893 -2971
rect -917 -2978 -913 -2975
rect -893 -2978 -889 -2975
rect -885 -2975 -873 -2971
rect -859 -2975 -851 -2971
rect -885 -2978 -881 -2975
rect -851 -2978 -847 -2975
rect -843 -2975 -831 -2971
rect -817 -2975 -805 -2971
rect -843 -2978 -839 -2975
rect -809 -2978 -805 -2975
rect -801 -2975 -789 -2971
rect -775 -2971 -771 -2954
rect -751 -2957 -747 -2910
rect -751 -2971 -747 -2961
rect -775 -2975 -763 -2971
rect -801 -2978 -797 -2975
rect -767 -2978 -763 -2975
rect -759 -2975 -747 -2971
rect -759 -2978 -755 -2975
rect -926 -2986 -922 -2982
rect -909 -2986 -905 -2982
rect -868 -2986 -864 -2982
rect -826 -2986 -822 -2982
rect -784 -2986 -780 -2982
rect -743 -2986 -739 -2982
rect -926 -3073 -922 -3069
rect -909 -3073 -905 -3069
rect -889 -3073 -885 -3069
rect -868 -3073 -864 -3069
rect -847 -3073 -843 -3069
rect -826 -3073 -822 -3069
rect -805 -3073 -801 -3069
rect -784 -3073 -780 -3069
rect -763 -3073 -759 -3069
rect -743 -3073 -739 -3069
rect -935 -3128 -931 -3081
rect -935 -3149 -931 -3132
rect -917 -3142 -913 -3081
rect -901 -3142 -897 -3081
rect -877 -3121 -873 -3081
rect -877 -3142 -873 -3125
rect -859 -3142 -855 -3081
rect -835 -3128 -831 -3081
rect -835 -3142 -831 -3132
rect -817 -3121 -813 -3081
rect -817 -3142 -813 -3125
rect -793 -3135 -789 -3081
rect -775 -3113 -771 -3081
rect -775 -3121 -771 -3117
rect -793 -3142 -789 -3139
rect -917 -3146 -908 -3142
rect -901 -3146 -893 -3142
rect -917 -3149 -913 -3146
rect -893 -3149 -889 -3146
rect -885 -3146 -873 -3142
rect -859 -3146 -851 -3142
rect -885 -3149 -881 -3146
rect -851 -3149 -847 -3146
rect -843 -3146 -831 -3142
rect -817 -3146 -805 -3142
rect -843 -3149 -839 -3146
rect -809 -3149 -805 -3146
rect -801 -3146 -789 -3142
rect -775 -3142 -771 -3125
rect -751 -3128 -747 -3081
rect -751 -3142 -747 -3132
rect -775 -3146 -763 -3142
rect -801 -3149 -797 -3146
rect -767 -3149 -763 -3146
rect -759 -3146 -747 -3142
rect -759 -3149 -755 -3146
rect -926 -3157 -922 -3153
rect -909 -3157 -905 -3153
rect -868 -3157 -864 -3153
rect -826 -3157 -822 -3153
rect -784 -3157 -780 -3153
rect -743 -3157 -739 -3153
rect -725 -3165 -721 -3117
rect -603 -3121 -599 -2878
rect -926 -3244 -922 -3240
rect -909 -3244 -905 -3240
rect -889 -3244 -885 -3240
rect -868 -3244 -864 -3240
rect -847 -3244 -843 -3240
rect -826 -3244 -822 -3240
rect -805 -3244 -801 -3240
rect -784 -3244 -780 -3240
rect -763 -3244 -759 -3240
rect -743 -3244 -739 -3240
rect -935 -3299 -931 -3252
rect -935 -3320 -931 -3303
rect -917 -3313 -913 -3252
rect -901 -3313 -897 -3252
rect -877 -3292 -873 -3252
rect -877 -3313 -873 -3296
rect -859 -3313 -855 -3252
rect -835 -3299 -831 -3252
rect -835 -3313 -831 -3303
rect -817 -3292 -813 -3252
rect -817 -3313 -813 -3296
rect -793 -3306 -789 -3252
rect -775 -3284 -771 -3252
rect -775 -3292 -771 -3288
rect -793 -3313 -789 -3310
rect -917 -3317 -908 -3313
rect -901 -3317 -893 -3313
rect -917 -3320 -913 -3317
rect -893 -3320 -889 -3317
rect -885 -3317 -873 -3313
rect -859 -3317 -851 -3313
rect -885 -3320 -881 -3317
rect -851 -3320 -847 -3317
rect -843 -3317 -831 -3313
rect -817 -3317 -805 -3313
rect -843 -3320 -839 -3317
rect -809 -3320 -805 -3317
rect -801 -3317 -789 -3313
rect -775 -3313 -771 -3296
rect -751 -3299 -747 -3252
rect -751 -3313 -747 -3303
rect -775 -3317 -763 -3313
rect -801 -3320 -797 -3317
rect -767 -3320 -763 -3317
rect -759 -3317 -747 -3313
rect -759 -3320 -755 -3317
rect -926 -3328 -922 -3324
rect -909 -3328 -905 -3324
rect -868 -3328 -864 -3324
rect -826 -3328 -822 -3324
rect -784 -3328 -780 -3324
rect -743 -3328 -739 -3324
rect -935 -3355 -931 -3351
rect -918 -3355 -914 -3351
rect -927 -3366 -923 -3363
rect -927 -3370 -912 -3366
rect -949 -3383 -934 -3379
rect -1225 -3598 -1221 -3594
rect -1181 -3598 -1177 -3594
rect -1147 -3598 -1143 -3594
rect -1257 -3863 -1253 -3609
rect -1113 -3612 -1109 -3580
rect -1246 -3692 -1242 -3616
rect -1225 -3644 -1221 -3640
rect -1208 -3644 -1204 -3640
rect -1188 -3644 -1184 -3640
rect -1167 -3644 -1163 -3640
rect -1146 -3644 -1142 -3640
rect -1125 -3644 -1121 -3640
rect -1104 -3644 -1100 -3640
rect -1083 -3644 -1079 -3640
rect -1062 -3644 -1058 -3640
rect -1042 -3644 -1038 -3640
rect -1234 -3699 -1230 -3652
rect -1234 -3720 -1230 -3703
rect -1216 -3713 -1212 -3652
rect -1200 -3713 -1196 -3652
rect -1176 -3692 -1172 -3652
rect -1176 -3713 -1172 -3696
rect -1158 -3713 -1154 -3652
rect -1134 -3699 -1130 -3652
rect -1134 -3713 -1130 -3703
rect -1116 -3692 -1112 -3652
rect -1116 -3713 -1112 -3696
rect -1092 -3706 -1088 -3652
rect -1074 -3684 -1070 -3652
rect -1074 -3692 -1070 -3688
rect -1092 -3713 -1088 -3710
rect -1216 -3717 -1207 -3713
rect -1200 -3717 -1192 -3713
rect -1216 -3720 -1212 -3717
rect -1192 -3720 -1188 -3717
rect -1184 -3717 -1172 -3713
rect -1158 -3717 -1150 -3713
rect -1184 -3720 -1180 -3717
rect -1150 -3720 -1146 -3717
rect -1142 -3717 -1130 -3713
rect -1116 -3717 -1104 -3713
rect -1142 -3720 -1138 -3717
rect -1108 -3720 -1104 -3717
rect -1100 -3717 -1088 -3713
rect -1074 -3713 -1070 -3696
rect -1050 -3699 -1046 -3652
rect -1050 -3713 -1046 -3703
rect -1074 -3717 -1062 -3713
rect -1100 -3720 -1096 -3717
rect -1066 -3720 -1062 -3717
rect -1058 -3717 -1046 -3713
rect -1058 -3720 -1054 -3717
rect -1225 -3728 -1221 -3724
rect -1208 -3728 -1204 -3724
rect -1167 -3728 -1163 -3724
rect -1125 -3728 -1121 -3724
rect -1083 -3728 -1079 -3724
rect -1042 -3728 -1038 -3724
rect -1225 -3815 -1221 -3811
rect -1208 -3815 -1204 -3811
rect -1188 -3815 -1184 -3811
rect -1167 -3815 -1163 -3811
rect -1146 -3815 -1142 -3811
rect -1125 -3815 -1121 -3811
rect -1104 -3815 -1100 -3811
rect -1083 -3815 -1079 -3811
rect -1062 -3815 -1058 -3811
rect -1042 -3815 -1038 -3811
rect -1234 -3870 -1230 -3823
rect -1234 -3891 -1230 -3874
rect -1216 -3884 -1212 -3823
rect -1200 -3884 -1196 -3823
rect -1176 -3863 -1172 -3823
rect -1176 -3884 -1172 -3867
rect -1158 -3884 -1154 -3823
rect -1134 -3870 -1130 -3823
rect -1134 -3884 -1130 -3874
rect -1116 -3863 -1112 -3823
rect -1116 -3884 -1112 -3867
rect -1092 -3877 -1088 -3823
rect -1074 -3855 -1070 -3823
rect -1074 -3863 -1070 -3859
rect -1092 -3884 -1088 -3881
rect -1216 -3888 -1207 -3884
rect -1200 -3888 -1192 -3884
rect -1216 -3891 -1212 -3888
rect -1192 -3891 -1188 -3888
rect -1184 -3888 -1172 -3884
rect -1158 -3888 -1150 -3884
rect -1184 -3891 -1180 -3888
rect -1150 -3891 -1146 -3888
rect -1142 -3888 -1130 -3884
rect -1116 -3888 -1104 -3884
rect -1142 -3891 -1138 -3888
rect -1108 -3891 -1104 -3888
rect -1100 -3888 -1088 -3884
rect -1074 -3884 -1070 -3867
rect -1050 -3870 -1046 -3823
rect -1050 -3884 -1046 -3874
rect -1074 -3888 -1062 -3884
rect -1100 -3891 -1096 -3888
rect -1066 -3891 -1062 -3888
rect -1058 -3888 -1046 -3884
rect -1058 -3891 -1054 -3888
rect -1225 -3899 -1221 -3895
rect -1208 -3899 -1204 -3895
rect -1167 -3899 -1163 -3895
rect -1125 -3899 -1121 -3895
rect -1083 -3899 -1079 -3895
rect -1042 -3899 -1038 -3895
rect -1028 -3906 -1024 -3859
rect -963 -3863 -959 -3616
rect -1309 -4105 -1305 -4101
rect -1292 -4105 -1288 -4101
rect -1301 -4116 -1297 -4113
rect -1301 -4120 -1286 -4116
rect -1319 -4133 -1308 -4129
rect -1805 -4387 -1801 -4383
rect -1788 -4387 -1784 -4383
rect -1768 -4387 -1764 -4383
rect -1747 -4387 -1743 -4383
rect -1726 -4387 -1722 -4383
rect -1705 -4387 -1701 -4383
rect -1684 -4387 -1680 -4383
rect -1663 -4387 -1659 -4383
rect -1642 -4387 -1638 -4383
rect -1622 -4387 -1618 -4383
rect -1542 -4387 -1538 -4383
rect -1525 -4387 -1521 -4383
rect -1505 -4387 -1501 -4383
rect -1484 -4387 -1480 -4383
rect -1463 -4387 -1459 -4383
rect -1442 -4387 -1438 -4383
rect -1421 -4387 -1417 -4383
rect -1400 -4387 -1396 -4383
rect -1379 -4387 -1375 -4383
rect -1359 -4387 -1355 -4383
rect -1814 -4442 -1810 -4395
rect -1814 -4463 -1810 -4446
rect -1796 -4456 -1792 -4395
rect -1780 -4456 -1776 -4395
rect -1756 -4435 -1752 -4395
rect -1756 -4456 -1752 -4439
rect -1738 -4456 -1734 -4395
rect -1714 -4442 -1710 -4395
rect -1714 -4456 -1710 -4446
rect -1696 -4435 -1692 -4395
rect -1696 -4456 -1692 -4439
rect -1672 -4449 -1668 -4395
rect -1654 -4427 -1650 -4395
rect -1654 -4435 -1650 -4431
rect -1672 -4456 -1668 -4453
rect -1796 -4460 -1787 -4456
rect -1780 -4460 -1772 -4456
rect -1796 -4463 -1792 -4460
rect -1772 -4463 -1768 -4460
rect -1764 -4460 -1752 -4456
rect -1738 -4460 -1730 -4456
rect -1764 -4463 -1760 -4460
rect -1730 -4463 -1726 -4460
rect -1722 -4460 -1710 -4456
rect -1696 -4460 -1684 -4456
rect -1722 -4463 -1718 -4460
rect -1688 -4463 -1684 -4460
rect -1680 -4460 -1668 -4456
rect -1654 -4456 -1650 -4439
rect -1630 -4442 -1626 -4395
rect -1630 -4456 -1626 -4446
rect -1654 -4460 -1642 -4456
rect -1680 -4463 -1676 -4460
rect -1646 -4463 -1642 -4460
rect -1638 -4460 -1626 -4456
rect -1551 -4442 -1547 -4395
rect -1638 -4463 -1634 -4460
rect -1551 -4463 -1547 -4446
rect -1533 -4456 -1529 -4395
rect -1517 -4456 -1513 -4395
rect -1493 -4435 -1489 -4395
rect -1493 -4456 -1489 -4439
rect -1475 -4456 -1471 -4395
rect -1451 -4442 -1447 -4395
rect -1451 -4456 -1447 -4446
rect -1433 -4435 -1429 -4395
rect -1433 -4456 -1429 -4439
rect -1409 -4449 -1405 -4395
rect -1391 -4427 -1387 -4395
rect -1391 -4435 -1387 -4431
rect -1409 -4456 -1405 -4453
rect -1533 -4460 -1524 -4456
rect -1517 -4460 -1509 -4456
rect -1533 -4463 -1529 -4460
rect -1509 -4463 -1505 -4460
rect -1501 -4460 -1489 -4456
rect -1475 -4460 -1467 -4456
rect -1501 -4463 -1497 -4460
rect -1467 -4463 -1463 -4460
rect -1459 -4460 -1447 -4456
rect -1433 -4460 -1421 -4456
rect -1459 -4463 -1455 -4460
rect -1425 -4463 -1421 -4460
rect -1417 -4460 -1405 -4456
rect -1391 -4456 -1387 -4439
rect -1367 -4442 -1363 -4395
rect -1367 -4456 -1363 -4446
rect -1391 -4460 -1379 -4456
rect -1417 -4463 -1413 -4460
rect -1383 -4463 -1379 -4460
rect -1375 -4460 -1363 -4456
rect -1375 -4463 -1371 -4460
rect -1805 -4471 -1801 -4467
rect -1788 -4471 -1784 -4467
rect -1747 -4471 -1743 -4467
rect -1705 -4471 -1701 -4467
rect -1663 -4471 -1659 -4467
rect -1622 -4471 -1618 -4467
rect -1542 -4471 -1538 -4467
rect -1525 -4471 -1521 -4467
rect -1484 -4471 -1480 -4467
rect -1442 -4471 -1438 -4467
rect -1400 -4471 -1396 -4467
rect -1359 -4471 -1355 -4467
rect -1346 -4478 -1342 -4431
rect -1831 -4606 -1827 -4482
rect -1805 -4558 -1801 -4554
rect -1788 -4558 -1784 -4554
rect -1768 -4558 -1764 -4554
rect -1747 -4558 -1743 -4554
rect -1726 -4558 -1722 -4554
rect -1705 -4558 -1701 -4554
rect -1684 -4558 -1680 -4554
rect -1663 -4558 -1659 -4554
rect -1642 -4558 -1638 -4554
rect -1622 -4558 -1618 -4554
rect -1542 -4558 -1538 -4554
rect -1525 -4558 -1521 -4554
rect -1505 -4558 -1501 -4554
rect -1484 -4558 -1480 -4554
rect -1463 -4558 -1459 -4554
rect -1442 -4558 -1438 -4554
rect -1421 -4558 -1417 -4554
rect -1400 -4558 -1396 -4554
rect -1379 -4558 -1375 -4554
rect -1359 -4558 -1355 -4554
rect -1814 -4613 -1810 -4566
rect -1814 -4634 -1810 -4617
rect -1796 -4627 -1792 -4566
rect -1780 -4627 -1776 -4566
rect -1756 -4606 -1752 -4566
rect -1756 -4627 -1752 -4610
rect -1738 -4627 -1734 -4566
rect -1714 -4613 -1710 -4566
rect -1714 -4627 -1710 -4617
rect -1696 -4606 -1692 -4566
rect -1696 -4627 -1692 -4610
rect -1672 -4620 -1668 -4566
rect -1654 -4598 -1650 -4566
rect -1654 -4606 -1650 -4602
rect -1672 -4627 -1668 -4624
rect -1796 -4631 -1787 -4627
rect -1780 -4631 -1772 -4627
rect -1796 -4634 -1792 -4631
rect -1772 -4634 -1768 -4631
rect -1764 -4631 -1752 -4627
rect -1738 -4631 -1730 -4627
rect -1764 -4634 -1760 -4631
rect -1730 -4634 -1726 -4631
rect -1722 -4631 -1710 -4627
rect -1696 -4631 -1684 -4627
rect -1722 -4634 -1718 -4631
rect -1688 -4634 -1684 -4631
rect -1680 -4631 -1668 -4627
rect -1654 -4627 -1650 -4610
rect -1630 -4613 -1626 -4566
rect -1630 -4627 -1626 -4617
rect -1654 -4631 -1642 -4627
rect -1680 -4634 -1676 -4631
rect -1646 -4634 -1642 -4631
rect -1638 -4631 -1626 -4627
rect -1551 -4613 -1547 -4566
rect -1638 -4634 -1634 -4631
rect -1551 -4634 -1547 -4617
rect -1533 -4627 -1529 -4566
rect -1517 -4627 -1513 -4566
rect -1493 -4606 -1489 -4566
rect -1493 -4627 -1489 -4610
rect -1475 -4627 -1471 -4566
rect -1451 -4613 -1447 -4566
rect -1451 -4627 -1447 -4617
rect -1433 -4606 -1429 -4566
rect -1433 -4627 -1429 -4610
rect -1409 -4620 -1405 -4566
rect -1391 -4598 -1387 -4566
rect -1391 -4606 -1387 -4602
rect -1409 -4627 -1405 -4624
rect -1533 -4631 -1524 -4627
rect -1517 -4631 -1509 -4627
rect -1533 -4634 -1529 -4631
rect -1509 -4634 -1505 -4631
rect -1501 -4631 -1489 -4627
rect -1475 -4631 -1467 -4627
rect -1501 -4634 -1497 -4631
rect -1467 -4634 -1463 -4631
rect -1459 -4631 -1447 -4627
rect -1433 -4631 -1421 -4627
rect -1459 -4634 -1455 -4631
rect -1425 -4634 -1421 -4631
rect -1417 -4631 -1405 -4627
rect -1391 -4627 -1387 -4610
rect -1367 -4613 -1363 -4566
rect -1367 -4627 -1363 -4617
rect -1391 -4631 -1379 -4627
rect -1417 -4634 -1413 -4631
rect -1383 -4634 -1379 -4631
rect -1375 -4631 -1363 -4627
rect -1375 -4634 -1371 -4631
rect -1805 -4642 -1801 -4638
rect -1788 -4642 -1784 -4638
rect -1747 -4642 -1743 -4638
rect -1705 -4642 -1701 -4638
rect -1663 -4642 -1659 -4638
rect -1622 -4642 -1618 -4638
rect -1542 -4642 -1538 -4638
rect -1525 -4642 -1521 -4638
rect -1484 -4642 -1480 -4638
rect -1442 -4642 -1438 -4638
rect -1400 -4642 -1396 -4638
rect -1359 -4642 -1355 -4638
rect -1347 -4650 -1343 -4602
rect -1566 -4777 -1562 -4654
rect -1542 -4729 -1538 -4725
rect -1525 -4729 -1521 -4725
rect -1505 -4729 -1501 -4725
rect -1484 -4729 -1480 -4725
rect -1463 -4729 -1459 -4725
rect -1442 -4729 -1438 -4725
rect -1421 -4729 -1417 -4725
rect -1400 -4729 -1396 -4725
rect -1379 -4729 -1375 -4725
rect -1359 -4729 -1355 -4725
rect -1551 -4784 -1547 -4737
rect -1551 -4805 -1547 -4788
rect -1533 -4798 -1529 -4737
rect -1517 -4798 -1513 -4737
rect -1493 -4777 -1489 -4737
rect -1493 -4798 -1489 -4781
rect -1475 -4798 -1471 -4737
rect -1451 -4784 -1447 -4737
rect -1451 -4798 -1447 -4788
rect -1433 -4777 -1429 -4737
rect -1433 -4798 -1429 -4781
rect -1409 -4791 -1405 -4737
rect -1391 -4769 -1387 -4737
rect -1391 -4777 -1387 -4773
rect -1409 -4798 -1405 -4795
rect -1533 -4802 -1524 -4798
rect -1517 -4802 -1509 -4798
rect -1533 -4805 -1529 -4802
rect -1509 -4805 -1505 -4802
rect -1501 -4802 -1489 -4798
rect -1475 -4802 -1467 -4798
rect -1501 -4805 -1497 -4802
rect -1467 -4805 -1463 -4802
rect -1459 -4802 -1447 -4798
rect -1433 -4802 -1421 -4798
rect -1459 -4805 -1455 -4802
rect -1425 -4805 -1421 -4802
rect -1417 -4802 -1405 -4798
rect -1391 -4798 -1387 -4781
rect -1367 -4784 -1363 -4737
rect -1367 -4798 -1363 -4788
rect -1391 -4802 -1379 -4798
rect -1417 -4805 -1413 -4802
rect -1383 -4805 -1379 -4802
rect -1375 -4802 -1363 -4798
rect -1375 -4805 -1371 -4802
rect -1542 -4813 -1538 -4809
rect -1525 -4813 -1521 -4809
rect -1484 -4813 -1480 -4809
rect -1442 -4813 -1438 -4809
rect -1400 -4813 -1396 -4809
rect -1359 -4813 -1355 -4809
rect -1346 -4876 -1342 -4773
rect -1319 -4777 -1315 -4133
rect -1290 -4159 -1286 -4120
rect -1290 -4174 -1286 -4163
rect -1309 -4178 -1286 -4174
rect -1309 -4181 -1305 -4178
rect -1283 -4181 -1279 -4113
rect -1292 -4189 -1288 -4185
rect -1283 -4319 -1279 -4185
rect -1257 -4312 -1253 -3910
rect -1225 -3990 -1221 -3986
rect -1208 -3990 -1204 -3986
rect -1188 -3990 -1184 -3986
rect -1167 -3990 -1163 -3986
rect -1146 -3990 -1142 -3986
rect -1125 -3990 -1121 -3986
rect -1104 -3990 -1100 -3986
rect -1083 -3990 -1079 -3986
rect -1062 -3990 -1058 -3986
rect -1042 -3990 -1038 -3986
rect -1234 -4045 -1230 -3998
rect -1234 -4066 -1230 -4049
rect -1216 -4059 -1212 -3998
rect -1200 -4059 -1196 -3998
rect -1176 -4038 -1172 -3998
rect -1176 -4059 -1172 -4042
rect -1158 -4059 -1154 -3998
rect -1134 -4045 -1130 -3998
rect -1134 -4059 -1130 -4049
rect -1116 -4038 -1112 -3998
rect -1116 -4059 -1112 -4042
rect -1092 -4052 -1088 -3998
rect -1074 -4030 -1070 -3998
rect -1074 -4038 -1070 -4034
rect -1092 -4059 -1088 -4056
rect -1216 -4063 -1207 -4059
rect -1200 -4063 -1192 -4059
rect -1216 -4066 -1212 -4063
rect -1192 -4066 -1188 -4063
rect -1184 -4063 -1172 -4059
rect -1158 -4063 -1150 -4059
rect -1184 -4066 -1180 -4063
rect -1150 -4066 -1146 -4063
rect -1142 -4063 -1130 -4059
rect -1116 -4063 -1104 -4059
rect -1142 -4066 -1138 -4063
rect -1108 -4066 -1104 -4063
rect -1100 -4063 -1088 -4059
rect -1074 -4059 -1070 -4042
rect -1050 -4045 -1046 -3998
rect -1050 -4059 -1046 -4049
rect -1074 -4063 -1062 -4059
rect -1100 -4066 -1096 -4063
rect -1066 -4066 -1062 -4063
rect -1058 -4063 -1046 -4059
rect -1058 -4066 -1054 -4063
rect -1225 -4074 -1221 -4070
rect -1208 -4074 -1204 -4070
rect -1167 -4074 -1163 -4070
rect -1125 -4074 -1121 -4070
rect -1083 -4074 -1079 -4070
rect -1042 -4074 -1038 -4070
rect -1024 -4129 -1020 -4034
rect -1225 -4264 -1221 -4260
rect -1208 -4264 -1204 -4260
rect -1168 -4264 -1164 -4260
rect -1147 -4264 -1143 -4260
rect -1234 -4305 -1230 -4272
rect -1234 -4340 -1230 -4309
rect -1216 -4299 -1212 -4272
rect -1216 -4303 -1207 -4299
rect -1216 -4340 -1212 -4303
rect -1190 -4326 -1186 -4272
rect -1190 -4333 -1186 -4330
rect -1156 -4333 -1152 -4272
rect -1138 -4304 -1134 -4272
rect -979 -4296 -975 -4154
rect -1208 -4340 -1204 -4337
rect -1199 -4337 -1186 -4333
rect -1199 -4340 -1195 -4337
rect -1172 -4340 -1168 -4337
rect -1164 -4337 -1145 -4333
rect -1164 -4340 -1160 -4337
rect -1138 -4340 -1134 -4308
rect -963 -4311 -959 -3911
rect -949 -4038 -945 -3383
rect -916 -3409 -912 -3370
rect -916 -3424 -912 -3413
rect -935 -3428 -912 -3424
rect -909 -3400 -905 -3363
rect -722 -3379 -718 -3288
rect -935 -3431 -931 -3428
rect -909 -3431 -905 -3404
rect -918 -3439 -914 -3435
rect -926 -3514 -922 -3510
rect -900 -3514 -896 -3510
rect -883 -3514 -879 -3510
rect -843 -3514 -839 -3510
rect -822 -3514 -818 -3510
rect -805 -3514 -801 -3510
rect -765 -3514 -761 -3510
rect -741 -3514 -737 -3510
rect -704 -3514 -700 -3510
rect -935 -3539 -931 -3522
rect -935 -3590 -931 -3543
rect -917 -3532 -913 -3522
rect -917 -3590 -913 -3536
rect -909 -3561 -905 -3522
rect -891 -3554 -887 -3522
rect -909 -3590 -905 -3565
rect -891 -3590 -887 -3558
rect -865 -3546 -861 -3522
rect -865 -3583 -861 -3550
rect -831 -3583 -827 -3522
rect -813 -3539 -809 -3522
rect -883 -3590 -879 -3587
rect -875 -3587 -861 -3583
rect -875 -3590 -871 -3587
rect -847 -3590 -843 -3587
rect -839 -3587 -820 -3583
rect -839 -3590 -835 -3587
rect -813 -3590 -809 -3543
rect -787 -3554 -783 -3522
rect -787 -3583 -783 -3558
rect -753 -3576 -749 -3522
rect -753 -3580 -736 -3576
rect -805 -3590 -801 -3587
rect -796 -3587 -783 -3583
rect -796 -3590 -792 -3587
rect -769 -3590 -765 -3587
rect -745 -3590 -741 -3580
rect -729 -3583 -725 -3522
rect -721 -3576 -717 -3522
rect -695 -3546 -691 -3522
rect -721 -3580 -702 -3576
rect -737 -3587 -720 -3583
rect -737 -3590 -733 -3587
rect -713 -3590 -709 -3580
rect -695 -3590 -691 -3550
rect -926 -3598 -922 -3594
rect -900 -3598 -896 -3594
rect -857 -3598 -853 -3594
rect -822 -3598 -818 -3594
rect -778 -3598 -774 -3594
rect -761 -3598 -757 -3594
rect -725 -3598 -721 -3594
rect -704 -3598 -700 -3594
rect -687 -3605 -683 -3558
rect -616 -3561 -612 -3404
rect -603 -3546 -599 -3168
rect -591 -3292 -587 -2652
rect -558 -2678 -554 -2639
rect -558 -2693 -554 -2682
rect -577 -2697 -554 -2693
rect -551 -2669 -547 -2632
rect -373 -2648 -369 -2563
rect -577 -2700 -573 -2697
rect -551 -2700 -547 -2673
rect -560 -2708 -556 -2704
rect -568 -2783 -564 -2779
rect -542 -2783 -538 -2779
rect -525 -2783 -521 -2779
rect -485 -2783 -481 -2779
rect -464 -2783 -460 -2779
rect -447 -2783 -443 -2779
rect -407 -2783 -403 -2779
rect -383 -2783 -379 -2779
rect -346 -2783 -342 -2779
rect -577 -2808 -573 -2791
rect -577 -2859 -573 -2812
rect -559 -2801 -555 -2791
rect -559 -2859 -555 -2805
rect -551 -2830 -547 -2791
rect -533 -2823 -529 -2791
rect -551 -2859 -547 -2834
rect -533 -2859 -529 -2827
rect -507 -2815 -503 -2791
rect -507 -2852 -503 -2819
rect -473 -2852 -469 -2791
rect -455 -2808 -451 -2791
rect -525 -2859 -521 -2856
rect -517 -2856 -503 -2852
rect -517 -2859 -513 -2856
rect -489 -2859 -485 -2856
rect -481 -2856 -462 -2852
rect -481 -2859 -477 -2856
rect -455 -2859 -451 -2812
rect -429 -2823 -425 -2791
rect -429 -2852 -425 -2827
rect -395 -2845 -391 -2791
rect -395 -2849 -378 -2845
rect -447 -2859 -443 -2856
rect -438 -2856 -425 -2852
rect -438 -2859 -434 -2856
rect -411 -2859 -407 -2856
rect -387 -2859 -383 -2849
rect -371 -2852 -367 -2791
rect -363 -2845 -359 -2791
rect -337 -2814 -333 -2791
rect -363 -2849 -344 -2845
rect -379 -2856 -362 -2852
rect -379 -2859 -375 -2856
rect -355 -2859 -351 -2849
rect -337 -2859 -333 -2818
rect -568 -2867 -564 -2863
rect -542 -2867 -538 -2863
rect -499 -2867 -495 -2863
rect -464 -2867 -460 -2863
rect -420 -2867 -416 -2863
rect -403 -2867 -399 -2863
rect -367 -2867 -363 -2863
rect -346 -2867 -342 -2863
rect -329 -2881 -325 -2827
rect -263 -2830 -259 -2673
rect -249 -2815 -245 -2444
rect -233 -2567 -229 -1902
rect -200 -1928 -196 -1889
rect -200 -1943 -196 -1932
rect -219 -1947 -196 -1943
rect -193 -1919 -189 -1882
rect -9 -1898 -5 -1811
rect -219 -1950 -215 -1947
rect -193 -1950 -189 -1923
rect -202 -1958 -198 -1954
rect -210 -2033 -206 -2029
rect -184 -2033 -180 -2029
rect -167 -2033 -163 -2029
rect -127 -2033 -123 -2029
rect -106 -2033 -102 -2029
rect -89 -2033 -85 -2029
rect -49 -2033 -45 -2029
rect -25 -2033 -21 -2029
rect 12 -2033 16 -2029
rect -219 -2058 -215 -2041
rect -219 -2109 -215 -2062
rect -201 -2051 -197 -2041
rect -201 -2109 -197 -2055
rect -193 -2080 -189 -2041
rect -175 -2073 -171 -2041
rect -193 -2109 -189 -2084
rect -175 -2109 -171 -2077
rect -149 -2065 -145 -2041
rect -149 -2102 -145 -2069
rect -115 -2102 -111 -2041
rect -97 -2058 -93 -2041
rect -167 -2109 -163 -2106
rect -159 -2106 -145 -2102
rect -159 -2109 -155 -2106
rect -131 -2109 -127 -2106
rect -123 -2106 -104 -2102
rect -123 -2109 -119 -2106
rect -97 -2109 -93 -2062
rect -71 -2073 -67 -2041
rect -71 -2102 -67 -2077
rect -37 -2095 -33 -2041
rect -37 -2099 -20 -2095
rect -89 -2109 -85 -2106
rect -80 -2106 -67 -2102
rect -80 -2109 -76 -2106
rect -53 -2109 -49 -2106
rect -29 -2109 -25 -2099
rect -13 -2102 -9 -2041
rect -5 -2095 -1 -2041
rect 21 -2065 25 -2041
rect -5 -2099 14 -2095
rect -21 -2106 -4 -2102
rect -21 -2109 -17 -2106
rect 3 -2109 7 -2099
rect 21 -2109 25 -2069
rect -210 -2117 -206 -2113
rect -184 -2117 -180 -2113
rect -141 -2117 -137 -2113
rect -106 -2117 -102 -2113
rect -62 -2117 -58 -2113
rect -45 -2117 -41 -2113
rect -9 -2117 -5 -2113
rect 12 -2117 16 -2113
rect 29 -2124 33 -2077
rect 93 -2080 97 -1923
rect 107 -2065 111 -1692
rect 125 -1815 129 -1166
rect 158 -1192 162 -1153
rect 158 -1207 162 -1196
rect 139 -1211 162 -1207
rect 165 -1183 169 -1146
rect 139 -1214 143 -1211
rect 165 -1214 169 -1187
rect 156 -1222 160 -1218
rect 148 -1302 152 -1298
rect 174 -1302 178 -1298
rect 191 -1302 195 -1298
rect 231 -1302 235 -1298
rect 252 -1302 256 -1298
rect 269 -1302 273 -1298
rect 309 -1302 313 -1298
rect 333 -1302 337 -1298
rect 370 -1302 374 -1298
rect 139 -1327 143 -1310
rect 139 -1378 143 -1331
rect 157 -1320 161 -1310
rect 157 -1378 161 -1324
rect 165 -1349 169 -1310
rect 183 -1342 187 -1310
rect 165 -1378 169 -1353
rect 183 -1378 187 -1346
rect 209 -1334 213 -1310
rect 209 -1371 213 -1338
rect 243 -1371 247 -1310
rect 261 -1327 265 -1310
rect 191 -1378 195 -1375
rect 199 -1375 213 -1371
rect 199 -1378 203 -1375
rect 227 -1378 231 -1375
rect 235 -1375 254 -1371
rect 235 -1378 239 -1375
rect 261 -1378 265 -1331
rect 287 -1342 291 -1310
rect 287 -1371 291 -1346
rect 321 -1364 325 -1310
rect 321 -1368 338 -1364
rect 269 -1378 273 -1375
rect 278 -1375 291 -1371
rect 278 -1378 282 -1375
rect 305 -1378 309 -1375
rect 329 -1378 333 -1368
rect 345 -1371 349 -1310
rect 353 -1364 357 -1310
rect 379 -1334 383 -1310
rect 353 -1368 372 -1364
rect 337 -1375 354 -1371
rect 337 -1378 341 -1375
rect 361 -1378 365 -1368
rect 379 -1378 383 -1338
rect 148 -1386 152 -1382
rect 174 -1386 178 -1382
rect 217 -1386 221 -1382
rect 252 -1386 256 -1382
rect 296 -1386 300 -1382
rect 313 -1386 317 -1382
rect 349 -1386 353 -1382
rect 370 -1386 374 -1382
rect 386 -1400 390 -1346
rect 447 -1349 451 -1187
rect 470 -1334 474 -832
rect 481 -1162 485 -816
rect 514 -857 518 -803
rect 495 -861 514 -857
rect 521 -836 525 -796
rect 839 -812 843 -748
rect 853 -788 857 -784
rect 870 -788 874 -784
rect 861 -799 865 -796
rect 861 -803 876 -799
rect 839 -816 854 -812
rect 495 -864 499 -861
rect 521 -864 525 -840
rect 512 -872 516 -868
rect 504 -1022 508 -1018
rect 521 -1022 525 -1018
rect 541 -1022 545 -1018
rect 562 -1022 566 -1018
rect 583 -1022 587 -1018
rect 604 -1022 608 -1018
rect 625 -1022 629 -1018
rect 646 -1022 650 -1018
rect 667 -1022 671 -1018
rect 687 -1022 691 -1018
rect 495 -1077 499 -1030
rect 495 -1098 499 -1081
rect 513 -1091 517 -1030
rect 529 -1091 533 -1030
rect 553 -1070 557 -1030
rect 553 -1091 557 -1074
rect 571 -1091 575 -1030
rect 595 -1077 599 -1030
rect 595 -1091 599 -1081
rect 613 -1070 617 -1030
rect 613 -1091 617 -1074
rect 637 -1084 641 -1030
rect 655 -1062 659 -1030
rect 655 -1070 659 -1066
rect 637 -1091 641 -1088
rect 513 -1095 522 -1091
rect 529 -1095 537 -1091
rect 513 -1098 517 -1095
rect 537 -1098 541 -1095
rect 545 -1095 557 -1091
rect 571 -1095 579 -1091
rect 545 -1098 549 -1095
rect 579 -1098 583 -1095
rect 587 -1095 599 -1091
rect 613 -1095 625 -1091
rect 587 -1098 591 -1095
rect 621 -1098 625 -1095
rect 629 -1095 641 -1091
rect 655 -1091 659 -1074
rect 679 -1077 683 -1030
rect 679 -1091 683 -1081
rect 655 -1095 667 -1091
rect 629 -1098 633 -1095
rect 663 -1098 667 -1095
rect 671 -1095 683 -1091
rect 671 -1098 675 -1095
rect 504 -1106 508 -1102
rect 521 -1106 525 -1102
rect 562 -1106 566 -1102
rect 604 -1106 608 -1102
rect 646 -1106 650 -1102
rect 687 -1106 691 -1102
rect 495 -1138 499 -1134
rect 512 -1138 516 -1134
rect 503 -1149 507 -1146
rect 503 -1153 518 -1149
rect 481 -1166 496 -1162
rect 148 -1425 152 -1421
rect 165 -1425 169 -1421
rect 185 -1425 189 -1421
rect 206 -1425 210 -1421
rect 227 -1425 231 -1421
rect 248 -1425 252 -1421
rect 269 -1425 273 -1421
rect 290 -1425 294 -1421
rect 311 -1425 315 -1421
rect 331 -1425 335 -1421
rect 139 -1480 143 -1433
rect 139 -1501 143 -1484
rect 157 -1494 161 -1433
rect 173 -1494 177 -1433
rect 197 -1473 201 -1433
rect 197 -1494 201 -1477
rect 215 -1494 219 -1433
rect 239 -1480 243 -1433
rect 239 -1494 243 -1484
rect 257 -1473 261 -1433
rect 257 -1494 261 -1477
rect 281 -1487 285 -1433
rect 299 -1465 303 -1433
rect 299 -1473 303 -1469
rect 281 -1494 285 -1491
rect 157 -1498 166 -1494
rect 173 -1498 181 -1494
rect 157 -1501 161 -1498
rect 181 -1501 185 -1498
rect 189 -1498 201 -1494
rect 215 -1498 223 -1494
rect 189 -1501 193 -1498
rect 223 -1501 227 -1498
rect 231 -1498 243 -1494
rect 257 -1498 269 -1494
rect 231 -1501 235 -1498
rect 265 -1501 269 -1498
rect 273 -1498 285 -1494
rect 299 -1494 303 -1477
rect 323 -1480 327 -1433
rect 323 -1494 327 -1484
rect 299 -1498 311 -1494
rect 273 -1501 277 -1498
rect 307 -1501 311 -1498
rect 315 -1498 327 -1494
rect 315 -1501 319 -1498
rect 148 -1509 152 -1505
rect 165 -1509 169 -1505
rect 206 -1509 210 -1505
rect 248 -1509 252 -1505
rect 290 -1509 294 -1505
rect 331 -1509 335 -1505
rect 148 -1596 152 -1592
rect 165 -1596 169 -1592
rect 185 -1596 189 -1592
rect 206 -1596 210 -1592
rect 227 -1596 231 -1592
rect 248 -1596 252 -1592
rect 269 -1596 273 -1592
rect 290 -1596 294 -1592
rect 311 -1596 315 -1592
rect 331 -1596 335 -1592
rect 139 -1651 143 -1604
rect 139 -1672 143 -1655
rect 157 -1665 161 -1604
rect 173 -1665 177 -1604
rect 197 -1644 201 -1604
rect 197 -1665 201 -1648
rect 215 -1665 219 -1604
rect 239 -1651 243 -1604
rect 239 -1665 243 -1655
rect 257 -1644 261 -1604
rect 257 -1665 261 -1648
rect 281 -1658 285 -1604
rect 299 -1636 303 -1604
rect 299 -1644 303 -1640
rect 281 -1665 285 -1662
rect 157 -1669 166 -1665
rect 173 -1669 181 -1665
rect 157 -1672 161 -1669
rect 181 -1672 185 -1669
rect 189 -1669 201 -1665
rect 215 -1669 223 -1665
rect 189 -1672 193 -1669
rect 223 -1672 227 -1669
rect 231 -1669 243 -1665
rect 257 -1669 269 -1665
rect 231 -1672 235 -1669
rect 265 -1672 269 -1669
rect 273 -1669 285 -1665
rect 299 -1665 303 -1648
rect 323 -1651 327 -1604
rect 323 -1665 327 -1655
rect 299 -1669 311 -1665
rect 273 -1672 277 -1669
rect 307 -1672 311 -1669
rect 315 -1669 327 -1665
rect 315 -1672 319 -1669
rect 148 -1680 152 -1676
rect 165 -1680 169 -1676
rect 206 -1680 210 -1676
rect 248 -1680 252 -1676
rect 290 -1680 294 -1676
rect 331 -1680 335 -1676
rect 346 -1688 350 -1640
rect 470 -1644 474 -1404
rect 148 -1767 152 -1763
rect 165 -1767 169 -1763
rect 185 -1767 189 -1763
rect 206 -1767 210 -1763
rect 227 -1767 231 -1763
rect 248 -1767 252 -1763
rect 269 -1767 273 -1763
rect 290 -1767 294 -1763
rect 311 -1767 315 -1763
rect 331 -1767 335 -1763
rect 139 -1822 143 -1775
rect 139 -1843 143 -1826
rect 157 -1836 161 -1775
rect 173 -1836 177 -1775
rect 197 -1815 201 -1775
rect 197 -1836 201 -1819
rect 215 -1836 219 -1775
rect 239 -1822 243 -1775
rect 239 -1836 243 -1826
rect 257 -1815 261 -1775
rect 257 -1836 261 -1819
rect 281 -1829 285 -1775
rect 299 -1807 303 -1775
rect 299 -1815 303 -1811
rect 281 -1836 285 -1833
rect 157 -1840 166 -1836
rect 173 -1840 181 -1836
rect 157 -1843 161 -1840
rect 181 -1843 185 -1840
rect 189 -1840 201 -1836
rect 215 -1840 223 -1836
rect 189 -1843 193 -1840
rect 223 -1843 227 -1840
rect 231 -1840 243 -1836
rect 257 -1840 269 -1836
rect 231 -1843 235 -1840
rect 265 -1843 269 -1840
rect 273 -1840 285 -1836
rect 299 -1836 303 -1819
rect 323 -1822 327 -1775
rect 323 -1836 327 -1826
rect 299 -1840 311 -1836
rect 273 -1843 277 -1840
rect 307 -1843 311 -1840
rect 315 -1840 327 -1836
rect 315 -1843 319 -1840
rect 148 -1851 152 -1847
rect 165 -1851 169 -1847
rect 206 -1851 210 -1847
rect 248 -1851 252 -1847
rect 290 -1851 294 -1847
rect 331 -1851 335 -1847
rect 139 -1874 143 -1870
rect 156 -1874 160 -1870
rect 147 -1885 151 -1882
rect 147 -1889 162 -1885
rect 125 -1902 140 -1898
rect -210 -2177 -206 -2173
rect -193 -2177 -189 -2173
rect -173 -2177 -169 -2173
rect -152 -2177 -148 -2173
rect -131 -2177 -127 -2173
rect -110 -2177 -106 -2173
rect -89 -2177 -85 -2173
rect -68 -2177 -64 -2173
rect -47 -2177 -43 -2173
rect -27 -2177 -23 -2173
rect -219 -2232 -215 -2185
rect -219 -2253 -215 -2236
rect -201 -2246 -197 -2185
rect -185 -2246 -181 -2185
rect -161 -2225 -157 -2185
rect -161 -2246 -157 -2229
rect -143 -2246 -139 -2185
rect -119 -2232 -115 -2185
rect -119 -2246 -115 -2236
rect -101 -2225 -97 -2185
rect -101 -2246 -97 -2229
rect -77 -2239 -73 -2185
rect -59 -2217 -55 -2185
rect -59 -2225 -55 -2221
rect -77 -2246 -73 -2243
rect -201 -2250 -192 -2246
rect -185 -2250 -177 -2246
rect -201 -2253 -197 -2250
rect -177 -2253 -173 -2250
rect -169 -2250 -157 -2246
rect -143 -2250 -135 -2246
rect -169 -2253 -165 -2250
rect -135 -2253 -131 -2250
rect -127 -2250 -115 -2246
rect -101 -2250 -89 -2246
rect -127 -2253 -123 -2250
rect -93 -2253 -89 -2250
rect -85 -2250 -73 -2246
rect -59 -2246 -55 -2229
rect -35 -2232 -31 -2185
rect -35 -2246 -31 -2236
rect -59 -2250 -47 -2246
rect -85 -2253 -81 -2250
rect -51 -2253 -47 -2250
rect -43 -2250 -31 -2246
rect -43 -2253 -39 -2250
rect -210 -2261 -206 -2257
rect -193 -2261 -189 -2257
rect -152 -2261 -148 -2257
rect -110 -2261 -106 -2257
rect -68 -2261 -64 -2257
rect -27 -2261 -23 -2257
rect -210 -2348 -206 -2344
rect -193 -2348 -189 -2344
rect -173 -2348 -169 -2344
rect -152 -2348 -148 -2344
rect -131 -2348 -127 -2344
rect -110 -2348 -106 -2344
rect -89 -2348 -85 -2344
rect -68 -2348 -64 -2344
rect -47 -2348 -43 -2344
rect -27 -2348 -23 -2344
rect -219 -2403 -215 -2356
rect -219 -2424 -215 -2407
rect -201 -2417 -197 -2356
rect -185 -2417 -181 -2356
rect -161 -2396 -157 -2356
rect -161 -2417 -157 -2400
rect -143 -2417 -139 -2356
rect -119 -2403 -115 -2356
rect -119 -2417 -115 -2407
rect -101 -2396 -97 -2356
rect -101 -2417 -97 -2400
rect -77 -2410 -73 -2356
rect -59 -2388 -55 -2356
rect -59 -2396 -55 -2392
rect -77 -2417 -73 -2414
rect -201 -2421 -192 -2417
rect -185 -2421 -177 -2417
rect -201 -2424 -197 -2421
rect -177 -2424 -173 -2421
rect -169 -2421 -157 -2417
rect -143 -2421 -135 -2417
rect -169 -2424 -165 -2421
rect -135 -2424 -131 -2421
rect -127 -2421 -115 -2417
rect -101 -2421 -89 -2417
rect -127 -2424 -123 -2421
rect -93 -2424 -89 -2421
rect -85 -2421 -73 -2417
rect -59 -2417 -55 -2400
rect -35 -2403 -31 -2356
rect -35 -2417 -31 -2407
rect -59 -2421 -47 -2417
rect -85 -2424 -81 -2421
rect -51 -2424 -47 -2421
rect -43 -2421 -31 -2417
rect -43 -2424 -39 -2421
rect -210 -2432 -206 -2428
rect -193 -2432 -189 -2428
rect -152 -2432 -148 -2428
rect -110 -2432 -106 -2428
rect -68 -2432 -64 -2428
rect -27 -2432 -23 -2428
rect -8 -2440 -4 -2392
rect 111 -2396 115 -2128
rect -211 -2519 -207 -2515
rect -194 -2519 -190 -2515
rect -174 -2519 -170 -2515
rect -153 -2519 -149 -2515
rect -132 -2519 -128 -2515
rect -111 -2519 -107 -2515
rect -90 -2519 -86 -2515
rect -69 -2519 -65 -2515
rect -48 -2519 -44 -2515
rect -28 -2519 -24 -2515
rect -220 -2574 -216 -2527
rect -220 -2595 -216 -2578
rect -202 -2588 -198 -2527
rect -186 -2588 -182 -2527
rect -162 -2567 -158 -2527
rect -162 -2588 -158 -2571
rect -144 -2588 -140 -2527
rect -120 -2574 -116 -2527
rect -120 -2588 -116 -2578
rect -102 -2567 -98 -2527
rect -102 -2588 -98 -2571
rect -78 -2581 -74 -2527
rect -60 -2559 -56 -2527
rect -60 -2567 -56 -2563
rect -78 -2588 -74 -2585
rect -202 -2592 -193 -2588
rect -186 -2592 -178 -2588
rect -202 -2595 -198 -2592
rect -178 -2595 -174 -2592
rect -170 -2592 -158 -2588
rect -144 -2592 -136 -2588
rect -170 -2595 -166 -2592
rect -136 -2595 -132 -2592
rect -128 -2592 -116 -2588
rect -102 -2592 -90 -2588
rect -128 -2595 -124 -2592
rect -94 -2595 -90 -2592
rect -86 -2592 -74 -2588
rect -60 -2588 -56 -2571
rect -36 -2574 -32 -2527
rect -36 -2588 -32 -2578
rect -60 -2592 -48 -2588
rect -86 -2595 -82 -2592
rect -52 -2595 -48 -2592
rect -44 -2592 -32 -2588
rect -44 -2595 -40 -2592
rect -211 -2603 -207 -2599
rect -194 -2603 -190 -2599
rect -153 -2603 -149 -2599
rect -111 -2603 -107 -2599
rect -69 -2603 -65 -2599
rect -28 -2603 -24 -2599
rect -219 -2624 -215 -2620
rect -202 -2624 -198 -2620
rect -211 -2635 -207 -2632
rect -211 -2639 -196 -2635
rect -233 -2652 -218 -2648
rect -568 -2902 -564 -2898
rect -551 -2902 -547 -2898
rect -531 -2902 -527 -2898
rect -510 -2902 -506 -2898
rect -489 -2902 -485 -2898
rect -468 -2902 -464 -2898
rect -447 -2902 -443 -2898
rect -426 -2902 -422 -2898
rect -405 -2902 -401 -2898
rect -385 -2902 -381 -2898
rect -577 -2957 -573 -2910
rect -577 -2978 -573 -2961
rect -559 -2971 -555 -2910
rect -543 -2971 -539 -2910
rect -519 -2950 -515 -2910
rect -519 -2971 -515 -2954
rect -501 -2971 -497 -2910
rect -477 -2957 -473 -2910
rect -477 -2971 -473 -2961
rect -459 -2950 -455 -2910
rect -459 -2971 -455 -2954
rect -435 -2964 -431 -2910
rect -417 -2942 -413 -2910
rect -417 -2950 -413 -2946
rect -435 -2971 -431 -2968
rect -559 -2975 -550 -2971
rect -543 -2975 -535 -2971
rect -559 -2978 -555 -2975
rect -535 -2978 -531 -2975
rect -527 -2975 -515 -2971
rect -501 -2975 -493 -2971
rect -527 -2978 -523 -2975
rect -493 -2978 -489 -2975
rect -485 -2975 -473 -2971
rect -459 -2975 -447 -2971
rect -485 -2978 -481 -2975
rect -451 -2978 -447 -2975
rect -443 -2975 -431 -2971
rect -417 -2971 -413 -2954
rect -393 -2957 -389 -2910
rect -393 -2971 -389 -2961
rect -417 -2975 -405 -2971
rect -443 -2978 -439 -2975
rect -409 -2978 -405 -2975
rect -401 -2975 -389 -2971
rect -401 -2978 -397 -2975
rect -568 -2986 -564 -2982
rect -551 -2986 -547 -2982
rect -510 -2986 -506 -2982
rect -468 -2986 -464 -2982
rect -426 -2986 -422 -2982
rect -385 -2986 -381 -2982
rect -568 -3073 -564 -3069
rect -551 -3073 -547 -3069
rect -531 -3073 -527 -3069
rect -510 -3073 -506 -3069
rect -489 -3073 -485 -3069
rect -468 -3073 -464 -3069
rect -447 -3073 -443 -3069
rect -426 -3073 -422 -3069
rect -405 -3073 -401 -3069
rect -385 -3073 -381 -3069
rect -577 -3128 -573 -3081
rect -577 -3149 -573 -3132
rect -559 -3142 -555 -3081
rect -543 -3142 -539 -3081
rect -519 -3121 -515 -3081
rect -519 -3142 -515 -3125
rect -501 -3142 -497 -3081
rect -477 -3128 -473 -3081
rect -477 -3142 -473 -3132
rect -459 -3121 -455 -3081
rect -459 -3142 -455 -3125
rect -435 -3135 -431 -3081
rect -417 -3113 -413 -3081
rect -417 -3121 -413 -3117
rect -435 -3142 -431 -3139
rect -559 -3146 -550 -3142
rect -543 -3146 -535 -3142
rect -559 -3149 -555 -3146
rect -535 -3149 -531 -3146
rect -527 -3146 -515 -3142
rect -501 -3146 -493 -3142
rect -527 -3149 -523 -3146
rect -493 -3149 -489 -3146
rect -485 -3146 -473 -3142
rect -459 -3146 -447 -3142
rect -485 -3149 -481 -3146
rect -451 -3149 -447 -3146
rect -443 -3146 -431 -3142
rect -417 -3142 -413 -3125
rect -393 -3128 -389 -3081
rect -393 -3142 -389 -3132
rect -417 -3146 -405 -3142
rect -443 -3149 -439 -3146
rect -409 -3149 -405 -3146
rect -401 -3146 -389 -3142
rect -401 -3149 -397 -3146
rect -568 -3157 -564 -3153
rect -551 -3157 -547 -3153
rect -510 -3157 -506 -3153
rect -468 -3157 -464 -3153
rect -426 -3157 -422 -3153
rect -385 -3157 -381 -3153
rect -367 -3164 -363 -3117
rect -249 -3121 -245 -2885
rect -568 -3244 -564 -3240
rect -551 -3244 -547 -3240
rect -531 -3244 -527 -3240
rect -510 -3244 -506 -3240
rect -489 -3244 -485 -3240
rect -468 -3244 -464 -3240
rect -447 -3244 -443 -3240
rect -426 -3244 -422 -3240
rect -405 -3244 -401 -3240
rect -385 -3244 -381 -3240
rect -577 -3299 -573 -3252
rect -577 -3320 -573 -3303
rect -559 -3313 -555 -3252
rect -543 -3313 -539 -3252
rect -519 -3292 -515 -3252
rect -519 -3313 -515 -3296
rect -501 -3313 -497 -3252
rect -477 -3299 -473 -3252
rect -477 -3313 -473 -3303
rect -459 -3292 -455 -3252
rect -459 -3313 -455 -3296
rect -435 -3306 -431 -3252
rect -417 -3284 -413 -3252
rect -417 -3292 -413 -3288
rect -435 -3313 -431 -3310
rect -559 -3317 -550 -3313
rect -543 -3317 -535 -3313
rect -559 -3320 -555 -3317
rect -535 -3320 -531 -3317
rect -527 -3317 -515 -3313
rect -501 -3317 -493 -3313
rect -527 -3320 -523 -3317
rect -493 -3320 -489 -3317
rect -485 -3317 -473 -3313
rect -459 -3317 -447 -3313
rect -485 -3320 -481 -3317
rect -451 -3320 -447 -3317
rect -443 -3317 -431 -3313
rect -417 -3313 -413 -3296
rect -393 -3299 -389 -3252
rect -393 -3313 -389 -3303
rect -417 -3317 -405 -3313
rect -443 -3320 -439 -3317
rect -409 -3320 -405 -3317
rect -401 -3317 -389 -3313
rect -401 -3320 -397 -3317
rect -568 -3328 -564 -3324
rect -551 -3328 -547 -3324
rect -510 -3328 -506 -3324
rect -468 -3328 -464 -3324
rect -426 -3328 -422 -3324
rect -385 -3328 -381 -3324
rect -577 -3355 -573 -3351
rect -560 -3355 -556 -3351
rect -569 -3366 -565 -3363
rect -569 -3370 -554 -3366
rect -591 -3383 -576 -3379
rect -925 -3644 -921 -3640
rect -908 -3644 -904 -3640
rect -888 -3644 -884 -3640
rect -867 -3644 -863 -3640
rect -846 -3644 -842 -3640
rect -825 -3644 -821 -3640
rect -804 -3644 -800 -3640
rect -783 -3644 -779 -3640
rect -762 -3644 -758 -3640
rect -742 -3644 -738 -3640
rect -934 -3699 -930 -3652
rect -934 -3720 -930 -3703
rect -916 -3713 -912 -3652
rect -900 -3713 -896 -3652
rect -876 -3692 -872 -3652
rect -876 -3713 -872 -3696
rect -858 -3713 -854 -3652
rect -834 -3699 -830 -3652
rect -834 -3713 -830 -3703
rect -816 -3692 -812 -3652
rect -816 -3713 -812 -3696
rect -792 -3706 -788 -3652
rect -774 -3684 -770 -3652
rect -774 -3692 -770 -3688
rect -792 -3713 -788 -3710
rect -916 -3717 -907 -3713
rect -900 -3717 -892 -3713
rect -916 -3720 -912 -3717
rect -892 -3720 -888 -3717
rect -884 -3717 -872 -3713
rect -858 -3717 -850 -3713
rect -884 -3720 -880 -3717
rect -850 -3720 -846 -3717
rect -842 -3717 -830 -3713
rect -816 -3717 -804 -3713
rect -842 -3720 -838 -3717
rect -808 -3720 -804 -3717
rect -800 -3717 -788 -3713
rect -774 -3713 -770 -3696
rect -750 -3699 -746 -3652
rect -750 -3713 -746 -3703
rect -774 -3717 -762 -3713
rect -800 -3720 -796 -3717
rect -766 -3720 -762 -3717
rect -758 -3717 -746 -3713
rect -758 -3720 -754 -3717
rect -925 -3728 -921 -3724
rect -908 -3728 -904 -3724
rect -867 -3728 -863 -3724
rect -825 -3728 -821 -3724
rect -783 -3728 -779 -3724
rect -742 -3728 -738 -3724
rect -925 -3815 -921 -3811
rect -908 -3815 -904 -3811
rect -888 -3815 -884 -3811
rect -867 -3815 -863 -3811
rect -846 -3815 -842 -3811
rect -825 -3815 -821 -3811
rect -804 -3815 -800 -3811
rect -783 -3815 -779 -3811
rect -762 -3815 -758 -3811
rect -742 -3815 -738 -3811
rect -934 -3870 -930 -3823
rect -934 -3891 -930 -3874
rect -916 -3884 -912 -3823
rect -900 -3884 -896 -3823
rect -876 -3863 -872 -3823
rect -876 -3884 -872 -3867
rect -858 -3884 -854 -3823
rect -834 -3870 -830 -3823
rect -834 -3884 -830 -3874
rect -816 -3863 -812 -3823
rect -816 -3884 -812 -3867
rect -792 -3877 -788 -3823
rect -774 -3855 -770 -3823
rect -774 -3863 -770 -3859
rect -792 -3884 -788 -3881
rect -916 -3888 -907 -3884
rect -900 -3888 -892 -3884
rect -916 -3891 -912 -3888
rect -892 -3891 -888 -3888
rect -884 -3888 -872 -3884
rect -858 -3888 -850 -3884
rect -884 -3891 -880 -3888
rect -850 -3891 -846 -3888
rect -842 -3888 -830 -3884
rect -816 -3888 -804 -3884
rect -842 -3891 -838 -3888
rect -808 -3891 -804 -3888
rect -800 -3888 -788 -3884
rect -774 -3884 -770 -3867
rect -750 -3870 -746 -3823
rect -750 -3884 -746 -3874
rect -774 -3888 -762 -3884
rect -800 -3891 -796 -3888
rect -766 -3891 -762 -3888
rect -758 -3888 -746 -3884
rect -758 -3891 -754 -3888
rect -925 -3899 -921 -3895
rect -908 -3899 -904 -3895
rect -867 -3899 -863 -3895
rect -825 -3899 -821 -3895
rect -783 -3899 -779 -3895
rect -742 -3899 -738 -3895
rect -723 -3907 -719 -3859
rect -603 -3863 -599 -3609
rect -926 -3990 -922 -3986
rect -909 -3990 -905 -3986
rect -889 -3990 -885 -3986
rect -868 -3990 -864 -3986
rect -847 -3990 -843 -3986
rect -826 -3990 -822 -3986
rect -805 -3990 -801 -3986
rect -784 -3990 -780 -3986
rect -763 -3990 -759 -3986
rect -743 -3990 -739 -3986
rect -935 -4045 -931 -3998
rect -935 -4066 -931 -4049
rect -917 -4059 -913 -3998
rect -901 -4059 -897 -3998
rect -877 -4038 -873 -3998
rect -877 -4059 -873 -4042
rect -859 -4059 -855 -3998
rect -835 -4045 -831 -3998
rect -835 -4059 -831 -4049
rect -817 -4038 -813 -3998
rect -817 -4059 -813 -4042
rect -793 -4052 -789 -3998
rect -775 -4030 -771 -3998
rect -775 -4038 -771 -4034
rect -793 -4059 -789 -4056
rect -917 -4063 -908 -4059
rect -901 -4063 -893 -4059
rect -917 -4066 -913 -4063
rect -893 -4066 -889 -4063
rect -885 -4063 -873 -4059
rect -859 -4063 -851 -4059
rect -885 -4066 -881 -4063
rect -851 -4066 -847 -4063
rect -843 -4063 -831 -4059
rect -817 -4063 -805 -4059
rect -843 -4066 -839 -4063
rect -809 -4066 -805 -4063
rect -801 -4063 -789 -4059
rect -775 -4059 -771 -4042
rect -751 -4045 -747 -3998
rect -751 -4059 -747 -4049
rect -775 -4063 -763 -4059
rect -801 -4066 -797 -4063
rect -767 -4066 -763 -4063
rect -759 -4063 -747 -4059
rect -759 -4066 -755 -4063
rect -926 -4074 -922 -4070
rect -909 -4074 -905 -4070
rect -868 -4074 -864 -4070
rect -826 -4074 -822 -4070
rect -784 -4074 -780 -4070
rect -743 -4074 -739 -4070
rect -935 -4105 -931 -4101
rect -918 -4105 -914 -4101
rect -927 -4116 -923 -4113
rect -927 -4120 -912 -4116
rect -949 -4133 -934 -4129
rect -1225 -4348 -1221 -4344
rect -1181 -4348 -1177 -4344
rect -1147 -4348 -1143 -4344
rect -1257 -4606 -1253 -4359
rect -1114 -4362 -1110 -4330
rect -1246 -4435 -1242 -4366
rect -1225 -4387 -1221 -4383
rect -1208 -4387 -1204 -4383
rect -1188 -4387 -1184 -4383
rect -1167 -4387 -1163 -4383
rect -1146 -4387 -1142 -4383
rect -1125 -4387 -1121 -4383
rect -1104 -4387 -1100 -4383
rect -1083 -4387 -1079 -4383
rect -1062 -4387 -1058 -4383
rect -1042 -4387 -1038 -4383
rect -1234 -4442 -1230 -4395
rect -1234 -4463 -1230 -4446
rect -1216 -4456 -1212 -4395
rect -1200 -4456 -1196 -4395
rect -1176 -4435 -1172 -4395
rect -1176 -4456 -1172 -4439
rect -1158 -4456 -1154 -4395
rect -1134 -4442 -1130 -4395
rect -1134 -4456 -1130 -4446
rect -1116 -4435 -1112 -4395
rect -1116 -4456 -1112 -4439
rect -1092 -4449 -1088 -4395
rect -1074 -4427 -1070 -4395
rect -1074 -4435 -1070 -4431
rect -1092 -4456 -1088 -4453
rect -1216 -4460 -1207 -4456
rect -1200 -4460 -1192 -4456
rect -1216 -4463 -1212 -4460
rect -1192 -4463 -1188 -4460
rect -1184 -4460 -1172 -4456
rect -1158 -4460 -1150 -4456
rect -1184 -4463 -1180 -4460
rect -1150 -4463 -1146 -4460
rect -1142 -4460 -1130 -4456
rect -1116 -4460 -1104 -4456
rect -1142 -4463 -1138 -4460
rect -1108 -4463 -1104 -4460
rect -1100 -4460 -1088 -4456
rect -1074 -4456 -1070 -4439
rect -1050 -4442 -1046 -4395
rect -1050 -4456 -1046 -4446
rect -1074 -4460 -1062 -4456
rect -1100 -4463 -1096 -4460
rect -1066 -4463 -1062 -4460
rect -1058 -4460 -1046 -4456
rect -1058 -4463 -1054 -4460
rect -1225 -4471 -1221 -4467
rect -1208 -4471 -1204 -4467
rect -1167 -4471 -1163 -4467
rect -1125 -4471 -1121 -4467
rect -1083 -4471 -1079 -4467
rect -1042 -4471 -1038 -4467
rect -1225 -4558 -1221 -4554
rect -1208 -4558 -1204 -4554
rect -1188 -4558 -1184 -4554
rect -1167 -4558 -1163 -4554
rect -1146 -4558 -1142 -4554
rect -1125 -4558 -1121 -4554
rect -1104 -4558 -1100 -4554
rect -1083 -4558 -1079 -4554
rect -1062 -4558 -1058 -4554
rect -1042 -4558 -1038 -4554
rect -1234 -4613 -1230 -4566
rect -1234 -4634 -1230 -4617
rect -1216 -4627 -1212 -4566
rect -1200 -4627 -1196 -4566
rect -1176 -4606 -1172 -4566
rect -1176 -4627 -1172 -4610
rect -1158 -4627 -1154 -4566
rect -1134 -4613 -1130 -4566
rect -1134 -4627 -1130 -4617
rect -1116 -4606 -1112 -4566
rect -1116 -4627 -1112 -4610
rect -1092 -4620 -1088 -4566
rect -1074 -4598 -1070 -4566
rect -1074 -4606 -1070 -4602
rect -1092 -4627 -1088 -4624
rect -1216 -4631 -1207 -4627
rect -1200 -4631 -1192 -4627
rect -1216 -4634 -1212 -4631
rect -1192 -4634 -1188 -4631
rect -1184 -4631 -1172 -4627
rect -1158 -4631 -1150 -4627
rect -1184 -4634 -1180 -4631
rect -1150 -4634 -1146 -4631
rect -1142 -4631 -1130 -4627
rect -1116 -4631 -1104 -4627
rect -1142 -4634 -1138 -4631
rect -1108 -4634 -1104 -4631
rect -1100 -4631 -1088 -4627
rect -1074 -4627 -1070 -4610
rect -1050 -4613 -1046 -4566
rect -1050 -4627 -1046 -4617
rect -1074 -4631 -1062 -4627
rect -1100 -4634 -1096 -4631
rect -1066 -4634 -1062 -4631
rect -1058 -4631 -1046 -4627
rect -1058 -4634 -1054 -4631
rect -1225 -4642 -1221 -4638
rect -1208 -4642 -1204 -4638
rect -1167 -4642 -1163 -4638
rect -1125 -4642 -1121 -4638
rect -1083 -4642 -1079 -4638
rect -1042 -4642 -1038 -4638
rect -1023 -4650 -1019 -4602
rect -963 -4606 -959 -4366
rect -1309 -4844 -1305 -4840
rect -1292 -4844 -1288 -4840
rect -1301 -4855 -1297 -4852
rect -1301 -4859 -1286 -4855
rect -1319 -4872 -1308 -4868
rect -1801 -5122 -1797 -5118
rect -1784 -5122 -1780 -5118
rect -1764 -5122 -1760 -5118
rect -1743 -5122 -1739 -5118
rect -1722 -5122 -1718 -5118
rect -1701 -5122 -1697 -5118
rect -1680 -5122 -1676 -5118
rect -1659 -5122 -1655 -5118
rect -1638 -5122 -1634 -5118
rect -1618 -5122 -1614 -5118
rect -1538 -5122 -1534 -5118
rect -1521 -5122 -1517 -5118
rect -1501 -5122 -1497 -5118
rect -1480 -5122 -1476 -5118
rect -1459 -5122 -1455 -5118
rect -1438 -5122 -1434 -5118
rect -1417 -5122 -1413 -5118
rect -1396 -5122 -1392 -5118
rect -1375 -5122 -1371 -5118
rect -1355 -5122 -1351 -5118
rect -1810 -5177 -1806 -5130
rect -1810 -5198 -1806 -5181
rect -1792 -5191 -1788 -5130
rect -1776 -5191 -1772 -5130
rect -1752 -5170 -1748 -5130
rect -1752 -5191 -1748 -5174
rect -1734 -5191 -1730 -5130
rect -1710 -5177 -1706 -5130
rect -1710 -5191 -1706 -5181
rect -1692 -5170 -1688 -5130
rect -1692 -5191 -1688 -5174
rect -1668 -5184 -1664 -5130
rect -1650 -5162 -1646 -5130
rect -1650 -5170 -1646 -5166
rect -1668 -5191 -1664 -5188
rect -1792 -5195 -1783 -5191
rect -1776 -5195 -1768 -5191
rect -1792 -5198 -1788 -5195
rect -1768 -5198 -1764 -5195
rect -1760 -5195 -1748 -5191
rect -1734 -5195 -1726 -5191
rect -1760 -5198 -1756 -5195
rect -1726 -5198 -1722 -5195
rect -1718 -5195 -1706 -5191
rect -1692 -5195 -1680 -5191
rect -1718 -5198 -1714 -5195
rect -1684 -5198 -1680 -5195
rect -1676 -5195 -1664 -5191
rect -1650 -5191 -1646 -5174
rect -1626 -5177 -1622 -5130
rect -1626 -5191 -1622 -5181
rect -1650 -5195 -1638 -5191
rect -1676 -5198 -1672 -5195
rect -1642 -5198 -1638 -5195
rect -1634 -5195 -1622 -5191
rect -1547 -5177 -1543 -5130
rect -1634 -5198 -1630 -5195
rect -1547 -5198 -1543 -5181
rect -1529 -5191 -1525 -5130
rect -1513 -5191 -1509 -5130
rect -1489 -5170 -1485 -5130
rect -1489 -5191 -1485 -5174
rect -1471 -5191 -1467 -5130
rect -1447 -5177 -1443 -5130
rect -1447 -5191 -1443 -5181
rect -1429 -5170 -1425 -5130
rect -1429 -5191 -1425 -5174
rect -1405 -5184 -1401 -5130
rect -1387 -5162 -1383 -5130
rect -1387 -5170 -1383 -5166
rect -1405 -5191 -1401 -5188
rect -1529 -5195 -1520 -5191
rect -1513 -5195 -1505 -5191
rect -1529 -5198 -1525 -5195
rect -1505 -5198 -1501 -5195
rect -1497 -5195 -1485 -5191
rect -1471 -5195 -1463 -5191
rect -1497 -5198 -1493 -5195
rect -1463 -5198 -1459 -5195
rect -1455 -5195 -1443 -5191
rect -1429 -5195 -1417 -5191
rect -1455 -5198 -1451 -5195
rect -1421 -5198 -1417 -5195
rect -1413 -5195 -1401 -5191
rect -1387 -5191 -1383 -5174
rect -1363 -5177 -1359 -5130
rect -1363 -5191 -1359 -5181
rect -1387 -5195 -1375 -5191
rect -1413 -5198 -1409 -5195
rect -1379 -5198 -1375 -5195
rect -1371 -5195 -1359 -5191
rect -1371 -5198 -1367 -5195
rect -1801 -5206 -1797 -5202
rect -1784 -5206 -1780 -5202
rect -1743 -5206 -1739 -5202
rect -1701 -5206 -1697 -5202
rect -1659 -5206 -1655 -5202
rect -1618 -5206 -1614 -5202
rect -1538 -5206 -1534 -5202
rect -1521 -5206 -1517 -5202
rect -1480 -5206 -1476 -5202
rect -1438 -5206 -1434 -5202
rect -1396 -5206 -1392 -5202
rect -1355 -5206 -1351 -5202
rect -1340 -5214 -1336 -5166
rect -1825 -5341 -1821 -5218
rect -1801 -5293 -1797 -5289
rect -1784 -5293 -1780 -5289
rect -1764 -5293 -1760 -5289
rect -1743 -5293 -1739 -5289
rect -1722 -5293 -1718 -5289
rect -1701 -5293 -1697 -5289
rect -1680 -5293 -1676 -5289
rect -1659 -5293 -1655 -5289
rect -1638 -5293 -1634 -5289
rect -1618 -5293 -1614 -5289
rect -1538 -5293 -1534 -5289
rect -1521 -5293 -1517 -5289
rect -1501 -5293 -1497 -5289
rect -1480 -5293 -1476 -5289
rect -1459 -5293 -1455 -5289
rect -1438 -5293 -1434 -5289
rect -1417 -5293 -1413 -5289
rect -1396 -5293 -1392 -5289
rect -1375 -5293 -1371 -5289
rect -1355 -5293 -1351 -5289
rect -1810 -5348 -1806 -5301
rect -1810 -5369 -1806 -5352
rect -1792 -5362 -1788 -5301
rect -1776 -5362 -1772 -5301
rect -1752 -5341 -1748 -5301
rect -1752 -5362 -1748 -5345
rect -1734 -5362 -1730 -5301
rect -1710 -5348 -1706 -5301
rect -1710 -5362 -1706 -5352
rect -1692 -5341 -1688 -5301
rect -1692 -5362 -1688 -5345
rect -1668 -5355 -1664 -5301
rect -1650 -5333 -1646 -5301
rect -1650 -5341 -1646 -5337
rect -1668 -5362 -1664 -5359
rect -1792 -5366 -1783 -5362
rect -1776 -5366 -1768 -5362
rect -1792 -5369 -1788 -5366
rect -1768 -5369 -1764 -5366
rect -1760 -5366 -1748 -5362
rect -1734 -5366 -1726 -5362
rect -1760 -5369 -1756 -5366
rect -1726 -5369 -1722 -5366
rect -1718 -5366 -1706 -5362
rect -1692 -5366 -1680 -5362
rect -1718 -5369 -1714 -5366
rect -1684 -5369 -1680 -5366
rect -1676 -5366 -1664 -5362
rect -1650 -5362 -1646 -5345
rect -1626 -5348 -1622 -5301
rect -1626 -5362 -1622 -5352
rect -1650 -5366 -1638 -5362
rect -1676 -5369 -1672 -5366
rect -1642 -5369 -1638 -5366
rect -1634 -5366 -1622 -5362
rect -1547 -5348 -1543 -5301
rect -1634 -5369 -1630 -5366
rect -1547 -5369 -1543 -5352
rect -1529 -5362 -1525 -5301
rect -1513 -5362 -1509 -5301
rect -1489 -5341 -1485 -5301
rect -1489 -5362 -1485 -5345
rect -1471 -5362 -1467 -5301
rect -1447 -5348 -1443 -5301
rect -1447 -5362 -1443 -5352
rect -1429 -5341 -1425 -5301
rect -1429 -5362 -1425 -5345
rect -1405 -5355 -1401 -5301
rect -1387 -5333 -1383 -5301
rect -1387 -5341 -1383 -5337
rect -1405 -5362 -1401 -5359
rect -1529 -5366 -1520 -5362
rect -1513 -5366 -1505 -5362
rect -1529 -5369 -1525 -5366
rect -1505 -5369 -1501 -5366
rect -1497 -5366 -1485 -5362
rect -1471 -5366 -1463 -5362
rect -1497 -5369 -1493 -5366
rect -1463 -5369 -1459 -5366
rect -1455 -5366 -1443 -5362
rect -1429 -5366 -1417 -5362
rect -1455 -5369 -1451 -5366
rect -1421 -5369 -1417 -5366
rect -1413 -5366 -1401 -5362
rect -1387 -5362 -1383 -5345
rect -1363 -5348 -1359 -5301
rect -1363 -5362 -1359 -5352
rect -1387 -5366 -1375 -5362
rect -1413 -5369 -1409 -5366
rect -1379 -5369 -1375 -5366
rect -1371 -5366 -1359 -5362
rect -1371 -5369 -1367 -5366
rect -1801 -5377 -1797 -5373
rect -1784 -5377 -1780 -5373
rect -1743 -5377 -1739 -5373
rect -1701 -5377 -1697 -5373
rect -1659 -5377 -1655 -5373
rect -1618 -5377 -1614 -5373
rect -1538 -5377 -1534 -5373
rect -1521 -5377 -1517 -5373
rect -1480 -5377 -1476 -5373
rect -1438 -5377 -1434 -5373
rect -1396 -5377 -1392 -5373
rect -1355 -5377 -1351 -5373
rect -1340 -5385 -1336 -5337
rect -1826 -5501 -1822 -5389
rect -1801 -5453 -1797 -5449
rect -1784 -5453 -1780 -5449
rect -1764 -5453 -1760 -5449
rect -1743 -5453 -1739 -5449
rect -1722 -5453 -1718 -5449
rect -1701 -5453 -1697 -5449
rect -1680 -5453 -1676 -5449
rect -1659 -5453 -1655 -5449
rect -1638 -5453 -1634 -5449
rect -1618 -5453 -1614 -5449
rect -1538 -5453 -1534 -5449
rect -1521 -5453 -1517 -5449
rect -1501 -5453 -1497 -5449
rect -1480 -5453 -1476 -5449
rect -1459 -5453 -1455 -5449
rect -1438 -5453 -1434 -5449
rect -1417 -5453 -1413 -5449
rect -1396 -5453 -1392 -5449
rect -1375 -5453 -1371 -5449
rect -1355 -5453 -1351 -5449
rect -1810 -5508 -1806 -5461
rect -1810 -5529 -1806 -5512
rect -1792 -5522 -1788 -5461
rect -1776 -5522 -1772 -5461
rect -1752 -5501 -1748 -5461
rect -1752 -5522 -1748 -5505
rect -1734 -5522 -1730 -5461
rect -1710 -5508 -1706 -5461
rect -1710 -5522 -1706 -5512
rect -1692 -5501 -1688 -5461
rect -1692 -5522 -1688 -5505
rect -1668 -5515 -1664 -5461
rect -1650 -5493 -1646 -5461
rect -1650 -5501 -1646 -5497
rect -1668 -5522 -1664 -5519
rect -1792 -5526 -1783 -5522
rect -1776 -5526 -1768 -5522
rect -1792 -5529 -1788 -5526
rect -1768 -5529 -1764 -5526
rect -1760 -5526 -1748 -5522
rect -1734 -5526 -1726 -5522
rect -1760 -5529 -1756 -5526
rect -1726 -5529 -1722 -5526
rect -1718 -5526 -1706 -5522
rect -1692 -5526 -1680 -5522
rect -1718 -5529 -1714 -5526
rect -1684 -5529 -1680 -5526
rect -1676 -5526 -1664 -5522
rect -1650 -5522 -1646 -5505
rect -1626 -5508 -1622 -5461
rect -1626 -5522 -1622 -5512
rect -1650 -5526 -1638 -5522
rect -1676 -5529 -1672 -5526
rect -1642 -5529 -1638 -5526
rect -1634 -5526 -1622 -5522
rect -1547 -5508 -1543 -5461
rect -1634 -5529 -1630 -5526
rect -1547 -5529 -1543 -5512
rect -1529 -5522 -1525 -5461
rect -1513 -5522 -1509 -5461
rect -1489 -5501 -1485 -5461
rect -1489 -5522 -1485 -5505
rect -1471 -5522 -1467 -5461
rect -1447 -5508 -1443 -5461
rect -1447 -5522 -1443 -5512
rect -1429 -5501 -1425 -5461
rect -1429 -5522 -1425 -5505
rect -1405 -5515 -1401 -5461
rect -1387 -5493 -1383 -5461
rect -1387 -5501 -1383 -5497
rect -1405 -5522 -1401 -5519
rect -1529 -5526 -1520 -5522
rect -1513 -5526 -1505 -5522
rect -1529 -5529 -1525 -5526
rect -1505 -5529 -1501 -5526
rect -1497 -5526 -1485 -5522
rect -1471 -5526 -1463 -5522
rect -1497 -5529 -1493 -5526
rect -1463 -5529 -1459 -5526
rect -1455 -5526 -1443 -5522
rect -1429 -5526 -1417 -5522
rect -1455 -5529 -1451 -5526
rect -1421 -5529 -1417 -5526
rect -1413 -5526 -1401 -5522
rect -1387 -5522 -1383 -5505
rect -1363 -5508 -1359 -5461
rect -1363 -5522 -1359 -5512
rect -1387 -5526 -1375 -5522
rect -1413 -5529 -1409 -5526
rect -1379 -5529 -1375 -5526
rect -1371 -5526 -1359 -5522
rect -1371 -5529 -1367 -5526
rect -1801 -5537 -1797 -5533
rect -1784 -5537 -1780 -5533
rect -1743 -5537 -1739 -5533
rect -1701 -5537 -1697 -5533
rect -1659 -5537 -1655 -5533
rect -1618 -5537 -1614 -5533
rect -1538 -5537 -1534 -5533
rect -1521 -5537 -1517 -5533
rect -1480 -5537 -1476 -5533
rect -1438 -5537 -1434 -5533
rect -1396 -5537 -1392 -5533
rect -1355 -5537 -1351 -5533
rect -1342 -5599 -1338 -5497
rect -1319 -5501 -1315 -4872
rect -1290 -4898 -1286 -4859
rect -1290 -4913 -1286 -4902
rect -1309 -4917 -1286 -4913
rect -1309 -4920 -1305 -4917
rect -1283 -4920 -1279 -4852
rect -1292 -4928 -1288 -4924
rect -1283 -5058 -1279 -4924
rect -1257 -5051 -1253 -4654
rect -1225 -4729 -1221 -4725
rect -1208 -4729 -1204 -4725
rect -1188 -4729 -1184 -4725
rect -1167 -4729 -1163 -4725
rect -1146 -4729 -1142 -4725
rect -1125 -4729 -1121 -4725
rect -1104 -4729 -1100 -4725
rect -1083 -4729 -1079 -4725
rect -1062 -4729 -1058 -4725
rect -1042 -4729 -1038 -4725
rect -1234 -4784 -1230 -4737
rect -1234 -4805 -1230 -4788
rect -1216 -4798 -1212 -4737
rect -1200 -4798 -1196 -4737
rect -1176 -4777 -1172 -4737
rect -1176 -4798 -1172 -4781
rect -1158 -4798 -1154 -4737
rect -1134 -4784 -1130 -4737
rect -1134 -4798 -1130 -4788
rect -1116 -4777 -1112 -4737
rect -1116 -4798 -1112 -4781
rect -1092 -4791 -1088 -4737
rect -1074 -4769 -1070 -4737
rect -1074 -4777 -1070 -4773
rect -1092 -4798 -1088 -4795
rect -1216 -4802 -1207 -4798
rect -1200 -4802 -1192 -4798
rect -1216 -4805 -1212 -4802
rect -1192 -4805 -1188 -4802
rect -1184 -4802 -1172 -4798
rect -1158 -4802 -1150 -4798
rect -1184 -4805 -1180 -4802
rect -1150 -4805 -1146 -4802
rect -1142 -4802 -1130 -4798
rect -1116 -4802 -1104 -4798
rect -1142 -4805 -1138 -4802
rect -1108 -4805 -1104 -4802
rect -1100 -4802 -1088 -4798
rect -1074 -4798 -1070 -4781
rect -1050 -4784 -1046 -4737
rect -1050 -4798 -1046 -4788
rect -1074 -4802 -1062 -4798
rect -1100 -4805 -1096 -4802
rect -1066 -4805 -1062 -4802
rect -1058 -4802 -1046 -4798
rect -1058 -4805 -1054 -4802
rect -1225 -4813 -1221 -4809
rect -1208 -4813 -1204 -4809
rect -1167 -4813 -1163 -4809
rect -1125 -4813 -1121 -4809
rect -1083 -4813 -1079 -4809
rect -1042 -4813 -1038 -4809
rect -1022 -4868 -1018 -4773
rect -1225 -5003 -1221 -4999
rect -1208 -5003 -1204 -4999
rect -1168 -5003 -1164 -4999
rect -1147 -5003 -1143 -4999
rect -1234 -5044 -1230 -5011
rect -1234 -5079 -1230 -5048
rect -1216 -5038 -1212 -5011
rect -1216 -5042 -1207 -5038
rect -1216 -5079 -1212 -5042
rect -1190 -5065 -1186 -5011
rect -1190 -5072 -1186 -5069
rect -1156 -5072 -1152 -5011
rect -1138 -5043 -1134 -5011
rect -979 -5035 -975 -4893
rect -1208 -5079 -1204 -5076
rect -1199 -5076 -1186 -5072
rect -1199 -5079 -1195 -5076
rect -1172 -5079 -1168 -5076
rect -1164 -5076 -1145 -5072
rect -1164 -5079 -1160 -5076
rect -1138 -5079 -1134 -5047
rect -963 -5050 -959 -4653
rect -949 -4777 -945 -4133
rect -916 -4159 -912 -4120
rect -916 -4174 -912 -4163
rect -935 -4178 -912 -4174
rect -909 -4150 -905 -4113
rect -719 -4129 -715 -4034
rect -935 -4181 -931 -4178
rect -909 -4181 -905 -4154
rect -918 -4189 -914 -4185
rect -926 -4264 -922 -4260
rect -900 -4264 -896 -4260
rect -883 -4264 -879 -4260
rect -843 -4264 -839 -4260
rect -822 -4264 -818 -4260
rect -805 -4264 -801 -4260
rect -765 -4264 -761 -4260
rect -741 -4264 -737 -4260
rect -704 -4264 -700 -4260
rect -935 -4289 -931 -4272
rect -935 -4340 -931 -4293
rect -917 -4282 -913 -4272
rect -917 -4340 -913 -4286
rect -909 -4311 -905 -4272
rect -891 -4304 -887 -4272
rect -909 -4340 -905 -4315
rect -891 -4340 -887 -4308
rect -865 -4296 -861 -4272
rect -865 -4333 -861 -4300
rect -831 -4333 -827 -4272
rect -813 -4289 -809 -4272
rect -883 -4340 -879 -4337
rect -875 -4337 -861 -4333
rect -875 -4340 -871 -4337
rect -847 -4340 -843 -4337
rect -839 -4337 -820 -4333
rect -839 -4340 -835 -4337
rect -813 -4340 -809 -4293
rect -787 -4304 -783 -4272
rect -787 -4333 -783 -4308
rect -753 -4326 -749 -4272
rect -753 -4330 -736 -4326
rect -805 -4340 -801 -4337
rect -796 -4337 -783 -4333
rect -796 -4340 -792 -4337
rect -769 -4340 -765 -4337
rect -745 -4340 -741 -4330
rect -729 -4333 -725 -4272
rect -721 -4326 -717 -4272
rect -695 -4296 -691 -4272
rect -721 -4330 -702 -4326
rect -737 -4337 -720 -4333
rect -737 -4340 -733 -4337
rect -713 -4340 -709 -4330
rect -695 -4340 -691 -4300
rect -926 -4348 -922 -4344
rect -900 -4348 -896 -4344
rect -857 -4348 -853 -4344
rect -822 -4348 -818 -4344
rect -778 -4348 -774 -4344
rect -761 -4348 -757 -4344
rect -725 -4348 -721 -4344
rect -704 -4348 -700 -4344
rect -687 -4355 -683 -4308
rect -616 -4311 -612 -4154
rect -603 -4296 -599 -3910
rect -591 -4038 -587 -3383
rect -558 -3409 -554 -3370
rect -558 -3424 -554 -3413
rect -577 -3428 -554 -3424
rect -551 -3400 -547 -3363
rect -369 -3379 -365 -3288
rect -577 -3431 -573 -3428
rect -551 -3431 -547 -3404
rect -560 -3439 -556 -3435
rect -568 -3514 -564 -3510
rect -542 -3514 -538 -3510
rect -525 -3514 -521 -3510
rect -485 -3514 -481 -3510
rect -464 -3514 -460 -3510
rect -447 -3514 -443 -3510
rect -407 -3514 -403 -3510
rect -383 -3514 -379 -3510
rect -346 -3514 -342 -3510
rect -577 -3539 -573 -3522
rect -577 -3590 -573 -3543
rect -559 -3532 -555 -3522
rect -559 -3590 -555 -3536
rect -551 -3561 -547 -3522
rect -533 -3554 -529 -3522
rect -551 -3590 -547 -3565
rect -533 -3590 -529 -3558
rect -507 -3546 -503 -3522
rect -507 -3583 -503 -3550
rect -473 -3583 -469 -3522
rect -455 -3539 -451 -3522
rect -525 -3590 -521 -3587
rect -517 -3587 -503 -3583
rect -517 -3590 -513 -3587
rect -489 -3590 -485 -3587
rect -481 -3587 -462 -3583
rect -481 -3590 -477 -3587
rect -455 -3590 -451 -3543
rect -429 -3554 -425 -3522
rect -429 -3583 -425 -3558
rect -395 -3576 -391 -3522
rect -395 -3580 -378 -3576
rect -447 -3590 -443 -3587
rect -438 -3587 -425 -3583
rect -438 -3590 -434 -3587
rect -411 -3590 -407 -3587
rect -387 -3590 -383 -3580
rect -371 -3583 -367 -3522
rect -363 -3576 -359 -3522
rect -337 -3545 -333 -3522
rect -363 -3580 -344 -3576
rect -379 -3587 -362 -3583
rect -379 -3590 -375 -3587
rect -355 -3590 -351 -3580
rect -337 -3590 -333 -3549
rect -568 -3598 -564 -3594
rect -542 -3598 -538 -3594
rect -499 -3598 -495 -3594
rect -464 -3598 -460 -3594
rect -420 -3598 -416 -3594
rect -403 -3598 -399 -3594
rect -367 -3598 -363 -3594
rect -346 -3598 -342 -3594
rect -328 -3612 -324 -3558
rect -263 -3561 -259 -3404
rect -249 -3546 -245 -3169
rect -233 -3292 -229 -2652
rect -200 -2678 -196 -2639
rect -200 -2693 -196 -2682
rect -219 -2697 -196 -2693
rect -193 -2669 -189 -2632
rect -12 -2648 -8 -2563
rect -219 -2700 -215 -2697
rect -193 -2700 -189 -2673
rect -202 -2708 -198 -2704
rect -210 -2783 -206 -2779
rect -184 -2783 -180 -2779
rect -167 -2783 -163 -2779
rect -127 -2783 -123 -2779
rect -106 -2783 -102 -2779
rect -89 -2783 -85 -2779
rect -49 -2783 -45 -2779
rect -25 -2783 -21 -2779
rect 12 -2783 16 -2779
rect -219 -2808 -215 -2791
rect -219 -2859 -215 -2812
rect -201 -2801 -197 -2791
rect -201 -2859 -197 -2805
rect -193 -2830 -189 -2791
rect -175 -2823 -171 -2791
rect -193 -2859 -189 -2834
rect -175 -2859 -171 -2827
rect -149 -2815 -145 -2791
rect -149 -2852 -145 -2819
rect -115 -2852 -111 -2791
rect -97 -2808 -93 -2791
rect -167 -2859 -163 -2856
rect -159 -2856 -145 -2852
rect -159 -2859 -155 -2856
rect -131 -2859 -127 -2856
rect -123 -2856 -104 -2852
rect -123 -2859 -119 -2856
rect -97 -2859 -93 -2812
rect -71 -2823 -67 -2791
rect -71 -2852 -67 -2827
rect -37 -2845 -33 -2791
rect -37 -2849 -20 -2845
rect -89 -2859 -85 -2856
rect -80 -2856 -67 -2852
rect -80 -2859 -76 -2856
rect -53 -2859 -49 -2856
rect -29 -2859 -25 -2849
rect -13 -2852 -9 -2791
rect -5 -2845 -1 -2791
rect 21 -2815 25 -2791
rect -5 -2849 14 -2845
rect -21 -2856 -4 -2852
rect -21 -2859 -17 -2856
rect 3 -2859 7 -2849
rect 21 -2859 25 -2819
rect -210 -2867 -206 -2863
rect -184 -2867 -180 -2863
rect -141 -2867 -137 -2863
rect -106 -2867 -102 -2863
rect -62 -2867 -58 -2863
rect -45 -2867 -41 -2863
rect -9 -2867 -5 -2863
rect 12 -2867 16 -2863
rect 28 -2874 32 -2827
rect 97 -2830 101 -2673
rect 111 -2815 115 -2443
rect 125 -2567 129 -1902
rect 158 -1928 162 -1889
rect 158 -1943 162 -1932
rect 139 -1947 162 -1943
rect 165 -1919 169 -1882
rect 350 -1898 354 -1811
rect 139 -1950 143 -1947
rect 165 -1950 169 -1923
rect 156 -1958 160 -1954
rect 148 -2033 152 -2029
rect 174 -2033 178 -2029
rect 191 -2033 195 -2029
rect 231 -2033 235 -2029
rect 252 -2033 256 -2029
rect 269 -2033 273 -2029
rect 309 -2033 313 -2029
rect 333 -2033 337 -2029
rect 370 -2033 374 -2029
rect 139 -2058 143 -2041
rect 139 -2109 143 -2062
rect 157 -2051 161 -2041
rect 157 -2109 161 -2055
rect 165 -2080 169 -2041
rect 183 -2073 187 -2041
rect 165 -2109 169 -2084
rect 183 -2109 187 -2077
rect 209 -2065 213 -2041
rect 209 -2102 213 -2069
rect 243 -2102 247 -2041
rect 261 -2058 265 -2041
rect 191 -2109 195 -2106
rect 199 -2106 213 -2102
rect 199 -2109 203 -2106
rect 227 -2109 231 -2106
rect 235 -2106 254 -2102
rect 235 -2109 239 -2106
rect 261 -2109 265 -2062
rect 287 -2073 291 -2041
rect 287 -2102 291 -2077
rect 321 -2095 325 -2041
rect 321 -2099 338 -2095
rect 269 -2109 273 -2106
rect 278 -2106 291 -2102
rect 278 -2109 282 -2106
rect 305 -2109 309 -2106
rect 329 -2109 333 -2099
rect 345 -2102 349 -2041
rect 353 -2095 357 -2041
rect 379 -2065 383 -2041
rect 353 -2099 372 -2095
rect 337 -2106 354 -2102
rect 337 -2109 341 -2106
rect 361 -2109 365 -2099
rect 379 -2109 383 -2069
rect 148 -2117 152 -2113
rect 174 -2117 178 -2113
rect 217 -2117 221 -2113
rect 252 -2117 256 -2113
rect 296 -2117 300 -2113
rect 313 -2117 317 -2113
rect 349 -2117 353 -2113
rect 370 -2117 374 -2113
rect 388 -2131 392 -2077
rect 451 -2080 455 -1923
rect 470 -2065 474 -1691
rect 481 -1815 485 -1166
rect 514 -1192 518 -1153
rect 514 -1207 518 -1196
rect 495 -1211 518 -1207
rect 521 -1183 525 -1146
rect 495 -1214 499 -1211
rect 521 -1214 525 -1187
rect 512 -1222 516 -1218
rect 504 -1302 508 -1298
rect 530 -1302 534 -1298
rect 547 -1302 551 -1298
rect 587 -1302 591 -1298
rect 608 -1302 612 -1298
rect 625 -1302 629 -1298
rect 665 -1302 669 -1298
rect 689 -1302 693 -1298
rect 726 -1302 730 -1298
rect 495 -1327 499 -1310
rect 495 -1378 499 -1331
rect 513 -1320 517 -1310
rect 513 -1378 517 -1324
rect 521 -1349 525 -1310
rect 539 -1342 543 -1310
rect 521 -1378 525 -1353
rect 539 -1378 543 -1346
rect 565 -1334 569 -1310
rect 565 -1371 569 -1338
rect 599 -1371 603 -1310
rect 617 -1327 621 -1310
rect 547 -1378 551 -1375
rect 555 -1375 569 -1371
rect 555 -1378 559 -1375
rect 583 -1378 587 -1375
rect 591 -1375 610 -1371
rect 591 -1378 595 -1375
rect 617 -1378 621 -1331
rect 643 -1342 647 -1310
rect 643 -1371 647 -1346
rect 677 -1364 681 -1310
rect 677 -1368 694 -1364
rect 625 -1378 629 -1375
rect 634 -1375 647 -1371
rect 634 -1378 638 -1375
rect 661 -1378 665 -1375
rect 685 -1378 689 -1368
rect 701 -1371 705 -1310
rect 709 -1364 713 -1310
rect 735 -1334 739 -1310
rect 709 -1368 728 -1364
rect 693 -1375 710 -1371
rect 693 -1378 697 -1375
rect 717 -1378 721 -1368
rect 735 -1378 739 -1338
rect 504 -1386 508 -1382
rect 530 -1386 534 -1382
rect 573 -1386 577 -1382
rect 608 -1386 612 -1382
rect 652 -1386 656 -1382
rect 669 -1386 673 -1382
rect 705 -1386 709 -1382
rect 726 -1386 730 -1382
rect 742 -1407 746 -1346
rect 805 -1349 809 -1187
rect 821 -1334 825 -840
rect 839 -1162 843 -816
rect 872 -857 876 -803
rect 853 -861 872 -857
rect 879 -828 883 -796
rect 853 -864 857 -861
rect 879 -864 883 -832
rect 1197 -812 1201 -748
rect 1211 -788 1215 -784
rect 1228 -788 1232 -784
rect 1219 -799 1223 -796
rect 1219 -803 1234 -799
rect 1197 -816 1212 -812
rect 870 -872 874 -868
rect 862 -1022 866 -1018
rect 879 -1022 883 -1018
rect 899 -1022 903 -1018
rect 920 -1022 924 -1018
rect 941 -1022 945 -1018
rect 962 -1022 966 -1018
rect 983 -1022 987 -1018
rect 1004 -1022 1008 -1018
rect 1025 -1022 1029 -1018
rect 1045 -1022 1049 -1018
rect 853 -1077 857 -1030
rect 853 -1098 857 -1081
rect 871 -1091 875 -1030
rect 887 -1091 891 -1030
rect 911 -1070 915 -1030
rect 911 -1091 915 -1074
rect 929 -1091 933 -1030
rect 953 -1077 957 -1030
rect 953 -1091 957 -1081
rect 971 -1070 975 -1030
rect 971 -1091 975 -1074
rect 995 -1084 999 -1030
rect 1013 -1062 1017 -1030
rect 1013 -1070 1017 -1066
rect 995 -1091 999 -1088
rect 871 -1095 880 -1091
rect 887 -1095 895 -1091
rect 871 -1098 875 -1095
rect 895 -1098 899 -1095
rect 903 -1095 915 -1091
rect 929 -1095 937 -1091
rect 903 -1098 907 -1095
rect 937 -1098 941 -1095
rect 945 -1095 957 -1091
rect 971 -1095 983 -1091
rect 945 -1098 949 -1095
rect 979 -1098 983 -1095
rect 987 -1095 999 -1091
rect 1013 -1091 1017 -1074
rect 1037 -1077 1041 -1030
rect 1037 -1091 1041 -1081
rect 1013 -1095 1025 -1091
rect 987 -1098 991 -1095
rect 1021 -1098 1025 -1095
rect 1029 -1095 1041 -1091
rect 1029 -1098 1033 -1095
rect 862 -1106 866 -1102
rect 879 -1106 883 -1102
rect 920 -1106 924 -1102
rect 962 -1106 966 -1102
rect 1004 -1106 1008 -1102
rect 1045 -1106 1049 -1102
rect 853 -1138 857 -1134
rect 870 -1138 874 -1134
rect 861 -1149 865 -1146
rect 861 -1153 876 -1149
rect 839 -1166 854 -1162
rect 504 -1425 508 -1421
rect 521 -1425 525 -1421
rect 541 -1425 545 -1421
rect 562 -1425 566 -1421
rect 583 -1425 587 -1421
rect 604 -1425 608 -1421
rect 625 -1425 629 -1421
rect 646 -1425 650 -1421
rect 667 -1425 671 -1421
rect 687 -1425 691 -1421
rect 495 -1480 499 -1433
rect 495 -1501 499 -1484
rect 513 -1494 517 -1433
rect 529 -1494 533 -1433
rect 553 -1473 557 -1433
rect 553 -1494 557 -1477
rect 571 -1494 575 -1433
rect 595 -1480 599 -1433
rect 595 -1494 599 -1484
rect 613 -1473 617 -1433
rect 613 -1494 617 -1477
rect 637 -1487 641 -1433
rect 655 -1465 659 -1433
rect 655 -1473 659 -1469
rect 637 -1494 641 -1491
rect 513 -1498 522 -1494
rect 529 -1498 537 -1494
rect 513 -1501 517 -1498
rect 537 -1501 541 -1498
rect 545 -1498 557 -1494
rect 571 -1498 579 -1494
rect 545 -1501 549 -1498
rect 579 -1501 583 -1498
rect 587 -1498 599 -1494
rect 613 -1498 625 -1494
rect 587 -1501 591 -1498
rect 621 -1501 625 -1498
rect 629 -1498 641 -1494
rect 655 -1494 659 -1477
rect 679 -1480 683 -1433
rect 679 -1494 683 -1484
rect 655 -1498 667 -1494
rect 629 -1501 633 -1498
rect 663 -1501 667 -1498
rect 671 -1498 683 -1494
rect 671 -1501 675 -1498
rect 504 -1509 508 -1505
rect 521 -1509 525 -1505
rect 562 -1509 566 -1505
rect 604 -1509 608 -1505
rect 646 -1509 650 -1505
rect 687 -1509 691 -1505
rect 504 -1596 508 -1592
rect 521 -1596 525 -1592
rect 541 -1596 545 -1592
rect 562 -1596 566 -1592
rect 583 -1596 587 -1592
rect 604 -1596 608 -1592
rect 625 -1596 629 -1592
rect 646 -1596 650 -1592
rect 667 -1596 671 -1592
rect 687 -1596 691 -1592
rect 495 -1651 499 -1604
rect 495 -1672 499 -1655
rect 513 -1665 517 -1604
rect 529 -1665 533 -1604
rect 553 -1644 557 -1604
rect 553 -1665 557 -1648
rect 571 -1665 575 -1604
rect 595 -1651 599 -1604
rect 595 -1665 599 -1655
rect 613 -1644 617 -1604
rect 613 -1665 617 -1648
rect 637 -1658 641 -1604
rect 655 -1636 659 -1604
rect 655 -1644 659 -1640
rect 637 -1665 641 -1662
rect 513 -1669 522 -1665
rect 529 -1669 537 -1665
rect 513 -1672 517 -1669
rect 537 -1672 541 -1669
rect 545 -1669 557 -1665
rect 571 -1669 579 -1665
rect 545 -1672 549 -1669
rect 579 -1672 583 -1669
rect 587 -1669 599 -1665
rect 613 -1669 625 -1665
rect 587 -1672 591 -1669
rect 621 -1672 625 -1669
rect 629 -1669 641 -1665
rect 655 -1665 659 -1648
rect 679 -1651 683 -1604
rect 679 -1665 683 -1655
rect 655 -1669 667 -1665
rect 629 -1672 633 -1669
rect 663 -1672 667 -1669
rect 671 -1669 683 -1665
rect 671 -1672 675 -1669
rect 504 -1680 508 -1676
rect 521 -1680 525 -1676
rect 562 -1680 566 -1676
rect 604 -1680 608 -1676
rect 646 -1680 650 -1676
rect 687 -1680 691 -1676
rect 704 -1687 708 -1640
rect 823 -1644 827 -1411
rect 504 -1767 508 -1763
rect 521 -1767 525 -1763
rect 541 -1767 545 -1763
rect 562 -1767 566 -1763
rect 583 -1767 587 -1763
rect 604 -1767 608 -1763
rect 625 -1767 629 -1763
rect 646 -1767 650 -1763
rect 667 -1767 671 -1763
rect 687 -1767 691 -1763
rect 495 -1822 499 -1775
rect 495 -1843 499 -1826
rect 513 -1836 517 -1775
rect 529 -1836 533 -1775
rect 553 -1815 557 -1775
rect 553 -1836 557 -1819
rect 571 -1836 575 -1775
rect 595 -1822 599 -1775
rect 595 -1836 599 -1826
rect 613 -1815 617 -1775
rect 613 -1836 617 -1819
rect 637 -1829 641 -1775
rect 655 -1807 659 -1775
rect 655 -1815 659 -1811
rect 637 -1836 641 -1833
rect 513 -1840 522 -1836
rect 529 -1840 537 -1836
rect 513 -1843 517 -1840
rect 537 -1843 541 -1840
rect 545 -1840 557 -1836
rect 571 -1840 579 -1836
rect 545 -1843 549 -1840
rect 579 -1843 583 -1840
rect 587 -1840 599 -1836
rect 613 -1840 625 -1836
rect 587 -1843 591 -1840
rect 621 -1843 625 -1840
rect 629 -1840 641 -1836
rect 655 -1836 659 -1819
rect 679 -1822 683 -1775
rect 679 -1836 683 -1826
rect 655 -1840 667 -1836
rect 629 -1843 633 -1840
rect 663 -1843 667 -1840
rect 671 -1840 683 -1836
rect 671 -1843 675 -1840
rect 504 -1851 508 -1847
rect 521 -1851 525 -1847
rect 562 -1851 566 -1847
rect 604 -1851 608 -1847
rect 646 -1851 650 -1847
rect 687 -1851 691 -1847
rect 495 -1874 499 -1870
rect 512 -1874 516 -1870
rect 503 -1885 507 -1882
rect 503 -1889 518 -1885
rect 481 -1902 496 -1898
rect 148 -2177 152 -2173
rect 165 -2177 169 -2173
rect 185 -2177 189 -2173
rect 206 -2177 210 -2173
rect 227 -2177 231 -2173
rect 248 -2177 252 -2173
rect 269 -2177 273 -2173
rect 290 -2177 294 -2173
rect 311 -2177 315 -2173
rect 331 -2177 335 -2173
rect 139 -2232 143 -2185
rect 139 -2253 143 -2236
rect 157 -2246 161 -2185
rect 173 -2246 177 -2185
rect 197 -2225 201 -2185
rect 197 -2246 201 -2229
rect 215 -2246 219 -2185
rect 239 -2232 243 -2185
rect 239 -2246 243 -2236
rect 257 -2225 261 -2185
rect 257 -2246 261 -2229
rect 281 -2239 285 -2185
rect 299 -2217 303 -2185
rect 299 -2225 303 -2221
rect 281 -2246 285 -2243
rect 157 -2250 166 -2246
rect 173 -2250 181 -2246
rect 157 -2253 161 -2250
rect 181 -2253 185 -2250
rect 189 -2250 201 -2246
rect 215 -2250 223 -2246
rect 189 -2253 193 -2250
rect 223 -2253 227 -2250
rect 231 -2250 243 -2246
rect 257 -2250 269 -2246
rect 231 -2253 235 -2250
rect 265 -2253 269 -2250
rect 273 -2250 285 -2246
rect 299 -2246 303 -2229
rect 323 -2232 327 -2185
rect 323 -2246 327 -2236
rect 299 -2250 311 -2246
rect 273 -2253 277 -2250
rect 307 -2253 311 -2250
rect 315 -2250 327 -2246
rect 315 -2253 319 -2250
rect 148 -2261 152 -2257
rect 165 -2261 169 -2257
rect 206 -2261 210 -2257
rect 248 -2261 252 -2257
rect 290 -2261 294 -2257
rect 331 -2261 335 -2257
rect 148 -2348 152 -2344
rect 165 -2348 169 -2344
rect 185 -2348 189 -2344
rect 206 -2348 210 -2344
rect 227 -2348 231 -2344
rect 248 -2348 252 -2344
rect 269 -2348 273 -2344
rect 290 -2348 294 -2344
rect 311 -2348 315 -2344
rect 331 -2348 335 -2344
rect 139 -2403 143 -2356
rect 139 -2424 143 -2407
rect 157 -2417 161 -2356
rect 173 -2417 177 -2356
rect 197 -2396 201 -2356
rect 197 -2417 201 -2400
rect 215 -2417 219 -2356
rect 239 -2403 243 -2356
rect 239 -2417 243 -2407
rect 257 -2396 261 -2356
rect 257 -2417 261 -2400
rect 281 -2410 285 -2356
rect 299 -2388 303 -2356
rect 299 -2396 303 -2392
rect 281 -2417 285 -2414
rect 157 -2421 166 -2417
rect 173 -2421 181 -2417
rect 157 -2424 161 -2421
rect 181 -2424 185 -2421
rect 189 -2421 201 -2417
rect 215 -2421 223 -2417
rect 189 -2424 193 -2421
rect 223 -2424 227 -2421
rect 231 -2421 243 -2417
rect 257 -2421 269 -2417
rect 231 -2424 235 -2421
rect 265 -2424 269 -2421
rect 273 -2421 285 -2417
rect 299 -2417 303 -2400
rect 323 -2403 327 -2356
rect 323 -2417 327 -2407
rect 299 -2421 311 -2417
rect 273 -2424 277 -2421
rect 307 -2424 311 -2421
rect 315 -2421 327 -2417
rect 315 -2424 319 -2421
rect 148 -2432 152 -2428
rect 165 -2432 169 -2428
rect 206 -2432 210 -2428
rect 248 -2432 252 -2428
rect 290 -2432 294 -2428
rect 331 -2432 335 -2428
rect 346 -2439 350 -2392
rect 465 -2396 469 -2135
rect 148 -2519 152 -2515
rect 165 -2519 169 -2515
rect 185 -2519 189 -2515
rect 206 -2519 210 -2515
rect 227 -2519 231 -2515
rect 248 -2519 252 -2515
rect 269 -2519 273 -2515
rect 290 -2519 294 -2515
rect 311 -2519 315 -2515
rect 331 -2519 335 -2515
rect 139 -2574 143 -2527
rect 139 -2595 143 -2578
rect 157 -2588 161 -2527
rect 173 -2588 177 -2527
rect 197 -2567 201 -2527
rect 197 -2588 201 -2571
rect 215 -2588 219 -2527
rect 239 -2574 243 -2527
rect 239 -2588 243 -2578
rect 257 -2567 261 -2527
rect 257 -2588 261 -2571
rect 281 -2581 285 -2527
rect 299 -2559 303 -2527
rect 299 -2567 303 -2563
rect 281 -2588 285 -2585
rect 157 -2592 166 -2588
rect 173 -2592 181 -2588
rect 157 -2595 161 -2592
rect 181 -2595 185 -2592
rect 189 -2592 201 -2588
rect 215 -2592 223 -2588
rect 189 -2595 193 -2592
rect 223 -2595 227 -2592
rect 231 -2592 243 -2588
rect 257 -2592 269 -2588
rect 231 -2595 235 -2592
rect 265 -2595 269 -2592
rect 273 -2592 285 -2588
rect 299 -2588 303 -2571
rect 323 -2574 327 -2527
rect 323 -2588 327 -2578
rect 299 -2592 311 -2588
rect 273 -2595 277 -2592
rect 307 -2595 311 -2592
rect 315 -2592 327 -2588
rect 315 -2595 319 -2592
rect 148 -2603 152 -2599
rect 165 -2603 169 -2599
rect 206 -2603 210 -2599
rect 248 -2603 252 -2599
rect 290 -2603 294 -2599
rect 331 -2603 335 -2599
rect 139 -2624 143 -2620
rect 156 -2624 160 -2620
rect 147 -2635 151 -2632
rect 147 -2639 162 -2635
rect 125 -2652 140 -2648
rect -210 -2902 -206 -2898
rect -193 -2902 -189 -2898
rect -173 -2902 -169 -2898
rect -152 -2902 -148 -2898
rect -131 -2902 -127 -2898
rect -110 -2902 -106 -2898
rect -89 -2902 -85 -2898
rect -68 -2902 -64 -2898
rect -47 -2902 -43 -2898
rect -27 -2902 -23 -2898
rect -219 -2957 -215 -2910
rect -219 -2978 -215 -2961
rect -201 -2971 -197 -2910
rect -185 -2971 -181 -2910
rect -161 -2950 -157 -2910
rect -161 -2971 -157 -2954
rect -143 -2971 -139 -2910
rect -119 -2957 -115 -2910
rect -119 -2971 -115 -2961
rect -101 -2950 -97 -2910
rect -101 -2971 -97 -2954
rect -77 -2964 -73 -2910
rect -59 -2942 -55 -2910
rect -59 -2950 -55 -2946
rect -77 -2971 -73 -2968
rect -201 -2975 -192 -2971
rect -185 -2975 -177 -2971
rect -201 -2978 -197 -2975
rect -177 -2978 -173 -2975
rect -169 -2975 -157 -2971
rect -143 -2975 -135 -2971
rect -169 -2978 -165 -2975
rect -135 -2978 -131 -2975
rect -127 -2975 -115 -2971
rect -101 -2975 -89 -2971
rect -127 -2978 -123 -2975
rect -93 -2978 -89 -2975
rect -85 -2975 -73 -2971
rect -59 -2971 -55 -2954
rect -35 -2957 -31 -2910
rect -35 -2971 -31 -2961
rect -59 -2975 -47 -2971
rect -85 -2978 -81 -2975
rect -51 -2978 -47 -2975
rect -43 -2975 -31 -2971
rect -43 -2978 -39 -2975
rect -210 -2986 -206 -2982
rect -193 -2986 -189 -2982
rect -152 -2986 -148 -2982
rect -110 -2986 -106 -2982
rect -68 -2986 -64 -2982
rect -27 -2986 -23 -2982
rect -210 -3073 -206 -3069
rect -193 -3073 -189 -3069
rect -173 -3073 -169 -3069
rect -152 -3073 -148 -3069
rect -131 -3073 -127 -3069
rect -110 -3073 -106 -3069
rect -89 -3073 -85 -3069
rect -68 -3073 -64 -3069
rect -47 -3073 -43 -3069
rect -27 -3073 -23 -3069
rect -219 -3128 -215 -3081
rect -219 -3149 -215 -3132
rect -201 -3142 -197 -3081
rect -185 -3142 -181 -3081
rect -161 -3121 -157 -3081
rect -161 -3142 -157 -3125
rect -143 -3142 -139 -3081
rect -119 -3128 -115 -3081
rect -119 -3142 -115 -3132
rect -101 -3121 -97 -3081
rect -101 -3142 -97 -3125
rect -77 -3135 -73 -3081
rect -59 -3113 -55 -3081
rect -59 -3121 -55 -3117
rect -77 -3142 -73 -3139
rect -201 -3146 -192 -3142
rect -185 -3146 -177 -3142
rect -201 -3149 -197 -3146
rect -177 -3149 -173 -3146
rect -169 -3146 -157 -3142
rect -143 -3146 -135 -3142
rect -169 -3149 -165 -3146
rect -135 -3149 -131 -3146
rect -127 -3146 -115 -3142
rect -101 -3146 -89 -3142
rect -127 -3149 -123 -3146
rect -93 -3149 -89 -3146
rect -85 -3146 -73 -3142
rect -59 -3142 -55 -3125
rect -35 -3128 -31 -3081
rect -35 -3142 -31 -3132
rect -59 -3146 -47 -3142
rect -85 -3149 -81 -3146
rect -51 -3149 -47 -3146
rect -43 -3146 -31 -3142
rect -43 -3149 -39 -3146
rect -210 -3157 -206 -3153
rect -193 -3157 -189 -3153
rect -152 -3157 -148 -3153
rect -110 -3157 -106 -3153
rect -68 -3157 -64 -3153
rect -27 -3157 -23 -3153
rect -13 -3165 -9 -3117
rect 111 -3121 115 -2878
rect -210 -3244 -206 -3240
rect -193 -3244 -189 -3240
rect -173 -3244 -169 -3240
rect -152 -3244 -148 -3240
rect -131 -3244 -127 -3240
rect -110 -3244 -106 -3240
rect -89 -3244 -85 -3240
rect -68 -3244 -64 -3240
rect -47 -3244 -43 -3240
rect -27 -3244 -23 -3240
rect -219 -3299 -215 -3252
rect -219 -3320 -215 -3303
rect -201 -3313 -197 -3252
rect -185 -3313 -181 -3252
rect -161 -3292 -157 -3252
rect -161 -3313 -157 -3296
rect -143 -3313 -139 -3252
rect -119 -3299 -115 -3252
rect -119 -3313 -115 -3303
rect -101 -3292 -97 -3252
rect -101 -3313 -97 -3296
rect -77 -3306 -73 -3252
rect -59 -3284 -55 -3252
rect -59 -3292 -55 -3288
rect -77 -3313 -73 -3310
rect -201 -3317 -192 -3313
rect -185 -3317 -177 -3313
rect -201 -3320 -197 -3317
rect -177 -3320 -173 -3317
rect -169 -3317 -157 -3313
rect -143 -3317 -135 -3313
rect -169 -3320 -165 -3317
rect -135 -3320 -131 -3317
rect -127 -3317 -115 -3313
rect -101 -3317 -89 -3313
rect -127 -3320 -123 -3317
rect -93 -3320 -89 -3317
rect -85 -3317 -73 -3313
rect -59 -3313 -55 -3296
rect -35 -3299 -31 -3252
rect -35 -3313 -31 -3303
rect -59 -3317 -47 -3313
rect -85 -3320 -81 -3317
rect -51 -3320 -47 -3317
rect -43 -3317 -31 -3313
rect -43 -3320 -39 -3317
rect -210 -3328 -206 -3324
rect -193 -3328 -189 -3324
rect -152 -3328 -148 -3324
rect -110 -3328 -106 -3324
rect -68 -3328 -64 -3324
rect -27 -3328 -23 -3324
rect -219 -3355 -215 -3351
rect -202 -3355 -198 -3351
rect -211 -3366 -207 -3363
rect -211 -3370 -196 -3366
rect -233 -3383 -218 -3379
rect -568 -3644 -564 -3640
rect -551 -3644 -547 -3640
rect -531 -3644 -527 -3640
rect -510 -3644 -506 -3640
rect -489 -3644 -485 -3640
rect -468 -3644 -464 -3640
rect -447 -3644 -443 -3640
rect -426 -3644 -422 -3640
rect -405 -3644 -401 -3640
rect -385 -3644 -381 -3640
rect -577 -3699 -573 -3652
rect -577 -3720 -573 -3703
rect -559 -3713 -555 -3652
rect -543 -3713 -539 -3652
rect -519 -3692 -515 -3652
rect -519 -3713 -515 -3696
rect -501 -3713 -497 -3652
rect -477 -3699 -473 -3652
rect -477 -3713 -473 -3703
rect -459 -3692 -455 -3652
rect -459 -3713 -455 -3696
rect -435 -3706 -431 -3652
rect -417 -3684 -413 -3652
rect -417 -3692 -413 -3688
rect -435 -3713 -431 -3710
rect -559 -3717 -550 -3713
rect -543 -3717 -535 -3713
rect -559 -3720 -555 -3717
rect -535 -3720 -531 -3717
rect -527 -3717 -515 -3713
rect -501 -3717 -493 -3713
rect -527 -3720 -523 -3717
rect -493 -3720 -489 -3717
rect -485 -3717 -473 -3713
rect -459 -3717 -447 -3713
rect -485 -3720 -481 -3717
rect -451 -3720 -447 -3717
rect -443 -3717 -431 -3713
rect -417 -3713 -413 -3696
rect -393 -3699 -389 -3652
rect -393 -3713 -389 -3703
rect -417 -3717 -405 -3713
rect -443 -3720 -439 -3717
rect -409 -3720 -405 -3717
rect -401 -3717 -389 -3713
rect -401 -3720 -397 -3717
rect -568 -3728 -564 -3724
rect -551 -3728 -547 -3724
rect -510 -3728 -506 -3724
rect -468 -3728 -464 -3724
rect -426 -3728 -422 -3724
rect -385 -3728 -381 -3724
rect -568 -3815 -564 -3811
rect -551 -3815 -547 -3811
rect -531 -3815 -527 -3811
rect -510 -3815 -506 -3811
rect -489 -3815 -485 -3811
rect -468 -3815 -464 -3811
rect -447 -3815 -443 -3811
rect -426 -3815 -422 -3811
rect -405 -3815 -401 -3811
rect -385 -3815 -381 -3811
rect -577 -3870 -573 -3823
rect -577 -3891 -573 -3874
rect -559 -3884 -555 -3823
rect -543 -3884 -539 -3823
rect -519 -3863 -515 -3823
rect -519 -3884 -515 -3867
rect -501 -3884 -497 -3823
rect -477 -3870 -473 -3823
rect -477 -3884 -473 -3874
rect -459 -3863 -455 -3823
rect -459 -3884 -455 -3867
rect -435 -3877 -431 -3823
rect -417 -3855 -413 -3823
rect -417 -3863 -413 -3859
rect -435 -3884 -431 -3881
rect -559 -3888 -550 -3884
rect -543 -3888 -535 -3884
rect -559 -3891 -555 -3888
rect -535 -3891 -531 -3888
rect -527 -3888 -515 -3884
rect -501 -3888 -493 -3884
rect -527 -3891 -523 -3888
rect -493 -3891 -489 -3888
rect -485 -3888 -473 -3884
rect -459 -3888 -447 -3884
rect -485 -3891 -481 -3888
rect -451 -3891 -447 -3888
rect -443 -3888 -431 -3884
rect -417 -3884 -413 -3867
rect -393 -3870 -389 -3823
rect -393 -3884 -389 -3874
rect -417 -3888 -405 -3884
rect -443 -3891 -439 -3888
rect -409 -3891 -405 -3888
rect -401 -3888 -389 -3884
rect -401 -3891 -397 -3888
rect -568 -3899 -564 -3895
rect -551 -3899 -547 -3895
rect -510 -3899 -506 -3895
rect -468 -3899 -464 -3895
rect -426 -3899 -422 -3895
rect -385 -3899 -381 -3895
rect -369 -3906 -365 -3859
rect -249 -3863 -245 -3616
rect -568 -3990 -564 -3986
rect -551 -3990 -547 -3986
rect -531 -3990 -527 -3986
rect -510 -3990 -506 -3986
rect -489 -3990 -485 -3986
rect -468 -3990 -464 -3986
rect -447 -3990 -443 -3986
rect -426 -3990 -422 -3986
rect -405 -3990 -401 -3986
rect -385 -3990 -381 -3986
rect -577 -4045 -573 -3998
rect -577 -4066 -573 -4049
rect -559 -4059 -555 -3998
rect -543 -4059 -539 -3998
rect -519 -4038 -515 -3998
rect -519 -4059 -515 -4042
rect -501 -4059 -497 -3998
rect -477 -4045 -473 -3998
rect -477 -4059 -473 -4049
rect -459 -4038 -455 -3998
rect -459 -4059 -455 -4042
rect -435 -4052 -431 -3998
rect -417 -4030 -413 -3998
rect -417 -4038 -413 -4034
rect -435 -4059 -431 -4056
rect -559 -4063 -550 -4059
rect -543 -4063 -535 -4059
rect -559 -4066 -555 -4063
rect -535 -4066 -531 -4063
rect -527 -4063 -515 -4059
rect -501 -4063 -493 -4059
rect -527 -4066 -523 -4063
rect -493 -4066 -489 -4063
rect -485 -4063 -473 -4059
rect -459 -4063 -447 -4059
rect -485 -4066 -481 -4063
rect -451 -4066 -447 -4063
rect -443 -4063 -431 -4059
rect -417 -4059 -413 -4042
rect -393 -4045 -389 -3998
rect -393 -4059 -389 -4049
rect -417 -4063 -405 -4059
rect -443 -4066 -439 -4063
rect -409 -4066 -405 -4063
rect -401 -4063 -389 -4059
rect -401 -4066 -397 -4063
rect -568 -4074 -564 -4070
rect -551 -4074 -547 -4070
rect -510 -4074 -506 -4070
rect -468 -4074 -464 -4070
rect -426 -4074 -422 -4070
rect -385 -4074 -381 -4070
rect -577 -4105 -573 -4101
rect -560 -4105 -556 -4101
rect -569 -4116 -565 -4113
rect -569 -4120 -554 -4116
rect -591 -4133 -576 -4129
rect -926 -4387 -922 -4383
rect -909 -4387 -905 -4383
rect -889 -4387 -885 -4383
rect -868 -4387 -864 -4383
rect -847 -4387 -843 -4383
rect -826 -4387 -822 -4383
rect -805 -4387 -801 -4383
rect -784 -4387 -780 -4383
rect -763 -4387 -759 -4383
rect -743 -4387 -739 -4383
rect -935 -4442 -931 -4395
rect -935 -4463 -931 -4446
rect -917 -4456 -913 -4395
rect -901 -4456 -897 -4395
rect -877 -4435 -873 -4395
rect -877 -4456 -873 -4439
rect -859 -4456 -855 -4395
rect -835 -4442 -831 -4395
rect -835 -4456 -831 -4446
rect -817 -4435 -813 -4395
rect -817 -4456 -813 -4439
rect -793 -4449 -789 -4395
rect -775 -4427 -771 -4395
rect -775 -4435 -771 -4431
rect -793 -4456 -789 -4453
rect -917 -4460 -908 -4456
rect -901 -4460 -893 -4456
rect -917 -4463 -913 -4460
rect -893 -4463 -889 -4460
rect -885 -4460 -873 -4456
rect -859 -4460 -851 -4456
rect -885 -4463 -881 -4460
rect -851 -4463 -847 -4460
rect -843 -4460 -831 -4456
rect -817 -4460 -805 -4456
rect -843 -4463 -839 -4460
rect -809 -4463 -805 -4460
rect -801 -4460 -789 -4456
rect -775 -4456 -771 -4439
rect -751 -4442 -747 -4395
rect -751 -4456 -747 -4446
rect -775 -4460 -763 -4456
rect -801 -4463 -797 -4460
rect -767 -4463 -763 -4460
rect -759 -4460 -747 -4456
rect -759 -4463 -755 -4460
rect -926 -4471 -922 -4467
rect -909 -4471 -905 -4467
rect -868 -4471 -864 -4467
rect -826 -4471 -822 -4467
rect -784 -4471 -780 -4467
rect -743 -4471 -739 -4467
rect -926 -4558 -922 -4554
rect -909 -4558 -905 -4554
rect -889 -4558 -885 -4554
rect -868 -4558 -864 -4554
rect -847 -4558 -843 -4554
rect -826 -4558 -822 -4554
rect -805 -4558 -801 -4554
rect -784 -4558 -780 -4554
rect -763 -4558 -759 -4554
rect -743 -4558 -739 -4554
rect -935 -4613 -931 -4566
rect -935 -4634 -931 -4617
rect -917 -4627 -913 -4566
rect -901 -4627 -897 -4566
rect -877 -4606 -873 -4566
rect -877 -4627 -873 -4610
rect -859 -4627 -855 -4566
rect -835 -4613 -831 -4566
rect -835 -4627 -831 -4617
rect -817 -4606 -813 -4566
rect -817 -4627 -813 -4610
rect -793 -4620 -789 -4566
rect -775 -4598 -771 -4566
rect -775 -4606 -771 -4602
rect -793 -4627 -789 -4624
rect -917 -4631 -908 -4627
rect -901 -4631 -893 -4627
rect -917 -4634 -913 -4631
rect -893 -4634 -889 -4631
rect -885 -4631 -873 -4627
rect -859 -4631 -851 -4627
rect -885 -4634 -881 -4631
rect -851 -4634 -847 -4631
rect -843 -4631 -831 -4627
rect -817 -4631 -805 -4627
rect -843 -4634 -839 -4631
rect -809 -4634 -805 -4631
rect -801 -4631 -789 -4627
rect -775 -4627 -771 -4610
rect -751 -4613 -747 -4566
rect -751 -4627 -747 -4617
rect -775 -4631 -763 -4627
rect -801 -4634 -797 -4631
rect -767 -4634 -763 -4631
rect -759 -4631 -747 -4627
rect -759 -4634 -755 -4631
rect -926 -4642 -922 -4638
rect -909 -4642 -905 -4638
rect -868 -4642 -864 -4638
rect -826 -4642 -822 -4638
rect -784 -4642 -780 -4638
rect -743 -4642 -739 -4638
rect -729 -4649 -725 -4602
rect -603 -4606 -599 -4359
rect -926 -4729 -922 -4725
rect -909 -4729 -905 -4725
rect -889 -4729 -885 -4725
rect -868 -4729 -864 -4725
rect -847 -4729 -843 -4725
rect -826 -4729 -822 -4725
rect -805 -4729 -801 -4725
rect -784 -4729 -780 -4725
rect -763 -4729 -759 -4725
rect -743 -4729 -739 -4725
rect -935 -4784 -931 -4737
rect -935 -4805 -931 -4788
rect -917 -4798 -913 -4737
rect -901 -4798 -897 -4737
rect -877 -4777 -873 -4737
rect -877 -4798 -873 -4781
rect -859 -4798 -855 -4737
rect -835 -4784 -831 -4737
rect -835 -4798 -831 -4788
rect -817 -4777 -813 -4737
rect -817 -4798 -813 -4781
rect -793 -4791 -789 -4737
rect -775 -4769 -771 -4737
rect -775 -4777 -771 -4773
rect -793 -4798 -789 -4795
rect -917 -4802 -908 -4798
rect -901 -4802 -893 -4798
rect -917 -4805 -913 -4802
rect -893 -4805 -889 -4802
rect -885 -4802 -873 -4798
rect -859 -4802 -851 -4798
rect -885 -4805 -881 -4802
rect -851 -4805 -847 -4802
rect -843 -4802 -831 -4798
rect -817 -4802 -805 -4798
rect -843 -4805 -839 -4802
rect -809 -4805 -805 -4802
rect -801 -4802 -789 -4798
rect -775 -4798 -771 -4781
rect -751 -4784 -747 -4737
rect -751 -4798 -747 -4788
rect -775 -4802 -763 -4798
rect -801 -4805 -797 -4802
rect -767 -4805 -763 -4802
rect -759 -4802 -747 -4798
rect -759 -4805 -755 -4802
rect -926 -4813 -922 -4809
rect -909 -4813 -905 -4809
rect -868 -4813 -864 -4809
rect -826 -4813 -822 -4809
rect -784 -4813 -780 -4809
rect -743 -4813 -739 -4809
rect -935 -4844 -931 -4840
rect -918 -4844 -914 -4840
rect -927 -4855 -923 -4852
rect -927 -4859 -912 -4855
rect -949 -4872 -934 -4868
rect -1225 -5087 -1221 -5083
rect -1181 -5087 -1177 -5083
rect -1147 -5087 -1143 -5083
rect -1257 -5341 -1253 -5098
rect -1102 -5102 -1098 -5069
rect -1246 -5170 -1242 -5106
rect -1225 -5122 -1221 -5118
rect -1208 -5122 -1204 -5118
rect -1188 -5122 -1184 -5118
rect -1167 -5122 -1163 -5118
rect -1146 -5122 -1142 -5118
rect -1125 -5122 -1121 -5118
rect -1104 -5122 -1100 -5118
rect -1083 -5122 -1079 -5118
rect -1062 -5122 -1058 -5118
rect -1042 -5122 -1038 -5118
rect -1234 -5177 -1230 -5130
rect -1234 -5198 -1230 -5181
rect -1216 -5191 -1212 -5130
rect -1200 -5191 -1196 -5130
rect -1176 -5170 -1172 -5130
rect -1176 -5191 -1172 -5174
rect -1158 -5191 -1154 -5130
rect -1134 -5177 -1130 -5130
rect -1134 -5191 -1130 -5181
rect -1116 -5170 -1112 -5130
rect -1116 -5191 -1112 -5174
rect -1092 -5184 -1088 -5130
rect -1074 -5162 -1070 -5130
rect -1074 -5170 -1070 -5166
rect -1092 -5191 -1088 -5188
rect -1216 -5195 -1207 -5191
rect -1200 -5195 -1192 -5191
rect -1216 -5198 -1212 -5195
rect -1192 -5198 -1188 -5195
rect -1184 -5195 -1172 -5191
rect -1158 -5195 -1150 -5191
rect -1184 -5198 -1180 -5195
rect -1150 -5198 -1146 -5195
rect -1142 -5195 -1130 -5191
rect -1116 -5195 -1104 -5191
rect -1142 -5198 -1138 -5195
rect -1108 -5198 -1104 -5195
rect -1100 -5195 -1088 -5191
rect -1074 -5191 -1070 -5174
rect -1050 -5177 -1046 -5130
rect -1050 -5191 -1046 -5181
rect -1074 -5195 -1062 -5191
rect -1100 -5198 -1096 -5195
rect -1066 -5198 -1062 -5195
rect -1058 -5195 -1046 -5191
rect -1058 -5198 -1054 -5195
rect -1225 -5206 -1221 -5202
rect -1208 -5206 -1204 -5202
rect -1167 -5206 -1163 -5202
rect -1125 -5206 -1121 -5202
rect -1083 -5206 -1079 -5202
rect -1042 -5206 -1038 -5202
rect -1225 -5293 -1221 -5289
rect -1208 -5293 -1204 -5289
rect -1188 -5293 -1184 -5289
rect -1167 -5293 -1163 -5289
rect -1146 -5293 -1142 -5289
rect -1125 -5293 -1121 -5289
rect -1104 -5293 -1100 -5289
rect -1083 -5293 -1079 -5289
rect -1062 -5293 -1058 -5289
rect -1042 -5293 -1038 -5289
rect -1234 -5348 -1230 -5301
rect -1234 -5369 -1230 -5352
rect -1216 -5362 -1212 -5301
rect -1200 -5362 -1196 -5301
rect -1176 -5341 -1172 -5301
rect -1176 -5362 -1172 -5345
rect -1158 -5362 -1154 -5301
rect -1134 -5348 -1130 -5301
rect -1134 -5362 -1130 -5352
rect -1116 -5341 -1112 -5301
rect -1116 -5362 -1112 -5345
rect -1092 -5355 -1088 -5301
rect -1074 -5333 -1070 -5301
rect -1074 -5341 -1070 -5337
rect -1092 -5362 -1088 -5359
rect -1216 -5366 -1207 -5362
rect -1200 -5366 -1192 -5362
rect -1216 -5369 -1212 -5366
rect -1192 -5369 -1188 -5366
rect -1184 -5366 -1172 -5362
rect -1158 -5366 -1150 -5362
rect -1184 -5369 -1180 -5366
rect -1150 -5369 -1146 -5366
rect -1142 -5366 -1130 -5362
rect -1116 -5366 -1104 -5362
rect -1142 -5369 -1138 -5366
rect -1108 -5369 -1104 -5366
rect -1100 -5366 -1088 -5362
rect -1074 -5362 -1070 -5345
rect -1050 -5348 -1046 -5301
rect -1050 -5362 -1046 -5352
rect -1074 -5366 -1062 -5362
rect -1100 -5369 -1096 -5366
rect -1066 -5369 -1062 -5366
rect -1058 -5366 -1046 -5362
rect -1058 -5369 -1054 -5366
rect -1225 -5377 -1221 -5373
rect -1208 -5377 -1204 -5373
rect -1167 -5377 -1163 -5373
rect -1125 -5377 -1121 -5373
rect -1083 -5377 -1079 -5373
rect -1042 -5377 -1038 -5373
rect -1024 -5384 -1020 -5337
rect -963 -5341 -959 -5105
rect -1309 -5567 -1305 -5563
rect -1292 -5567 -1288 -5563
rect -1301 -5578 -1297 -5575
rect -1301 -5582 -1286 -5578
rect -1290 -5621 -1286 -5582
rect -1290 -5636 -1286 -5625
rect -1309 -5640 -1286 -5636
rect -1309 -5643 -1305 -5640
rect -1283 -5643 -1279 -5575
rect -1292 -5651 -1288 -5647
rect -1283 -5781 -1279 -5647
rect -1257 -5774 -1253 -5388
rect -1225 -5453 -1221 -5449
rect -1208 -5453 -1204 -5449
rect -1188 -5453 -1184 -5449
rect -1167 -5453 -1163 -5449
rect -1146 -5453 -1142 -5449
rect -1125 -5453 -1121 -5449
rect -1104 -5453 -1100 -5449
rect -1083 -5453 -1079 -5449
rect -1062 -5453 -1058 -5449
rect -1042 -5453 -1038 -5449
rect -1234 -5508 -1230 -5461
rect -1234 -5529 -1230 -5512
rect -1216 -5522 -1212 -5461
rect -1200 -5522 -1196 -5461
rect -1176 -5501 -1172 -5461
rect -1176 -5522 -1172 -5505
rect -1158 -5522 -1154 -5461
rect -1134 -5508 -1130 -5461
rect -1134 -5522 -1130 -5512
rect -1116 -5501 -1112 -5461
rect -1116 -5522 -1112 -5505
rect -1092 -5515 -1088 -5461
rect -1074 -5493 -1070 -5461
rect -1074 -5501 -1070 -5497
rect -1092 -5522 -1088 -5519
rect -1216 -5526 -1207 -5522
rect -1200 -5526 -1192 -5522
rect -1216 -5529 -1212 -5526
rect -1192 -5529 -1188 -5526
rect -1184 -5526 -1172 -5522
rect -1158 -5526 -1150 -5522
rect -1184 -5529 -1180 -5526
rect -1150 -5529 -1146 -5526
rect -1142 -5526 -1130 -5522
rect -1116 -5526 -1104 -5522
rect -1142 -5529 -1138 -5526
rect -1108 -5529 -1104 -5526
rect -1100 -5526 -1088 -5522
rect -1074 -5522 -1070 -5505
rect -1050 -5508 -1046 -5461
rect -1050 -5522 -1046 -5512
rect -1074 -5526 -1062 -5522
rect -1100 -5529 -1096 -5526
rect -1066 -5529 -1062 -5526
rect -1058 -5526 -1046 -5522
rect -1058 -5529 -1054 -5526
rect -1225 -5537 -1221 -5533
rect -1208 -5537 -1204 -5533
rect -1167 -5537 -1163 -5533
rect -1125 -5537 -1121 -5533
rect -1083 -5537 -1079 -5533
rect -1042 -5537 -1038 -5533
rect -1020 -5591 -1016 -5497
rect -1225 -5726 -1221 -5722
rect -1208 -5726 -1204 -5722
rect -1168 -5726 -1164 -5722
rect -1147 -5726 -1143 -5722
rect -1234 -5767 -1230 -5734
rect -1234 -5802 -1230 -5771
rect -1216 -5761 -1212 -5734
rect -1216 -5765 -1207 -5761
rect -1216 -5802 -1212 -5765
rect -1190 -5788 -1186 -5734
rect -1190 -5795 -1186 -5792
rect -1156 -5795 -1152 -5734
rect -1138 -5766 -1134 -5734
rect -979 -5758 -975 -5616
rect -1208 -5802 -1204 -5799
rect -1199 -5799 -1186 -5795
rect -1199 -5802 -1195 -5799
rect -1172 -5802 -1168 -5799
rect -1164 -5799 -1145 -5795
rect -1164 -5802 -1160 -5799
rect -1138 -5802 -1134 -5770
rect -963 -5773 -959 -5388
rect -949 -5501 -945 -4872
rect -916 -4898 -912 -4859
rect -916 -4913 -912 -4902
rect -935 -4917 -912 -4913
rect -909 -4889 -905 -4852
rect -722 -4868 -718 -4773
rect -935 -4920 -931 -4917
rect -909 -4920 -905 -4893
rect -918 -4928 -914 -4924
rect -926 -5003 -922 -4999
rect -900 -5003 -896 -4999
rect -883 -5003 -879 -4999
rect -843 -5003 -839 -4999
rect -822 -5003 -818 -4999
rect -805 -5003 -801 -4999
rect -765 -5003 -761 -4999
rect -741 -5003 -737 -4999
rect -704 -5003 -700 -4999
rect -935 -5028 -931 -5011
rect -935 -5079 -931 -5032
rect -917 -5021 -913 -5011
rect -917 -5079 -913 -5025
rect -909 -5050 -905 -5011
rect -891 -5043 -887 -5011
rect -909 -5079 -905 -5054
rect -891 -5079 -887 -5047
rect -865 -5035 -861 -5011
rect -865 -5072 -861 -5039
rect -831 -5072 -827 -5011
rect -813 -5028 -809 -5011
rect -883 -5079 -879 -5076
rect -875 -5076 -861 -5072
rect -875 -5079 -871 -5076
rect -847 -5079 -843 -5076
rect -839 -5076 -820 -5072
rect -839 -5079 -835 -5076
rect -813 -5079 -809 -5032
rect -787 -5043 -783 -5011
rect -787 -5072 -783 -5047
rect -753 -5065 -749 -5011
rect -753 -5069 -736 -5065
rect -805 -5079 -801 -5076
rect -796 -5076 -783 -5072
rect -796 -5079 -792 -5076
rect -769 -5079 -765 -5076
rect -745 -5079 -741 -5069
rect -729 -5072 -725 -5011
rect -721 -5065 -717 -5011
rect -695 -5035 -691 -5011
rect -721 -5069 -702 -5065
rect -737 -5076 -720 -5072
rect -737 -5079 -733 -5076
rect -713 -5079 -709 -5069
rect -695 -5079 -691 -5039
rect -926 -5087 -922 -5083
rect -900 -5087 -896 -5083
rect -857 -5087 -853 -5083
rect -822 -5087 -818 -5083
rect -778 -5087 -774 -5083
rect -761 -5087 -757 -5083
rect -725 -5087 -721 -5083
rect -704 -5087 -700 -5083
rect -687 -5094 -683 -5047
rect -616 -5050 -612 -4893
rect -603 -5035 -599 -4653
rect -591 -4777 -587 -4133
rect -558 -4159 -554 -4120
rect -558 -4174 -554 -4163
rect -577 -4178 -554 -4174
rect -551 -4150 -547 -4113
rect -369 -4129 -365 -4034
rect -577 -4181 -573 -4178
rect -551 -4181 -547 -4154
rect -560 -4189 -556 -4185
rect -568 -4264 -564 -4260
rect -542 -4264 -538 -4260
rect -525 -4264 -521 -4260
rect -485 -4264 -481 -4260
rect -464 -4264 -460 -4260
rect -447 -4264 -443 -4260
rect -407 -4264 -403 -4260
rect -383 -4264 -379 -4260
rect -346 -4264 -342 -4260
rect -577 -4289 -573 -4272
rect -577 -4340 -573 -4293
rect -559 -4282 -555 -4272
rect -559 -4340 -555 -4286
rect -551 -4311 -547 -4272
rect -533 -4304 -529 -4272
rect -551 -4340 -547 -4315
rect -533 -4340 -529 -4308
rect -507 -4296 -503 -4272
rect -507 -4333 -503 -4300
rect -473 -4333 -469 -4272
rect -455 -4289 -451 -4272
rect -525 -4340 -521 -4337
rect -517 -4337 -503 -4333
rect -517 -4340 -513 -4337
rect -489 -4340 -485 -4337
rect -481 -4337 -462 -4333
rect -481 -4340 -477 -4337
rect -455 -4340 -451 -4293
rect -429 -4304 -425 -4272
rect -429 -4333 -425 -4308
rect -395 -4326 -391 -4272
rect -395 -4330 -378 -4326
rect -447 -4340 -443 -4337
rect -438 -4337 -425 -4333
rect -438 -4340 -434 -4337
rect -411 -4340 -407 -4337
rect -387 -4340 -383 -4330
rect -371 -4333 -367 -4272
rect -363 -4326 -359 -4272
rect -337 -4295 -333 -4272
rect -363 -4330 -344 -4326
rect -379 -4337 -362 -4333
rect -379 -4340 -375 -4337
rect -355 -4340 -351 -4330
rect -337 -4340 -333 -4299
rect -568 -4348 -564 -4344
rect -542 -4348 -538 -4344
rect -499 -4348 -495 -4344
rect -464 -4348 -460 -4344
rect -420 -4348 -416 -4344
rect -403 -4348 -399 -4344
rect -367 -4348 -363 -4344
rect -346 -4348 -342 -4344
rect -328 -4362 -324 -4308
rect -263 -4311 -259 -4154
rect -249 -4296 -245 -3910
rect -233 -4038 -229 -3383
rect -200 -3409 -196 -3370
rect -200 -3424 -196 -3413
rect -219 -3428 -196 -3424
rect -193 -3400 -189 -3363
rect -13 -3379 -9 -3288
rect -219 -3431 -215 -3428
rect -193 -3431 -189 -3404
rect -202 -3439 -198 -3435
rect -210 -3514 -206 -3510
rect -184 -3514 -180 -3510
rect -167 -3514 -163 -3510
rect -127 -3514 -123 -3510
rect -106 -3514 -102 -3510
rect -89 -3514 -85 -3510
rect -49 -3514 -45 -3510
rect -25 -3514 -21 -3510
rect 12 -3514 16 -3510
rect -219 -3539 -215 -3522
rect -219 -3590 -215 -3543
rect -201 -3532 -197 -3522
rect -201 -3590 -197 -3536
rect -193 -3561 -189 -3522
rect -175 -3554 -171 -3522
rect -193 -3590 -189 -3565
rect -175 -3590 -171 -3558
rect -149 -3546 -145 -3522
rect -149 -3583 -145 -3550
rect -115 -3583 -111 -3522
rect -97 -3539 -93 -3522
rect -167 -3590 -163 -3587
rect -159 -3587 -145 -3583
rect -159 -3590 -155 -3587
rect -131 -3590 -127 -3587
rect -123 -3587 -104 -3583
rect -123 -3590 -119 -3587
rect -97 -3590 -93 -3543
rect -71 -3554 -67 -3522
rect -71 -3583 -67 -3558
rect -37 -3576 -33 -3522
rect -37 -3580 -20 -3576
rect -89 -3590 -85 -3587
rect -80 -3587 -67 -3583
rect -80 -3590 -76 -3587
rect -53 -3590 -49 -3587
rect -29 -3590 -25 -3580
rect -13 -3583 -9 -3522
rect -5 -3576 -1 -3522
rect 21 -3546 25 -3522
rect -5 -3580 14 -3576
rect -21 -3587 -4 -3583
rect -21 -3590 -17 -3587
rect 3 -3590 7 -3580
rect 21 -3590 25 -3550
rect -210 -3598 -206 -3594
rect -184 -3598 -180 -3594
rect -141 -3598 -137 -3594
rect -106 -3598 -102 -3594
rect -62 -3598 -58 -3594
rect -45 -3598 -41 -3594
rect -9 -3598 -5 -3594
rect 12 -3598 16 -3594
rect 29 -3605 33 -3558
rect 97 -3561 101 -3404
rect 111 -3546 115 -3168
rect 125 -3292 129 -2652
rect 158 -2678 162 -2639
rect 158 -2693 162 -2682
rect 139 -2697 162 -2693
rect 165 -2669 169 -2632
rect 347 -2648 351 -2563
rect 139 -2700 143 -2697
rect 165 -2700 169 -2673
rect 156 -2708 160 -2704
rect 148 -2783 152 -2779
rect 174 -2783 178 -2779
rect 191 -2783 195 -2779
rect 231 -2783 235 -2779
rect 252 -2783 256 -2779
rect 269 -2783 273 -2779
rect 309 -2783 313 -2779
rect 333 -2783 337 -2779
rect 370 -2783 374 -2779
rect 139 -2808 143 -2791
rect 139 -2859 143 -2812
rect 157 -2801 161 -2791
rect 157 -2859 161 -2805
rect 165 -2830 169 -2791
rect 183 -2823 187 -2791
rect 165 -2859 169 -2834
rect 183 -2859 187 -2827
rect 209 -2815 213 -2791
rect 209 -2852 213 -2819
rect 243 -2852 247 -2791
rect 261 -2808 265 -2791
rect 191 -2859 195 -2856
rect 199 -2856 213 -2852
rect 199 -2859 203 -2856
rect 227 -2859 231 -2856
rect 235 -2856 254 -2852
rect 235 -2859 239 -2856
rect 261 -2859 265 -2812
rect 287 -2823 291 -2791
rect 287 -2852 291 -2827
rect 321 -2845 325 -2791
rect 321 -2849 338 -2845
rect 269 -2859 273 -2856
rect 278 -2856 291 -2852
rect 278 -2859 282 -2856
rect 305 -2859 309 -2856
rect 329 -2859 333 -2849
rect 345 -2852 349 -2791
rect 353 -2845 357 -2791
rect 379 -2815 383 -2791
rect 353 -2849 372 -2845
rect 337 -2856 354 -2852
rect 337 -2859 341 -2856
rect 361 -2859 365 -2849
rect 379 -2859 383 -2819
rect 148 -2867 152 -2863
rect 174 -2867 178 -2863
rect 217 -2867 221 -2863
rect 252 -2867 256 -2863
rect 296 -2867 300 -2863
rect 313 -2867 317 -2863
rect 349 -2867 353 -2863
rect 370 -2867 374 -2863
rect 389 -2881 393 -2827
rect 451 -2830 455 -2673
rect 465 -2815 469 -2443
rect 481 -2567 485 -1902
rect 514 -1928 518 -1889
rect 514 -1943 518 -1932
rect 495 -1947 518 -1943
rect 521 -1919 525 -1882
rect 703 -1898 707 -1811
rect 495 -1950 499 -1947
rect 521 -1950 525 -1923
rect 512 -1958 516 -1954
rect 504 -2033 508 -2029
rect 530 -2033 534 -2029
rect 547 -2033 551 -2029
rect 587 -2033 591 -2029
rect 608 -2033 612 -2029
rect 625 -2033 629 -2029
rect 665 -2033 669 -2029
rect 689 -2033 693 -2029
rect 726 -2033 730 -2029
rect 495 -2058 499 -2041
rect 495 -2109 499 -2062
rect 513 -2051 517 -2041
rect 513 -2109 517 -2055
rect 521 -2080 525 -2041
rect 539 -2073 543 -2041
rect 521 -2109 525 -2084
rect 539 -2109 543 -2077
rect 565 -2065 569 -2041
rect 565 -2102 569 -2069
rect 599 -2102 603 -2041
rect 617 -2058 621 -2041
rect 547 -2109 551 -2106
rect 555 -2106 569 -2102
rect 555 -2109 559 -2106
rect 583 -2109 587 -2106
rect 591 -2106 610 -2102
rect 591 -2109 595 -2106
rect 617 -2109 621 -2062
rect 643 -2073 647 -2041
rect 643 -2102 647 -2077
rect 677 -2095 681 -2041
rect 677 -2099 694 -2095
rect 625 -2109 629 -2106
rect 634 -2106 647 -2102
rect 634 -2109 638 -2106
rect 661 -2109 665 -2106
rect 685 -2109 689 -2099
rect 701 -2102 705 -2041
rect 709 -2095 713 -2041
rect 735 -2065 739 -2041
rect 709 -2099 728 -2095
rect 693 -2106 710 -2102
rect 693 -2109 697 -2106
rect 717 -2109 721 -2099
rect 735 -2109 739 -2069
rect 504 -2117 508 -2113
rect 530 -2117 534 -2113
rect 573 -2117 577 -2113
rect 608 -2117 612 -2113
rect 652 -2117 656 -2113
rect 669 -2117 673 -2113
rect 705 -2117 709 -2113
rect 726 -2117 730 -2113
rect 743 -2124 747 -2077
rect 809 -2080 813 -1923
rect 823 -2065 827 -1691
rect 839 -1815 843 -1166
rect 872 -1192 876 -1153
rect 872 -1207 876 -1196
rect 853 -1211 876 -1207
rect 879 -1183 883 -1146
rect 1197 -1162 1201 -816
rect 1230 -857 1234 -803
rect 1211 -861 1230 -857
rect 1237 -836 1241 -796
rect 1211 -864 1215 -861
rect 1237 -864 1241 -840
rect 1228 -872 1232 -868
rect 1211 -1138 1215 -1134
rect 1228 -1138 1232 -1134
rect 1219 -1149 1223 -1146
rect 1219 -1153 1234 -1149
rect 1197 -1166 1212 -1162
rect 853 -1214 857 -1211
rect 879 -1214 883 -1187
rect 870 -1222 874 -1218
rect 862 -1302 866 -1298
rect 888 -1302 892 -1298
rect 905 -1302 909 -1298
rect 945 -1302 949 -1298
rect 966 -1302 970 -1298
rect 983 -1302 987 -1298
rect 1023 -1302 1027 -1298
rect 1047 -1302 1051 -1298
rect 1084 -1302 1088 -1298
rect 853 -1327 857 -1310
rect 853 -1378 857 -1331
rect 871 -1320 875 -1310
rect 871 -1378 875 -1324
rect 879 -1349 883 -1310
rect 897 -1342 901 -1310
rect 879 -1378 883 -1353
rect 897 -1378 901 -1346
rect 923 -1334 927 -1310
rect 923 -1371 927 -1338
rect 957 -1371 961 -1310
rect 975 -1327 979 -1310
rect 905 -1378 909 -1375
rect 913 -1375 927 -1371
rect 913 -1378 917 -1375
rect 941 -1378 945 -1375
rect 949 -1375 968 -1371
rect 949 -1378 953 -1375
rect 975 -1378 979 -1331
rect 1001 -1342 1005 -1310
rect 1001 -1371 1005 -1346
rect 1035 -1364 1039 -1310
rect 1035 -1368 1052 -1364
rect 983 -1378 987 -1375
rect 992 -1375 1005 -1371
rect 992 -1378 996 -1375
rect 1019 -1378 1023 -1375
rect 1043 -1378 1047 -1368
rect 1059 -1371 1063 -1310
rect 1067 -1364 1071 -1310
rect 1093 -1350 1097 -1310
rect 1067 -1368 1086 -1364
rect 1051 -1375 1068 -1371
rect 1051 -1378 1055 -1375
rect 1075 -1378 1079 -1368
rect 1093 -1378 1097 -1354
rect 862 -1386 866 -1382
rect 888 -1386 892 -1382
rect 931 -1386 935 -1382
rect 966 -1386 970 -1382
rect 1010 -1386 1014 -1382
rect 1027 -1386 1031 -1382
rect 1063 -1386 1067 -1382
rect 1084 -1386 1088 -1382
rect 1100 -1400 1104 -1346
rect 1163 -1357 1167 -1187
rect 862 -1425 866 -1421
rect 879 -1425 883 -1421
rect 899 -1425 903 -1421
rect 920 -1425 924 -1421
rect 941 -1425 945 -1421
rect 962 -1425 966 -1421
rect 983 -1425 987 -1421
rect 1004 -1425 1008 -1421
rect 1025 -1425 1029 -1421
rect 1045 -1425 1049 -1421
rect 853 -1480 857 -1433
rect 853 -1501 857 -1484
rect 871 -1494 875 -1433
rect 887 -1494 891 -1433
rect 911 -1473 915 -1433
rect 911 -1494 915 -1477
rect 929 -1494 933 -1433
rect 953 -1480 957 -1433
rect 953 -1494 957 -1484
rect 971 -1473 975 -1433
rect 971 -1494 975 -1477
rect 995 -1487 999 -1433
rect 1013 -1465 1017 -1433
rect 1013 -1473 1017 -1469
rect 995 -1494 999 -1491
rect 871 -1498 880 -1494
rect 887 -1498 895 -1494
rect 871 -1501 875 -1498
rect 895 -1501 899 -1498
rect 903 -1498 915 -1494
rect 929 -1498 937 -1494
rect 903 -1501 907 -1498
rect 937 -1501 941 -1498
rect 945 -1498 957 -1494
rect 971 -1498 983 -1494
rect 945 -1501 949 -1498
rect 979 -1501 983 -1498
rect 987 -1498 999 -1494
rect 1013 -1494 1017 -1477
rect 1037 -1480 1041 -1433
rect 1037 -1494 1041 -1484
rect 1013 -1498 1025 -1494
rect 987 -1501 991 -1498
rect 1021 -1501 1025 -1498
rect 1029 -1498 1041 -1494
rect 1029 -1501 1033 -1498
rect 862 -1509 866 -1505
rect 879 -1509 883 -1505
rect 920 -1509 924 -1505
rect 962 -1509 966 -1505
rect 1004 -1509 1008 -1505
rect 1045 -1509 1049 -1505
rect 862 -1596 866 -1592
rect 879 -1596 883 -1592
rect 899 -1596 903 -1592
rect 920 -1596 924 -1592
rect 941 -1596 945 -1592
rect 962 -1596 966 -1592
rect 983 -1596 987 -1592
rect 1004 -1596 1008 -1592
rect 1025 -1596 1029 -1592
rect 1045 -1596 1049 -1592
rect 853 -1651 857 -1604
rect 853 -1672 857 -1655
rect 871 -1665 875 -1604
rect 887 -1665 891 -1604
rect 911 -1644 915 -1604
rect 911 -1665 915 -1648
rect 929 -1665 933 -1604
rect 953 -1651 957 -1604
rect 953 -1665 957 -1655
rect 971 -1644 975 -1604
rect 971 -1665 975 -1648
rect 995 -1658 999 -1604
rect 1013 -1636 1017 -1604
rect 1013 -1644 1017 -1640
rect 995 -1665 999 -1662
rect 871 -1669 880 -1665
rect 887 -1669 895 -1665
rect 871 -1672 875 -1669
rect 895 -1672 899 -1669
rect 903 -1669 915 -1665
rect 929 -1669 937 -1665
rect 903 -1672 907 -1669
rect 937 -1672 941 -1669
rect 945 -1669 957 -1665
rect 971 -1669 983 -1665
rect 945 -1672 949 -1669
rect 979 -1672 983 -1669
rect 987 -1669 999 -1665
rect 1013 -1665 1017 -1648
rect 1037 -1651 1041 -1604
rect 1037 -1665 1041 -1655
rect 1013 -1669 1025 -1665
rect 987 -1672 991 -1669
rect 1021 -1672 1025 -1669
rect 1029 -1669 1041 -1665
rect 1029 -1672 1033 -1669
rect 862 -1680 866 -1676
rect 879 -1680 883 -1676
rect 920 -1680 924 -1676
rect 962 -1680 966 -1676
rect 1004 -1680 1008 -1676
rect 1045 -1680 1049 -1676
rect 1063 -1687 1067 -1640
rect 1184 -1644 1188 -1404
rect 862 -1767 866 -1763
rect 879 -1767 883 -1763
rect 899 -1767 903 -1763
rect 920 -1767 924 -1763
rect 941 -1767 945 -1763
rect 962 -1767 966 -1763
rect 983 -1767 987 -1763
rect 1004 -1767 1008 -1763
rect 1025 -1767 1029 -1763
rect 1045 -1767 1049 -1763
rect 853 -1822 857 -1775
rect 853 -1843 857 -1826
rect 871 -1836 875 -1775
rect 887 -1836 891 -1775
rect 911 -1815 915 -1775
rect 911 -1836 915 -1819
rect 929 -1836 933 -1775
rect 953 -1822 957 -1775
rect 953 -1836 957 -1826
rect 971 -1815 975 -1775
rect 971 -1836 975 -1819
rect 995 -1829 999 -1775
rect 1013 -1807 1017 -1775
rect 1013 -1815 1017 -1811
rect 995 -1836 999 -1833
rect 871 -1840 880 -1836
rect 887 -1840 895 -1836
rect 871 -1843 875 -1840
rect 895 -1843 899 -1840
rect 903 -1840 915 -1836
rect 929 -1840 937 -1836
rect 903 -1843 907 -1840
rect 937 -1843 941 -1840
rect 945 -1840 957 -1836
rect 971 -1840 983 -1836
rect 945 -1843 949 -1840
rect 979 -1843 983 -1840
rect 987 -1840 999 -1836
rect 1013 -1836 1017 -1819
rect 1037 -1822 1041 -1775
rect 1037 -1836 1041 -1826
rect 1013 -1840 1025 -1836
rect 987 -1843 991 -1840
rect 1021 -1843 1025 -1840
rect 1029 -1840 1041 -1836
rect 1029 -1843 1033 -1840
rect 862 -1851 866 -1847
rect 879 -1851 883 -1847
rect 920 -1851 924 -1847
rect 962 -1851 966 -1847
rect 1004 -1851 1008 -1847
rect 1045 -1851 1049 -1847
rect 853 -1874 857 -1870
rect 870 -1874 874 -1870
rect 861 -1885 865 -1882
rect 861 -1889 876 -1885
rect 839 -1902 854 -1898
rect 504 -2177 508 -2173
rect 521 -2177 525 -2173
rect 541 -2177 545 -2173
rect 562 -2177 566 -2173
rect 583 -2177 587 -2173
rect 604 -2177 608 -2173
rect 625 -2177 629 -2173
rect 646 -2177 650 -2173
rect 667 -2177 671 -2173
rect 687 -2177 691 -2173
rect 495 -2232 499 -2185
rect 495 -2253 499 -2236
rect 513 -2246 517 -2185
rect 529 -2246 533 -2185
rect 553 -2225 557 -2185
rect 553 -2246 557 -2229
rect 571 -2246 575 -2185
rect 595 -2232 599 -2185
rect 595 -2246 599 -2236
rect 613 -2225 617 -2185
rect 613 -2246 617 -2229
rect 637 -2239 641 -2185
rect 655 -2217 659 -2185
rect 655 -2225 659 -2221
rect 637 -2246 641 -2243
rect 513 -2250 522 -2246
rect 529 -2250 537 -2246
rect 513 -2253 517 -2250
rect 537 -2253 541 -2250
rect 545 -2250 557 -2246
rect 571 -2250 579 -2246
rect 545 -2253 549 -2250
rect 579 -2253 583 -2250
rect 587 -2250 599 -2246
rect 613 -2250 625 -2246
rect 587 -2253 591 -2250
rect 621 -2253 625 -2250
rect 629 -2250 641 -2246
rect 655 -2246 659 -2229
rect 679 -2232 683 -2185
rect 679 -2246 683 -2236
rect 655 -2250 667 -2246
rect 629 -2253 633 -2250
rect 663 -2253 667 -2250
rect 671 -2250 683 -2246
rect 671 -2253 675 -2250
rect 504 -2261 508 -2257
rect 521 -2261 525 -2257
rect 562 -2261 566 -2257
rect 604 -2261 608 -2257
rect 646 -2261 650 -2257
rect 687 -2261 691 -2257
rect 504 -2348 508 -2344
rect 521 -2348 525 -2344
rect 541 -2348 545 -2344
rect 562 -2348 566 -2344
rect 583 -2348 587 -2344
rect 604 -2348 608 -2344
rect 625 -2348 629 -2344
rect 646 -2348 650 -2344
rect 667 -2348 671 -2344
rect 687 -2348 691 -2344
rect 495 -2403 499 -2356
rect 495 -2424 499 -2407
rect 513 -2417 517 -2356
rect 529 -2417 533 -2356
rect 553 -2396 557 -2356
rect 553 -2417 557 -2400
rect 571 -2417 575 -2356
rect 595 -2403 599 -2356
rect 595 -2417 599 -2407
rect 613 -2396 617 -2356
rect 613 -2417 617 -2400
rect 637 -2410 641 -2356
rect 655 -2388 659 -2356
rect 655 -2396 659 -2392
rect 637 -2417 641 -2414
rect 513 -2421 522 -2417
rect 529 -2421 537 -2417
rect 513 -2424 517 -2421
rect 537 -2424 541 -2421
rect 545 -2421 557 -2417
rect 571 -2421 579 -2417
rect 545 -2424 549 -2421
rect 579 -2424 583 -2421
rect 587 -2421 599 -2417
rect 613 -2421 625 -2417
rect 587 -2424 591 -2421
rect 621 -2424 625 -2421
rect 629 -2421 641 -2417
rect 655 -2417 659 -2400
rect 679 -2403 683 -2356
rect 679 -2417 683 -2407
rect 655 -2421 667 -2417
rect 629 -2424 633 -2421
rect 663 -2424 667 -2421
rect 671 -2421 683 -2417
rect 671 -2424 675 -2421
rect 504 -2432 508 -2428
rect 521 -2432 525 -2428
rect 562 -2432 566 -2428
rect 604 -2432 608 -2428
rect 646 -2432 650 -2428
rect 687 -2432 691 -2428
rect 705 -2439 709 -2392
rect 824 -2396 828 -2128
rect 504 -2519 508 -2515
rect 521 -2519 525 -2515
rect 541 -2519 545 -2515
rect 562 -2519 566 -2515
rect 583 -2519 587 -2515
rect 604 -2519 608 -2515
rect 625 -2519 629 -2515
rect 646 -2519 650 -2515
rect 667 -2519 671 -2515
rect 687 -2519 691 -2515
rect 495 -2574 499 -2527
rect 495 -2595 499 -2578
rect 513 -2588 517 -2527
rect 529 -2588 533 -2527
rect 553 -2567 557 -2527
rect 553 -2588 557 -2571
rect 571 -2588 575 -2527
rect 595 -2574 599 -2527
rect 595 -2588 599 -2578
rect 613 -2567 617 -2527
rect 613 -2588 617 -2571
rect 637 -2581 641 -2527
rect 655 -2559 659 -2527
rect 655 -2567 659 -2563
rect 637 -2588 641 -2585
rect 513 -2592 522 -2588
rect 529 -2592 537 -2588
rect 513 -2595 517 -2592
rect 537 -2595 541 -2592
rect 545 -2592 557 -2588
rect 571 -2592 579 -2588
rect 545 -2595 549 -2592
rect 579 -2595 583 -2592
rect 587 -2592 599 -2588
rect 613 -2592 625 -2588
rect 587 -2595 591 -2592
rect 621 -2595 625 -2592
rect 629 -2592 641 -2588
rect 655 -2588 659 -2571
rect 679 -2574 683 -2527
rect 679 -2588 683 -2578
rect 655 -2592 667 -2588
rect 629 -2595 633 -2592
rect 663 -2595 667 -2592
rect 671 -2592 683 -2588
rect 671 -2595 675 -2592
rect 504 -2603 508 -2599
rect 521 -2603 525 -2599
rect 562 -2603 566 -2599
rect 604 -2603 608 -2599
rect 646 -2603 650 -2599
rect 687 -2603 691 -2599
rect 495 -2624 499 -2620
rect 512 -2624 516 -2620
rect 503 -2635 507 -2632
rect 503 -2639 518 -2635
rect 481 -2652 496 -2648
rect 148 -2902 152 -2898
rect 165 -2902 169 -2898
rect 185 -2902 189 -2898
rect 206 -2902 210 -2898
rect 227 -2902 231 -2898
rect 248 -2902 252 -2898
rect 269 -2902 273 -2898
rect 290 -2902 294 -2898
rect 311 -2902 315 -2898
rect 331 -2902 335 -2898
rect 139 -2957 143 -2910
rect 139 -2978 143 -2961
rect 157 -2971 161 -2910
rect 173 -2971 177 -2910
rect 197 -2950 201 -2910
rect 197 -2971 201 -2954
rect 215 -2971 219 -2910
rect 239 -2957 243 -2910
rect 239 -2971 243 -2961
rect 257 -2950 261 -2910
rect 257 -2971 261 -2954
rect 281 -2964 285 -2910
rect 299 -2942 303 -2910
rect 299 -2950 303 -2946
rect 281 -2971 285 -2968
rect 157 -2975 166 -2971
rect 173 -2975 181 -2971
rect 157 -2978 161 -2975
rect 181 -2978 185 -2975
rect 189 -2975 201 -2971
rect 215 -2975 223 -2971
rect 189 -2978 193 -2975
rect 223 -2978 227 -2975
rect 231 -2975 243 -2971
rect 257 -2975 269 -2971
rect 231 -2978 235 -2975
rect 265 -2978 269 -2975
rect 273 -2975 285 -2971
rect 299 -2971 303 -2954
rect 323 -2957 327 -2910
rect 323 -2971 327 -2961
rect 299 -2975 311 -2971
rect 273 -2978 277 -2975
rect 307 -2978 311 -2975
rect 315 -2975 327 -2971
rect 315 -2978 319 -2975
rect 148 -2986 152 -2982
rect 165 -2986 169 -2982
rect 206 -2986 210 -2982
rect 248 -2986 252 -2982
rect 290 -2986 294 -2982
rect 331 -2986 335 -2982
rect 148 -3073 152 -3069
rect 165 -3073 169 -3069
rect 185 -3073 189 -3069
rect 206 -3073 210 -3069
rect 227 -3073 231 -3069
rect 248 -3073 252 -3069
rect 269 -3073 273 -3069
rect 290 -3073 294 -3069
rect 311 -3073 315 -3069
rect 331 -3073 335 -3069
rect 139 -3128 143 -3081
rect 139 -3149 143 -3132
rect 157 -3142 161 -3081
rect 173 -3142 177 -3081
rect 197 -3121 201 -3081
rect 197 -3142 201 -3125
rect 215 -3142 219 -3081
rect 239 -3128 243 -3081
rect 239 -3142 243 -3132
rect 257 -3121 261 -3081
rect 257 -3142 261 -3125
rect 281 -3135 285 -3081
rect 299 -3113 303 -3081
rect 299 -3121 303 -3117
rect 281 -3142 285 -3139
rect 157 -3146 166 -3142
rect 173 -3146 181 -3142
rect 157 -3149 161 -3146
rect 181 -3149 185 -3146
rect 189 -3146 201 -3142
rect 215 -3146 223 -3142
rect 189 -3149 193 -3146
rect 223 -3149 227 -3146
rect 231 -3146 243 -3142
rect 257 -3146 269 -3142
rect 231 -3149 235 -3146
rect 265 -3149 269 -3146
rect 273 -3146 285 -3142
rect 299 -3142 303 -3125
rect 323 -3128 327 -3081
rect 323 -3142 327 -3132
rect 299 -3146 311 -3142
rect 273 -3149 277 -3146
rect 307 -3149 311 -3146
rect 315 -3146 327 -3142
rect 315 -3149 319 -3146
rect 148 -3157 152 -3153
rect 165 -3157 169 -3153
rect 206 -3157 210 -3153
rect 248 -3157 252 -3153
rect 290 -3157 294 -3153
rect 331 -3157 335 -3153
rect 345 -3164 349 -3117
rect 465 -3121 469 -2885
rect 148 -3244 152 -3240
rect 165 -3244 169 -3240
rect 185 -3244 189 -3240
rect 206 -3244 210 -3240
rect 227 -3244 231 -3240
rect 248 -3244 252 -3240
rect 269 -3244 273 -3240
rect 290 -3244 294 -3240
rect 311 -3244 315 -3240
rect 331 -3244 335 -3240
rect 139 -3299 143 -3252
rect 139 -3320 143 -3303
rect 157 -3313 161 -3252
rect 173 -3313 177 -3252
rect 197 -3292 201 -3252
rect 197 -3313 201 -3296
rect 215 -3313 219 -3252
rect 239 -3299 243 -3252
rect 239 -3313 243 -3303
rect 257 -3292 261 -3252
rect 257 -3313 261 -3296
rect 281 -3306 285 -3252
rect 299 -3284 303 -3252
rect 299 -3292 303 -3288
rect 281 -3313 285 -3310
rect 157 -3317 166 -3313
rect 173 -3317 181 -3313
rect 157 -3320 161 -3317
rect 181 -3320 185 -3317
rect 189 -3317 201 -3313
rect 215 -3317 223 -3313
rect 189 -3320 193 -3317
rect 223 -3320 227 -3317
rect 231 -3317 243 -3313
rect 257 -3317 269 -3313
rect 231 -3320 235 -3317
rect 265 -3320 269 -3317
rect 273 -3317 285 -3313
rect 299 -3313 303 -3296
rect 323 -3299 327 -3252
rect 323 -3313 327 -3303
rect 299 -3317 311 -3313
rect 273 -3320 277 -3317
rect 307 -3320 311 -3317
rect 315 -3317 327 -3313
rect 315 -3320 319 -3317
rect 148 -3328 152 -3324
rect 165 -3328 169 -3324
rect 206 -3328 210 -3324
rect 248 -3328 252 -3324
rect 290 -3328 294 -3324
rect 331 -3328 335 -3324
rect 139 -3355 143 -3351
rect 156 -3355 160 -3351
rect 147 -3366 151 -3363
rect 147 -3370 162 -3366
rect 125 -3383 140 -3379
rect -210 -3644 -206 -3640
rect -193 -3644 -189 -3640
rect -173 -3644 -169 -3640
rect -152 -3644 -148 -3640
rect -131 -3644 -127 -3640
rect -110 -3644 -106 -3640
rect -89 -3644 -85 -3640
rect -68 -3644 -64 -3640
rect -47 -3644 -43 -3640
rect -27 -3644 -23 -3640
rect -219 -3699 -215 -3652
rect -219 -3720 -215 -3703
rect -201 -3713 -197 -3652
rect -185 -3713 -181 -3652
rect -161 -3692 -157 -3652
rect -161 -3713 -157 -3696
rect -143 -3713 -139 -3652
rect -119 -3699 -115 -3652
rect -119 -3713 -115 -3703
rect -101 -3692 -97 -3652
rect -101 -3713 -97 -3696
rect -77 -3706 -73 -3652
rect -59 -3684 -55 -3652
rect -59 -3692 -55 -3688
rect -77 -3713 -73 -3710
rect -201 -3717 -192 -3713
rect -185 -3717 -177 -3713
rect -201 -3720 -197 -3717
rect -177 -3720 -173 -3717
rect -169 -3717 -157 -3713
rect -143 -3717 -135 -3713
rect -169 -3720 -165 -3717
rect -135 -3720 -131 -3717
rect -127 -3717 -115 -3713
rect -101 -3717 -89 -3713
rect -127 -3720 -123 -3717
rect -93 -3720 -89 -3717
rect -85 -3717 -73 -3713
rect -59 -3713 -55 -3696
rect -35 -3699 -31 -3652
rect -35 -3713 -31 -3703
rect -59 -3717 -47 -3713
rect -85 -3720 -81 -3717
rect -51 -3720 -47 -3717
rect -43 -3717 -31 -3713
rect -43 -3720 -39 -3717
rect -210 -3728 -206 -3724
rect -193 -3728 -189 -3724
rect -152 -3728 -148 -3724
rect -110 -3728 -106 -3724
rect -68 -3728 -64 -3724
rect -27 -3728 -23 -3724
rect -210 -3815 -206 -3811
rect -193 -3815 -189 -3811
rect -173 -3815 -169 -3811
rect -152 -3815 -148 -3811
rect -131 -3815 -127 -3811
rect -110 -3815 -106 -3811
rect -89 -3815 -85 -3811
rect -68 -3815 -64 -3811
rect -47 -3815 -43 -3811
rect -27 -3815 -23 -3811
rect -219 -3870 -215 -3823
rect -219 -3891 -215 -3874
rect -201 -3884 -197 -3823
rect -185 -3884 -181 -3823
rect -161 -3863 -157 -3823
rect -161 -3884 -157 -3867
rect -143 -3884 -139 -3823
rect -119 -3870 -115 -3823
rect -119 -3884 -115 -3874
rect -101 -3863 -97 -3823
rect -101 -3884 -97 -3867
rect -77 -3877 -73 -3823
rect -59 -3855 -55 -3823
rect -59 -3863 -55 -3859
rect -77 -3884 -73 -3881
rect -201 -3888 -192 -3884
rect -185 -3888 -177 -3884
rect -201 -3891 -197 -3888
rect -177 -3891 -173 -3888
rect -169 -3888 -157 -3884
rect -143 -3888 -135 -3884
rect -169 -3891 -165 -3888
rect -135 -3891 -131 -3888
rect -127 -3888 -115 -3884
rect -101 -3888 -89 -3884
rect -127 -3891 -123 -3888
rect -93 -3891 -89 -3888
rect -85 -3888 -73 -3884
rect -59 -3884 -55 -3867
rect -35 -3870 -31 -3823
rect -35 -3884 -31 -3874
rect -59 -3888 -47 -3884
rect -85 -3891 -81 -3888
rect -51 -3891 -47 -3888
rect -43 -3888 -31 -3884
rect -43 -3891 -39 -3888
rect -210 -3899 -206 -3895
rect -193 -3899 -189 -3895
rect -152 -3899 -148 -3895
rect -110 -3899 -106 -3895
rect -68 -3899 -64 -3895
rect -27 -3899 -23 -3895
rect -9 -3906 -5 -3859
rect 111 -3863 115 -3609
rect -210 -3990 -206 -3986
rect -193 -3990 -189 -3986
rect -173 -3990 -169 -3986
rect -152 -3990 -148 -3986
rect -131 -3990 -127 -3986
rect -110 -3990 -106 -3986
rect -89 -3990 -85 -3986
rect -68 -3990 -64 -3986
rect -47 -3990 -43 -3986
rect -27 -3990 -23 -3986
rect -219 -4045 -215 -3998
rect -219 -4066 -215 -4049
rect -201 -4059 -197 -3998
rect -185 -4059 -181 -3998
rect -161 -4038 -157 -3998
rect -161 -4059 -157 -4042
rect -143 -4059 -139 -3998
rect -119 -4045 -115 -3998
rect -119 -4059 -115 -4049
rect -101 -4038 -97 -3998
rect -101 -4059 -97 -4042
rect -77 -4052 -73 -3998
rect -59 -4030 -55 -3998
rect -59 -4038 -55 -4034
rect -77 -4059 -73 -4056
rect -201 -4063 -192 -4059
rect -185 -4063 -177 -4059
rect -201 -4066 -197 -4063
rect -177 -4066 -173 -4063
rect -169 -4063 -157 -4059
rect -143 -4063 -135 -4059
rect -169 -4066 -165 -4063
rect -135 -4066 -131 -4063
rect -127 -4063 -115 -4059
rect -101 -4063 -89 -4059
rect -127 -4066 -123 -4063
rect -93 -4066 -89 -4063
rect -85 -4063 -73 -4059
rect -59 -4059 -55 -4042
rect -35 -4045 -31 -3998
rect -35 -4059 -31 -4049
rect -59 -4063 -47 -4059
rect -85 -4066 -81 -4063
rect -51 -4066 -47 -4063
rect -43 -4063 -31 -4059
rect -43 -4066 -39 -4063
rect -210 -4074 -206 -4070
rect -193 -4074 -189 -4070
rect -152 -4074 -148 -4070
rect -110 -4074 -106 -4070
rect -68 -4074 -64 -4070
rect -27 -4074 -23 -4070
rect -219 -4105 -215 -4101
rect -202 -4105 -198 -4101
rect -211 -4116 -207 -4113
rect -211 -4120 -196 -4116
rect -233 -4133 -218 -4129
rect -568 -4387 -564 -4383
rect -551 -4387 -547 -4383
rect -531 -4387 -527 -4383
rect -510 -4387 -506 -4383
rect -489 -4387 -485 -4383
rect -468 -4387 -464 -4383
rect -447 -4387 -443 -4383
rect -426 -4387 -422 -4383
rect -405 -4387 -401 -4383
rect -385 -4387 -381 -4383
rect -577 -4442 -573 -4395
rect -577 -4463 -573 -4446
rect -559 -4456 -555 -4395
rect -543 -4456 -539 -4395
rect -519 -4435 -515 -4395
rect -519 -4456 -515 -4439
rect -501 -4456 -497 -4395
rect -477 -4442 -473 -4395
rect -477 -4456 -473 -4446
rect -459 -4435 -455 -4395
rect -459 -4456 -455 -4439
rect -435 -4449 -431 -4395
rect -417 -4427 -413 -4395
rect -417 -4435 -413 -4431
rect -435 -4456 -431 -4453
rect -559 -4460 -550 -4456
rect -543 -4460 -535 -4456
rect -559 -4463 -555 -4460
rect -535 -4463 -531 -4460
rect -527 -4460 -515 -4456
rect -501 -4460 -493 -4456
rect -527 -4463 -523 -4460
rect -493 -4463 -489 -4460
rect -485 -4460 -473 -4456
rect -459 -4460 -447 -4456
rect -485 -4463 -481 -4460
rect -451 -4463 -447 -4460
rect -443 -4460 -431 -4456
rect -417 -4456 -413 -4439
rect -393 -4442 -389 -4395
rect -393 -4456 -389 -4446
rect -417 -4460 -405 -4456
rect -443 -4463 -439 -4460
rect -409 -4463 -405 -4460
rect -401 -4460 -389 -4456
rect -401 -4463 -397 -4460
rect -568 -4471 -564 -4467
rect -551 -4471 -547 -4467
rect -510 -4471 -506 -4467
rect -468 -4471 -464 -4467
rect -426 -4471 -422 -4467
rect -385 -4471 -381 -4467
rect -568 -4558 -564 -4554
rect -551 -4558 -547 -4554
rect -531 -4558 -527 -4554
rect -510 -4558 -506 -4554
rect -489 -4558 -485 -4554
rect -468 -4558 -464 -4554
rect -447 -4558 -443 -4554
rect -426 -4558 -422 -4554
rect -405 -4558 -401 -4554
rect -385 -4558 -381 -4554
rect -577 -4613 -573 -4566
rect -577 -4634 -573 -4617
rect -559 -4627 -555 -4566
rect -543 -4627 -539 -4566
rect -519 -4606 -515 -4566
rect -519 -4627 -515 -4610
rect -501 -4627 -497 -4566
rect -477 -4613 -473 -4566
rect -477 -4627 -473 -4617
rect -459 -4606 -455 -4566
rect -459 -4627 -455 -4610
rect -435 -4620 -431 -4566
rect -417 -4598 -413 -4566
rect -417 -4606 -413 -4602
rect -435 -4627 -431 -4624
rect -559 -4631 -550 -4627
rect -543 -4631 -535 -4627
rect -559 -4634 -555 -4631
rect -535 -4634 -531 -4631
rect -527 -4631 -515 -4627
rect -501 -4631 -493 -4627
rect -527 -4634 -523 -4631
rect -493 -4634 -489 -4631
rect -485 -4631 -473 -4627
rect -459 -4631 -447 -4627
rect -485 -4634 -481 -4631
rect -451 -4634 -447 -4631
rect -443 -4631 -431 -4627
rect -417 -4627 -413 -4610
rect -393 -4613 -389 -4566
rect -393 -4627 -389 -4617
rect -417 -4631 -405 -4627
rect -443 -4634 -439 -4631
rect -409 -4634 -405 -4631
rect -401 -4631 -389 -4627
rect -401 -4634 -397 -4631
rect -568 -4642 -564 -4638
rect -551 -4642 -547 -4638
rect -510 -4642 -506 -4638
rect -468 -4642 -464 -4638
rect -426 -4642 -422 -4638
rect -385 -4642 -381 -4638
rect -370 -4649 -366 -4602
rect -249 -4606 -245 -4366
rect -568 -4729 -564 -4725
rect -551 -4729 -547 -4725
rect -531 -4729 -527 -4725
rect -510 -4729 -506 -4725
rect -489 -4729 -485 -4725
rect -468 -4729 -464 -4725
rect -447 -4729 -443 -4725
rect -426 -4729 -422 -4725
rect -405 -4729 -401 -4725
rect -385 -4729 -381 -4725
rect -577 -4784 -573 -4737
rect -577 -4805 -573 -4788
rect -559 -4798 -555 -4737
rect -543 -4798 -539 -4737
rect -519 -4777 -515 -4737
rect -519 -4798 -515 -4781
rect -501 -4798 -497 -4737
rect -477 -4784 -473 -4737
rect -477 -4798 -473 -4788
rect -459 -4777 -455 -4737
rect -459 -4798 -455 -4781
rect -435 -4791 -431 -4737
rect -417 -4769 -413 -4737
rect -417 -4777 -413 -4773
rect -435 -4798 -431 -4795
rect -559 -4802 -550 -4798
rect -543 -4802 -535 -4798
rect -559 -4805 -555 -4802
rect -535 -4805 -531 -4802
rect -527 -4802 -515 -4798
rect -501 -4802 -493 -4798
rect -527 -4805 -523 -4802
rect -493 -4805 -489 -4802
rect -485 -4802 -473 -4798
rect -459 -4802 -447 -4798
rect -485 -4805 -481 -4802
rect -451 -4805 -447 -4802
rect -443 -4802 -431 -4798
rect -417 -4798 -413 -4781
rect -393 -4784 -389 -4737
rect -393 -4798 -389 -4788
rect -417 -4802 -405 -4798
rect -443 -4805 -439 -4802
rect -409 -4805 -405 -4802
rect -401 -4802 -389 -4798
rect -401 -4805 -397 -4802
rect -568 -4813 -564 -4809
rect -551 -4813 -547 -4809
rect -510 -4813 -506 -4809
rect -468 -4813 -464 -4809
rect -426 -4813 -422 -4809
rect -385 -4813 -381 -4809
rect -577 -4844 -573 -4840
rect -560 -4844 -556 -4840
rect -569 -4855 -565 -4852
rect -569 -4859 -554 -4855
rect -591 -4872 -576 -4868
rect -926 -5122 -922 -5118
rect -909 -5122 -905 -5118
rect -889 -5122 -885 -5118
rect -868 -5122 -864 -5118
rect -847 -5122 -843 -5118
rect -826 -5122 -822 -5118
rect -805 -5122 -801 -5118
rect -784 -5122 -780 -5118
rect -763 -5122 -759 -5118
rect -743 -5122 -739 -5118
rect -935 -5177 -931 -5130
rect -935 -5198 -931 -5181
rect -917 -5191 -913 -5130
rect -901 -5191 -897 -5130
rect -877 -5170 -873 -5130
rect -877 -5191 -873 -5174
rect -859 -5191 -855 -5130
rect -835 -5177 -831 -5130
rect -835 -5191 -831 -5181
rect -817 -5170 -813 -5130
rect -817 -5191 -813 -5174
rect -793 -5184 -789 -5130
rect -775 -5162 -771 -5130
rect -775 -5170 -771 -5166
rect -793 -5191 -789 -5188
rect -917 -5195 -908 -5191
rect -901 -5195 -893 -5191
rect -917 -5198 -913 -5195
rect -893 -5198 -889 -5195
rect -885 -5195 -873 -5191
rect -859 -5195 -851 -5191
rect -885 -5198 -881 -5195
rect -851 -5198 -847 -5195
rect -843 -5195 -831 -5191
rect -817 -5195 -805 -5191
rect -843 -5198 -839 -5195
rect -809 -5198 -805 -5195
rect -801 -5195 -789 -5191
rect -775 -5191 -771 -5174
rect -751 -5177 -747 -5130
rect -751 -5191 -747 -5181
rect -775 -5195 -763 -5191
rect -801 -5198 -797 -5195
rect -767 -5198 -763 -5195
rect -759 -5195 -747 -5191
rect -759 -5198 -755 -5195
rect -926 -5206 -922 -5202
rect -909 -5206 -905 -5202
rect -868 -5206 -864 -5202
rect -826 -5206 -822 -5202
rect -784 -5206 -780 -5202
rect -743 -5206 -739 -5202
rect -926 -5293 -922 -5289
rect -909 -5293 -905 -5289
rect -889 -5293 -885 -5289
rect -868 -5293 -864 -5289
rect -847 -5293 -843 -5289
rect -826 -5293 -822 -5289
rect -805 -5293 -801 -5289
rect -784 -5293 -780 -5289
rect -763 -5293 -759 -5289
rect -743 -5293 -739 -5289
rect -935 -5348 -931 -5301
rect -935 -5369 -931 -5352
rect -917 -5362 -913 -5301
rect -901 -5362 -897 -5301
rect -877 -5341 -873 -5301
rect -877 -5362 -873 -5345
rect -859 -5362 -855 -5301
rect -835 -5348 -831 -5301
rect -835 -5362 -831 -5352
rect -817 -5341 -813 -5301
rect -817 -5362 -813 -5345
rect -793 -5355 -789 -5301
rect -775 -5333 -771 -5301
rect -775 -5341 -771 -5337
rect -793 -5362 -789 -5359
rect -917 -5366 -908 -5362
rect -901 -5366 -893 -5362
rect -917 -5369 -913 -5366
rect -893 -5369 -889 -5366
rect -885 -5366 -873 -5362
rect -859 -5366 -851 -5362
rect -885 -5369 -881 -5366
rect -851 -5369 -847 -5366
rect -843 -5366 -831 -5362
rect -817 -5366 -805 -5362
rect -843 -5369 -839 -5366
rect -809 -5369 -805 -5366
rect -801 -5366 -789 -5362
rect -775 -5362 -771 -5345
rect -751 -5348 -747 -5301
rect -751 -5362 -747 -5352
rect -775 -5366 -763 -5362
rect -801 -5369 -797 -5366
rect -767 -5369 -763 -5366
rect -759 -5366 -747 -5362
rect -759 -5369 -755 -5366
rect -926 -5377 -922 -5373
rect -909 -5377 -905 -5373
rect -868 -5377 -864 -5373
rect -826 -5377 -822 -5373
rect -784 -5377 -780 -5373
rect -743 -5377 -739 -5373
rect -725 -5384 -721 -5337
rect -603 -5341 -599 -5098
rect -926 -5453 -922 -5449
rect -909 -5453 -905 -5449
rect -889 -5453 -885 -5449
rect -868 -5453 -864 -5449
rect -847 -5453 -843 -5449
rect -826 -5453 -822 -5449
rect -805 -5453 -801 -5449
rect -784 -5453 -780 -5449
rect -763 -5453 -759 -5449
rect -743 -5453 -739 -5449
rect -935 -5508 -931 -5461
rect -935 -5529 -931 -5512
rect -917 -5522 -913 -5461
rect -901 -5522 -897 -5461
rect -877 -5501 -873 -5461
rect -877 -5522 -873 -5505
rect -859 -5522 -855 -5461
rect -835 -5508 -831 -5461
rect -835 -5522 -831 -5512
rect -817 -5501 -813 -5461
rect -817 -5522 -813 -5505
rect -793 -5515 -789 -5461
rect -775 -5493 -771 -5461
rect -775 -5501 -771 -5497
rect -793 -5522 -789 -5519
rect -917 -5526 -908 -5522
rect -901 -5526 -893 -5522
rect -917 -5529 -913 -5526
rect -893 -5529 -889 -5526
rect -885 -5526 -873 -5522
rect -859 -5526 -851 -5522
rect -885 -5529 -881 -5526
rect -851 -5529 -847 -5526
rect -843 -5526 -831 -5522
rect -817 -5526 -805 -5522
rect -843 -5529 -839 -5526
rect -809 -5529 -805 -5526
rect -801 -5526 -789 -5522
rect -775 -5522 -771 -5505
rect -751 -5508 -747 -5461
rect -751 -5522 -747 -5512
rect -775 -5526 -763 -5522
rect -801 -5529 -797 -5526
rect -767 -5529 -763 -5526
rect -759 -5526 -747 -5522
rect -759 -5529 -755 -5526
rect -926 -5537 -922 -5533
rect -909 -5537 -905 -5533
rect -868 -5537 -864 -5533
rect -826 -5537 -822 -5533
rect -784 -5537 -780 -5533
rect -743 -5537 -739 -5533
rect -935 -5567 -931 -5563
rect -918 -5567 -914 -5563
rect -927 -5578 -923 -5575
rect -927 -5582 -912 -5578
rect -916 -5621 -912 -5582
rect -916 -5636 -912 -5625
rect -935 -5640 -912 -5636
rect -909 -5612 -905 -5575
rect -725 -5591 -721 -5497
rect -935 -5643 -931 -5640
rect -909 -5643 -905 -5616
rect -918 -5651 -914 -5647
rect -926 -5726 -922 -5722
rect -900 -5726 -896 -5722
rect -883 -5726 -879 -5722
rect -843 -5726 -839 -5722
rect -822 -5726 -818 -5722
rect -805 -5726 -801 -5722
rect -765 -5726 -761 -5722
rect -741 -5726 -737 -5722
rect -704 -5726 -700 -5722
rect -935 -5751 -931 -5734
rect -1225 -5810 -1221 -5806
rect -1181 -5810 -1177 -5806
rect -1147 -5810 -1143 -5806
rect -1103 -5820 -1099 -5792
rect -935 -5802 -931 -5755
rect -917 -5744 -913 -5734
rect -917 -5802 -913 -5748
rect -909 -5773 -905 -5734
rect -891 -5766 -887 -5734
rect -909 -5802 -905 -5777
rect -891 -5802 -887 -5770
rect -865 -5758 -861 -5734
rect -865 -5795 -861 -5762
rect -831 -5795 -827 -5734
rect -813 -5751 -809 -5734
rect -883 -5802 -879 -5799
rect -875 -5799 -861 -5795
rect -875 -5802 -871 -5799
rect -847 -5802 -843 -5799
rect -839 -5799 -820 -5795
rect -839 -5802 -835 -5799
rect -813 -5802 -809 -5755
rect -787 -5766 -783 -5734
rect -787 -5795 -783 -5770
rect -753 -5788 -749 -5734
rect -753 -5792 -736 -5788
rect -805 -5802 -801 -5799
rect -796 -5799 -783 -5795
rect -796 -5802 -792 -5799
rect -769 -5802 -765 -5799
rect -745 -5802 -741 -5792
rect -729 -5795 -725 -5734
rect -721 -5788 -717 -5734
rect -695 -5758 -691 -5734
rect -721 -5792 -702 -5788
rect -737 -5799 -720 -5795
rect -737 -5802 -733 -5799
rect -713 -5802 -709 -5792
rect -695 -5802 -691 -5762
rect -926 -5810 -922 -5806
rect -900 -5810 -896 -5806
rect -857 -5810 -853 -5806
rect -822 -5810 -818 -5806
rect -778 -5810 -774 -5806
rect -761 -5810 -757 -5806
rect -725 -5810 -721 -5806
rect -704 -5810 -700 -5806
rect -683 -5817 -679 -5770
rect -616 -5773 -612 -5616
rect -603 -5758 -599 -5389
rect -591 -5501 -587 -4872
rect -558 -4898 -554 -4859
rect -558 -4913 -554 -4902
rect -577 -4917 -554 -4913
rect -551 -4889 -547 -4852
rect -369 -4868 -365 -4773
rect -577 -4920 -573 -4917
rect -551 -4920 -547 -4893
rect -560 -4928 -556 -4924
rect -568 -5003 -564 -4999
rect -542 -5003 -538 -4999
rect -525 -5003 -521 -4999
rect -485 -5003 -481 -4999
rect -464 -5003 -460 -4999
rect -447 -5003 -443 -4999
rect -407 -5003 -403 -4999
rect -383 -5003 -379 -4999
rect -346 -5003 -342 -4999
rect -577 -5028 -573 -5011
rect -577 -5079 -573 -5032
rect -559 -5021 -555 -5011
rect -559 -5079 -555 -5025
rect -551 -5050 -547 -5011
rect -533 -5043 -529 -5011
rect -551 -5079 -547 -5054
rect -533 -5079 -529 -5047
rect -507 -5035 -503 -5011
rect -507 -5072 -503 -5039
rect -473 -5072 -469 -5011
rect -455 -5028 -451 -5011
rect -525 -5079 -521 -5076
rect -517 -5076 -503 -5072
rect -517 -5079 -513 -5076
rect -489 -5079 -485 -5076
rect -481 -5076 -462 -5072
rect -481 -5079 -477 -5076
rect -455 -5079 -451 -5032
rect -429 -5043 -425 -5011
rect -429 -5072 -425 -5047
rect -395 -5065 -391 -5011
rect -395 -5069 -378 -5065
rect -447 -5079 -443 -5076
rect -438 -5076 -425 -5072
rect -438 -5079 -434 -5076
rect -411 -5079 -407 -5076
rect -387 -5079 -383 -5069
rect -371 -5072 -367 -5011
rect -363 -5065 -359 -5011
rect -337 -5034 -333 -5011
rect -363 -5069 -344 -5065
rect -379 -5076 -362 -5072
rect -379 -5079 -375 -5076
rect -355 -5079 -351 -5069
rect -337 -5079 -333 -5038
rect -568 -5087 -564 -5083
rect -542 -5087 -538 -5083
rect -499 -5087 -495 -5083
rect -464 -5087 -460 -5083
rect -420 -5087 -416 -5083
rect -403 -5087 -399 -5083
rect -367 -5087 -363 -5083
rect -346 -5087 -342 -5083
rect -328 -5101 -324 -5047
rect -263 -5050 -259 -4893
rect -249 -5035 -245 -4653
rect -233 -4777 -229 -4133
rect -200 -4159 -196 -4120
rect -200 -4174 -196 -4163
rect -219 -4178 -196 -4174
rect -193 -4150 -189 -4113
rect -9 -4129 -5 -4034
rect -219 -4181 -215 -4178
rect -193 -4181 -189 -4154
rect -202 -4189 -198 -4185
rect -210 -4264 -206 -4260
rect -184 -4264 -180 -4260
rect -167 -4264 -163 -4260
rect -127 -4264 -123 -4260
rect -106 -4264 -102 -4260
rect -89 -4264 -85 -4260
rect -49 -4264 -45 -4260
rect -25 -4264 -21 -4260
rect 12 -4264 16 -4260
rect -219 -4289 -215 -4272
rect -219 -4340 -215 -4293
rect -201 -4282 -197 -4272
rect -201 -4340 -197 -4286
rect -193 -4311 -189 -4272
rect -175 -4304 -171 -4272
rect -193 -4340 -189 -4315
rect -175 -4340 -171 -4308
rect -149 -4296 -145 -4272
rect -149 -4333 -145 -4300
rect -115 -4333 -111 -4272
rect -97 -4289 -93 -4272
rect -167 -4340 -163 -4337
rect -159 -4337 -145 -4333
rect -159 -4340 -155 -4337
rect -131 -4340 -127 -4337
rect -123 -4337 -104 -4333
rect -123 -4340 -119 -4337
rect -97 -4340 -93 -4293
rect -71 -4304 -67 -4272
rect -71 -4333 -67 -4308
rect -37 -4326 -33 -4272
rect -37 -4330 -20 -4326
rect -89 -4340 -85 -4337
rect -80 -4337 -67 -4333
rect -80 -4340 -76 -4337
rect -53 -4340 -49 -4337
rect -29 -4340 -25 -4330
rect -13 -4333 -9 -4272
rect -5 -4326 -1 -4272
rect 21 -4296 25 -4272
rect -5 -4330 14 -4326
rect -21 -4337 -4 -4333
rect -21 -4340 -17 -4337
rect 3 -4340 7 -4330
rect 21 -4340 25 -4300
rect -210 -4348 -206 -4344
rect -184 -4348 -180 -4344
rect -141 -4348 -137 -4344
rect -106 -4348 -102 -4344
rect -62 -4348 -58 -4344
rect -45 -4348 -41 -4344
rect -9 -4348 -5 -4344
rect 12 -4348 16 -4344
rect 29 -4355 33 -4308
rect 97 -4311 101 -4154
rect 111 -4296 115 -3910
rect 125 -4038 129 -3383
rect 158 -3409 162 -3370
rect 158 -3424 162 -3413
rect 139 -3428 162 -3424
rect 165 -3400 169 -3363
rect 347 -3379 351 -3288
rect 139 -3431 143 -3428
rect 165 -3431 169 -3404
rect 156 -3439 160 -3435
rect 148 -3514 152 -3510
rect 174 -3514 178 -3510
rect 191 -3514 195 -3510
rect 231 -3514 235 -3510
rect 252 -3514 256 -3510
rect 269 -3514 273 -3510
rect 309 -3514 313 -3510
rect 333 -3514 337 -3510
rect 370 -3514 374 -3510
rect 139 -3539 143 -3522
rect 139 -3590 143 -3543
rect 157 -3532 161 -3522
rect 157 -3590 161 -3536
rect 165 -3561 169 -3522
rect 183 -3554 187 -3522
rect 165 -3590 169 -3565
rect 183 -3590 187 -3558
rect 209 -3546 213 -3522
rect 209 -3583 213 -3550
rect 243 -3583 247 -3522
rect 261 -3539 265 -3522
rect 191 -3590 195 -3587
rect 199 -3587 213 -3583
rect 199 -3590 203 -3587
rect 227 -3590 231 -3587
rect 235 -3587 254 -3583
rect 235 -3590 239 -3587
rect 261 -3590 265 -3543
rect 287 -3554 291 -3522
rect 287 -3583 291 -3558
rect 321 -3576 325 -3522
rect 321 -3580 338 -3576
rect 269 -3590 273 -3587
rect 278 -3587 291 -3583
rect 278 -3590 282 -3587
rect 305 -3590 309 -3587
rect 329 -3590 333 -3580
rect 345 -3583 349 -3522
rect 353 -3576 357 -3522
rect 379 -3546 383 -3522
rect 353 -3580 372 -3576
rect 337 -3587 354 -3583
rect 337 -3590 341 -3587
rect 361 -3590 365 -3580
rect 379 -3590 383 -3550
rect 148 -3598 152 -3594
rect 174 -3598 178 -3594
rect 217 -3598 221 -3594
rect 252 -3598 256 -3594
rect 296 -3598 300 -3594
rect 313 -3598 317 -3594
rect 349 -3598 353 -3594
rect 370 -3598 374 -3594
rect 388 -3612 392 -3558
rect 451 -3561 455 -3404
rect 465 -3546 469 -3168
rect 481 -3292 485 -2652
rect 514 -2678 518 -2639
rect 514 -2693 518 -2682
rect 495 -2697 518 -2693
rect 521 -2669 525 -2632
rect 703 -2648 707 -2563
rect 495 -2700 499 -2697
rect 521 -2700 525 -2673
rect 512 -2708 516 -2704
rect 504 -2783 508 -2779
rect 530 -2783 534 -2779
rect 547 -2783 551 -2779
rect 587 -2783 591 -2779
rect 608 -2783 612 -2779
rect 625 -2783 629 -2779
rect 665 -2783 669 -2779
rect 689 -2783 693 -2779
rect 726 -2783 730 -2779
rect 495 -2808 499 -2791
rect 495 -2859 499 -2812
rect 513 -2801 517 -2791
rect 513 -2859 517 -2805
rect 521 -2830 525 -2791
rect 539 -2823 543 -2791
rect 521 -2859 525 -2834
rect 539 -2859 543 -2827
rect 565 -2815 569 -2791
rect 565 -2852 569 -2819
rect 599 -2852 603 -2791
rect 617 -2808 621 -2791
rect 547 -2859 551 -2856
rect 555 -2856 569 -2852
rect 555 -2859 559 -2856
rect 583 -2859 587 -2856
rect 591 -2856 610 -2852
rect 591 -2859 595 -2856
rect 617 -2859 621 -2812
rect 643 -2823 647 -2791
rect 643 -2852 647 -2827
rect 677 -2845 681 -2791
rect 677 -2849 694 -2845
rect 625 -2859 629 -2856
rect 634 -2856 647 -2852
rect 634 -2859 638 -2856
rect 661 -2859 665 -2856
rect 685 -2859 689 -2849
rect 701 -2852 705 -2791
rect 709 -2845 713 -2791
rect 735 -2815 739 -2791
rect 709 -2849 728 -2845
rect 693 -2856 710 -2852
rect 693 -2859 697 -2856
rect 717 -2859 721 -2849
rect 735 -2859 739 -2819
rect 504 -2867 508 -2863
rect 530 -2867 534 -2863
rect 573 -2867 577 -2863
rect 608 -2867 612 -2863
rect 652 -2867 656 -2863
rect 669 -2867 673 -2863
rect 705 -2867 709 -2863
rect 726 -2867 730 -2863
rect 742 -2874 746 -2827
rect 810 -2830 814 -2673
rect 824 -2815 828 -2444
rect 839 -2567 843 -1902
rect 872 -1928 876 -1889
rect 872 -1943 876 -1932
rect 853 -1947 876 -1943
rect 879 -1919 883 -1882
rect 1060 -1898 1064 -1811
rect 853 -1950 857 -1947
rect 879 -1950 883 -1923
rect 870 -1958 874 -1954
rect 862 -2033 866 -2029
rect 888 -2033 892 -2029
rect 905 -2033 909 -2029
rect 945 -2033 949 -2029
rect 966 -2033 970 -2029
rect 983 -2033 987 -2029
rect 1023 -2033 1027 -2029
rect 1047 -2033 1051 -2029
rect 1084 -2033 1088 -2029
rect 853 -2058 857 -2041
rect 853 -2109 857 -2062
rect 871 -2051 875 -2041
rect 871 -2109 875 -2055
rect 879 -2080 883 -2041
rect 897 -2073 901 -2041
rect 879 -2109 883 -2084
rect 897 -2109 901 -2077
rect 923 -2065 927 -2041
rect 923 -2102 927 -2069
rect 957 -2102 961 -2041
rect 975 -2058 979 -2041
rect 905 -2109 909 -2106
rect 913 -2106 927 -2102
rect 913 -2109 917 -2106
rect 941 -2109 945 -2106
rect 949 -2106 968 -2102
rect 949 -2109 953 -2106
rect 975 -2109 979 -2062
rect 1001 -2073 1005 -2041
rect 1001 -2102 1005 -2077
rect 1035 -2095 1039 -2041
rect 1035 -2099 1052 -2095
rect 983 -2109 987 -2106
rect 992 -2106 1005 -2102
rect 992 -2109 996 -2106
rect 1019 -2109 1023 -2106
rect 1043 -2109 1047 -2099
rect 1059 -2102 1063 -2041
rect 1067 -2095 1071 -2041
rect 1093 -2063 1097 -2041
rect 1093 -2081 1097 -2067
rect 1167 -2065 1171 -1923
rect 1067 -2099 1086 -2095
rect 1051 -2106 1068 -2102
rect 1051 -2109 1055 -2106
rect 1075 -2109 1079 -2099
rect 1093 -2109 1097 -2085
rect 862 -2117 866 -2113
rect 888 -2117 892 -2113
rect 931 -2117 935 -2113
rect 966 -2117 970 -2113
rect 1010 -2117 1014 -2113
rect 1027 -2117 1031 -2113
rect 1063 -2117 1067 -2113
rect 1084 -2117 1088 -2113
rect 1101 -2131 1105 -2077
rect 1184 -2080 1188 -1692
rect 1197 -1815 1201 -1166
rect 1230 -1192 1234 -1153
rect 1230 -1207 1234 -1196
rect 1211 -1211 1234 -1207
rect 1237 -1183 1241 -1146
rect 1211 -1214 1215 -1211
rect 1237 -1214 1241 -1187
rect 1228 -1222 1232 -1218
rect 1220 -1302 1224 -1298
rect 1237 -1302 1241 -1298
rect 1277 -1302 1281 -1298
rect 1298 -1302 1302 -1298
rect 1211 -1343 1215 -1310
rect 1211 -1378 1215 -1347
rect 1229 -1337 1233 -1310
rect 1229 -1341 1238 -1337
rect 1229 -1378 1233 -1341
rect 1255 -1364 1259 -1310
rect 1255 -1371 1259 -1368
rect 1289 -1371 1293 -1310
rect 1307 -1342 1311 -1310
rect 1311 -1346 1333 -1342
rect 1237 -1378 1241 -1375
rect 1246 -1375 1259 -1371
rect 1246 -1378 1250 -1375
rect 1273 -1378 1277 -1375
rect 1281 -1375 1300 -1371
rect 1281 -1378 1285 -1375
rect 1307 -1378 1311 -1346
rect 1220 -1386 1224 -1382
rect 1264 -1386 1268 -1382
rect 1298 -1386 1302 -1382
rect 1322 -1407 1326 -1368
rect 1329 -1400 1333 -1346
rect 1220 -1596 1224 -1592
rect 1237 -1596 1241 -1592
rect 1257 -1596 1261 -1592
rect 1278 -1596 1282 -1592
rect 1299 -1596 1303 -1592
rect 1320 -1596 1324 -1592
rect 1341 -1596 1345 -1592
rect 1362 -1596 1366 -1592
rect 1383 -1596 1387 -1592
rect 1403 -1596 1407 -1592
rect 1211 -1651 1215 -1604
rect 1211 -1672 1215 -1655
rect 1229 -1665 1233 -1604
rect 1245 -1665 1249 -1604
rect 1269 -1644 1273 -1604
rect 1269 -1665 1273 -1648
rect 1287 -1665 1291 -1604
rect 1311 -1651 1315 -1604
rect 1311 -1665 1315 -1655
rect 1329 -1644 1333 -1604
rect 1329 -1665 1333 -1648
rect 1353 -1658 1357 -1604
rect 1371 -1636 1375 -1604
rect 1371 -1644 1375 -1640
rect 1353 -1665 1357 -1662
rect 1229 -1669 1238 -1665
rect 1245 -1669 1253 -1665
rect 1229 -1672 1233 -1669
rect 1253 -1672 1257 -1669
rect 1261 -1669 1273 -1665
rect 1287 -1669 1295 -1665
rect 1261 -1672 1265 -1669
rect 1295 -1672 1299 -1669
rect 1303 -1669 1315 -1665
rect 1329 -1669 1341 -1665
rect 1303 -1672 1307 -1669
rect 1337 -1672 1341 -1669
rect 1345 -1669 1357 -1665
rect 1371 -1665 1375 -1648
rect 1395 -1651 1399 -1604
rect 1395 -1665 1399 -1655
rect 1371 -1669 1383 -1665
rect 1345 -1672 1349 -1669
rect 1379 -1672 1383 -1669
rect 1387 -1669 1399 -1665
rect 1387 -1672 1391 -1669
rect 1220 -1680 1224 -1676
rect 1237 -1680 1241 -1676
rect 1278 -1680 1282 -1676
rect 1320 -1680 1324 -1676
rect 1362 -1680 1366 -1676
rect 1403 -1680 1407 -1676
rect 1424 -1688 1428 -1640
rect 1220 -1767 1224 -1763
rect 1237 -1767 1241 -1763
rect 1257 -1767 1261 -1763
rect 1278 -1767 1282 -1763
rect 1299 -1767 1303 -1763
rect 1320 -1767 1324 -1763
rect 1341 -1767 1345 -1763
rect 1362 -1767 1366 -1763
rect 1383 -1767 1387 -1763
rect 1403 -1767 1407 -1763
rect 1211 -1822 1215 -1775
rect 1211 -1843 1215 -1826
rect 1229 -1836 1233 -1775
rect 1245 -1836 1249 -1775
rect 1269 -1815 1273 -1775
rect 1269 -1836 1273 -1819
rect 1287 -1836 1291 -1775
rect 1311 -1822 1315 -1775
rect 1311 -1836 1315 -1826
rect 1329 -1815 1333 -1775
rect 1329 -1836 1333 -1819
rect 1353 -1829 1357 -1775
rect 1371 -1807 1375 -1775
rect 1371 -1815 1375 -1811
rect 1353 -1836 1357 -1833
rect 1229 -1840 1238 -1836
rect 1245 -1840 1253 -1836
rect 1229 -1843 1233 -1840
rect 1253 -1843 1257 -1840
rect 1261 -1840 1273 -1836
rect 1287 -1840 1295 -1836
rect 1261 -1843 1265 -1840
rect 1295 -1843 1299 -1840
rect 1303 -1840 1315 -1836
rect 1329 -1840 1341 -1836
rect 1303 -1843 1307 -1840
rect 1337 -1843 1341 -1840
rect 1345 -1840 1357 -1836
rect 1371 -1836 1375 -1819
rect 1395 -1822 1399 -1775
rect 1395 -1836 1399 -1826
rect 1371 -1840 1383 -1836
rect 1345 -1843 1349 -1840
rect 1379 -1843 1383 -1840
rect 1387 -1840 1399 -1836
rect 1387 -1843 1391 -1840
rect 1220 -1851 1224 -1847
rect 1237 -1851 1241 -1847
rect 1278 -1851 1282 -1847
rect 1320 -1851 1324 -1847
rect 1362 -1851 1366 -1847
rect 1403 -1851 1407 -1847
rect 1211 -1874 1215 -1870
rect 1228 -1874 1232 -1870
rect 1219 -1885 1223 -1882
rect 1219 -1889 1234 -1885
rect 1197 -1902 1212 -1898
rect 862 -2348 866 -2344
rect 879 -2348 883 -2344
rect 899 -2348 903 -2344
rect 920 -2348 924 -2344
rect 941 -2348 945 -2344
rect 962 -2348 966 -2344
rect 983 -2348 987 -2344
rect 1004 -2348 1008 -2344
rect 1025 -2348 1029 -2344
rect 1045 -2348 1049 -2344
rect 853 -2403 857 -2356
rect 853 -2424 857 -2407
rect 871 -2417 875 -2356
rect 887 -2417 891 -2356
rect 911 -2396 915 -2356
rect 911 -2417 915 -2400
rect 929 -2417 933 -2356
rect 953 -2403 957 -2356
rect 953 -2417 957 -2407
rect 971 -2396 975 -2356
rect 971 -2417 975 -2400
rect 995 -2410 999 -2356
rect 1013 -2388 1017 -2356
rect 1013 -2396 1017 -2392
rect 995 -2417 999 -2414
rect 871 -2421 880 -2417
rect 887 -2421 895 -2417
rect 871 -2424 875 -2421
rect 895 -2424 899 -2421
rect 903 -2421 915 -2417
rect 929 -2421 937 -2417
rect 903 -2424 907 -2421
rect 937 -2424 941 -2421
rect 945 -2421 957 -2417
rect 971 -2421 983 -2417
rect 945 -2424 949 -2421
rect 979 -2424 983 -2421
rect 987 -2421 999 -2417
rect 1013 -2417 1017 -2400
rect 1037 -2403 1041 -2356
rect 1037 -2417 1041 -2407
rect 1013 -2421 1025 -2417
rect 987 -2424 991 -2421
rect 1021 -2424 1025 -2421
rect 1029 -2421 1041 -2417
rect 1029 -2424 1033 -2421
rect 862 -2432 866 -2428
rect 879 -2432 883 -2428
rect 920 -2432 924 -2428
rect 962 -2432 966 -2428
rect 1004 -2432 1008 -2428
rect 1045 -2432 1049 -2428
rect 1062 -2440 1066 -2392
rect 1184 -2396 1188 -2135
rect 862 -2519 866 -2515
rect 879 -2519 883 -2515
rect 899 -2519 903 -2515
rect 920 -2519 924 -2515
rect 941 -2519 945 -2515
rect 962 -2519 966 -2515
rect 983 -2519 987 -2515
rect 1004 -2519 1008 -2515
rect 1025 -2519 1029 -2515
rect 1045 -2519 1049 -2515
rect 853 -2574 857 -2527
rect 853 -2595 857 -2578
rect 871 -2588 875 -2527
rect 887 -2588 891 -2527
rect 911 -2567 915 -2527
rect 911 -2588 915 -2571
rect 929 -2588 933 -2527
rect 953 -2574 957 -2527
rect 953 -2588 957 -2578
rect 971 -2567 975 -2527
rect 971 -2588 975 -2571
rect 995 -2581 999 -2527
rect 1013 -2559 1017 -2527
rect 1013 -2567 1017 -2563
rect 995 -2588 999 -2585
rect 871 -2592 880 -2588
rect 887 -2592 895 -2588
rect 871 -2595 875 -2592
rect 895 -2595 899 -2592
rect 903 -2592 915 -2588
rect 929 -2592 937 -2588
rect 903 -2595 907 -2592
rect 937 -2595 941 -2592
rect 945 -2592 957 -2588
rect 971 -2592 983 -2588
rect 945 -2595 949 -2592
rect 979 -2595 983 -2592
rect 987 -2592 999 -2588
rect 1013 -2588 1017 -2571
rect 1037 -2574 1041 -2527
rect 1037 -2588 1041 -2578
rect 1013 -2592 1025 -2588
rect 987 -2595 991 -2592
rect 1021 -2595 1025 -2592
rect 1029 -2592 1041 -2588
rect 1029 -2595 1033 -2592
rect 862 -2603 866 -2599
rect 879 -2603 883 -2599
rect 920 -2603 924 -2599
rect 962 -2603 966 -2599
rect 1004 -2603 1008 -2599
rect 1045 -2603 1049 -2599
rect 853 -2624 857 -2620
rect 870 -2624 874 -2620
rect 861 -2635 865 -2632
rect 861 -2639 876 -2635
rect 839 -2652 854 -2648
rect 504 -3073 508 -3069
rect 521 -3073 525 -3069
rect 541 -3073 545 -3069
rect 562 -3073 566 -3069
rect 583 -3073 587 -3069
rect 604 -3073 608 -3069
rect 625 -3073 629 -3069
rect 646 -3073 650 -3069
rect 667 -3073 671 -3069
rect 687 -3073 691 -3069
rect 495 -3128 499 -3081
rect 495 -3149 499 -3132
rect 513 -3142 517 -3081
rect 529 -3142 533 -3081
rect 553 -3121 557 -3081
rect 553 -3142 557 -3125
rect 571 -3142 575 -3081
rect 595 -3128 599 -3081
rect 595 -3142 599 -3132
rect 613 -3121 617 -3081
rect 613 -3142 617 -3125
rect 637 -3135 641 -3081
rect 655 -3113 659 -3081
rect 655 -3121 659 -3117
rect 637 -3142 641 -3139
rect 513 -3146 522 -3142
rect 529 -3146 537 -3142
rect 513 -3149 517 -3146
rect 537 -3149 541 -3146
rect 545 -3146 557 -3142
rect 571 -3146 579 -3142
rect 545 -3149 549 -3146
rect 579 -3149 583 -3146
rect 587 -3146 599 -3142
rect 613 -3146 625 -3142
rect 587 -3149 591 -3146
rect 621 -3149 625 -3146
rect 629 -3146 641 -3142
rect 655 -3142 659 -3125
rect 679 -3128 683 -3081
rect 679 -3142 683 -3132
rect 655 -3146 667 -3142
rect 629 -3149 633 -3146
rect 663 -3149 667 -3146
rect 671 -3146 683 -3142
rect 671 -3149 675 -3146
rect 504 -3157 508 -3153
rect 521 -3157 525 -3153
rect 562 -3157 566 -3153
rect 604 -3157 608 -3153
rect 646 -3157 650 -3153
rect 687 -3157 691 -3153
rect 701 -3164 705 -3117
rect 823 -3121 827 -2878
rect 504 -3244 508 -3240
rect 521 -3244 525 -3240
rect 541 -3244 545 -3240
rect 562 -3244 566 -3240
rect 583 -3244 587 -3240
rect 604 -3244 608 -3240
rect 625 -3244 629 -3240
rect 646 -3244 650 -3240
rect 667 -3244 671 -3240
rect 687 -3244 691 -3240
rect 495 -3299 499 -3252
rect 495 -3320 499 -3303
rect 513 -3313 517 -3252
rect 529 -3313 533 -3252
rect 553 -3292 557 -3252
rect 553 -3313 557 -3296
rect 571 -3313 575 -3252
rect 595 -3299 599 -3252
rect 595 -3313 599 -3303
rect 613 -3292 617 -3252
rect 613 -3313 617 -3296
rect 637 -3306 641 -3252
rect 655 -3284 659 -3252
rect 655 -3292 659 -3288
rect 637 -3313 641 -3310
rect 513 -3317 522 -3313
rect 529 -3317 537 -3313
rect 513 -3320 517 -3317
rect 537 -3320 541 -3317
rect 545 -3317 557 -3313
rect 571 -3317 579 -3313
rect 545 -3320 549 -3317
rect 579 -3320 583 -3317
rect 587 -3317 599 -3313
rect 613 -3317 625 -3313
rect 587 -3320 591 -3317
rect 621 -3320 625 -3317
rect 629 -3317 641 -3313
rect 655 -3313 659 -3296
rect 679 -3299 683 -3252
rect 679 -3313 683 -3303
rect 655 -3317 667 -3313
rect 629 -3320 633 -3317
rect 663 -3320 667 -3317
rect 671 -3317 683 -3313
rect 671 -3320 675 -3317
rect 504 -3328 508 -3324
rect 521 -3328 525 -3324
rect 562 -3328 566 -3324
rect 604 -3328 608 -3324
rect 646 -3328 650 -3324
rect 687 -3328 691 -3324
rect 495 -3355 499 -3351
rect 512 -3355 516 -3351
rect 503 -3366 507 -3363
rect 503 -3370 518 -3366
rect 481 -3383 496 -3379
rect 148 -3815 152 -3811
rect 165 -3815 169 -3811
rect 185 -3815 189 -3811
rect 206 -3815 210 -3811
rect 227 -3815 231 -3811
rect 248 -3815 252 -3811
rect 269 -3815 273 -3811
rect 290 -3815 294 -3811
rect 311 -3815 315 -3811
rect 331 -3815 335 -3811
rect 139 -3870 143 -3823
rect 139 -3891 143 -3874
rect 157 -3884 161 -3823
rect 173 -3884 177 -3823
rect 197 -3863 201 -3823
rect 197 -3884 201 -3867
rect 215 -3884 219 -3823
rect 239 -3870 243 -3823
rect 239 -3884 243 -3874
rect 257 -3863 261 -3823
rect 257 -3884 261 -3867
rect 281 -3877 285 -3823
rect 299 -3855 303 -3823
rect 299 -3863 303 -3859
rect 281 -3884 285 -3881
rect 157 -3888 166 -3884
rect 173 -3888 181 -3884
rect 157 -3891 161 -3888
rect 181 -3891 185 -3888
rect 189 -3888 201 -3884
rect 215 -3888 223 -3884
rect 189 -3891 193 -3888
rect 223 -3891 227 -3888
rect 231 -3888 243 -3884
rect 257 -3888 269 -3884
rect 231 -3891 235 -3888
rect 265 -3891 269 -3888
rect 273 -3888 285 -3884
rect 299 -3884 303 -3867
rect 323 -3870 327 -3823
rect 323 -3884 327 -3874
rect 299 -3888 311 -3884
rect 273 -3891 277 -3888
rect 307 -3891 311 -3888
rect 315 -3888 327 -3884
rect 315 -3891 319 -3888
rect 148 -3899 152 -3895
rect 165 -3899 169 -3895
rect 206 -3899 210 -3895
rect 248 -3899 252 -3895
rect 290 -3899 294 -3895
rect 331 -3899 335 -3895
rect 349 -3906 353 -3859
rect 465 -3863 469 -3616
rect 148 -3990 152 -3986
rect 165 -3990 169 -3986
rect 185 -3990 189 -3986
rect 206 -3990 210 -3986
rect 227 -3990 231 -3986
rect 248 -3990 252 -3986
rect 269 -3990 273 -3986
rect 290 -3990 294 -3986
rect 311 -3990 315 -3986
rect 331 -3990 335 -3986
rect 139 -4045 143 -3998
rect 139 -4066 143 -4049
rect 157 -4059 161 -3998
rect 173 -4059 177 -3998
rect 197 -4038 201 -3998
rect 197 -4059 201 -4042
rect 215 -4059 219 -3998
rect 239 -4045 243 -3998
rect 239 -4059 243 -4049
rect 257 -4038 261 -3998
rect 257 -4059 261 -4042
rect 281 -4052 285 -3998
rect 299 -4030 303 -3998
rect 299 -4038 303 -4034
rect 281 -4059 285 -4056
rect 157 -4063 166 -4059
rect 173 -4063 181 -4059
rect 157 -4066 161 -4063
rect 181 -4066 185 -4063
rect 189 -4063 201 -4059
rect 215 -4063 223 -4059
rect 189 -4066 193 -4063
rect 223 -4066 227 -4063
rect 231 -4063 243 -4059
rect 257 -4063 269 -4059
rect 231 -4066 235 -4063
rect 265 -4066 269 -4063
rect 273 -4063 285 -4059
rect 299 -4059 303 -4042
rect 323 -4045 327 -3998
rect 323 -4059 327 -4049
rect 299 -4063 311 -4059
rect 273 -4066 277 -4063
rect 307 -4066 311 -4063
rect 315 -4063 327 -4059
rect 315 -4066 319 -4063
rect 148 -4074 152 -4070
rect 165 -4074 169 -4070
rect 206 -4074 210 -4070
rect 248 -4074 252 -4070
rect 290 -4074 294 -4070
rect 331 -4074 335 -4070
rect 139 -4105 143 -4101
rect 156 -4105 160 -4101
rect 147 -4116 151 -4113
rect 147 -4120 162 -4116
rect 125 -4133 140 -4129
rect -210 -4558 -206 -4554
rect -193 -4558 -189 -4554
rect -173 -4558 -169 -4554
rect -152 -4558 -148 -4554
rect -131 -4558 -127 -4554
rect -110 -4558 -106 -4554
rect -89 -4558 -85 -4554
rect -68 -4558 -64 -4554
rect -47 -4558 -43 -4554
rect -27 -4558 -23 -4554
rect -219 -4613 -215 -4566
rect -219 -4634 -215 -4617
rect -201 -4627 -197 -4566
rect -185 -4627 -181 -4566
rect -161 -4606 -157 -4566
rect -161 -4627 -157 -4610
rect -143 -4627 -139 -4566
rect -119 -4613 -115 -4566
rect -119 -4627 -115 -4617
rect -101 -4606 -97 -4566
rect -101 -4627 -97 -4610
rect -77 -4620 -73 -4566
rect -59 -4598 -55 -4566
rect -59 -4606 -55 -4602
rect -77 -4627 -73 -4624
rect -201 -4631 -192 -4627
rect -185 -4631 -177 -4627
rect -201 -4634 -197 -4631
rect -177 -4634 -173 -4631
rect -169 -4631 -157 -4627
rect -143 -4631 -135 -4627
rect -169 -4634 -165 -4631
rect -135 -4634 -131 -4631
rect -127 -4631 -115 -4627
rect -101 -4631 -89 -4627
rect -127 -4634 -123 -4631
rect -93 -4634 -89 -4631
rect -85 -4631 -73 -4627
rect -59 -4627 -55 -4610
rect -35 -4613 -31 -4566
rect -35 -4627 -31 -4617
rect -59 -4631 -47 -4627
rect -85 -4634 -81 -4631
rect -51 -4634 -47 -4631
rect -43 -4631 -31 -4627
rect -43 -4634 -39 -4631
rect -210 -4642 -206 -4638
rect -193 -4642 -189 -4638
rect -152 -4642 -148 -4638
rect -110 -4642 -106 -4638
rect -68 -4642 -64 -4638
rect -27 -4642 -23 -4638
rect -9 -4649 -5 -4602
rect 111 -4606 115 -4359
rect -210 -4729 -206 -4725
rect -193 -4729 -189 -4725
rect -173 -4729 -169 -4725
rect -152 -4729 -148 -4725
rect -131 -4729 -127 -4725
rect -110 -4729 -106 -4725
rect -89 -4729 -85 -4725
rect -68 -4729 -64 -4725
rect -47 -4729 -43 -4725
rect -27 -4729 -23 -4725
rect -219 -4784 -215 -4737
rect -219 -4805 -215 -4788
rect -201 -4798 -197 -4737
rect -185 -4798 -181 -4737
rect -161 -4777 -157 -4737
rect -161 -4798 -157 -4781
rect -143 -4798 -139 -4737
rect -119 -4784 -115 -4737
rect -119 -4798 -115 -4788
rect -101 -4777 -97 -4737
rect -101 -4798 -97 -4781
rect -77 -4791 -73 -4737
rect -59 -4769 -55 -4737
rect -59 -4777 -55 -4773
rect -77 -4798 -73 -4795
rect -201 -4802 -192 -4798
rect -185 -4802 -177 -4798
rect -201 -4805 -197 -4802
rect -177 -4805 -173 -4802
rect -169 -4802 -157 -4798
rect -143 -4802 -135 -4798
rect -169 -4805 -165 -4802
rect -135 -4805 -131 -4802
rect -127 -4802 -115 -4798
rect -101 -4802 -89 -4798
rect -127 -4805 -123 -4802
rect -93 -4805 -89 -4802
rect -85 -4802 -73 -4798
rect -59 -4798 -55 -4781
rect -35 -4784 -31 -4737
rect -35 -4798 -31 -4788
rect -59 -4802 -47 -4798
rect -85 -4805 -81 -4802
rect -51 -4805 -47 -4802
rect -43 -4802 -31 -4798
rect -43 -4805 -39 -4802
rect -210 -4813 -206 -4809
rect -193 -4813 -189 -4809
rect -152 -4813 -148 -4809
rect -110 -4813 -106 -4809
rect -68 -4813 -64 -4809
rect -27 -4813 -23 -4809
rect -219 -4844 -215 -4840
rect -202 -4844 -198 -4840
rect -211 -4855 -207 -4852
rect -211 -4859 -196 -4855
rect -233 -4872 -218 -4868
rect -568 -5293 -564 -5289
rect -551 -5293 -547 -5289
rect -531 -5293 -527 -5289
rect -510 -5293 -506 -5289
rect -489 -5293 -485 -5289
rect -468 -5293 -464 -5289
rect -447 -5293 -443 -5289
rect -426 -5293 -422 -5289
rect -405 -5293 -401 -5289
rect -385 -5293 -381 -5289
rect -577 -5348 -573 -5301
rect -577 -5369 -573 -5352
rect -559 -5362 -555 -5301
rect -543 -5362 -539 -5301
rect -519 -5341 -515 -5301
rect -519 -5362 -515 -5345
rect -501 -5362 -497 -5301
rect -477 -5348 -473 -5301
rect -477 -5362 -473 -5352
rect -459 -5341 -455 -5301
rect -459 -5362 -455 -5345
rect -435 -5355 -431 -5301
rect -417 -5333 -413 -5301
rect -417 -5341 -413 -5337
rect -435 -5362 -431 -5359
rect -559 -5366 -550 -5362
rect -543 -5366 -535 -5362
rect -559 -5369 -555 -5366
rect -535 -5369 -531 -5366
rect -527 -5366 -515 -5362
rect -501 -5366 -493 -5362
rect -527 -5369 -523 -5366
rect -493 -5369 -489 -5366
rect -485 -5366 -473 -5362
rect -459 -5366 -447 -5362
rect -485 -5369 -481 -5366
rect -451 -5369 -447 -5366
rect -443 -5366 -431 -5362
rect -417 -5362 -413 -5345
rect -393 -5348 -389 -5301
rect -393 -5362 -389 -5352
rect -417 -5366 -405 -5362
rect -443 -5369 -439 -5366
rect -409 -5369 -405 -5366
rect -401 -5366 -389 -5362
rect -401 -5369 -397 -5366
rect -568 -5377 -564 -5373
rect -551 -5377 -547 -5373
rect -510 -5377 -506 -5373
rect -468 -5377 -464 -5373
rect -426 -5377 -422 -5373
rect -385 -5377 -381 -5373
rect -369 -5385 -365 -5337
rect -249 -5341 -245 -5105
rect -568 -5453 -564 -5449
rect -551 -5453 -547 -5449
rect -531 -5453 -527 -5449
rect -510 -5453 -506 -5449
rect -489 -5453 -485 -5449
rect -468 -5453 -464 -5449
rect -447 -5453 -443 -5449
rect -426 -5453 -422 -5449
rect -405 -5453 -401 -5449
rect -385 -5453 -381 -5449
rect -577 -5508 -573 -5461
rect -577 -5529 -573 -5512
rect -559 -5522 -555 -5461
rect -543 -5522 -539 -5461
rect -519 -5501 -515 -5461
rect -519 -5522 -515 -5505
rect -501 -5522 -497 -5461
rect -477 -5508 -473 -5461
rect -477 -5522 -473 -5512
rect -459 -5501 -455 -5461
rect -459 -5522 -455 -5505
rect -435 -5515 -431 -5461
rect -417 -5493 -413 -5461
rect -417 -5501 -413 -5497
rect -435 -5522 -431 -5519
rect -559 -5526 -550 -5522
rect -543 -5526 -535 -5522
rect -559 -5529 -555 -5526
rect -535 -5529 -531 -5526
rect -527 -5526 -515 -5522
rect -501 -5526 -493 -5522
rect -527 -5529 -523 -5526
rect -493 -5529 -489 -5526
rect -485 -5526 -473 -5522
rect -459 -5526 -447 -5522
rect -485 -5529 -481 -5526
rect -451 -5529 -447 -5526
rect -443 -5526 -431 -5522
rect -417 -5522 -413 -5505
rect -393 -5508 -389 -5461
rect -393 -5522 -389 -5512
rect -417 -5526 -405 -5522
rect -443 -5529 -439 -5526
rect -409 -5529 -405 -5526
rect -401 -5526 -389 -5522
rect -401 -5529 -397 -5526
rect -568 -5537 -564 -5533
rect -551 -5537 -547 -5533
rect -510 -5537 -506 -5533
rect -468 -5537 -464 -5533
rect -426 -5537 -422 -5533
rect -385 -5537 -381 -5533
rect -577 -5567 -573 -5563
rect -560 -5567 -556 -5563
rect -569 -5578 -565 -5575
rect -569 -5582 -554 -5578
rect -558 -5621 -554 -5582
rect -558 -5636 -554 -5625
rect -577 -5640 -554 -5636
rect -551 -5612 -547 -5575
rect -368 -5591 -364 -5497
rect -577 -5643 -573 -5640
rect -551 -5643 -547 -5616
rect -560 -5651 -556 -5647
rect -568 -5726 -564 -5722
rect -542 -5726 -538 -5722
rect -525 -5726 -521 -5722
rect -485 -5726 -481 -5722
rect -464 -5726 -460 -5722
rect -447 -5726 -443 -5722
rect -407 -5726 -403 -5722
rect -383 -5726 -379 -5722
rect -346 -5726 -342 -5722
rect -577 -5751 -573 -5734
rect -577 -5802 -573 -5755
rect -559 -5744 -555 -5734
rect -559 -5802 -555 -5748
rect -551 -5773 -547 -5734
rect -533 -5766 -529 -5734
rect -551 -5802 -547 -5777
rect -533 -5802 -529 -5770
rect -507 -5758 -503 -5734
rect -507 -5795 -503 -5762
rect -473 -5795 -469 -5734
rect -455 -5751 -451 -5734
rect -525 -5802 -521 -5799
rect -517 -5799 -503 -5795
rect -517 -5802 -513 -5799
rect -489 -5802 -485 -5799
rect -481 -5799 -462 -5795
rect -481 -5802 -477 -5799
rect -455 -5802 -451 -5755
rect -429 -5766 -425 -5734
rect -429 -5795 -425 -5770
rect -395 -5788 -391 -5734
rect -395 -5792 -378 -5788
rect -447 -5802 -443 -5799
rect -438 -5799 -425 -5795
rect -438 -5802 -434 -5799
rect -411 -5802 -407 -5799
rect -387 -5802 -383 -5792
rect -371 -5795 -367 -5734
rect -363 -5788 -359 -5734
rect -337 -5757 -333 -5734
rect -363 -5792 -344 -5788
rect -379 -5799 -362 -5795
rect -379 -5802 -375 -5799
rect -355 -5802 -351 -5792
rect -337 -5802 -333 -5761
rect -568 -5810 -564 -5806
rect -542 -5810 -538 -5806
rect -499 -5810 -495 -5806
rect -464 -5810 -460 -5806
rect -420 -5810 -416 -5806
rect -403 -5810 -399 -5806
rect -367 -5810 -363 -5806
rect -346 -5810 -342 -5806
rect -326 -5817 -322 -5770
rect -263 -5773 -259 -5616
rect -249 -5758 -245 -5388
rect -233 -5501 -229 -4872
rect -200 -4898 -196 -4859
rect -200 -4913 -196 -4902
rect -219 -4917 -196 -4913
rect -193 -4889 -189 -4852
rect -11 -4868 -7 -4773
rect -219 -4920 -215 -4917
rect -193 -4920 -189 -4893
rect -202 -4928 -198 -4924
rect -210 -5003 -206 -4999
rect -184 -5003 -180 -4999
rect -167 -5003 -163 -4999
rect -127 -5003 -123 -4999
rect -106 -5003 -102 -4999
rect -89 -5003 -85 -4999
rect -49 -5003 -45 -4999
rect -25 -5003 -21 -4999
rect 12 -5003 16 -4999
rect -219 -5028 -215 -5011
rect -219 -5079 -215 -5032
rect -201 -5021 -197 -5011
rect -201 -5079 -197 -5025
rect -193 -5050 -189 -5011
rect -175 -5043 -171 -5011
rect -193 -5079 -189 -5054
rect -175 -5079 -171 -5047
rect -149 -5035 -145 -5011
rect -149 -5072 -145 -5039
rect -115 -5072 -111 -5011
rect -97 -5028 -93 -5011
rect -167 -5079 -163 -5076
rect -159 -5076 -145 -5072
rect -159 -5079 -155 -5076
rect -131 -5079 -127 -5076
rect -123 -5076 -104 -5072
rect -123 -5079 -119 -5076
rect -97 -5079 -93 -5032
rect -71 -5043 -67 -5011
rect -71 -5072 -67 -5047
rect -37 -5065 -33 -5011
rect -37 -5069 -20 -5065
rect -89 -5079 -85 -5076
rect -80 -5076 -67 -5072
rect -80 -5079 -76 -5076
rect -53 -5079 -49 -5076
rect -29 -5079 -25 -5069
rect -13 -5072 -9 -5011
rect -5 -5065 -1 -5011
rect 21 -5035 25 -5011
rect -5 -5069 14 -5065
rect -21 -5076 -4 -5072
rect -21 -5079 -17 -5076
rect 3 -5079 7 -5069
rect 21 -5079 25 -5039
rect -210 -5087 -206 -5083
rect -184 -5087 -180 -5083
rect -141 -5087 -137 -5083
rect -106 -5087 -102 -5083
rect -62 -5087 -58 -5083
rect -45 -5087 -41 -5083
rect -9 -5087 -5 -5083
rect 12 -5087 16 -5083
rect 29 -5094 33 -5047
rect 97 -5050 101 -4893
rect 111 -5035 115 -4655
rect 125 -4777 129 -4133
rect 158 -4159 162 -4120
rect 158 -4174 162 -4163
rect 139 -4178 162 -4174
rect 165 -4150 169 -4113
rect 348 -4129 352 -4034
rect 139 -4181 143 -4178
rect 165 -4181 169 -4154
rect 156 -4189 160 -4185
rect 148 -4264 152 -4260
rect 174 -4264 178 -4260
rect 191 -4264 195 -4260
rect 231 -4264 235 -4260
rect 252 -4264 256 -4260
rect 269 -4264 273 -4260
rect 309 -4264 313 -4260
rect 333 -4264 337 -4260
rect 370 -4264 374 -4260
rect 139 -4289 143 -4272
rect 139 -4340 143 -4293
rect 157 -4282 161 -4272
rect 157 -4340 161 -4286
rect 165 -4311 169 -4272
rect 183 -4304 187 -4272
rect 165 -4340 169 -4315
rect 183 -4340 187 -4308
rect 209 -4296 213 -4272
rect 209 -4333 213 -4300
rect 243 -4333 247 -4272
rect 261 -4289 265 -4272
rect 191 -4340 195 -4337
rect 199 -4337 213 -4333
rect 199 -4340 203 -4337
rect 227 -4340 231 -4337
rect 235 -4337 254 -4333
rect 235 -4340 239 -4337
rect 261 -4340 265 -4293
rect 287 -4304 291 -4272
rect 287 -4333 291 -4308
rect 321 -4326 325 -4272
rect 321 -4330 338 -4326
rect 269 -4340 273 -4337
rect 278 -4337 291 -4333
rect 278 -4340 282 -4337
rect 305 -4340 309 -4337
rect 329 -4340 333 -4330
rect 345 -4333 349 -4272
rect 353 -4326 357 -4272
rect 379 -4296 383 -4272
rect 353 -4330 372 -4326
rect 337 -4337 354 -4333
rect 337 -4340 341 -4337
rect 361 -4340 365 -4330
rect 379 -4340 383 -4300
rect 148 -4348 152 -4344
rect 174 -4348 178 -4344
rect 217 -4348 221 -4344
rect 252 -4348 256 -4344
rect 296 -4348 300 -4344
rect 313 -4348 317 -4344
rect 349 -4348 353 -4344
rect 370 -4348 374 -4344
rect 388 -4362 392 -4308
rect 451 -4311 455 -4154
rect 465 -4296 469 -3911
rect 481 -4038 485 -3383
rect 514 -3409 518 -3370
rect 514 -3424 518 -3413
rect 495 -3428 518 -3424
rect 521 -3400 525 -3363
rect 705 -3379 709 -3288
rect 495 -3431 499 -3428
rect 521 -3431 525 -3404
rect 512 -3439 516 -3435
rect 809 -3506 813 -3404
rect 823 -3506 827 -3168
rect 839 -3292 843 -2652
rect 872 -2678 876 -2639
rect 872 -2693 876 -2682
rect 853 -2697 876 -2693
rect 879 -2669 883 -2632
rect 1062 -2648 1066 -2563
rect 853 -2700 857 -2697
rect 879 -2700 883 -2673
rect 870 -2708 874 -2704
rect 862 -2783 866 -2779
rect 888 -2783 892 -2779
rect 905 -2783 909 -2779
rect 945 -2783 949 -2779
rect 966 -2783 970 -2779
rect 983 -2783 987 -2779
rect 1023 -2783 1027 -2779
rect 1047 -2783 1051 -2779
rect 1084 -2783 1088 -2779
rect 853 -2808 857 -2791
rect 853 -2859 857 -2812
rect 871 -2801 875 -2791
rect 871 -2859 875 -2805
rect 879 -2830 883 -2791
rect 897 -2823 901 -2791
rect 879 -2859 883 -2834
rect 897 -2859 901 -2827
rect 923 -2815 927 -2791
rect 923 -2852 927 -2819
rect 957 -2852 961 -2791
rect 975 -2808 979 -2791
rect 905 -2859 909 -2856
rect 913 -2856 927 -2852
rect 913 -2859 917 -2856
rect 941 -2859 945 -2856
rect 949 -2856 968 -2852
rect 949 -2859 953 -2856
rect 975 -2859 979 -2812
rect 1001 -2823 1005 -2791
rect 1001 -2852 1005 -2827
rect 1035 -2845 1039 -2791
rect 1035 -2849 1052 -2845
rect 983 -2859 987 -2856
rect 992 -2856 1005 -2852
rect 992 -2859 996 -2856
rect 1019 -2859 1023 -2856
rect 1043 -2859 1047 -2849
rect 1059 -2852 1063 -2791
rect 1067 -2845 1071 -2791
rect 1093 -2813 1097 -2791
rect 1093 -2831 1097 -2817
rect 1167 -2815 1171 -2673
rect 1067 -2849 1086 -2845
rect 1051 -2856 1068 -2852
rect 1051 -2859 1055 -2856
rect 1075 -2859 1079 -2849
rect 1093 -2859 1097 -2835
rect 862 -2867 866 -2863
rect 888 -2867 892 -2863
rect 931 -2867 935 -2863
rect 966 -2867 970 -2863
rect 1010 -2867 1014 -2863
rect 1027 -2867 1031 -2863
rect 1063 -2867 1067 -2863
rect 1084 -2867 1088 -2863
rect 1103 -2881 1107 -2827
rect 1184 -2830 1188 -2444
rect 1197 -2567 1201 -1902
rect 1230 -1928 1234 -1889
rect 1230 -1943 1234 -1932
rect 1211 -1947 1234 -1943
rect 1237 -1919 1241 -1882
rect 1419 -1898 1423 -1811
rect 1211 -1950 1215 -1947
rect 1237 -1950 1241 -1923
rect 1228 -1958 1232 -1954
rect 1220 -2033 1224 -2029
rect 1246 -2033 1250 -2029
rect 1263 -2033 1267 -2029
rect 1303 -2033 1307 -2029
rect 1324 -2033 1328 -2029
rect 1341 -2033 1345 -2029
rect 1381 -2033 1385 -2029
rect 1405 -2033 1409 -2029
rect 1442 -2033 1446 -2029
rect 1211 -2058 1215 -2041
rect 1211 -2109 1215 -2062
rect 1229 -2051 1233 -2041
rect 1229 -2109 1233 -2055
rect 1237 -2080 1241 -2041
rect 1255 -2073 1259 -2041
rect 1237 -2109 1241 -2084
rect 1255 -2109 1259 -2077
rect 1281 -2065 1285 -2041
rect 1281 -2102 1285 -2069
rect 1315 -2102 1319 -2041
rect 1333 -2058 1337 -2041
rect 1263 -2109 1267 -2106
rect 1271 -2106 1285 -2102
rect 1271 -2109 1275 -2106
rect 1299 -2109 1303 -2106
rect 1307 -2106 1326 -2102
rect 1307 -2109 1311 -2106
rect 1333 -2109 1337 -2062
rect 1359 -2073 1363 -2041
rect 1359 -2102 1363 -2077
rect 1393 -2095 1397 -2041
rect 1393 -2099 1410 -2095
rect 1341 -2109 1345 -2106
rect 1350 -2106 1363 -2102
rect 1350 -2109 1354 -2106
rect 1377 -2109 1381 -2106
rect 1401 -2109 1405 -2099
rect 1417 -2102 1421 -2041
rect 1425 -2095 1429 -2041
rect 1425 -2099 1444 -2095
rect 1409 -2106 1426 -2102
rect 1409 -2109 1413 -2106
rect 1433 -2109 1437 -2099
rect 1451 -2109 1455 -2041
rect 1220 -2117 1224 -2113
rect 1246 -2117 1250 -2113
rect 1289 -2117 1293 -2113
rect 1324 -2117 1328 -2113
rect 1368 -2117 1372 -2113
rect 1385 -2117 1389 -2113
rect 1421 -2117 1425 -2113
rect 1442 -2117 1446 -2113
rect 1451 -2131 1455 -2113
rect 1466 -2124 1470 -2077
rect 1220 -2348 1224 -2344
rect 1237 -2348 1241 -2344
rect 1257 -2348 1261 -2344
rect 1278 -2348 1282 -2344
rect 1299 -2348 1303 -2344
rect 1320 -2348 1324 -2344
rect 1341 -2348 1345 -2344
rect 1362 -2348 1366 -2344
rect 1383 -2348 1387 -2344
rect 1403 -2348 1407 -2344
rect 1211 -2403 1215 -2356
rect 1211 -2424 1215 -2407
rect 1229 -2417 1233 -2356
rect 1245 -2417 1249 -2356
rect 1269 -2396 1273 -2356
rect 1269 -2417 1273 -2400
rect 1287 -2417 1291 -2356
rect 1311 -2403 1315 -2356
rect 1311 -2417 1315 -2407
rect 1329 -2396 1333 -2356
rect 1329 -2417 1333 -2400
rect 1353 -2410 1357 -2356
rect 1371 -2388 1375 -2356
rect 1371 -2396 1375 -2392
rect 1353 -2417 1357 -2414
rect 1229 -2421 1238 -2417
rect 1245 -2421 1253 -2417
rect 1229 -2424 1233 -2421
rect 1253 -2424 1257 -2421
rect 1261 -2421 1273 -2417
rect 1287 -2421 1295 -2417
rect 1261 -2424 1265 -2421
rect 1295 -2424 1299 -2421
rect 1303 -2421 1315 -2417
rect 1329 -2421 1341 -2417
rect 1303 -2424 1307 -2421
rect 1337 -2424 1341 -2421
rect 1345 -2421 1357 -2417
rect 1371 -2417 1375 -2400
rect 1395 -2403 1399 -2356
rect 1395 -2417 1399 -2407
rect 1371 -2421 1383 -2417
rect 1345 -2424 1349 -2421
rect 1379 -2424 1383 -2421
rect 1387 -2421 1399 -2417
rect 1387 -2424 1391 -2421
rect 1220 -2432 1224 -2428
rect 1237 -2432 1241 -2428
rect 1278 -2432 1282 -2428
rect 1320 -2432 1324 -2428
rect 1362 -2432 1366 -2428
rect 1403 -2432 1407 -2428
rect 1421 -2440 1425 -2392
rect 1220 -2519 1224 -2515
rect 1237 -2519 1241 -2515
rect 1257 -2519 1261 -2515
rect 1278 -2519 1282 -2515
rect 1299 -2519 1303 -2515
rect 1320 -2519 1324 -2515
rect 1341 -2519 1345 -2515
rect 1362 -2519 1366 -2515
rect 1383 -2519 1387 -2515
rect 1403 -2519 1407 -2515
rect 1211 -2574 1215 -2527
rect 1211 -2595 1215 -2578
rect 1229 -2588 1233 -2527
rect 1245 -2588 1249 -2527
rect 1269 -2567 1273 -2527
rect 1269 -2588 1273 -2571
rect 1287 -2588 1291 -2527
rect 1311 -2574 1315 -2527
rect 1311 -2588 1315 -2578
rect 1329 -2567 1333 -2527
rect 1329 -2588 1333 -2571
rect 1353 -2581 1357 -2527
rect 1371 -2559 1375 -2527
rect 1371 -2567 1375 -2563
rect 1353 -2588 1357 -2585
rect 1229 -2592 1238 -2588
rect 1245 -2592 1253 -2588
rect 1229 -2595 1233 -2592
rect 1253 -2595 1257 -2592
rect 1261 -2592 1273 -2588
rect 1287 -2592 1295 -2588
rect 1261 -2595 1265 -2592
rect 1295 -2595 1299 -2592
rect 1303 -2592 1315 -2588
rect 1329 -2592 1341 -2588
rect 1303 -2595 1307 -2592
rect 1337 -2595 1341 -2592
rect 1345 -2592 1357 -2588
rect 1371 -2588 1375 -2571
rect 1395 -2574 1399 -2527
rect 1395 -2588 1399 -2578
rect 1371 -2592 1383 -2588
rect 1345 -2595 1349 -2592
rect 1379 -2595 1383 -2592
rect 1387 -2592 1399 -2588
rect 1387 -2595 1391 -2592
rect 1220 -2603 1224 -2599
rect 1237 -2603 1241 -2599
rect 1278 -2603 1282 -2599
rect 1320 -2603 1324 -2599
rect 1362 -2603 1366 -2599
rect 1403 -2603 1407 -2599
rect 1211 -2624 1215 -2620
rect 1228 -2624 1232 -2620
rect 1219 -2635 1223 -2632
rect 1219 -2639 1234 -2635
rect 1197 -2652 1212 -2648
rect 862 -3073 866 -3069
rect 879 -3073 883 -3069
rect 899 -3073 903 -3069
rect 920 -3073 924 -3069
rect 941 -3073 945 -3069
rect 962 -3073 966 -3069
rect 983 -3073 987 -3069
rect 1004 -3073 1008 -3069
rect 1025 -3073 1029 -3069
rect 1045 -3073 1049 -3069
rect 853 -3128 857 -3081
rect 853 -3149 857 -3132
rect 871 -3142 875 -3081
rect 887 -3142 891 -3081
rect 911 -3121 915 -3081
rect 911 -3142 915 -3125
rect 929 -3142 933 -3081
rect 953 -3128 957 -3081
rect 953 -3142 957 -3132
rect 971 -3121 975 -3081
rect 971 -3142 975 -3125
rect 995 -3135 999 -3081
rect 1013 -3113 1017 -3081
rect 1013 -3121 1017 -3117
rect 995 -3142 999 -3139
rect 871 -3146 880 -3142
rect 887 -3146 895 -3142
rect 871 -3149 875 -3146
rect 895 -3149 899 -3146
rect 903 -3146 915 -3142
rect 929 -3146 937 -3142
rect 903 -3149 907 -3146
rect 937 -3149 941 -3146
rect 945 -3146 957 -3142
rect 971 -3146 983 -3142
rect 945 -3149 949 -3146
rect 979 -3149 983 -3146
rect 987 -3146 999 -3142
rect 1013 -3142 1017 -3125
rect 1037 -3128 1041 -3081
rect 1037 -3142 1041 -3132
rect 1013 -3146 1025 -3142
rect 987 -3149 991 -3146
rect 1021 -3149 1025 -3146
rect 1029 -3146 1041 -3142
rect 1029 -3149 1033 -3146
rect 862 -3157 866 -3153
rect 879 -3157 883 -3153
rect 920 -3157 924 -3153
rect 962 -3157 966 -3153
rect 1004 -3157 1008 -3153
rect 1045 -3157 1049 -3153
rect 1060 -3164 1064 -3117
rect 1184 -3121 1188 -2885
rect 862 -3244 866 -3240
rect 879 -3244 883 -3240
rect 899 -3244 903 -3240
rect 920 -3244 924 -3240
rect 941 -3244 945 -3240
rect 962 -3244 966 -3240
rect 983 -3244 987 -3240
rect 1004 -3244 1008 -3240
rect 1025 -3244 1029 -3240
rect 1045 -3244 1049 -3240
rect 853 -3299 857 -3252
rect 853 -3320 857 -3303
rect 871 -3313 875 -3252
rect 887 -3313 891 -3252
rect 911 -3292 915 -3252
rect 911 -3313 915 -3296
rect 929 -3313 933 -3252
rect 953 -3299 957 -3252
rect 953 -3313 957 -3303
rect 971 -3292 975 -3252
rect 971 -3313 975 -3296
rect 995 -3306 999 -3252
rect 1013 -3284 1017 -3252
rect 1013 -3292 1017 -3288
rect 995 -3313 999 -3310
rect 871 -3317 880 -3313
rect 887 -3317 895 -3313
rect 871 -3320 875 -3317
rect 895 -3320 899 -3317
rect 903 -3317 915 -3313
rect 929 -3317 937 -3313
rect 903 -3320 907 -3317
rect 937 -3320 941 -3317
rect 945 -3317 957 -3313
rect 971 -3317 983 -3313
rect 945 -3320 949 -3317
rect 979 -3320 983 -3317
rect 987 -3317 999 -3313
rect 1013 -3313 1017 -3296
rect 1037 -3299 1041 -3252
rect 1037 -3313 1041 -3303
rect 1013 -3317 1025 -3313
rect 987 -3320 991 -3317
rect 1021 -3320 1025 -3317
rect 1029 -3317 1041 -3313
rect 1029 -3320 1033 -3317
rect 862 -3328 866 -3324
rect 879 -3328 883 -3324
rect 920 -3328 924 -3324
rect 962 -3328 966 -3324
rect 1004 -3328 1008 -3324
rect 1045 -3328 1049 -3324
rect 853 -3355 857 -3351
rect 870 -3355 874 -3351
rect 861 -3366 865 -3363
rect 861 -3370 876 -3366
rect 839 -3383 854 -3379
rect 504 -3514 508 -3510
rect 530 -3514 534 -3510
rect 547 -3514 551 -3510
rect 587 -3514 591 -3510
rect 608 -3514 612 -3510
rect 625 -3514 629 -3510
rect 665 -3514 669 -3510
rect 689 -3514 693 -3510
rect 726 -3514 730 -3510
rect 495 -3539 499 -3522
rect 495 -3590 499 -3543
rect 513 -3532 517 -3522
rect 513 -3590 517 -3536
rect 521 -3561 525 -3522
rect 539 -3554 543 -3522
rect 521 -3590 525 -3565
rect 539 -3590 543 -3558
rect 565 -3546 569 -3522
rect 565 -3583 569 -3550
rect 599 -3583 603 -3522
rect 617 -3539 621 -3522
rect 547 -3590 551 -3587
rect 555 -3587 569 -3583
rect 555 -3590 559 -3587
rect 583 -3590 587 -3587
rect 591 -3587 610 -3583
rect 591 -3590 595 -3587
rect 617 -3590 621 -3543
rect 643 -3554 647 -3522
rect 643 -3583 647 -3558
rect 677 -3576 681 -3522
rect 677 -3580 694 -3576
rect 625 -3590 629 -3587
rect 634 -3587 647 -3583
rect 634 -3590 638 -3587
rect 661 -3590 665 -3587
rect 685 -3590 689 -3580
rect 701 -3583 705 -3522
rect 709 -3576 713 -3522
rect 735 -3546 739 -3522
rect 709 -3580 728 -3576
rect 693 -3587 710 -3583
rect 693 -3590 697 -3587
rect 717 -3590 721 -3580
rect 735 -3590 739 -3550
rect 504 -3598 508 -3594
rect 530 -3598 534 -3594
rect 573 -3598 577 -3594
rect 608 -3598 612 -3594
rect 652 -3598 656 -3594
rect 669 -3598 673 -3594
rect 705 -3598 709 -3594
rect 726 -3598 730 -3594
rect 743 -3605 747 -3558
rect 810 -3561 814 -3506
rect 824 -3546 828 -3506
rect 504 -3815 508 -3811
rect 521 -3815 525 -3811
rect 541 -3815 545 -3811
rect 562 -3815 566 -3811
rect 583 -3815 587 -3811
rect 604 -3815 608 -3811
rect 625 -3815 629 -3811
rect 646 -3815 650 -3811
rect 667 -3815 671 -3811
rect 687 -3815 691 -3811
rect 495 -3870 499 -3823
rect 495 -3891 499 -3874
rect 513 -3884 517 -3823
rect 529 -3884 533 -3823
rect 553 -3863 557 -3823
rect 553 -3884 557 -3867
rect 571 -3884 575 -3823
rect 595 -3870 599 -3823
rect 595 -3884 599 -3874
rect 613 -3863 617 -3823
rect 613 -3884 617 -3867
rect 637 -3877 641 -3823
rect 655 -3855 659 -3823
rect 655 -3863 659 -3859
rect 637 -3884 641 -3881
rect 513 -3888 522 -3884
rect 529 -3888 537 -3884
rect 513 -3891 517 -3888
rect 537 -3891 541 -3888
rect 545 -3888 557 -3884
rect 571 -3888 579 -3884
rect 545 -3891 549 -3888
rect 579 -3891 583 -3888
rect 587 -3888 599 -3884
rect 613 -3888 625 -3884
rect 587 -3891 591 -3888
rect 621 -3891 625 -3888
rect 629 -3888 641 -3884
rect 655 -3884 659 -3867
rect 679 -3870 683 -3823
rect 679 -3884 683 -3874
rect 655 -3888 667 -3884
rect 629 -3891 633 -3888
rect 663 -3891 667 -3888
rect 671 -3888 683 -3884
rect 671 -3891 675 -3888
rect 504 -3899 508 -3895
rect 521 -3899 525 -3895
rect 562 -3899 566 -3895
rect 604 -3899 608 -3895
rect 646 -3899 650 -3895
rect 687 -3899 691 -3895
rect 702 -3907 706 -3859
rect 824 -3863 828 -3609
rect 504 -3990 508 -3986
rect 521 -3990 525 -3986
rect 541 -3990 545 -3986
rect 562 -3990 566 -3986
rect 583 -3990 587 -3986
rect 604 -3990 608 -3986
rect 625 -3990 629 -3986
rect 646 -3990 650 -3986
rect 667 -3990 671 -3986
rect 687 -3990 691 -3986
rect 495 -4045 499 -3998
rect 495 -4066 499 -4049
rect 513 -4059 517 -3998
rect 529 -4059 533 -3998
rect 553 -4038 557 -3998
rect 553 -4059 557 -4042
rect 571 -4059 575 -3998
rect 595 -4045 599 -3998
rect 595 -4059 599 -4049
rect 613 -4038 617 -3998
rect 613 -4059 617 -4042
rect 637 -4052 641 -3998
rect 655 -4030 659 -3998
rect 655 -4038 659 -4034
rect 637 -4059 641 -4056
rect 513 -4063 522 -4059
rect 529 -4063 537 -4059
rect 513 -4066 517 -4063
rect 537 -4066 541 -4063
rect 545 -4063 557 -4059
rect 571 -4063 579 -4059
rect 545 -4066 549 -4063
rect 579 -4066 583 -4063
rect 587 -4063 599 -4059
rect 613 -4063 625 -4059
rect 587 -4066 591 -4063
rect 621 -4066 625 -4063
rect 629 -4063 641 -4059
rect 655 -4059 659 -4042
rect 679 -4045 683 -3998
rect 679 -4059 683 -4049
rect 655 -4063 667 -4059
rect 629 -4066 633 -4063
rect 663 -4066 667 -4063
rect 671 -4063 683 -4059
rect 671 -4066 675 -4063
rect 504 -4074 508 -4070
rect 521 -4074 525 -4070
rect 562 -4074 566 -4070
rect 604 -4074 608 -4070
rect 646 -4074 650 -4070
rect 687 -4074 691 -4070
rect 495 -4105 499 -4101
rect 512 -4105 516 -4101
rect 503 -4116 507 -4113
rect 503 -4120 518 -4116
rect 481 -4133 496 -4129
rect 148 -4558 152 -4554
rect 165 -4558 169 -4554
rect 185 -4558 189 -4554
rect 206 -4558 210 -4554
rect 227 -4558 231 -4554
rect 248 -4558 252 -4554
rect 269 -4558 273 -4554
rect 290 -4558 294 -4554
rect 311 -4558 315 -4554
rect 331 -4558 335 -4554
rect 139 -4613 143 -4566
rect 139 -4634 143 -4617
rect 157 -4627 161 -4566
rect 173 -4627 177 -4566
rect 197 -4606 201 -4566
rect 197 -4627 201 -4610
rect 215 -4627 219 -4566
rect 239 -4613 243 -4566
rect 239 -4627 243 -4617
rect 257 -4606 261 -4566
rect 257 -4627 261 -4610
rect 281 -4620 285 -4566
rect 299 -4598 303 -4566
rect 299 -4606 303 -4602
rect 281 -4627 285 -4624
rect 157 -4631 166 -4627
rect 173 -4631 181 -4627
rect 157 -4634 161 -4631
rect 181 -4634 185 -4631
rect 189 -4631 201 -4627
rect 215 -4631 223 -4627
rect 189 -4634 193 -4631
rect 223 -4634 227 -4631
rect 231 -4631 243 -4627
rect 257 -4631 269 -4627
rect 231 -4634 235 -4631
rect 265 -4634 269 -4631
rect 273 -4631 285 -4627
rect 299 -4627 303 -4610
rect 323 -4613 327 -4566
rect 323 -4627 327 -4617
rect 299 -4631 311 -4627
rect 273 -4634 277 -4631
rect 307 -4634 311 -4631
rect 315 -4631 327 -4627
rect 315 -4634 319 -4631
rect 148 -4642 152 -4638
rect 165 -4642 169 -4638
rect 206 -4642 210 -4638
rect 248 -4642 252 -4638
rect 290 -4642 294 -4638
rect 331 -4642 335 -4638
rect 348 -4651 352 -4602
rect 465 -4606 469 -4366
rect 148 -4729 152 -4725
rect 165 -4729 169 -4725
rect 185 -4729 189 -4725
rect 206 -4729 210 -4725
rect 227 -4729 231 -4725
rect 248 -4729 252 -4725
rect 269 -4729 273 -4725
rect 290 -4729 294 -4725
rect 311 -4729 315 -4725
rect 331 -4729 335 -4725
rect 139 -4784 143 -4737
rect 139 -4805 143 -4788
rect 157 -4798 161 -4737
rect 173 -4798 177 -4737
rect 197 -4777 201 -4737
rect 197 -4798 201 -4781
rect 215 -4798 219 -4737
rect 239 -4784 243 -4737
rect 239 -4798 243 -4788
rect 257 -4777 261 -4737
rect 257 -4798 261 -4781
rect 281 -4791 285 -4737
rect 299 -4769 303 -4737
rect 299 -4777 303 -4773
rect 281 -4798 285 -4795
rect 157 -4802 166 -4798
rect 173 -4802 181 -4798
rect 157 -4805 161 -4802
rect 181 -4805 185 -4802
rect 189 -4802 201 -4798
rect 215 -4802 223 -4798
rect 189 -4805 193 -4802
rect 223 -4805 227 -4802
rect 231 -4802 243 -4798
rect 257 -4802 269 -4798
rect 231 -4805 235 -4802
rect 265 -4805 269 -4802
rect 273 -4802 285 -4798
rect 299 -4798 303 -4781
rect 323 -4784 327 -4737
rect 323 -4798 327 -4788
rect 299 -4802 311 -4798
rect 273 -4805 277 -4802
rect 307 -4805 311 -4802
rect 315 -4802 327 -4798
rect 315 -4805 319 -4802
rect 148 -4813 152 -4809
rect 165 -4813 169 -4809
rect 206 -4813 210 -4809
rect 248 -4813 252 -4809
rect 290 -4813 294 -4809
rect 331 -4813 335 -4809
rect 139 -4844 143 -4840
rect 156 -4844 160 -4840
rect 147 -4855 151 -4852
rect 147 -4859 162 -4855
rect 125 -4872 140 -4868
rect -210 -5293 -206 -5289
rect -193 -5293 -189 -5289
rect -173 -5293 -169 -5289
rect -152 -5293 -148 -5289
rect -131 -5293 -127 -5289
rect -110 -5293 -106 -5289
rect -89 -5293 -85 -5289
rect -68 -5293 -64 -5289
rect -47 -5293 -43 -5289
rect -27 -5293 -23 -5289
rect -219 -5348 -215 -5301
rect -219 -5369 -215 -5352
rect -201 -5362 -197 -5301
rect -185 -5362 -181 -5301
rect -161 -5341 -157 -5301
rect -161 -5362 -157 -5345
rect -143 -5362 -139 -5301
rect -119 -5348 -115 -5301
rect -119 -5362 -115 -5352
rect -101 -5341 -97 -5301
rect -101 -5362 -97 -5345
rect -77 -5355 -73 -5301
rect -59 -5333 -55 -5301
rect -59 -5341 -55 -5337
rect -77 -5362 -73 -5359
rect -201 -5366 -192 -5362
rect -185 -5366 -177 -5362
rect -201 -5369 -197 -5366
rect -177 -5369 -173 -5366
rect -169 -5366 -157 -5362
rect -143 -5366 -135 -5362
rect -169 -5369 -165 -5366
rect -135 -5369 -131 -5366
rect -127 -5366 -115 -5362
rect -101 -5366 -89 -5362
rect -127 -5369 -123 -5366
rect -93 -5369 -89 -5366
rect -85 -5366 -73 -5362
rect -59 -5362 -55 -5345
rect -35 -5348 -31 -5301
rect -35 -5362 -31 -5352
rect -59 -5366 -47 -5362
rect -85 -5369 -81 -5366
rect -51 -5369 -47 -5366
rect -43 -5366 -31 -5362
rect -43 -5369 -39 -5366
rect -210 -5377 -206 -5373
rect -193 -5377 -189 -5373
rect -152 -5377 -148 -5373
rect -110 -5377 -106 -5373
rect -68 -5377 -64 -5373
rect -27 -5377 -23 -5373
rect -7 -5384 -3 -5337
rect 108 -5341 112 -5098
rect -210 -5453 -206 -5449
rect -193 -5453 -189 -5449
rect -173 -5453 -169 -5449
rect -152 -5453 -148 -5449
rect -131 -5453 -127 -5449
rect -110 -5453 -106 -5449
rect -89 -5453 -85 -5449
rect -68 -5453 -64 -5449
rect -47 -5453 -43 -5449
rect -27 -5453 -23 -5449
rect -219 -5508 -215 -5461
rect -219 -5529 -215 -5512
rect -201 -5522 -197 -5461
rect -185 -5522 -181 -5461
rect -161 -5501 -157 -5461
rect -161 -5522 -157 -5505
rect -143 -5522 -139 -5461
rect -119 -5508 -115 -5461
rect -119 -5522 -115 -5512
rect -101 -5501 -97 -5461
rect -101 -5522 -97 -5505
rect -77 -5515 -73 -5461
rect -59 -5493 -55 -5461
rect -59 -5501 -55 -5497
rect -77 -5522 -73 -5519
rect -201 -5526 -192 -5522
rect -185 -5526 -177 -5522
rect -201 -5529 -197 -5526
rect -177 -5529 -173 -5526
rect -169 -5526 -157 -5522
rect -143 -5526 -135 -5522
rect -169 -5529 -165 -5526
rect -135 -5529 -131 -5526
rect -127 -5526 -115 -5522
rect -101 -5526 -89 -5522
rect -127 -5529 -123 -5526
rect -93 -5529 -89 -5526
rect -85 -5526 -73 -5522
rect -59 -5522 -55 -5505
rect -35 -5508 -31 -5461
rect -35 -5522 -31 -5512
rect -59 -5526 -47 -5522
rect -85 -5529 -81 -5526
rect -51 -5529 -47 -5526
rect -43 -5526 -31 -5522
rect -43 -5529 -39 -5526
rect -210 -5537 -206 -5533
rect -193 -5537 -189 -5533
rect -152 -5537 -148 -5533
rect -110 -5537 -106 -5533
rect -68 -5537 -64 -5533
rect -27 -5537 -23 -5533
rect -219 -5567 -215 -5563
rect -202 -5567 -198 -5563
rect -211 -5578 -207 -5575
rect -211 -5582 -196 -5578
rect -200 -5621 -196 -5582
rect -200 -5636 -196 -5625
rect -219 -5640 -196 -5636
rect -193 -5612 -189 -5575
rect -12 -5591 -8 -5497
rect -219 -5643 -215 -5640
rect -193 -5643 -189 -5616
rect -202 -5651 -198 -5647
rect -210 -5726 -206 -5722
rect -184 -5726 -180 -5722
rect -167 -5726 -163 -5722
rect -127 -5726 -123 -5722
rect -106 -5726 -102 -5722
rect -89 -5726 -85 -5722
rect -49 -5726 -45 -5722
rect -25 -5726 -21 -5722
rect 12 -5726 16 -5722
rect -219 -5751 -215 -5734
rect -219 -5802 -215 -5755
rect -201 -5744 -197 -5734
rect -201 -5802 -197 -5748
rect -193 -5773 -189 -5734
rect -175 -5766 -171 -5734
rect -193 -5802 -189 -5777
rect -175 -5802 -171 -5770
rect -149 -5758 -145 -5734
rect -149 -5795 -145 -5762
rect -115 -5795 -111 -5734
rect -97 -5751 -93 -5734
rect -167 -5802 -163 -5799
rect -159 -5799 -145 -5795
rect -159 -5802 -155 -5799
rect -131 -5802 -127 -5799
rect -123 -5799 -104 -5795
rect -123 -5802 -119 -5799
rect -97 -5802 -93 -5755
rect -71 -5766 -67 -5734
rect -71 -5795 -67 -5770
rect -37 -5788 -33 -5734
rect -37 -5792 -20 -5788
rect -89 -5802 -85 -5799
rect -80 -5799 -67 -5795
rect -80 -5802 -76 -5799
rect -53 -5802 -49 -5799
rect -29 -5802 -25 -5792
rect -13 -5795 -9 -5734
rect -5 -5788 -1 -5734
rect 21 -5758 25 -5734
rect -5 -5792 14 -5788
rect -21 -5799 -4 -5795
rect -21 -5802 -17 -5799
rect 3 -5802 7 -5792
rect 21 -5802 25 -5762
rect -210 -5810 -206 -5806
rect -184 -5810 -180 -5806
rect -141 -5810 -137 -5806
rect -106 -5810 -102 -5806
rect -62 -5810 -58 -5806
rect -45 -5810 -41 -5806
rect -9 -5810 -5 -5806
rect 12 -5810 16 -5806
rect 33 -5817 37 -5770
rect 97 -5773 101 -5616
rect 108 -5758 112 -5388
rect 125 -5501 129 -4872
rect 158 -4898 162 -4859
rect 158 -4913 162 -4902
rect 139 -4917 162 -4913
rect 165 -4889 169 -4852
rect 347 -4868 351 -4773
rect 139 -4920 143 -4917
rect 165 -4920 169 -4893
rect 156 -4928 160 -4924
rect 148 -5003 152 -4999
rect 174 -5003 178 -4999
rect 191 -5003 195 -4999
rect 231 -5003 235 -4999
rect 252 -5003 256 -4999
rect 269 -5003 273 -4999
rect 309 -5003 313 -4999
rect 333 -5003 337 -4999
rect 370 -5003 374 -4999
rect 139 -5028 143 -5011
rect 139 -5079 143 -5032
rect 157 -5021 161 -5011
rect 157 -5079 161 -5025
rect 165 -5050 169 -5011
rect 183 -5043 187 -5011
rect 165 -5079 169 -5054
rect 183 -5079 187 -5047
rect 209 -5035 213 -5011
rect 209 -5072 213 -5039
rect 243 -5072 247 -5011
rect 261 -5028 265 -5011
rect 191 -5079 195 -5076
rect 199 -5076 213 -5072
rect 199 -5079 203 -5076
rect 227 -5079 231 -5076
rect 235 -5076 254 -5072
rect 235 -5079 239 -5076
rect 261 -5079 265 -5032
rect 287 -5043 291 -5011
rect 287 -5072 291 -5047
rect 321 -5065 325 -5011
rect 321 -5069 338 -5065
rect 269 -5079 273 -5076
rect 278 -5076 291 -5072
rect 278 -5079 282 -5076
rect 305 -5079 309 -5076
rect 329 -5079 333 -5069
rect 345 -5072 349 -5011
rect 353 -5065 357 -5011
rect 379 -5035 383 -5011
rect 353 -5069 372 -5065
rect 337 -5076 354 -5072
rect 337 -5079 341 -5076
rect 361 -5079 365 -5069
rect 379 -5079 383 -5039
rect 148 -5087 152 -5083
rect 174 -5087 178 -5083
rect 217 -5087 221 -5083
rect 252 -5087 256 -5083
rect 296 -5087 300 -5083
rect 313 -5087 317 -5083
rect 349 -5087 353 -5083
rect 370 -5087 374 -5083
rect 388 -5101 392 -5047
rect 451 -5050 455 -4893
rect 465 -5035 469 -4654
rect 481 -4777 485 -4133
rect 514 -4159 518 -4120
rect 514 -4174 518 -4163
rect 495 -4178 518 -4174
rect 521 -4150 525 -4113
rect 705 -4129 709 -4034
rect 495 -4181 499 -4178
rect 521 -4181 525 -4154
rect 512 -4189 516 -4185
rect 504 -4264 508 -4260
rect 530 -4264 534 -4260
rect 547 -4264 551 -4260
rect 587 -4264 591 -4260
rect 608 -4264 612 -4260
rect 625 -4264 629 -4260
rect 665 -4264 669 -4260
rect 689 -4264 693 -4260
rect 726 -4264 730 -4260
rect 495 -4289 499 -4272
rect 495 -4340 499 -4293
rect 513 -4282 517 -4272
rect 513 -4340 517 -4286
rect 521 -4311 525 -4272
rect 539 -4304 543 -4272
rect 521 -4340 525 -4315
rect 539 -4340 543 -4308
rect 565 -4296 569 -4272
rect 565 -4333 569 -4300
rect 599 -4333 603 -4272
rect 617 -4289 621 -4272
rect 547 -4340 551 -4337
rect 555 -4337 569 -4333
rect 555 -4340 559 -4337
rect 583 -4340 587 -4337
rect 591 -4337 610 -4333
rect 591 -4340 595 -4337
rect 617 -4340 621 -4293
rect 643 -4304 647 -4272
rect 643 -4333 647 -4308
rect 677 -4326 681 -4272
rect 677 -4330 694 -4326
rect 625 -4340 629 -4337
rect 634 -4337 647 -4333
rect 634 -4340 638 -4337
rect 661 -4340 665 -4337
rect 685 -4340 689 -4330
rect 701 -4333 705 -4272
rect 709 -4326 713 -4272
rect 735 -4296 739 -4272
rect 709 -4330 728 -4326
rect 693 -4337 710 -4333
rect 693 -4340 697 -4337
rect 717 -4340 721 -4330
rect 735 -4340 739 -4300
rect 504 -4348 508 -4344
rect 530 -4348 534 -4344
rect 573 -4348 577 -4344
rect 608 -4348 612 -4344
rect 652 -4348 656 -4344
rect 669 -4348 673 -4344
rect 705 -4348 709 -4344
rect 726 -4348 730 -4344
rect 743 -4355 747 -4308
rect 810 -4311 814 -4154
rect 824 -4296 828 -3910
rect 839 -4038 843 -3383
rect 872 -3409 876 -3370
rect 872 -3424 876 -3413
rect 853 -3428 876 -3424
rect 879 -3400 883 -3363
rect 1066 -3379 1070 -3288
rect 853 -3431 857 -3428
rect 879 -3431 883 -3404
rect 870 -3439 874 -3435
rect 862 -3514 866 -3510
rect 888 -3514 892 -3510
rect 905 -3514 909 -3510
rect 945 -3514 949 -3510
rect 966 -3514 970 -3510
rect 983 -3514 987 -3510
rect 1023 -3514 1027 -3510
rect 1047 -3514 1051 -3510
rect 1084 -3514 1088 -3510
rect 853 -3539 857 -3522
rect 853 -3590 857 -3543
rect 871 -3532 875 -3522
rect 871 -3590 875 -3536
rect 879 -3561 883 -3522
rect 897 -3554 901 -3522
rect 879 -3590 883 -3565
rect 897 -3590 901 -3558
rect 923 -3546 927 -3522
rect 923 -3583 927 -3550
rect 957 -3583 961 -3522
rect 975 -3539 979 -3522
rect 905 -3590 909 -3587
rect 913 -3587 927 -3583
rect 913 -3590 917 -3587
rect 941 -3590 945 -3587
rect 949 -3587 968 -3583
rect 949 -3590 953 -3587
rect 975 -3590 979 -3543
rect 1001 -3554 1005 -3522
rect 1001 -3583 1005 -3558
rect 1035 -3576 1039 -3522
rect 1035 -3580 1052 -3576
rect 983 -3590 987 -3587
rect 992 -3587 1005 -3583
rect 992 -3590 996 -3587
rect 1019 -3590 1023 -3587
rect 1043 -3590 1047 -3580
rect 1059 -3583 1063 -3522
rect 1067 -3576 1071 -3522
rect 1093 -3544 1097 -3522
rect 1067 -3580 1086 -3576
rect 1051 -3587 1068 -3583
rect 1051 -3590 1055 -3587
rect 1075 -3590 1079 -3580
rect 1093 -3590 1097 -3548
rect 1167 -3546 1171 -3404
rect 862 -3598 866 -3594
rect 888 -3598 892 -3594
rect 931 -3598 935 -3594
rect 966 -3598 970 -3594
rect 1010 -3598 1014 -3594
rect 1027 -3598 1031 -3594
rect 1063 -3598 1067 -3594
rect 1084 -3598 1088 -3594
rect 1101 -3612 1105 -3558
rect 1184 -3561 1188 -3169
rect 1197 -3292 1201 -2652
rect 1230 -2678 1234 -2639
rect 1230 -2693 1234 -2682
rect 1211 -2697 1234 -2693
rect 1237 -2669 1241 -2632
rect 1419 -2648 1423 -2563
rect 1211 -2700 1215 -2697
rect 1237 -2700 1241 -2673
rect 1228 -2708 1232 -2704
rect 1220 -2783 1224 -2779
rect 1246 -2783 1250 -2779
rect 1263 -2783 1267 -2779
rect 1303 -2783 1307 -2779
rect 1324 -2783 1328 -2779
rect 1341 -2783 1345 -2779
rect 1381 -2783 1385 -2779
rect 1405 -2783 1409 -2779
rect 1442 -2783 1446 -2779
rect 1211 -2808 1215 -2791
rect 1211 -2859 1215 -2812
rect 1229 -2801 1233 -2791
rect 1229 -2859 1233 -2805
rect 1237 -2830 1241 -2791
rect 1255 -2823 1259 -2791
rect 1237 -2859 1241 -2834
rect 1255 -2859 1259 -2827
rect 1281 -2815 1285 -2791
rect 1281 -2852 1285 -2819
rect 1315 -2852 1319 -2791
rect 1333 -2808 1337 -2791
rect 1263 -2859 1267 -2856
rect 1271 -2856 1285 -2852
rect 1271 -2859 1275 -2856
rect 1299 -2859 1303 -2856
rect 1307 -2856 1326 -2852
rect 1307 -2859 1311 -2856
rect 1333 -2859 1337 -2812
rect 1359 -2823 1363 -2791
rect 1359 -2852 1363 -2827
rect 1393 -2845 1397 -2791
rect 1393 -2849 1410 -2845
rect 1341 -2859 1345 -2856
rect 1350 -2856 1363 -2852
rect 1350 -2859 1354 -2856
rect 1377 -2859 1381 -2856
rect 1401 -2859 1405 -2849
rect 1417 -2852 1421 -2791
rect 1425 -2845 1429 -2791
rect 1425 -2849 1444 -2845
rect 1409 -2856 1426 -2852
rect 1409 -2859 1413 -2856
rect 1433 -2859 1437 -2849
rect 1451 -2859 1455 -2791
rect 1220 -2867 1224 -2863
rect 1246 -2867 1250 -2863
rect 1289 -2867 1293 -2863
rect 1324 -2867 1328 -2863
rect 1368 -2867 1372 -2863
rect 1385 -2867 1389 -2863
rect 1421 -2867 1425 -2863
rect 1442 -2867 1446 -2863
rect 1451 -2881 1455 -2863
rect 1467 -2874 1471 -2827
rect 1220 -3073 1224 -3069
rect 1237 -3073 1241 -3069
rect 1257 -3073 1261 -3069
rect 1278 -3073 1282 -3069
rect 1299 -3073 1303 -3069
rect 1320 -3073 1324 -3069
rect 1341 -3073 1345 -3069
rect 1362 -3073 1366 -3069
rect 1383 -3073 1387 -3069
rect 1403 -3073 1407 -3069
rect 1211 -3128 1215 -3081
rect 1211 -3149 1215 -3132
rect 1229 -3142 1233 -3081
rect 1245 -3142 1249 -3081
rect 1269 -3121 1273 -3081
rect 1269 -3142 1273 -3125
rect 1287 -3142 1291 -3081
rect 1311 -3128 1315 -3081
rect 1311 -3142 1315 -3132
rect 1329 -3121 1333 -3081
rect 1329 -3142 1333 -3125
rect 1353 -3135 1357 -3081
rect 1371 -3113 1375 -3081
rect 1371 -3121 1375 -3117
rect 1353 -3142 1357 -3139
rect 1229 -3146 1238 -3142
rect 1245 -3146 1253 -3142
rect 1229 -3149 1233 -3146
rect 1253 -3149 1257 -3146
rect 1261 -3146 1273 -3142
rect 1287 -3146 1295 -3142
rect 1261 -3149 1265 -3146
rect 1295 -3149 1299 -3146
rect 1303 -3146 1315 -3142
rect 1329 -3146 1341 -3142
rect 1303 -3149 1307 -3146
rect 1337 -3149 1341 -3146
rect 1345 -3146 1357 -3142
rect 1371 -3142 1375 -3125
rect 1395 -3128 1399 -3081
rect 1395 -3142 1399 -3132
rect 1371 -3146 1383 -3142
rect 1345 -3149 1349 -3146
rect 1379 -3149 1383 -3146
rect 1387 -3146 1399 -3142
rect 1387 -3149 1391 -3146
rect 1220 -3157 1224 -3153
rect 1237 -3157 1241 -3153
rect 1278 -3157 1282 -3153
rect 1320 -3157 1324 -3153
rect 1362 -3157 1366 -3153
rect 1403 -3157 1407 -3153
rect 1419 -3165 1423 -3117
rect 1220 -3244 1224 -3240
rect 1237 -3244 1241 -3240
rect 1257 -3244 1261 -3240
rect 1278 -3244 1282 -3240
rect 1299 -3244 1303 -3240
rect 1320 -3244 1324 -3240
rect 1341 -3244 1345 -3240
rect 1362 -3244 1366 -3240
rect 1383 -3244 1387 -3240
rect 1403 -3244 1407 -3240
rect 1211 -3299 1215 -3252
rect 1211 -3320 1215 -3303
rect 1229 -3313 1233 -3252
rect 1245 -3313 1249 -3252
rect 1269 -3292 1273 -3252
rect 1269 -3313 1273 -3296
rect 1287 -3313 1291 -3252
rect 1311 -3299 1315 -3252
rect 1311 -3313 1315 -3303
rect 1329 -3292 1333 -3252
rect 1329 -3313 1333 -3296
rect 1353 -3306 1357 -3252
rect 1371 -3284 1375 -3252
rect 1371 -3292 1375 -3288
rect 1353 -3313 1357 -3310
rect 1229 -3317 1238 -3313
rect 1245 -3317 1253 -3313
rect 1229 -3320 1233 -3317
rect 1253 -3320 1257 -3317
rect 1261 -3317 1273 -3313
rect 1287 -3317 1295 -3313
rect 1261 -3320 1265 -3317
rect 1295 -3320 1299 -3317
rect 1303 -3317 1315 -3313
rect 1329 -3317 1341 -3313
rect 1303 -3320 1307 -3317
rect 1337 -3320 1341 -3317
rect 1345 -3317 1357 -3313
rect 1371 -3313 1375 -3296
rect 1395 -3299 1399 -3252
rect 1395 -3313 1399 -3303
rect 1371 -3317 1383 -3313
rect 1345 -3320 1349 -3317
rect 1379 -3320 1383 -3317
rect 1387 -3317 1399 -3313
rect 1387 -3320 1391 -3317
rect 1220 -3328 1224 -3324
rect 1237 -3328 1241 -3324
rect 1278 -3328 1282 -3324
rect 1320 -3328 1324 -3324
rect 1362 -3328 1366 -3324
rect 1403 -3328 1407 -3324
rect 1211 -3355 1215 -3351
rect 1228 -3355 1232 -3351
rect 1219 -3366 1223 -3363
rect 1219 -3370 1234 -3366
rect 1197 -3383 1212 -3379
rect 862 -3815 866 -3811
rect 879 -3815 883 -3811
rect 899 -3815 903 -3811
rect 920 -3815 924 -3811
rect 941 -3815 945 -3811
rect 962 -3815 966 -3811
rect 983 -3815 987 -3811
rect 1004 -3815 1008 -3811
rect 1025 -3815 1029 -3811
rect 1045 -3815 1049 -3811
rect 853 -3870 857 -3823
rect 853 -3891 857 -3874
rect 871 -3884 875 -3823
rect 887 -3884 891 -3823
rect 911 -3863 915 -3823
rect 911 -3884 915 -3867
rect 929 -3884 933 -3823
rect 953 -3870 957 -3823
rect 953 -3884 957 -3874
rect 971 -3863 975 -3823
rect 971 -3884 975 -3867
rect 995 -3877 999 -3823
rect 1013 -3855 1017 -3823
rect 1013 -3863 1017 -3859
rect 995 -3884 999 -3881
rect 871 -3888 880 -3884
rect 887 -3888 895 -3884
rect 871 -3891 875 -3888
rect 895 -3891 899 -3888
rect 903 -3888 915 -3884
rect 929 -3888 937 -3884
rect 903 -3891 907 -3888
rect 937 -3891 941 -3888
rect 945 -3888 957 -3884
rect 971 -3888 983 -3884
rect 945 -3891 949 -3888
rect 979 -3891 983 -3888
rect 987 -3888 999 -3884
rect 1013 -3884 1017 -3867
rect 1037 -3870 1041 -3823
rect 1037 -3884 1041 -3874
rect 1013 -3888 1025 -3884
rect 987 -3891 991 -3888
rect 1021 -3891 1025 -3888
rect 1029 -3888 1041 -3884
rect 1029 -3891 1033 -3888
rect 862 -3899 866 -3895
rect 879 -3899 883 -3895
rect 920 -3899 924 -3895
rect 962 -3899 966 -3895
rect 1004 -3899 1008 -3895
rect 1045 -3899 1049 -3895
rect 1060 -3906 1064 -3859
rect 1184 -3863 1188 -3616
rect 862 -3990 866 -3986
rect 879 -3990 883 -3986
rect 899 -3990 903 -3986
rect 920 -3990 924 -3986
rect 941 -3990 945 -3986
rect 962 -3990 966 -3986
rect 983 -3990 987 -3986
rect 1004 -3990 1008 -3986
rect 1025 -3990 1029 -3986
rect 1045 -3990 1049 -3986
rect 853 -4045 857 -3998
rect 853 -4066 857 -4049
rect 871 -4059 875 -3998
rect 887 -4059 891 -3998
rect 911 -4038 915 -3998
rect 911 -4059 915 -4042
rect 929 -4059 933 -3998
rect 953 -4045 957 -3998
rect 953 -4059 957 -4049
rect 971 -4038 975 -3998
rect 971 -4059 975 -4042
rect 995 -4052 999 -3998
rect 1013 -4030 1017 -3998
rect 1013 -4038 1017 -4034
rect 995 -4059 999 -4056
rect 871 -4063 880 -4059
rect 887 -4063 895 -4059
rect 871 -4066 875 -4063
rect 895 -4066 899 -4063
rect 903 -4063 915 -4059
rect 929 -4063 937 -4059
rect 903 -4066 907 -4063
rect 937 -4066 941 -4063
rect 945 -4063 957 -4059
rect 971 -4063 983 -4059
rect 945 -4066 949 -4063
rect 979 -4066 983 -4063
rect 987 -4063 999 -4059
rect 1013 -4059 1017 -4042
rect 1037 -4045 1041 -3998
rect 1037 -4059 1041 -4049
rect 1013 -4063 1025 -4059
rect 987 -4066 991 -4063
rect 1021 -4066 1025 -4063
rect 1029 -4063 1041 -4059
rect 1029 -4066 1033 -4063
rect 862 -4074 866 -4070
rect 879 -4074 883 -4070
rect 920 -4074 924 -4070
rect 962 -4074 966 -4070
rect 1004 -4074 1008 -4070
rect 1045 -4074 1049 -4070
rect 853 -4105 857 -4101
rect 870 -4105 874 -4101
rect 861 -4116 865 -4113
rect 861 -4120 876 -4116
rect 839 -4133 854 -4129
rect 504 -4558 508 -4554
rect 521 -4558 525 -4554
rect 541 -4558 545 -4554
rect 562 -4558 566 -4554
rect 583 -4558 587 -4554
rect 604 -4558 608 -4554
rect 625 -4558 629 -4554
rect 646 -4558 650 -4554
rect 667 -4558 671 -4554
rect 687 -4558 691 -4554
rect 495 -4613 499 -4566
rect 495 -4634 499 -4617
rect 513 -4627 517 -4566
rect 529 -4627 533 -4566
rect 553 -4606 557 -4566
rect 553 -4627 557 -4610
rect 571 -4627 575 -4566
rect 595 -4613 599 -4566
rect 595 -4627 599 -4617
rect 613 -4606 617 -4566
rect 613 -4627 617 -4610
rect 637 -4620 641 -4566
rect 655 -4598 659 -4566
rect 655 -4606 659 -4602
rect 637 -4627 641 -4624
rect 513 -4631 522 -4627
rect 529 -4631 537 -4627
rect 513 -4634 517 -4631
rect 537 -4634 541 -4631
rect 545 -4631 557 -4627
rect 571 -4631 579 -4627
rect 545 -4634 549 -4631
rect 579 -4634 583 -4631
rect 587 -4631 599 -4627
rect 613 -4631 625 -4627
rect 587 -4634 591 -4631
rect 621 -4634 625 -4631
rect 629 -4631 641 -4627
rect 655 -4627 659 -4610
rect 679 -4613 683 -4566
rect 679 -4627 683 -4617
rect 655 -4631 667 -4627
rect 629 -4634 633 -4631
rect 663 -4634 667 -4631
rect 671 -4631 683 -4627
rect 671 -4634 675 -4631
rect 504 -4642 508 -4638
rect 521 -4642 525 -4638
rect 562 -4642 566 -4638
rect 604 -4642 608 -4638
rect 646 -4642 650 -4638
rect 687 -4642 691 -4638
rect 700 -4650 704 -4602
rect 824 -4606 828 -4359
rect 504 -4729 508 -4725
rect 521 -4729 525 -4725
rect 541 -4729 545 -4725
rect 562 -4729 566 -4725
rect 583 -4729 587 -4725
rect 604 -4729 608 -4725
rect 625 -4729 629 -4725
rect 646 -4729 650 -4725
rect 667 -4729 671 -4725
rect 687 -4729 691 -4725
rect 495 -4784 499 -4737
rect 495 -4805 499 -4788
rect 513 -4798 517 -4737
rect 529 -4798 533 -4737
rect 553 -4777 557 -4737
rect 553 -4798 557 -4781
rect 571 -4798 575 -4737
rect 595 -4784 599 -4737
rect 595 -4798 599 -4788
rect 613 -4777 617 -4737
rect 613 -4798 617 -4781
rect 637 -4791 641 -4737
rect 655 -4769 659 -4737
rect 655 -4777 659 -4773
rect 637 -4798 641 -4795
rect 513 -4802 522 -4798
rect 529 -4802 537 -4798
rect 513 -4805 517 -4802
rect 537 -4805 541 -4802
rect 545 -4802 557 -4798
rect 571 -4802 579 -4798
rect 545 -4805 549 -4802
rect 579 -4805 583 -4802
rect 587 -4802 599 -4798
rect 613 -4802 625 -4798
rect 587 -4805 591 -4802
rect 621 -4805 625 -4802
rect 629 -4802 641 -4798
rect 655 -4798 659 -4781
rect 679 -4784 683 -4737
rect 679 -4798 683 -4788
rect 655 -4802 667 -4798
rect 629 -4805 633 -4802
rect 663 -4805 667 -4802
rect 671 -4802 683 -4798
rect 671 -4805 675 -4802
rect 504 -4813 508 -4809
rect 521 -4813 525 -4809
rect 562 -4813 566 -4809
rect 604 -4813 608 -4809
rect 646 -4813 650 -4809
rect 687 -4813 691 -4809
rect 495 -4844 499 -4840
rect 512 -4844 516 -4840
rect 503 -4855 507 -4852
rect 503 -4859 518 -4855
rect 481 -4872 496 -4868
rect 148 -5293 152 -5289
rect 165 -5293 169 -5289
rect 185 -5293 189 -5289
rect 206 -5293 210 -5289
rect 227 -5293 231 -5289
rect 248 -5293 252 -5289
rect 269 -5293 273 -5289
rect 290 -5293 294 -5289
rect 311 -5293 315 -5289
rect 331 -5293 335 -5289
rect 139 -5348 143 -5301
rect 139 -5369 143 -5352
rect 157 -5362 161 -5301
rect 173 -5362 177 -5301
rect 197 -5341 201 -5301
rect 197 -5362 201 -5345
rect 215 -5362 219 -5301
rect 239 -5348 243 -5301
rect 239 -5362 243 -5352
rect 257 -5341 261 -5301
rect 257 -5362 261 -5345
rect 281 -5355 285 -5301
rect 299 -5333 303 -5301
rect 299 -5341 303 -5337
rect 281 -5362 285 -5359
rect 157 -5366 166 -5362
rect 173 -5366 181 -5362
rect 157 -5369 161 -5366
rect 181 -5369 185 -5366
rect 189 -5366 201 -5362
rect 215 -5366 223 -5362
rect 189 -5369 193 -5366
rect 223 -5369 227 -5366
rect 231 -5366 243 -5362
rect 257 -5366 269 -5362
rect 231 -5369 235 -5366
rect 265 -5369 269 -5366
rect 273 -5366 285 -5362
rect 299 -5362 303 -5345
rect 323 -5348 327 -5301
rect 323 -5362 327 -5352
rect 299 -5366 311 -5362
rect 273 -5369 277 -5366
rect 307 -5369 311 -5366
rect 315 -5366 327 -5362
rect 315 -5369 319 -5366
rect 148 -5377 152 -5373
rect 165 -5377 169 -5373
rect 206 -5377 210 -5373
rect 248 -5377 252 -5373
rect 290 -5377 294 -5373
rect 331 -5377 335 -5373
rect 349 -5384 353 -5337
rect 464 -5341 468 -5105
rect 148 -5453 152 -5449
rect 165 -5453 169 -5449
rect 185 -5453 189 -5449
rect 206 -5453 210 -5449
rect 227 -5453 231 -5449
rect 248 -5453 252 -5449
rect 269 -5453 273 -5449
rect 290 -5453 294 -5449
rect 311 -5453 315 -5449
rect 331 -5453 335 -5449
rect 139 -5508 143 -5461
rect 139 -5529 143 -5512
rect 157 -5522 161 -5461
rect 173 -5522 177 -5461
rect 197 -5501 201 -5461
rect 197 -5522 201 -5505
rect 215 -5522 219 -5461
rect 239 -5508 243 -5461
rect 239 -5522 243 -5512
rect 257 -5501 261 -5461
rect 257 -5522 261 -5505
rect 281 -5515 285 -5461
rect 299 -5493 303 -5461
rect 299 -5501 303 -5497
rect 281 -5522 285 -5519
rect 157 -5526 166 -5522
rect 173 -5526 181 -5522
rect 157 -5529 161 -5526
rect 181 -5529 185 -5526
rect 189 -5526 201 -5522
rect 215 -5526 223 -5522
rect 189 -5529 193 -5526
rect 223 -5529 227 -5526
rect 231 -5526 243 -5522
rect 257 -5526 269 -5522
rect 231 -5529 235 -5526
rect 265 -5529 269 -5526
rect 273 -5526 285 -5522
rect 299 -5522 303 -5505
rect 323 -5508 327 -5461
rect 323 -5522 327 -5512
rect 299 -5526 311 -5522
rect 273 -5529 277 -5526
rect 307 -5529 311 -5526
rect 315 -5526 327 -5522
rect 315 -5529 319 -5526
rect 148 -5537 152 -5533
rect 165 -5537 169 -5533
rect 206 -5537 210 -5533
rect 248 -5537 252 -5533
rect 290 -5537 294 -5533
rect 331 -5537 335 -5533
rect 139 -5567 143 -5563
rect 156 -5567 160 -5563
rect 147 -5578 151 -5575
rect 147 -5582 162 -5578
rect 158 -5621 162 -5582
rect 158 -5636 162 -5625
rect 139 -5640 162 -5636
rect 165 -5612 169 -5575
rect 348 -5591 352 -5497
rect 139 -5643 143 -5640
rect 165 -5643 169 -5616
rect 156 -5651 160 -5647
rect 148 -5726 152 -5722
rect 174 -5726 178 -5722
rect 191 -5726 195 -5722
rect 231 -5726 235 -5722
rect 252 -5726 256 -5722
rect 269 -5726 273 -5722
rect 309 -5726 313 -5722
rect 333 -5726 337 -5722
rect 370 -5726 374 -5722
rect 139 -5751 143 -5734
rect 139 -5802 143 -5755
rect 157 -5744 161 -5734
rect 157 -5802 161 -5748
rect 165 -5773 169 -5734
rect 183 -5766 187 -5734
rect 165 -5802 169 -5777
rect 183 -5802 187 -5770
rect 209 -5758 213 -5734
rect 209 -5795 213 -5762
rect 243 -5795 247 -5734
rect 261 -5751 265 -5734
rect 191 -5802 195 -5799
rect 199 -5799 213 -5795
rect 199 -5802 203 -5799
rect 227 -5802 231 -5799
rect 235 -5799 254 -5795
rect 235 -5802 239 -5799
rect 261 -5802 265 -5755
rect 287 -5766 291 -5734
rect 287 -5795 291 -5770
rect 321 -5788 325 -5734
rect 321 -5792 338 -5788
rect 269 -5802 273 -5799
rect 278 -5799 291 -5795
rect 278 -5802 282 -5799
rect 305 -5802 309 -5799
rect 329 -5802 333 -5792
rect 345 -5795 349 -5734
rect 353 -5788 357 -5734
rect 379 -5758 383 -5734
rect 353 -5792 372 -5788
rect 337 -5799 354 -5795
rect 337 -5802 341 -5799
rect 361 -5802 365 -5792
rect 379 -5802 383 -5762
rect 148 -5810 152 -5806
rect 174 -5810 178 -5806
rect 217 -5810 221 -5806
rect 252 -5810 256 -5806
rect 296 -5810 300 -5806
rect 313 -5810 317 -5806
rect 349 -5810 353 -5806
rect 370 -5810 374 -5806
rect 392 -5818 396 -5770
rect 451 -5773 455 -5616
rect 464 -5758 468 -5390
rect 481 -5501 485 -4872
rect 514 -4898 518 -4859
rect 514 -4913 518 -4902
rect 495 -4917 518 -4913
rect 521 -4889 525 -4852
rect 706 -4868 710 -4773
rect 495 -4920 499 -4917
rect 521 -4920 525 -4893
rect 512 -4928 516 -4924
rect 504 -5003 508 -4999
rect 530 -5003 534 -4999
rect 547 -5003 551 -4999
rect 587 -5003 591 -4999
rect 608 -5003 612 -4999
rect 625 -5003 629 -4999
rect 665 -5003 669 -4999
rect 689 -5003 693 -4999
rect 726 -5003 730 -4999
rect 495 -5028 499 -5011
rect 495 -5079 499 -5032
rect 513 -5021 517 -5011
rect 513 -5079 517 -5025
rect 521 -5050 525 -5011
rect 539 -5043 543 -5011
rect 521 -5079 525 -5054
rect 539 -5079 543 -5047
rect 565 -5035 569 -5011
rect 565 -5072 569 -5039
rect 599 -5072 603 -5011
rect 617 -5028 621 -5011
rect 547 -5079 551 -5076
rect 555 -5076 569 -5072
rect 555 -5079 559 -5076
rect 583 -5079 587 -5076
rect 591 -5076 610 -5072
rect 591 -5079 595 -5076
rect 617 -5079 621 -5032
rect 643 -5043 647 -5011
rect 643 -5072 647 -5047
rect 677 -5065 681 -5011
rect 677 -5069 694 -5065
rect 625 -5079 629 -5076
rect 634 -5076 647 -5072
rect 634 -5079 638 -5076
rect 661 -5079 665 -5076
rect 685 -5079 689 -5069
rect 701 -5072 705 -5011
rect 709 -5065 713 -5011
rect 735 -5035 739 -5011
rect 709 -5069 728 -5065
rect 693 -5076 710 -5072
rect 693 -5079 697 -5076
rect 717 -5079 721 -5069
rect 735 -5079 739 -5039
rect 504 -5087 508 -5083
rect 530 -5087 534 -5083
rect 573 -5087 577 -5083
rect 608 -5087 612 -5083
rect 652 -5087 656 -5083
rect 669 -5087 673 -5083
rect 705 -5087 709 -5083
rect 726 -5087 730 -5083
rect 743 -5094 747 -5047
rect 810 -5050 814 -4893
rect 824 -5035 828 -4653
rect 839 -4777 843 -4133
rect 872 -4159 876 -4120
rect 872 -4174 876 -4163
rect 853 -4178 876 -4174
rect 879 -4150 883 -4113
rect 1063 -4129 1067 -4034
rect 853 -4181 857 -4178
rect 879 -4181 883 -4154
rect 870 -4189 874 -4185
rect 862 -4264 866 -4260
rect 888 -4264 892 -4260
rect 905 -4264 909 -4260
rect 945 -4264 949 -4260
rect 966 -4264 970 -4260
rect 983 -4264 987 -4260
rect 1023 -4264 1027 -4260
rect 1047 -4264 1051 -4260
rect 1084 -4264 1088 -4260
rect 853 -4289 857 -4272
rect 853 -4340 857 -4293
rect 871 -4282 875 -4272
rect 871 -4340 875 -4286
rect 879 -4311 883 -4272
rect 897 -4304 901 -4272
rect 879 -4340 883 -4315
rect 897 -4340 901 -4308
rect 923 -4296 927 -4272
rect 923 -4333 927 -4300
rect 957 -4333 961 -4272
rect 975 -4289 979 -4272
rect 905 -4340 909 -4337
rect 913 -4337 927 -4333
rect 913 -4340 917 -4337
rect 941 -4340 945 -4337
rect 949 -4337 968 -4333
rect 949 -4340 953 -4337
rect 975 -4340 979 -4293
rect 1001 -4304 1005 -4272
rect 1001 -4333 1005 -4308
rect 1035 -4326 1039 -4272
rect 1035 -4330 1052 -4326
rect 983 -4340 987 -4337
rect 992 -4337 1005 -4333
rect 992 -4340 996 -4337
rect 1019 -4340 1023 -4337
rect 1043 -4340 1047 -4330
rect 1059 -4333 1063 -4272
rect 1067 -4326 1071 -4272
rect 1093 -4294 1097 -4272
rect 1067 -4330 1086 -4326
rect 1051 -4337 1068 -4333
rect 1051 -4340 1055 -4337
rect 1075 -4340 1079 -4330
rect 1093 -4340 1097 -4298
rect 1167 -4296 1171 -4154
rect 862 -4348 866 -4344
rect 888 -4348 892 -4344
rect 931 -4348 935 -4344
rect 966 -4348 970 -4344
rect 1010 -4348 1014 -4344
rect 1027 -4348 1031 -4344
rect 1063 -4348 1067 -4344
rect 1084 -4348 1088 -4344
rect 1101 -4362 1105 -4308
rect 1184 -4311 1188 -3910
rect 1197 -4038 1201 -3383
rect 1230 -3409 1234 -3370
rect 1230 -3424 1234 -3413
rect 1211 -3428 1234 -3424
rect 1237 -3400 1241 -3363
rect 1422 -3379 1426 -3288
rect 1211 -3431 1215 -3428
rect 1237 -3431 1241 -3404
rect 1228 -3439 1232 -3435
rect 1220 -3514 1224 -3510
rect 1246 -3514 1250 -3510
rect 1263 -3514 1267 -3510
rect 1303 -3514 1307 -3510
rect 1324 -3514 1328 -3510
rect 1341 -3514 1345 -3510
rect 1381 -3514 1385 -3510
rect 1405 -3514 1409 -3510
rect 1442 -3514 1446 -3510
rect 1211 -3539 1215 -3522
rect 1211 -3590 1215 -3543
rect 1229 -3532 1233 -3522
rect 1229 -3590 1233 -3536
rect 1237 -3561 1241 -3522
rect 1255 -3554 1259 -3522
rect 1237 -3590 1241 -3565
rect 1255 -3590 1259 -3558
rect 1281 -3546 1285 -3522
rect 1281 -3583 1285 -3550
rect 1315 -3583 1319 -3522
rect 1333 -3539 1337 -3522
rect 1263 -3590 1267 -3587
rect 1271 -3587 1285 -3583
rect 1271 -3590 1275 -3587
rect 1299 -3590 1303 -3587
rect 1307 -3587 1326 -3583
rect 1307 -3590 1311 -3587
rect 1333 -3590 1337 -3543
rect 1359 -3554 1363 -3522
rect 1359 -3583 1363 -3558
rect 1393 -3576 1397 -3522
rect 1393 -3580 1410 -3576
rect 1341 -3590 1345 -3587
rect 1350 -3587 1363 -3583
rect 1350 -3590 1354 -3587
rect 1377 -3590 1381 -3587
rect 1401 -3590 1405 -3580
rect 1417 -3583 1421 -3522
rect 1425 -3576 1429 -3522
rect 1425 -3580 1444 -3576
rect 1409 -3587 1426 -3583
rect 1409 -3590 1413 -3587
rect 1433 -3590 1437 -3580
rect 1451 -3590 1455 -3522
rect 1220 -3598 1224 -3594
rect 1246 -3598 1250 -3594
rect 1289 -3598 1293 -3594
rect 1324 -3598 1328 -3594
rect 1368 -3598 1372 -3594
rect 1385 -3598 1389 -3594
rect 1421 -3598 1425 -3594
rect 1442 -3598 1446 -3594
rect 1451 -3612 1455 -3594
rect 1464 -3605 1468 -3558
rect 1220 -3815 1224 -3811
rect 1237 -3815 1241 -3811
rect 1257 -3815 1261 -3811
rect 1278 -3815 1282 -3811
rect 1299 -3815 1303 -3811
rect 1320 -3815 1324 -3811
rect 1341 -3815 1345 -3811
rect 1362 -3815 1366 -3811
rect 1383 -3815 1387 -3811
rect 1403 -3815 1407 -3811
rect 1211 -3870 1215 -3823
rect 1211 -3891 1215 -3874
rect 1229 -3884 1233 -3823
rect 1245 -3884 1249 -3823
rect 1269 -3863 1273 -3823
rect 1269 -3884 1273 -3867
rect 1287 -3884 1291 -3823
rect 1311 -3870 1315 -3823
rect 1311 -3884 1315 -3874
rect 1329 -3863 1333 -3823
rect 1329 -3884 1333 -3867
rect 1353 -3877 1357 -3823
rect 1371 -3855 1375 -3823
rect 1371 -3863 1375 -3859
rect 1353 -3884 1357 -3881
rect 1229 -3888 1238 -3884
rect 1245 -3888 1253 -3884
rect 1229 -3891 1233 -3888
rect 1253 -3891 1257 -3888
rect 1261 -3888 1273 -3884
rect 1287 -3888 1295 -3884
rect 1261 -3891 1265 -3888
rect 1295 -3891 1299 -3888
rect 1303 -3888 1315 -3884
rect 1329 -3888 1341 -3884
rect 1303 -3891 1307 -3888
rect 1337 -3891 1341 -3888
rect 1345 -3888 1357 -3884
rect 1371 -3884 1375 -3867
rect 1395 -3870 1399 -3823
rect 1395 -3884 1399 -3874
rect 1371 -3888 1383 -3884
rect 1345 -3891 1349 -3888
rect 1379 -3891 1383 -3888
rect 1387 -3888 1399 -3884
rect 1387 -3891 1391 -3888
rect 1220 -3899 1224 -3895
rect 1237 -3899 1241 -3895
rect 1278 -3899 1282 -3895
rect 1320 -3899 1324 -3895
rect 1362 -3899 1366 -3895
rect 1403 -3899 1407 -3895
rect 1424 -3906 1428 -3859
rect 1220 -3990 1224 -3986
rect 1237 -3990 1241 -3986
rect 1257 -3990 1261 -3986
rect 1278 -3990 1282 -3986
rect 1299 -3990 1303 -3986
rect 1320 -3990 1324 -3986
rect 1341 -3990 1345 -3986
rect 1362 -3990 1366 -3986
rect 1383 -3990 1387 -3986
rect 1403 -3990 1407 -3986
rect 1211 -4045 1215 -3998
rect 1211 -4066 1215 -4049
rect 1229 -4059 1233 -3998
rect 1245 -4059 1249 -3998
rect 1269 -4038 1273 -3998
rect 1269 -4059 1273 -4042
rect 1287 -4059 1291 -3998
rect 1311 -4045 1315 -3998
rect 1311 -4059 1315 -4049
rect 1329 -4038 1333 -3998
rect 1329 -4059 1333 -4042
rect 1353 -4052 1357 -3998
rect 1371 -4030 1375 -3998
rect 1371 -4038 1375 -4034
rect 1353 -4059 1357 -4056
rect 1229 -4063 1238 -4059
rect 1245 -4063 1253 -4059
rect 1229 -4066 1233 -4063
rect 1253 -4066 1257 -4063
rect 1261 -4063 1273 -4059
rect 1287 -4063 1295 -4059
rect 1261 -4066 1265 -4063
rect 1295 -4066 1299 -4063
rect 1303 -4063 1315 -4059
rect 1329 -4063 1341 -4059
rect 1303 -4066 1307 -4063
rect 1337 -4066 1341 -4063
rect 1345 -4063 1357 -4059
rect 1371 -4059 1375 -4042
rect 1395 -4045 1399 -3998
rect 1395 -4059 1399 -4049
rect 1371 -4063 1383 -4059
rect 1345 -4066 1349 -4063
rect 1379 -4066 1383 -4063
rect 1387 -4063 1399 -4059
rect 1387 -4066 1391 -4063
rect 1220 -4074 1224 -4070
rect 1237 -4074 1241 -4070
rect 1278 -4074 1282 -4070
rect 1320 -4074 1324 -4070
rect 1362 -4074 1366 -4070
rect 1403 -4074 1407 -4070
rect 1211 -4105 1215 -4101
rect 1228 -4105 1232 -4101
rect 1219 -4116 1223 -4113
rect 1219 -4120 1234 -4116
rect 1197 -4133 1212 -4129
rect 862 -4558 866 -4554
rect 879 -4558 883 -4554
rect 899 -4558 903 -4554
rect 920 -4558 924 -4554
rect 941 -4558 945 -4554
rect 962 -4558 966 -4554
rect 983 -4558 987 -4554
rect 1004 -4558 1008 -4554
rect 1025 -4558 1029 -4554
rect 1045 -4558 1049 -4554
rect 853 -4613 857 -4566
rect 853 -4634 857 -4617
rect 871 -4627 875 -4566
rect 887 -4627 891 -4566
rect 911 -4606 915 -4566
rect 911 -4627 915 -4610
rect 929 -4627 933 -4566
rect 953 -4613 957 -4566
rect 953 -4627 957 -4617
rect 971 -4606 975 -4566
rect 971 -4627 975 -4610
rect 995 -4620 999 -4566
rect 1013 -4598 1017 -4566
rect 1013 -4606 1017 -4602
rect 995 -4627 999 -4624
rect 871 -4631 880 -4627
rect 887 -4631 895 -4627
rect 871 -4634 875 -4631
rect 895 -4634 899 -4631
rect 903 -4631 915 -4627
rect 929 -4631 937 -4627
rect 903 -4634 907 -4631
rect 937 -4634 941 -4631
rect 945 -4631 957 -4627
rect 971 -4631 983 -4627
rect 945 -4634 949 -4631
rect 979 -4634 983 -4631
rect 987 -4631 999 -4627
rect 1013 -4627 1017 -4610
rect 1037 -4613 1041 -4566
rect 1037 -4627 1041 -4617
rect 1013 -4631 1025 -4627
rect 987 -4634 991 -4631
rect 1021 -4634 1025 -4631
rect 1029 -4631 1041 -4627
rect 1029 -4634 1033 -4631
rect 862 -4642 866 -4638
rect 879 -4642 883 -4638
rect 920 -4642 924 -4638
rect 962 -4642 966 -4638
rect 1004 -4642 1008 -4638
rect 1045 -4642 1049 -4638
rect 1059 -4649 1063 -4602
rect 1184 -4606 1188 -4366
rect 862 -4729 866 -4725
rect 879 -4729 883 -4725
rect 899 -4729 903 -4725
rect 920 -4729 924 -4725
rect 941 -4729 945 -4725
rect 962 -4729 966 -4725
rect 983 -4729 987 -4725
rect 1004 -4729 1008 -4725
rect 1025 -4729 1029 -4725
rect 1045 -4729 1049 -4725
rect 853 -4784 857 -4737
rect 853 -4805 857 -4788
rect 871 -4798 875 -4737
rect 887 -4798 891 -4737
rect 911 -4777 915 -4737
rect 911 -4798 915 -4781
rect 929 -4798 933 -4737
rect 953 -4784 957 -4737
rect 953 -4798 957 -4788
rect 971 -4777 975 -4737
rect 971 -4798 975 -4781
rect 995 -4791 999 -4737
rect 1013 -4769 1017 -4737
rect 1013 -4777 1017 -4773
rect 995 -4798 999 -4795
rect 871 -4802 880 -4798
rect 887 -4802 895 -4798
rect 871 -4805 875 -4802
rect 895 -4805 899 -4802
rect 903 -4802 915 -4798
rect 929 -4802 937 -4798
rect 903 -4805 907 -4802
rect 937 -4805 941 -4802
rect 945 -4802 957 -4798
rect 971 -4802 983 -4798
rect 945 -4805 949 -4802
rect 979 -4805 983 -4802
rect 987 -4802 999 -4798
rect 1013 -4798 1017 -4781
rect 1037 -4784 1041 -4737
rect 1037 -4798 1041 -4788
rect 1013 -4802 1025 -4798
rect 987 -4805 991 -4802
rect 1021 -4805 1025 -4802
rect 1029 -4802 1041 -4798
rect 1029 -4805 1033 -4802
rect 862 -4813 866 -4809
rect 879 -4813 883 -4809
rect 920 -4813 924 -4809
rect 962 -4813 966 -4809
rect 1004 -4813 1008 -4809
rect 1045 -4813 1049 -4809
rect 853 -4844 857 -4840
rect 870 -4844 874 -4840
rect 861 -4855 865 -4852
rect 861 -4859 876 -4855
rect 839 -4872 854 -4868
rect 504 -5293 508 -5289
rect 521 -5293 525 -5289
rect 541 -5293 545 -5289
rect 562 -5293 566 -5289
rect 583 -5293 587 -5289
rect 604 -5293 608 -5289
rect 625 -5293 629 -5289
rect 646 -5293 650 -5289
rect 667 -5293 671 -5289
rect 687 -5293 691 -5289
rect 495 -5348 499 -5301
rect 495 -5369 499 -5352
rect 513 -5362 517 -5301
rect 529 -5362 533 -5301
rect 553 -5341 557 -5301
rect 553 -5362 557 -5345
rect 571 -5362 575 -5301
rect 595 -5348 599 -5301
rect 595 -5362 599 -5352
rect 613 -5341 617 -5301
rect 613 -5362 617 -5345
rect 637 -5355 641 -5301
rect 655 -5333 659 -5301
rect 655 -5341 659 -5337
rect 637 -5362 641 -5359
rect 513 -5366 522 -5362
rect 529 -5366 537 -5362
rect 513 -5369 517 -5366
rect 537 -5369 541 -5366
rect 545 -5366 557 -5362
rect 571 -5366 579 -5362
rect 545 -5369 549 -5366
rect 579 -5369 583 -5366
rect 587 -5366 599 -5362
rect 613 -5366 625 -5362
rect 587 -5369 591 -5366
rect 621 -5369 625 -5366
rect 629 -5366 641 -5362
rect 655 -5362 659 -5345
rect 679 -5348 683 -5301
rect 679 -5362 683 -5352
rect 655 -5366 667 -5362
rect 629 -5369 633 -5366
rect 663 -5369 667 -5366
rect 671 -5366 683 -5362
rect 671 -5369 675 -5366
rect 504 -5377 508 -5373
rect 521 -5377 525 -5373
rect 562 -5377 566 -5373
rect 604 -5377 608 -5373
rect 646 -5377 650 -5373
rect 687 -5377 691 -5373
rect 705 -5386 709 -5337
rect 822 -5341 826 -5098
rect 504 -5453 508 -5449
rect 521 -5453 525 -5449
rect 541 -5453 545 -5449
rect 562 -5453 566 -5449
rect 583 -5453 587 -5449
rect 604 -5453 608 -5449
rect 625 -5453 629 -5449
rect 646 -5453 650 -5449
rect 667 -5453 671 -5449
rect 687 -5453 691 -5449
rect 495 -5508 499 -5461
rect 495 -5529 499 -5512
rect 513 -5522 517 -5461
rect 529 -5522 533 -5461
rect 553 -5501 557 -5461
rect 553 -5522 557 -5505
rect 571 -5522 575 -5461
rect 595 -5508 599 -5461
rect 595 -5522 599 -5512
rect 613 -5501 617 -5461
rect 613 -5522 617 -5505
rect 637 -5515 641 -5461
rect 655 -5493 659 -5461
rect 655 -5501 659 -5497
rect 637 -5522 641 -5519
rect 513 -5526 522 -5522
rect 529 -5526 537 -5522
rect 513 -5529 517 -5526
rect 537 -5529 541 -5526
rect 545 -5526 557 -5522
rect 571 -5526 579 -5522
rect 545 -5529 549 -5526
rect 579 -5529 583 -5526
rect 587 -5526 599 -5522
rect 613 -5526 625 -5522
rect 587 -5529 591 -5526
rect 621 -5529 625 -5526
rect 629 -5526 641 -5522
rect 655 -5522 659 -5505
rect 679 -5508 683 -5461
rect 679 -5522 683 -5512
rect 655 -5526 667 -5522
rect 629 -5529 633 -5526
rect 663 -5529 667 -5526
rect 671 -5526 683 -5522
rect 671 -5529 675 -5526
rect 504 -5537 508 -5533
rect 521 -5537 525 -5533
rect 562 -5537 566 -5533
rect 604 -5537 608 -5533
rect 646 -5537 650 -5533
rect 687 -5537 691 -5533
rect 495 -5567 499 -5563
rect 512 -5567 516 -5563
rect 503 -5578 507 -5575
rect 503 -5582 518 -5578
rect 514 -5621 518 -5582
rect 514 -5636 518 -5625
rect 495 -5640 518 -5636
rect 521 -5612 525 -5575
rect 705 -5591 709 -5497
rect 495 -5643 499 -5640
rect 521 -5643 525 -5616
rect 512 -5651 516 -5647
rect 504 -5726 508 -5722
rect 530 -5726 534 -5722
rect 547 -5726 551 -5722
rect 587 -5726 591 -5722
rect 608 -5726 612 -5722
rect 625 -5726 629 -5722
rect 665 -5726 669 -5722
rect 689 -5726 693 -5722
rect 726 -5726 730 -5722
rect 495 -5751 499 -5734
rect 495 -5802 499 -5755
rect 513 -5744 517 -5734
rect 513 -5802 517 -5748
rect 521 -5773 525 -5734
rect 539 -5766 543 -5734
rect 521 -5802 525 -5777
rect 539 -5802 543 -5770
rect 565 -5758 569 -5734
rect 565 -5795 569 -5762
rect 599 -5795 603 -5734
rect 617 -5751 621 -5734
rect 547 -5802 551 -5799
rect 555 -5799 569 -5795
rect 555 -5802 559 -5799
rect 583 -5802 587 -5799
rect 591 -5799 610 -5795
rect 591 -5802 595 -5799
rect 617 -5802 621 -5755
rect 643 -5766 647 -5734
rect 643 -5795 647 -5770
rect 677 -5788 681 -5734
rect 677 -5792 694 -5788
rect 625 -5802 629 -5799
rect 634 -5799 647 -5795
rect 634 -5802 638 -5799
rect 661 -5802 665 -5799
rect 685 -5802 689 -5792
rect 701 -5795 705 -5734
rect 709 -5788 713 -5734
rect 735 -5758 739 -5734
rect 709 -5792 728 -5788
rect 693 -5799 710 -5795
rect 693 -5802 697 -5799
rect 717 -5802 721 -5792
rect 735 -5802 739 -5762
rect 504 -5810 508 -5806
rect 530 -5810 534 -5806
rect 573 -5810 577 -5806
rect 608 -5810 612 -5806
rect 652 -5810 656 -5806
rect 669 -5810 673 -5806
rect 705 -5810 709 -5806
rect 726 -5810 730 -5806
rect 748 -5817 752 -5770
rect 810 -5773 814 -5616
rect 822 -5758 826 -5389
rect 839 -5501 843 -4872
rect 872 -4898 876 -4859
rect 872 -4913 876 -4902
rect 853 -4917 876 -4913
rect 879 -4889 883 -4852
rect 1062 -4868 1066 -4773
rect 853 -4920 857 -4917
rect 879 -4920 883 -4893
rect 870 -4928 874 -4924
rect 862 -5003 866 -4999
rect 888 -5003 892 -4999
rect 905 -5003 909 -4999
rect 945 -5003 949 -4999
rect 966 -5003 970 -4999
rect 983 -5003 987 -4999
rect 1023 -5003 1027 -4999
rect 1047 -5003 1051 -4999
rect 1084 -5003 1088 -4999
rect 853 -5028 857 -5011
rect 853 -5079 857 -5032
rect 871 -5021 875 -5011
rect 871 -5079 875 -5025
rect 879 -5050 883 -5011
rect 897 -5043 901 -5011
rect 879 -5079 883 -5054
rect 897 -5079 901 -5047
rect 923 -5035 927 -5011
rect 923 -5072 927 -5039
rect 957 -5072 961 -5011
rect 975 -5028 979 -5011
rect 905 -5079 909 -5076
rect 913 -5076 927 -5072
rect 913 -5079 917 -5076
rect 941 -5079 945 -5076
rect 949 -5076 968 -5072
rect 949 -5079 953 -5076
rect 975 -5079 979 -5032
rect 1001 -5043 1005 -5011
rect 1001 -5072 1005 -5047
rect 1035 -5065 1039 -5011
rect 1035 -5069 1052 -5065
rect 983 -5079 987 -5076
rect 992 -5076 1005 -5072
rect 992 -5079 996 -5076
rect 1019 -5079 1023 -5076
rect 1043 -5079 1047 -5069
rect 1059 -5072 1063 -5011
rect 1067 -5065 1071 -5011
rect 1093 -5033 1097 -5011
rect 1067 -5069 1086 -5065
rect 1051 -5076 1068 -5072
rect 1051 -5079 1055 -5076
rect 1075 -5079 1079 -5069
rect 1093 -5079 1097 -5037
rect 1167 -5035 1171 -4893
rect 862 -5087 866 -5083
rect 888 -5087 892 -5083
rect 931 -5087 935 -5083
rect 966 -5087 970 -5083
rect 1010 -5087 1014 -5083
rect 1027 -5087 1031 -5083
rect 1063 -5087 1067 -5083
rect 1084 -5087 1088 -5083
rect 1101 -5101 1105 -5047
rect 1184 -5050 1188 -4653
rect 1197 -4777 1201 -4133
rect 1230 -4159 1234 -4120
rect 1230 -4174 1234 -4163
rect 1211 -4178 1234 -4174
rect 1237 -4150 1241 -4113
rect 1418 -4129 1422 -4034
rect 1211 -4181 1215 -4178
rect 1237 -4181 1241 -4154
rect 1228 -4189 1232 -4185
rect 1220 -4264 1224 -4260
rect 1246 -4264 1250 -4260
rect 1263 -4264 1267 -4260
rect 1303 -4264 1307 -4260
rect 1324 -4264 1328 -4260
rect 1341 -4264 1345 -4260
rect 1381 -4264 1385 -4260
rect 1405 -4264 1409 -4260
rect 1442 -4264 1446 -4260
rect 1211 -4289 1215 -4272
rect 1211 -4340 1215 -4293
rect 1229 -4282 1233 -4272
rect 1229 -4340 1233 -4286
rect 1237 -4311 1241 -4272
rect 1255 -4304 1259 -4272
rect 1237 -4340 1241 -4315
rect 1255 -4340 1259 -4308
rect 1281 -4296 1285 -4272
rect 1281 -4333 1285 -4300
rect 1315 -4333 1319 -4272
rect 1333 -4289 1337 -4272
rect 1263 -4340 1267 -4337
rect 1271 -4337 1285 -4333
rect 1271 -4340 1275 -4337
rect 1299 -4340 1303 -4337
rect 1307 -4337 1326 -4333
rect 1307 -4340 1311 -4337
rect 1333 -4340 1337 -4293
rect 1359 -4304 1363 -4272
rect 1359 -4333 1363 -4308
rect 1393 -4326 1397 -4272
rect 1393 -4330 1410 -4326
rect 1341 -4340 1345 -4337
rect 1350 -4337 1363 -4333
rect 1350 -4340 1354 -4337
rect 1377 -4340 1381 -4337
rect 1401 -4340 1405 -4330
rect 1417 -4333 1421 -4272
rect 1425 -4326 1429 -4272
rect 1425 -4330 1444 -4326
rect 1409 -4337 1426 -4333
rect 1409 -4340 1413 -4337
rect 1433 -4340 1437 -4330
rect 1451 -4340 1455 -4272
rect 1220 -4348 1224 -4344
rect 1246 -4348 1250 -4344
rect 1289 -4348 1293 -4344
rect 1324 -4348 1328 -4344
rect 1368 -4348 1372 -4344
rect 1385 -4348 1389 -4344
rect 1421 -4348 1425 -4344
rect 1442 -4348 1446 -4344
rect 1451 -4362 1455 -4344
rect 1464 -4355 1468 -4308
rect 1220 -4558 1224 -4554
rect 1237 -4558 1241 -4554
rect 1257 -4558 1261 -4554
rect 1278 -4558 1282 -4554
rect 1299 -4558 1303 -4554
rect 1320 -4558 1324 -4554
rect 1341 -4558 1345 -4554
rect 1362 -4558 1366 -4554
rect 1383 -4558 1387 -4554
rect 1403 -4558 1407 -4554
rect 1211 -4613 1215 -4566
rect 1211 -4634 1215 -4617
rect 1229 -4627 1233 -4566
rect 1245 -4627 1249 -4566
rect 1269 -4606 1273 -4566
rect 1269 -4627 1273 -4610
rect 1287 -4627 1291 -4566
rect 1311 -4613 1315 -4566
rect 1311 -4627 1315 -4617
rect 1329 -4606 1333 -4566
rect 1329 -4627 1333 -4610
rect 1353 -4620 1357 -4566
rect 1371 -4598 1375 -4566
rect 1371 -4606 1375 -4602
rect 1353 -4627 1357 -4624
rect 1229 -4631 1238 -4627
rect 1245 -4631 1253 -4627
rect 1229 -4634 1233 -4631
rect 1253 -4634 1257 -4631
rect 1261 -4631 1273 -4627
rect 1287 -4631 1295 -4627
rect 1261 -4634 1265 -4631
rect 1295 -4634 1299 -4631
rect 1303 -4631 1315 -4627
rect 1329 -4631 1341 -4627
rect 1303 -4634 1307 -4631
rect 1337 -4634 1341 -4631
rect 1345 -4631 1357 -4627
rect 1371 -4627 1375 -4610
rect 1395 -4613 1399 -4566
rect 1395 -4627 1399 -4617
rect 1371 -4631 1383 -4627
rect 1345 -4634 1349 -4631
rect 1379 -4634 1383 -4631
rect 1387 -4631 1399 -4627
rect 1387 -4634 1391 -4631
rect 1220 -4642 1224 -4638
rect 1237 -4642 1241 -4638
rect 1278 -4642 1282 -4638
rect 1320 -4642 1324 -4638
rect 1362 -4642 1366 -4638
rect 1403 -4642 1407 -4638
rect 1419 -4649 1423 -4602
rect 1220 -4729 1224 -4725
rect 1237 -4729 1241 -4725
rect 1257 -4729 1261 -4725
rect 1278 -4729 1282 -4725
rect 1299 -4729 1303 -4725
rect 1320 -4729 1324 -4725
rect 1341 -4729 1345 -4725
rect 1362 -4729 1366 -4725
rect 1383 -4729 1387 -4725
rect 1403 -4729 1407 -4725
rect 1211 -4784 1215 -4737
rect 1211 -4805 1215 -4788
rect 1229 -4798 1233 -4737
rect 1245 -4798 1249 -4737
rect 1269 -4777 1273 -4737
rect 1269 -4798 1273 -4781
rect 1287 -4798 1291 -4737
rect 1311 -4784 1315 -4737
rect 1311 -4798 1315 -4788
rect 1329 -4777 1333 -4737
rect 1329 -4798 1333 -4781
rect 1353 -4791 1357 -4737
rect 1371 -4769 1375 -4737
rect 1371 -4777 1375 -4773
rect 1353 -4798 1357 -4795
rect 1229 -4802 1238 -4798
rect 1245 -4802 1253 -4798
rect 1229 -4805 1233 -4802
rect 1253 -4805 1257 -4802
rect 1261 -4802 1273 -4798
rect 1287 -4802 1295 -4798
rect 1261 -4805 1265 -4802
rect 1295 -4805 1299 -4802
rect 1303 -4802 1315 -4798
rect 1329 -4802 1341 -4798
rect 1303 -4805 1307 -4802
rect 1337 -4805 1341 -4802
rect 1345 -4802 1357 -4798
rect 1371 -4798 1375 -4781
rect 1395 -4784 1399 -4737
rect 1395 -4798 1399 -4788
rect 1371 -4802 1383 -4798
rect 1345 -4805 1349 -4802
rect 1379 -4805 1383 -4802
rect 1387 -4802 1399 -4798
rect 1387 -4805 1391 -4802
rect 1220 -4813 1224 -4809
rect 1237 -4813 1241 -4809
rect 1278 -4813 1282 -4809
rect 1320 -4813 1324 -4809
rect 1362 -4813 1366 -4809
rect 1403 -4813 1407 -4809
rect 1211 -4844 1215 -4840
rect 1228 -4844 1232 -4840
rect 1219 -4855 1223 -4852
rect 1219 -4859 1234 -4855
rect 1197 -4872 1212 -4868
rect 862 -5293 866 -5289
rect 879 -5293 883 -5289
rect 899 -5293 903 -5289
rect 920 -5293 924 -5289
rect 941 -5293 945 -5289
rect 962 -5293 966 -5289
rect 983 -5293 987 -5289
rect 1004 -5293 1008 -5289
rect 1025 -5293 1029 -5289
rect 1045 -5293 1049 -5289
rect 853 -5348 857 -5301
rect 853 -5369 857 -5352
rect 871 -5362 875 -5301
rect 887 -5362 891 -5301
rect 911 -5341 915 -5301
rect 911 -5362 915 -5345
rect 929 -5362 933 -5301
rect 953 -5348 957 -5301
rect 953 -5362 957 -5352
rect 971 -5341 975 -5301
rect 971 -5362 975 -5345
rect 995 -5355 999 -5301
rect 1013 -5333 1017 -5301
rect 1013 -5341 1017 -5337
rect 995 -5362 999 -5359
rect 871 -5366 880 -5362
rect 887 -5366 895 -5362
rect 871 -5369 875 -5366
rect 895 -5369 899 -5366
rect 903 -5366 915 -5362
rect 929 -5366 937 -5362
rect 903 -5369 907 -5366
rect 937 -5369 941 -5366
rect 945 -5366 957 -5362
rect 971 -5366 983 -5362
rect 945 -5369 949 -5366
rect 979 -5369 983 -5366
rect 987 -5366 999 -5362
rect 1013 -5362 1017 -5345
rect 1037 -5348 1041 -5301
rect 1037 -5362 1041 -5352
rect 1013 -5366 1025 -5362
rect 987 -5369 991 -5366
rect 1021 -5369 1025 -5366
rect 1029 -5366 1041 -5362
rect 1029 -5369 1033 -5366
rect 862 -5377 866 -5373
rect 879 -5377 883 -5373
rect 920 -5377 924 -5373
rect 962 -5377 966 -5373
rect 1004 -5377 1008 -5373
rect 1045 -5377 1049 -5373
rect 1061 -5385 1065 -5337
rect 1177 -5341 1181 -5105
rect 862 -5453 866 -5449
rect 879 -5453 883 -5449
rect 899 -5453 903 -5449
rect 920 -5453 924 -5449
rect 941 -5453 945 -5449
rect 962 -5453 966 -5449
rect 983 -5453 987 -5449
rect 1004 -5453 1008 -5449
rect 1025 -5453 1029 -5449
rect 1045 -5453 1049 -5449
rect 853 -5508 857 -5461
rect 853 -5529 857 -5512
rect 871 -5522 875 -5461
rect 887 -5522 891 -5461
rect 911 -5501 915 -5461
rect 911 -5522 915 -5505
rect 929 -5522 933 -5461
rect 953 -5508 957 -5461
rect 953 -5522 957 -5512
rect 971 -5501 975 -5461
rect 971 -5522 975 -5505
rect 995 -5515 999 -5461
rect 1013 -5493 1017 -5461
rect 1013 -5501 1017 -5497
rect 995 -5522 999 -5519
rect 871 -5526 880 -5522
rect 887 -5526 895 -5522
rect 871 -5529 875 -5526
rect 895 -5529 899 -5526
rect 903 -5526 915 -5522
rect 929 -5526 937 -5522
rect 903 -5529 907 -5526
rect 937 -5529 941 -5526
rect 945 -5526 957 -5522
rect 971 -5526 983 -5522
rect 945 -5529 949 -5526
rect 979 -5529 983 -5526
rect 987 -5526 999 -5522
rect 1013 -5522 1017 -5505
rect 1037 -5508 1041 -5461
rect 1037 -5522 1041 -5512
rect 1013 -5526 1025 -5522
rect 987 -5529 991 -5526
rect 1021 -5529 1025 -5526
rect 1029 -5526 1041 -5522
rect 1029 -5529 1033 -5526
rect 862 -5537 866 -5533
rect 879 -5537 883 -5533
rect 920 -5537 924 -5533
rect 962 -5537 966 -5533
rect 1004 -5537 1008 -5533
rect 1045 -5537 1049 -5533
rect 853 -5567 857 -5563
rect 870 -5567 874 -5563
rect 861 -5578 865 -5575
rect 861 -5582 876 -5578
rect 872 -5621 876 -5582
rect 872 -5636 876 -5625
rect 853 -5640 876 -5636
rect 879 -5612 883 -5575
rect 1062 -5591 1066 -5497
rect 853 -5643 857 -5640
rect 879 -5643 883 -5616
rect 870 -5651 874 -5647
rect 862 -5726 866 -5722
rect 888 -5726 892 -5722
rect 905 -5726 909 -5722
rect 945 -5726 949 -5722
rect 966 -5726 970 -5722
rect 983 -5726 987 -5722
rect 1023 -5726 1027 -5722
rect 1047 -5726 1051 -5722
rect 1084 -5726 1088 -5722
rect 853 -5751 857 -5734
rect 853 -5802 857 -5755
rect 871 -5744 875 -5734
rect 871 -5802 875 -5748
rect 879 -5773 883 -5734
rect 897 -5766 901 -5734
rect 879 -5802 883 -5777
rect 897 -5802 901 -5770
rect 923 -5758 927 -5734
rect 923 -5795 927 -5762
rect 957 -5795 961 -5734
rect 975 -5751 979 -5734
rect 905 -5802 909 -5799
rect 913 -5799 927 -5795
rect 913 -5802 917 -5799
rect 941 -5802 945 -5799
rect 949 -5799 968 -5795
rect 949 -5802 953 -5799
rect 975 -5802 979 -5755
rect 1001 -5766 1005 -5734
rect 1001 -5795 1005 -5770
rect 1035 -5788 1039 -5734
rect 1035 -5792 1052 -5788
rect 983 -5802 987 -5799
rect 992 -5799 1005 -5795
rect 992 -5802 996 -5799
rect 1019 -5802 1023 -5799
rect 1043 -5802 1047 -5792
rect 1059 -5795 1063 -5734
rect 1067 -5788 1071 -5734
rect 1093 -5756 1097 -5734
rect 1067 -5792 1086 -5788
rect 1051 -5799 1068 -5795
rect 1051 -5802 1055 -5799
rect 1075 -5802 1079 -5792
rect 1093 -5802 1097 -5760
rect 1167 -5758 1171 -5616
rect 862 -5810 866 -5806
rect 888 -5810 892 -5806
rect 931 -5810 935 -5806
rect 966 -5810 970 -5806
rect 1010 -5810 1014 -5806
rect 1027 -5810 1031 -5806
rect 1063 -5810 1067 -5806
rect 1084 -5810 1088 -5806
rect 1106 -5817 1110 -5770
rect 1177 -5773 1181 -5388
rect 1197 -5501 1201 -4872
rect 1230 -4898 1234 -4859
rect 1230 -4913 1234 -4902
rect 1211 -4917 1234 -4913
rect 1237 -4889 1241 -4852
rect 1420 -4868 1424 -4773
rect 1211 -4920 1215 -4917
rect 1237 -4920 1241 -4893
rect 1228 -4928 1232 -4924
rect 1220 -5003 1224 -4999
rect 1246 -5003 1250 -4999
rect 1263 -5003 1267 -4999
rect 1303 -5003 1307 -4999
rect 1324 -5003 1328 -4999
rect 1341 -5003 1345 -4999
rect 1381 -5003 1385 -4999
rect 1405 -5003 1409 -4999
rect 1442 -5003 1446 -4999
rect 1211 -5028 1215 -5011
rect 1211 -5079 1215 -5032
rect 1229 -5021 1233 -5011
rect 1229 -5079 1233 -5025
rect 1237 -5050 1241 -5011
rect 1255 -5043 1259 -5011
rect 1237 -5079 1241 -5054
rect 1255 -5079 1259 -5047
rect 1281 -5035 1285 -5011
rect 1281 -5072 1285 -5039
rect 1315 -5072 1319 -5011
rect 1333 -5028 1337 -5011
rect 1263 -5079 1267 -5076
rect 1271 -5076 1285 -5072
rect 1271 -5079 1275 -5076
rect 1299 -5079 1303 -5076
rect 1307 -5076 1326 -5072
rect 1307 -5079 1311 -5076
rect 1333 -5079 1337 -5032
rect 1359 -5043 1363 -5011
rect 1359 -5072 1363 -5047
rect 1393 -5065 1397 -5011
rect 1393 -5069 1410 -5065
rect 1341 -5079 1345 -5076
rect 1350 -5076 1363 -5072
rect 1350 -5079 1354 -5076
rect 1377 -5079 1381 -5076
rect 1401 -5079 1405 -5069
rect 1417 -5072 1421 -5011
rect 1425 -5065 1429 -5011
rect 1425 -5069 1444 -5065
rect 1409 -5076 1426 -5072
rect 1409 -5079 1413 -5076
rect 1433 -5079 1437 -5069
rect 1451 -5079 1455 -5011
rect 1220 -5087 1224 -5083
rect 1246 -5087 1250 -5083
rect 1289 -5087 1293 -5083
rect 1324 -5087 1328 -5083
rect 1368 -5087 1372 -5083
rect 1385 -5087 1389 -5083
rect 1421 -5087 1425 -5083
rect 1442 -5087 1446 -5083
rect 1451 -5101 1455 -5083
rect 1464 -5094 1468 -5047
rect 1220 -5293 1224 -5289
rect 1237 -5293 1241 -5289
rect 1257 -5293 1261 -5289
rect 1278 -5293 1282 -5289
rect 1299 -5293 1303 -5289
rect 1320 -5293 1324 -5289
rect 1341 -5293 1345 -5289
rect 1362 -5293 1366 -5289
rect 1383 -5293 1387 -5289
rect 1403 -5293 1407 -5289
rect 1211 -5348 1215 -5301
rect 1211 -5369 1215 -5352
rect 1229 -5362 1233 -5301
rect 1245 -5362 1249 -5301
rect 1269 -5341 1273 -5301
rect 1269 -5362 1273 -5345
rect 1287 -5362 1291 -5301
rect 1311 -5348 1315 -5301
rect 1311 -5362 1315 -5352
rect 1329 -5341 1333 -5301
rect 1329 -5362 1333 -5345
rect 1353 -5355 1357 -5301
rect 1371 -5333 1375 -5301
rect 1371 -5341 1375 -5337
rect 1353 -5362 1357 -5359
rect 1229 -5366 1238 -5362
rect 1245 -5366 1253 -5362
rect 1229 -5369 1233 -5366
rect 1253 -5369 1257 -5366
rect 1261 -5366 1273 -5362
rect 1287 -5366 1295 -5362
rect 1261 -5369 1265 -5366
rect 1295 -5369 1299 -5366
rect 1303 -5366 1315 -5362
rect 1329 -5366 1341 -5362
rect 1303 -5369 1307 -5366
rect 1337 -5369 1341 -5366
rect 1345 -5366 1357 -5362
rect 1371 -5362 1375 -5345
rect 1395 -5348 1399 -5301
rect 1395 -5362 1399 -5352
rect 1371 -5366 1383 -5362
rect 1345 -5369 1349 -5366
rect 1379 -5369 1383 -5366
rect 1387 -5366 1399 -5362
rect 1387 -5369 1391 -5366
rect 1220 -5377 1224 -5373
rect 1237 -5377 1241 -5373
rect 1278 -5377 1282 -5373
rect 1320 -5377 1324 -5373
rect 1362 -5377 1366 -5373
rect 1403 -5377 1407 -5373
rect 1423 -5384 1427 -5337
rect 1220 -5453 1224 -5449
rect 1237 -5453 1241 -5449
rect 1257 -5453 1261 -5449
rect 1278 -5453 1282 -5449
rect 1299 -5453 1303 -5449
rect 1320 -5453 1324 -5449
rect 1341 -5453 1345 -5449
rect 1362 -5453 1366 -5449
rect 1383 -5453 1387 -5449
rect 1403 -5453 1407 -5449
rect 1211 -5508 1215 -5461
rect 1211 -5529 1215 -5512
rect 1229 -5522 1233 -5461
rect 1245 -5522 1249 -5461
rect 1269 -5501 1273 -5461
rect 1269 -5522 1273 -5505
rect 1287 -5522 1291 -5461
rect 1311 -5508 1315 -5461
rect 1311 -5522 1315 -5512
rect 1329 -5501 1333 -5461
rect 1329 -5522 1333 -5505
rect 1353 -5515 1357 -5461
rect 1371 -5493 1375 -5461
rect 1371 -5501 1375 -5497
rect 1353 -5522 1357 -5519
rect 1229 -5526 1238 -5522
rect 1245 -5526 1253 -5522
rect 1229 -5529 1233 -5526
rect 1253 -5529 1257 -5526
rect 1261 -5526 1273 -5522
rect 1287 -5526 1295 -5522
rect 1261 -5529 1265 -5526
rect 1295 -5529 1299 -5526
rect 1303 -5526 1315 -5522
rect 1329 -5526 1341 -5522
rect 1303 -5529 1307 -5526
rect 1337 -5529 1341 -5526
rect 1345 -5526 1357 -5522
rect 1371 -5522 1375 -5505
rect 1395 -5508 1399 -5461
rect 1395 -5522 1399 -5512
rect 1371 -5526 1383 -5522
rect 1345 -5529 1349 -5526
rect 1379 -5529 1383 -5526
rect 1387 -5526 1399 -5522
rect 1387 -5529 1391 -5526
rect 1220 -5537 1224 -5533
rect 1237 -5537 1241 -5533
rect 1278 -5537 1282 -5533
rect 1320 -5537 1324 -5533
rect 1362 -5537 1366 -5533
rect 1403 -5537 1407 -5533
rect 1211 -5567 1215 -5563
rect 1228 -5567 1232 -5563
rect 1219 -5578 1223 -5575
rect 1219 -5582 1234 -5578
rect 1230 -5621 1234 -5582
rect 1230 -5636 1234 -5625
rect 1211 -5640 1234 -5636
rect 1237 -5612 1241 -5575
rect 1423 -5591 1427 -5497
rect 1211 -5643 1215 -5640
rect 1237 -5643 1241 -5616
rect 1228 -5651 1232 -5647
rect 1220 -5726 1224 -5722
rect 1246 -5726 1250 -5722
rect 1263 -5726 1267 -5722
rect 1303 -5726 1307 -5722
rect 1324 -5726 1328 -5722
rect 1341 -5726 1345 -5722
rect 1381 -5726 1385 -5722
rect 1405 -5726 1409 -5722
rect 1442 -5726 1446 -5722
rect 1211 -5751 1215 -5734
rect 1211 -5802 1215 -5755
rect 1229 -5744 1233 -5734
rect 1229 -5802 1233 -5748
rect 1237 -5773 1241 -5734
rect 1255 -5766 1259 -5734
rect 1237 -5802 1241 -5777
rect 1255 -5802 1259 -5770
rect 1281 -5758 1285 -5734
rect 1281 -5795 1285 -5762
rect 1315 -5795 1319 -5734
rect 1333 -5751 1337 -5734
rect 1263 -5802 1267 -5799
rect 1271 -5799 1285 -5795
rect 1271 -5802 1275 -5799
rect 1299 -5802 1303 -5799
rect 1307 -5799 1326 -5795
rect 1307 -5802 1311 -5799
rect 1333 -5802 1337 -5755
rect 1359 -5766 1363 -5734
rect 1359 -5795 1363 -5770
rect 1393 -5788 1397 -5734
rect 1393 -5792 1410 -5788
rect 1341 -5802 1345 -5799
rect 1350 -5799 1363 -5795
rect 1350 -5802 1354 -5799
rect 1377 -5802 1381 -5799
rect 1401 -5802 1405 -5792
rect 1417 -5795 1421 -5734
rect 1425 -5788 1429 -5734
rect 1425 -5792 1444 -5788
rect 1409 -5799 1426 -5795
rect 1409 -5802 1413 -5799
rect 1433 -5802 1437 -5792
rect 1451 -5802 1455 -5734
rect 1220 -5810 1224 -5806
rect 1246 -5810 1250 -5806
rect 1289 -5810 1293 -5806
rect 1324 -5810 1328 -5806
rect 1368 -5810 1372 -5806
rect 1385 -5810 1389 -5806
rect 1421 -5810 1425 -5806
rect 1442 -5810 1446 -5806
rect -1246 -5897 -1242 -5824
rect -1225 -5849 -1221 -5845
rect -1208 -5849 -1204 -5845
rect -1188 -5849 -1184 -5845
rect -1167 -5849 -1163 -5845
rect -1146 -5849 -1142 -5845
rect -1125 -5849 -1121 -5845
rect -1104 -5849 -1100 -5845
rect -1083 -5849 -1079 -5845
rect -1062 -5849 -1058 -5845
rect -1042 -5849 -1038 -5845
rect -1234 -5904 -1230 -5857
rect -1234 -5925 -1230 -5908
rect -1216 -5918 -1212 -5857
rect -1200 -5918 -1196 -5857
rect -1176 -5897 -1172 -5857
rect -1176 -5918 -1172 -5901
rect -1158 -5918 -1154 -5857
rect -1134 -5904 -1130 -5857
rect -1134 -5918 -1130 -5908
rect -1116 -5897 -1112 -5857
rect -1116 -5918 -1112 -5901
rect -1092 -5911 -1088 -5857
rect -1074 -5889 -1070 -5857
rect -1074 -5897 -1070 -5893
rect -1092 -5918 -1088 -5915
rect -1216 -5922 -1207 -5918
rect -1200 -5922 -1192 -5918
rect -1216 -5925 -1212 -5922
rect -1192 -5925 -1188 -5922
rect -1184 -5922 -1172 -5918
rect -1158 -5922 -1150 -5918
rect -1184 -5925 -1180 -5922
rect -1150 -5925 -1146 -5922
rect -1142 -5922 -1130 -5918
rect -1116 -5922 -1104 -5918
rect -1142 -5925 -1138 -5922
rect -1108 -5925 -1104 -5922
rect -1100 -5922 -1088 -5918
rect -1074 -5918 -1070 -5901
rect -1050 -5904 -1046 -5857
rect -949 -5897 -945 -5821
rect -926 -5849 -922 -5845
rect -909 -5849 -905 -5845
rect -889 -5849 -885 -5845
rect -868 -5849 -864 -5845
rect -847 -5849 -843 -5845
rect -826 -5849 -822 -5845
rect -805 -5849 -801 -5845
rect -784 -5849 -780 -5845
rect -763 -5849 -759 -5845
rect -743 -5849 -739 -5845
rect -1050 -5918 -1046 -5908
rect -1074 -5922 -1062 -5918
rect -1100 -5925 -1096 -5922
rect -1066 -5925 -1062 -5922
rect -1058 -5922 -1046 -5918
rect -935 -5904 -931 -5857
rect -1058 -5925 -1054 -5922
rect -935 -5925 -931 -5908
rect -917 -5918 -913 -5857
rect -901 -5918 -897 -5857
rect -877 -5897 -873 -5857
rect -877 -5918 -873 -5901
rect -859 -5918 -855 -5857
rect -835 -5904 -831 -5857
rect -835 -5918 -831 -5908
rect -817 -5897 -813 -5857
rect -817 -5918 -813 -5901
rect -793 -5911 -789 -5857
rect -775 -5889 -771 -5857
rect -775 -5897 -771 -5893
rect -793 -5918 -789 -5915
rect -917 -5922 -908 -5918
rect -901 -5922 -893 -5918
rect -917 -5925 -913 -5922
rect -893 -5925 -889 -5922
rect -885 -5922 -873 -5918
rect -859 -5922 -851 -5918
rect -885 -5925 -881 -5922
rect -851 -5925 -847 -5922
rect -843 -5922 -831 -5918
rect -817 -5922 -805 -5918
rect -843 -5925 -839 -5922
rect -809 -5925 -805 -5922
rect -801 -5922 -789 -5918
rect -775 -5918 -771 -5901
rect -751 -5904 -747 -5857
rect -586 -5897 -582 -5821
rect -568 -5849 -564 -5845
rect -551 -5849 -547 -5845
rect -531 -5849 -527 -5845
rect -510 -5849 -506 -5845
rect -489 -5849 -485 -5845
rect -468 -5849 -464 -5845
rect -447 -5849 -443 -5845
rect -426 -5849 -422 -5845
rect -405 -5849 -401 -5845
rect -385 -5849 -381 -5845
rect -751 -5918 -747 -5908
rect -775 -5922 -763 -5918
rect -801 -5925 -797 -5922
rect -767 -5925 -763 -5922
rect -759 -5922 -747 -5918
rect -577 -5904 -573 -5857
rect -759 -5925 -755 -5922
rect -577 -5925 -573 -5908
rect -559 -5918 -555 -5857
rect -543 -5918 -539 -5857
rect -519 -5897 -515 -5857
rect -519 -5918 -515 -5901
rect -501 -5918 -497 -5857
rect -477 -5904 -473 -5857
rect -477 -5918 -473 -5908
rect -459 -5897 -455 -5857
rect -459 -5918 -455 -5901
rect -435 -5911 -431 -5857
rect -417 -5889 -413 -5857
rect -417 -5897 -413 -5893
rect -435 -5918 -431 -5915
rect -559 -5922 -550 -5918
rect -543 -5922 -535 -5918
rect -559 -5925 -555 -5922
rect -535 -5925 -531 -5922
rect -527 -5922 -515 -5918
rect -501 -5922 -493 -5918
rect -527 -5925 -523 -5922
rect -493 -5925 -489 -5922
rect -485 -5922 -473 -5918
rect -459 -5922 -447 -5918
rect -485 -5925 -481 -5922
rect -451 -5925 -447 -5922
rect -443 -5922 -431 -5918
rect -417 -5918 -413 -5901
rect -393 -5904 -389 -5857
rect -233 -5897 -229 -5821
rect -210 -5849 -206 -5845
rect -193 -5849 -189 -5845
rect -173 -5849 -169 -5845
rect -152 -5849 -148 -5845
rect -131 -5849 -127 -5845
rect -110 -5849 -106 -5845
rect -89 -5849 -85 -5845
rect -68 -5849 -64 -5845
rect -47 -5849 -43 -5845
rect -27 -5849 -23 -5845
rect -393 -5918 -389 -5908
rect -417 -5922 -405 -5918
rect -443 -5925 -439 -5922
rect -409 -5925 -405 -5922
rect -401 -5922 -389 -5918
rect -219 -5904 -215 -5857
rect -401 -5925 -397 -5922
rect -219 -5925 -215 -5908
rect -201 -5918 -197 -5857
rect -185 -5918 -181 -5857
rect -161 -5897 -157 -5857
rect -161 -5918 -157 -5901
rect -143 -5918 -139 -5857
rect -119 -5904 -115 -5857
rect -119 -5918 -115 -5908
rect -101 -5897 -97 -5857
rect -101 -5918 -97 -5901
rect -77 -5911 -73 -5857
rect -59 -5889 -55 -5857
rect -59 -5897 -55 -5893
rect -77 -5918 -73 -5915
rect -201 -5922 -192 -5918
rect -185 -5922 -177 -5918
rect -201 -5925 -197 -5922
rect -177 -5925 -173 -5922
rect -169 -5922 -157 -5918
rect -143 -5922 -135 -5918
rect -169 -5925 -165 -5922
rect -135 -5925 -131 -5922
rect -127 -5922 -115 -5918
rect -101 -5922 -89 -5918
rect -127 -5925 -123 -5922
rect -93 -5925 -89 -5922
rect -85 -5922 -73 -5918
rect -59 -5918 -55 -5901
rect -35 -5904 -31 -5857
rect 129 -5897 133 -5822
rect 148 -5849 152 -5845
rect 165 -5849 169 -5845
rect 185 -5849 189 -5845
rect 206 -5849 210 -5845
rect 227 -5849 231 -5845
rect 248 -5849 252 -5845
rect 269 -5849 273 -5845
rect 290 -5849 294 -5845
rect 311 -5849 315 -5845
rect 331 -5849 335 -5845
rect -35 -5918 -31 -5908
rect -59 -5922 -47 -5918
rect -85 -5925 -81 -5922
rect -51 -5925 -47 -5922
rect -43 -5922 -31 -5918
rect 139 -5904 143 -5857
rect -43 -5925 -39 -5922
rect 139 -5925 143 -5908
rect 157 -5918 161 -5857
rect 173 -5918 177 -5857
rect 197 -5897 201 -5857
rect 197 -5918 201 -5901
rect 215 -5918 219 -5857
rect 239 -5904 243 -5857
rect 239 -5918 243 -5908
rect 257 -5897 261 -5857
rect 257 -5918 261 -5901
rect 281 -5911 285 -5857
rect 299 -5889 303 -5857
rect 299 -5897 303 -5893
rect 281 -5918 285 -5915
rect 157 -5922 166 -5918
rect 173 -5922 181 -5918
rect 157 -5925 161 -5922
rect 181 -5925 185 -5922
rect 189 -5922 201 -5918
rect 215 -5922 223 -5918
rect 189 -5925 193 -5922
rect 223 -5925 227 -5922
rect 231 -5922 243 -5918
rect 257 -5922 269 -5918
rect 231 -5925 235 -5922
rect 265 -5925 269 -5922
rect 273 -5922 285 -5918
rect 299 -5918 303 -5901
rect 323 -5904 327 -5857
rect 484 -5897 488 -5821
rect 504 -5849 508 -5845
rect 521 -5849 525 -5845
rect 541 -5849 545 -5845
rect 562 -5849 566 -5845
rect 583 -5849 587 -5845
rect 604 -5849 608 -5845
rect 625 -5849 629 -5845
rect 646 -5849 650 -5845
rect 667 -5849 671 -5845
rect 687 -5849 691 -5845
rect 323 -5918 327 -5908
rect 299 -5922 311 -5918
rect 273 -5925 277 -5922
rect 307 -5925 311 -5922
rect 315 -5922 327 -5918
rect 495 -5904 499 -5857
rect 315 -5925 319 -5922
rect 495 -5925 499 -5908
rect 513 -5918 517 -5857
rect 529 -5918 533 -5857
rect 553 -5897 557 -5857
rect 553 -5918 557 -5901
rect 571 -5918 575 -5857
rect 595 -5904 599 -5857
rect 595 -5918 599 -5908
rect 613 -5897 617 -5857
rect 613 -5918 617 -5901
rect 637 -5911 641 -5857
rect 655 -5889 659 -5857
rect 655 -5897 659 -5893
rect 637 -5918 641 -5915
rect 513 -5922 522 -5918
rect 529 -5922 537 -5918
rect 513 -5925 517 -5922
rect 537 -5925 541 -5922
rect 545 -5922 557 -5918
rect 571 -5922 579 -5918
rect 545 -5925 549 -5922
rect 579 -5925 583 -5922
rect 587 -5922 599 -5918
rect 613 -5922 625 -5918
rect 587 -5925 591 -5922
rect 621 -5925 625 -5922
rect 629 -5922 641 -5918
rect 655 -5918 659 -5901
rect 679 -5904 683 -5857
rect 842 -5897 846 -5821
rect 862 -5849 866 -5845
rect 879 -5849 883 -5845
rect 899 -5849 903 -5845
rect 920 -5849 924 -5845
rect 941 -5849 945 -5845
rect 962 -5849 966 -5845
rect 983 -5849 987 -5845
rect 1004 -5849 1008 -5845
rect 1025 -5849 1029 -5845
rect 1045 -5849 1049 -5845
rect 679 -5918 683 -5908
rect 655 -5922 667 -5918
rect 629 -5925 633 -5922
rect 663 -5925 667 -5922
rect 671 -5922 683 -5918
rect 853 -5904 857 -5857
rect 671 -5925 675 -5922
rect 853 -5925 857 -5908
rect 871 -5918 875 -5857
rect 887 -5918 891 -5857
rect 911 -5897 915 -5857
rect 911 -5918 915 -5901
rect 929 -5918 933 -5857
rect 953 -5904 957 -5857
rect 953 -5918 957 -5908
rect 971 -5897 975 -5857
rect 971 -5918 975 -5901
rect 995 -5911 999 -5857
rect 1013 -5889 1017 -5857
rect 1013 -5897 1017 -5893
rect 995 -5918 999 -5915
rect 871 -5922 880 -5918
rect 887 -5922 895 -5918
rect 871 -5925 875 -5922
rect 895 -5925 899 -5922
rect 903 -5922 915 -5918
rect 929 -5922 937 -5918
rect 903 -5925 907 -5922
rect 937 -5925 941 -5922
rect 945 -5922 957 -5918
rect 971 -5922 983 -5918
rect 945 -5925 949 -5922
rect 979 -5925 983 -5922
rect 987 -5922 999 -5918
rect 1013 -5918 1017 -5901
rect 1037 -5904 1041 -5857
rect 1199 -5897 1203 -5821
rect 1220 -5849 1224 -5845
rect 1237 -5849 1241 -5845
rect 1257 -5849 1261 -5845
rect 1278 -5849 1282 -5845
rect 1299 -5849 1303 -5845
rect 1320 -5849 1324 -5845
rect 1341 -5849 1345 -5845
rect 1362 -5849 1366 -5845
rect 1383 -5849 1387 -5845
rect 1403 -5849 1407 -5845
rect 1037 -5918 1041 -5908
rect 1013 -5922 1025 -5918
rect 987 -5925 991 -5922
rect 1021 -5925 1025 -5922
rect 1029 -5922 1041 -5918
rect 1211 -5904 1215 -5857
rect 1029 -5925 1033 -5922
rect 1211 -5925 1215 -5908
rect 1229 -5918 1233 -5857
rect 1245 -5918 1249 -5857
rect 1269 -5897 1273 -5857
rect 1269 -5918 1273 -5901
rect 1287 -5918 1291 -5857
rect 1311 -5904 1315 -5857
rect 1311 -5918 1315 -5908
rect 1329 -5897 1333 -5857
rect 1329 -5918 1333 -5901
rect 1353 -5911 1357 -5857
rect 1371 -5889 1375 -5857
rect 1371 -5897 1375 -5893
rect 1353 -5918 1357 -5915
rect 1229 -5922 1238 -5918
rect 1245 -5922 1253 -5918
rect 1229 -5925 1233 -5922
rect 1253 -5925 1257 -5922
rect 1261 -5922 1273 -5918
rect 1287 -5922 1295 -5918
rect 1261 -5925 1265 -5922
rect 1295 -5925 1299 -5922
rect 1303 -5922 1315 -5918
rect 1329 -5922 1341 -5918
rect 1303 -5925 1307 -5922
rect 1337 -5925 1341 -5922
rect 1345 -5922 1357 -5918
rect 1371 -5918 1375 -5901
rect 1395 -5904 1399 -5857
rect 1451 -5897 1455 -5806
rect 1466 -5817 1470 -5770
rect 1564 -5849 1568 -5845
rect 1581 -5849 1585 -5845
rect 1601 -5849 1605 -5845
rect 1622 -5849 1626 -5845
rect 1643 -5849 1647 -5845
rect 1664 -5849 1668 -5845
rect 1685 -5849 1689 -5845
rect 1706 -5849 1710 -5845
rect 1727 -5849 1731 -5845
rect 1747 -5849 1751 -5845
rect 1395 -5918 1399 -5908
rect 1371 -5922 1383 -5918
rect 1345 -5925 1349 -5922
rect 1379 -5925 1383 -5922
rect 1387 -5922 1399 -5918
rect 1555 -5904 1559 -5857
rect 1387 -5925 1391 -5922
rect 1555 -5925 1559 -5908
rect 1573 -5918 1577 -5857
rect 1589 -5918 1593 -5857
rect 1613 -5897 1617 -5857
rect 1613 -5918 1617 -5901
rect 1631 -5918 1635 -5857
rect 1655 -5904 1659 -5857
rect 1655 -5918 1659 -5908
rect 1673 -5897 1677 -5857
rect 1673 -5918 1677 -5901
rect 1697 -5911 1701 -5857
rect 1715 -5889 1719 -5857
rect 1715 -5897 1719 -5893
rect 1697 -5918 1701 -5915
rect 1573 -5922 1582 -5918
rect 1589 -5922 1597 -5918
rect 1573 -5925 1577 -5922
rect 1597 -5925 1601 -5922
rect 1605 -5922 1617 -5918
rect 1631 -5922 1639 -5918
rect 1605 -5925 1609 -5922
rect 1639 -5925 1643 -5922
rect 1647 -5922 1659 -5918
rect 1673 -5922 1685 -5918
rect 1647 -5925 1651 -5922
rect 1681 -5925 1685 -5922
rect 1689 -5922 1701 -5918
rect 1715 -5918 1719 -5901
rect 1739 -5904 1743 -5857
rect 1739 -5918 1743 -5908
rect 1715 -5922 1727 -5918
rect 1689 -5925 1693 -5922
rect 1723 -5925 1727 -5922
rect 1731 -5922 1743 -5918
rect 1731 -5925 1735 -5922
rect -1225 -5933 -1221 -5929
rect -1208 -5933 -1204 -5929
rect -1167 -5933 -1163 -5929
rect -1125 -5933 -1121 -5929
rect -1083 -5933 -1079 -5929
rect -1042 -5933 -1038 -5929
rect -926 -5933 -922 -5929
rect -909 -5933 -905 -5929
rect -868 -5933 -864 -5929
rect -826 -5933 -822 -5929
rect -784 -5933 -780 -5929
rect -743 -5933 -739 -5929
rect -568 -5933 -564 -5929
rect -551 -5933 -547 -5929
rect -510 -5933 -506 -5929
rect -468 -5933 -464 -5929
rect -426 -5933 -422 -5929
rect -385 -5933 -381 -5929
rect -210 -5933 -206 -5929
rect -193 -5933 -189 -5929
rect -152 -5933 -148 -5929
rect -110 -5933 -106 -5929
rect -68 -5933 -64 -5929
rect -27 -5933 -23 -5929
rect 148 -5933 152 -5929
rect 165 -5933 169 -5929
rect 206 -5933 210 -5929
rect 248 -5933 252 -5929
rect 290 -5933 294 -5929
rect 331 -5933 335 -5929
rect 504 -5933 508 -5929
rect 521 -5933 525 -5929
rect 562 -5933 566 -5929
rect 604 -5933 608 -5929
rect 646 -5933 650 -5929
rect 687 -5933 691 -5929
rect 862 -5933 866 -5929
rect 879 -5933 883 -5929
rect 920 -5933 924 -5929
rect 962 -5933 966 -5929
rect 1004 -5933 1008 -5929
rect 1045 -5933 1049 -5929
rect 1220 -5933 1224 -5929
rect 1237 -5933 1241 -5929
rect 1278 -5933 1282 -5929
rect 1320 -5933 1324 -5929
rect 1362 -5933 1366 -5929
rect 1403 -5933 1407 -5929
rect 1564 -5933 1568 -5929
rect 1581 -5933 1585 -5929
rect 1622 -5933 1626 -5929
rect 1664 -5933 1668 -5929
rect 1706 -5933 1710 -5929
rect 1747 -5933 1751 -5929
<< metal2 >>
rect -2054 -784 -1307 -780
rect -1303 -784 -1290 -780
rect -1286 -784 -936 -780
rect -932 -784 -919 -780
rect -915 -784 -577 -780
rect -573 -784 -560 -780
rect -556 -784 -219 -780
rect -215 -784 -202 -780
rect -198 -784 138 -780
rect 142 -784 155 -780
rect 159 -784 495 -780
rect 499 -784 512 -780
rect 516 -784 853 -780
rect 857 -784 870 -780
rect 874 -784 1211 -780
rect 1215 -784 1228 -780
rect 1232 -784 1589 -780
rect -2054 -1014 -2027 -784
rect -1411 -824 -1295 -820
rect -1291 -824 -924 -820
rect -920 -824 -565 -820
rect -561 -824 -207 -820
rect -203 -824 150 -820
rect 154 -824 507 -820
rect 511 -824 865 -820
rect 869 -824 1223 -820
rect 1227 -824 1589 -820
rect -960 -832 -551 -828
rect -240 -832 164 -828
rect 474 -832 879 -828
rect -1247 -840 -910 -836
rect -601 -840 -193 -836
rect 111 -840 521 -836
rect 825 -840 1237 -836
rect -1411 -876 -1290 -872
rect -1286 -876 -919 -872
rect -915 -876 -560 -872
rect -556 -876 -202 -872
rect -198 -876 155 -872
rect 159 -876 512 -872
rect 516 -876 870 -872
rect 874 -876 1228 -872
rect 1232 -876 1831 -872
rect -2054 -1018 -1221 -1014
rect -1217 -1018 -1204 -1014
rect -1200 -1018 -1184 -1014
rect -1180 -1018 -1163 -1014
rect -1159 -1018 -1142 -1014
rect -1138 -1018 -1121 -1014
rect -1117 -1018 -1100 -1014
rect -1096 -1018 -1079 -1014
rect -1075 -1018 -1058 -1014
rect -1054 -1018 -1038 -1014
rect -1034 -1018 -926 -1014
rect -922 -1018 -909 -1014
rect -905 -1018 -889 -1014
rect -885 -1018 -868 -1014
rect -864 -1018 -847 -1014
rect -843 -1018 -826 -1014
rect -822 -1018 -805 -1014
rect -801 -1018 -784 -1014
rect -780 -1018 -763 -1014
rect -759 -1018 -743 -1014
rect -739 -1018 -568 -1014
rect -564 -1018 -551 -1014
rect -547 -1018 -531 -1014
rect -527 -1018 -510 -1014
rect -506 -1018 -489 -1014
rect -485 -1018 -468 -1014
rect -464 -1018 -447 -1014
rect -443 -1018 -426 -1014
rect -422 -1018 -405 -1014
rect -401 -1018 -385 -1014
rect -381 -1018 -210 -1014
rect -206 -1018 -193 -1014
rect -189 -1018 -173 -1014
rect -169 -1018 -152 -1014
rect -148 -1018 -131 -1014
rect -127 -1018 -110 -1014
rect -106 -1018 -89 -1014
rect -85 -1018 -68 -1014
rect -64 -1018 -47 -1014
rect -43 -1018 -27 -1014
rect -23 -1018 148 -1014
rect 152 -1018 165 -1014
rect 169 -1018 185 -1014
rect 189 -1018 206 -1014
rect 210 -1018 227 -1014
rect 231 -1018 248 -1014
rect 252 -1018 269 -1014
rect 273 -1018 290 -1014
rect 294 -1018 311 -1014
rect 315 -1018 331 -1014
rect 335 -1018 504 -1014
rect 508 -1018 521 -1014
rect 525 -1018 541 -1014
rect 545 -1018 562 -1014
rect 566 -1018 583 -1014
rect 587 -1018 604 -1014
rect 608 -1018 625 -1014
rect 629 -1018 646 -1014
rect 650 -1018 667 -1014
rect 671 -1018 687 -1014
rect 691 -1018 862 -1014
rect 866 -1018 879 -1014
rect 883 -1018 899 -1014
rect 903 -1018 920 -1014
rect 924 -1018 941 -1014
rect 945 -1018 962 -1014
rect 966 -1018 983 -1014
rect 987 -1018 1004 -1014
rect 1008 -1018 1025 -1014
rect 1029 -1018 1045 -1014
rect 1049 -1018 1368 -1014
rect -2054 -1130 -2027 -1018
rect -1199 -1066 -1165 -1062
rect -1101 -1066 -1081 -1062
rect -1066 -1066 -931 -1062
rect -904 -1066 -870 -1062
rect -806 -1066 -786 -1062
rect -771 -1066 -573 -1062
rect -546 -1066 -512 -1062
rect -448 -1066 -428 -1062
rect -413 -1066 -215 -1062
rect -188 -1066 -154 -1062
rect -90 -1066 -70 -1062
rect -55 -1066 143 -1062
rect 170 -1066 204 -1062
rect 268 -1066 288 -1062
rect 303 -1066 499 -1062
rect 526 -1066 560 -1062
rect 624 -1066 644 -1062
rect 659 -1066 857 -1062
rect 884 -1066 918 -1062
rect 982 -1066 1002 -1062
rect 1017 -1066 1053 -1062
rect -935 -1070 -931 -1066
rect -577 -1070 -573 -1066
rect -219 -1070 -215 -1066
rect 139 -1070 143 -1066
rect 495 -1070 499 -1066
rect 853 -1070 857 -1066
rect -1277 -1074 -1223 -1070
rect -1219 -1074 -1189 -1070
rect -1168 -1074 -1137 -1070
rect -1108 -1074 -1077 -1070
rect -1066 -1074 -1039 -1070
rect -935 -1074 -928 -1070
rect -924 -1074 -894 -1070
rect -873 -1074 -842 -1070
rect -813 -1074 -782 -1070
rect -771 -1074 -744 -1070
rect -577 -1074 -570 -1070
rect -566 -1074 -536 -1070
rect -515 -1074 -484 -1070
rect -455 -1074 -424 -1070
rect -413 -1074 -386 -1070
rect -219 -1074 -212 -1070
rect -208 -1074 -178 -1070
rect -157 -1074 -126 -1070
rect -97 -1074 -66 -1070
rect -55 -1074 -28 -1070
rect 139 -1074 146 -1070
rect 150 -1074 180 -1070
rect 201 -1074 232 -1070
rect 261 -1074 292 -1070
rect 303 -1074 330 -1070
rect 495 -1074 502 -1070
rect 506 -1074 536 -1070
rect 557 -1074 588 -1070
rect 617 -1074 648 -1070
rect 659 -1074 686 -1070
rect 853 -1074 860 -1070
rect 864 -1074 894 -1070
rect 915 -1074 946 -1070
rect 975 -1074 1006 -1070
rect 1017 -1074 1044 -1070
rect -1226 -1081 -1179 -1077
rect -1143 -1081 -1130 -1077
rect -1126 -1081 -1095 -1077
rect -1059 -1081 -1046 -1077
rect -1042 -1081 -1030 -1077
rect -931 -1081 -884 -1077
rect -848 -1081 -835 -1077
rect -831 -1081 -800 -1077
rect -764 -1081 -751 -1077
rect -747 -1081 -735 -1077
rect -573 -1081 -526 -1077
rect -490 -1081 -477 -1077
rect -473 -1081 -442 -1077
rect -406 -1081 -393 -1077
rect -389 -1081 -377 -1077
rect -215 -1081 -168 -1077
rect -132 -1081 -119 -1077
rect -115 -1081 -84 -1077
rect -48 -1081 -35 -1077
rect -31 -1081 -19 -1077
rect 143 -1081 190 -1077
rect 226 -1081 239 -1077
rect 243 -1081 274 -1077
rect 310 -1081 323 -1077
rect 327 -1081 339 -1077
rect 499 -1081 546 -1077
rect 582 -1081 595 -1077
rect 599 -1081 630 -1077
rect 666 -1081 679 -1077
rect 683 -1081 695 -1077
rect 857 -1081 904 -1077
rect 940 -1081 953 -1077
rect 957 -1081 988 -1077
rect 1024 -1081 1037 -1077
rect 1041 -1081 1053 -1077
rect -1234 -1088 -1219 -1084
rect -1215 -1088 -1105 -1084
rect -1084 -1088 -1053 -1084
rect -939 -1088 -924 -1084
rect -920 -1088 -810 -1084
rect -789 -1088 -758 -1084
rect -581 -1088 -566 -1084
rect -562 -1088 -452 -1084
rect -431 -1088 -400 -1084
rect -223 -1088 -208 -1084
rect -204 -1088 -94 -1084
rect -73 -1088 -42 -1084
rect 135 -1088 150 -1084
rect 154 -1088 264 -1084
rect 285 -1088 316 -1084
rect 491 -1088 506 -1084
rect 510 -1088 620 -1084
rect 641 -1088 672 -1084
rect 849 -1088 864 -1084
rect 868 -1088 978 -1084
rect 999 -1088 1030 -1084
rect -1184 -1095 -1161 -1091
rect -1142 -1095 -1123 -1091
rect -889 -1095 -866 -1091
rect -847 -1095 -828 -1091
rect -531 -1095 -508 -1091
rect -489 -1095 -470 -1091
rect -173 -1095 -150 -1091
rect -131 -1095 -112 -1091
rect 185 -1095 208 -1091
rect 227 -1095 246 -1091
rect 541 -1095 564 -1091
rect 583 -1095 602 -1091
rect 899 -1095 922 -1091
rect 941 -1095 960 -1091
rect 1804 -1106 1831 -876
rect -1636 -1110 -1221 -1106
rect -1217 -1110 -1204 -1106
rect -1200 -1110 -1163 -1106
rect -1159 -1110 -1121 -1106
rect -1117 -1110 -1079 -1106
rect -1075 -1110 -1038 -1106
rect -1034 -1110 -926 -1106
rect -922 -1110 -909 -1106
rect -905 -1110 -868 -1106
rect -864 -1110 -826 -1106
rect -822 -1110 -784 -1106
rect -780 -1110 -743 -1106
rect -739 -1110 -568 -1106
rect -564 -1110 -551 -1106
rect -547 -1110 -510 -1106
rect -506 -1110 -468 -1106
rect -464 -1110 -426 -1106
rect -422 -1110 -385 -1106
rect -381 -1110 -210 -1106
rect -206 -1110 -193 -1106
rect -189 -1110 -152 -1106
rect -148 -1110 -110 -1106
rect -106 -1110 -68 -1106
rect -64 -1110 -27 -1106
rect -23 -1110 148 -1106
rect 152 -1110 165 -1106
rect 169 -1110 206 -1106
rect 210 -1110 248 -1106
rect 252 -1110 290 -1106
rect 294 -1110 331 -1106
rect 335 -1110 504 -1106
rect 508 -1110 521 -1106
rect 525 -1110 562 -1106
rect 566 -1110 604 -1106
rect 608 -1110 646 -1106
rect 650 -1110 687 -1106
rect 691 -1110 862 -1106
rect 866 -1110 879 -1106
rect 883 -1110 920 -1106
rect 924 -1110 962 -1106
rect 966 -1110 1004 -1106
rect 1008 -1110 1045 -1106
rect 1049 -1110 1831 -1106
rect -2054 -1134 -1309 -1130
rect -1305 -1134 -1292 -1130
rect -1288 -1134 -935 -1130
rect -931 -1134 -918 -1130
rect -914 -1134 -577 -1130
rect -573 -1134 -560 -1130
rect -556 -1134 -219 -1130
rect -215 -1134 -202 -1130
rect -198 -1134 139 -1130
rect 143 -1134 156 -1130
rect 160 -1134 495 -1130
rect 499 -1134 512 -1130
rect 516 -1134 853 -1130
rect 857 -1134 870 -1130
rect 874 -1134 1211 -1130
rect 1215 -1134 1228 -1130
rect 1232 -1134 1589 -1130
rect -2054 -1294 -2027 -1134
rect -1411 -1174 -1297 -1170
rect -1293 -1174 -923 -1170
rect -919 -1174 -565 -1170
rect -561 -1174 -207 -1170
rect -203 -1174 151 -1170
rect 155 -1174 507 -1170
rect 511 -1174 865 -1170
rect 869 -1174 1223 -1170
rect 1227 -1174 1589 -1170
rect -972 -1187 -909 -1183
rect -614 -1187 -551 -1183
rect -263 -1187 -193 -1183
rect 95 -1187 165 -1183
rect 451 -1187 521 -1183
rect 809 -1187 879 -1183
rect 1167 -1187 1237 -1183
rect 1804 -1222 1831 -1110
rect -1411 -1226 -1292 -1222
rect -1288 -1226 -918 -1222
rect -914 -1226 -560 -1222
rect -556 -1226 -202 -1222
rect -198 -1226 156 -1222
rect 160 -1226 512 -1222
rect 516 -1226 870 -1222
rect 874 -1226 1228 -1222
rect 1232 -1226 1831 -1222
rect -2054 -1298 -1221 -1294
rect -1217 -1298 -1204 -1294
rect -1200 -1298 -1164 -1294
rect -1160 -1298 -1143 -1294
rect -1139 -1298 -926 -1294
rect -922 -1298 -900 -1294
rect -896 -1298 -883 -1294
rect -879 -1298 -843 -1294
rect -839 -1298 -822 -1294
rect -818 -1298 -805 -1294
rect -801 -1298 -765 -1294
rect -761 -1298 -741 -1294
rect -737 -1298 -704 -1294
rect -700 -1298 -568 -1294
rect -564 -1298 -542 -1294
rect -538 -1298 -525 -1294
rect -521 -1298 -485 -1294
rect -481 -1298 -464 -1294
rect -460 -1298 -447 -1294
rect -443 -1298 -407 -1294
rect -403 -1298 -383 -1294
rect -379 -1298 -346 -1294
rect -342 -1298 -210 -1294
rect -206 -1298 -184 -1294
rect -180 -1298 -167 -1294
rect -163 -1298 -127 -1294
rect -123 -1298 -106 -1294
rect -102 -1298 -89 -1294
rect -85 -1298 -49 -1294
rect -45 -1298 -25 -1294
rect -21 -1298 12 -1294
rect 16 -1298 148 -1294
rect 152 -1298 174 -1294
rect 178 -1298 191 -1294
rect 195 -1298 231 -1294
rect 235 -1298 252 -1294
rect 256 -1298 269 -1294
rect 273 -1298 309 -1294
rect 313 -1298 333 -1294
rect 337 -1298 370 -1294
rect 374 -1298 504 -1294
rect 508 -1298 530 -1294
rect 534 -1298 547 -1294
rect 551 -1298 587 -1294
rect 591 -1298 608 -1294
rect 612 -1298 625 -1294
rect 629 -1298 665 -1294
rect 669 -1298 689 -1294
rect 693 -1298 726 -1294
rect 730 -1298 862 -1294
rect 866 -1298 888 -1294
rect 892 -1298 905 -1294
rect 909 -1298 945 -1294
rect 949 -1298 966 -1294
rect 970 -1298 983 -1294
rect 987 -1298 1023 -1294
rect 1027 -1298 1047 -1294
rect 1051 -1298 1084 -1294
rect 1088 -1298 1220 -1294
rect 1224 -1298 1237 -1294
rect 1241 -1298 1277 -1294
rect 1281 -1298 1298 -1294
rect 1302 -1298 1589 -1294
rect -2054 -1417 -2027 -1298
rect -210 -1302 -206 -1298
rect -184 -1302 -180 -1298
rect -167 -1302 -163 -1298
rect -127 -1302 -123 -1298
rect -106 -1302 -102 -1298
rect -89 -1302 -85 -1298
rect -49 -1302 -45 -1298
rect -25 -1302 -21 -1298
rect 12 -1302 16 -1298
rect 148 -1302 152 -1298
rect 174 -1302 178 -1298
rect 191 -1302 195 -1298
rect 231 -1302 235 -1298
rect 252 -1302 256 -1298
rect 269 -1302 273 -1298
rect 309 -1302 313 -1298
rect 333 -1302 337 -1298
rect 370 -1302 374 -1298
rect 504 -1302 508 -1298
rect 530 -1302 534 -1298
rect 547 -1302 551 -1298
rect 587 -1302 591 -1298
rect 608 -1302 612 -1298
rect 625 -1302 629 -1298
rect 665 -1302 669 -1298
rect 689 -1302 693 -1298
rect 726 -1302 730 -1298
rect 862 -1302 866 -1298
rect 888 -1302 892 -1298
rect 905 -1302 909 -1298
rect 945 -1302 949 -1298
rect 966 -1302 970 -1298
rect 983 -1302 987 -1298
rect 1023 -1302 1027 -1298
rect 1047 -1302 1051 -1298
rect 1084 -1302 1088 -1298
rect -920 -1317 -858 -1313
rect -854 -1317 -824 -1313
rect -776 -1317 -746 -1313
rect -562 -1317 -500 -1313
rect -496 -1317 -466 -1313
rect -418 -1317 -388 -1313
rect -204 -1317 -142 -1313
rect -138 -1317 -108 -1313
rect -60 -1317 -30 -1313
rect 154 -1317 216 -1313
rect 220 -1317 250 -1313
rect 298 -1317 328 -1313
rect 510 -1317 572 -1313
rect 576 -1317 606 -1313
rect 654 -1317 684 -1313
rect 868 -1317 930 -1313
rect 934 -1317 964 -1313
rect 1012 -1317 1042 -1313
rect -913 -1324 -882 -1320
rect -555 -1324 -524 -1320
rect -197 -1324 -166 -1320
rect 161 -1324 192 -1320
rect 517 -1324 548 -1320
rect 875 -1324 906 -1320
rect -931 -1331 -848 -1327
rect -809 -1331 -706 -1327
rect -573 -1331 -490 -1327
rect -451 -1331 -348 -1327
rect -215 -1331 -132 -1327
rect -93 -1331 10 -1327
rect 143 -1331 226 -1327
rect 265 -1331 368 -1327
rect 499 -1331 582 -1327
rect 621 -1331 724 -1327
rect 857 -1331 940 -1327
rect 979 -1331 1082 -1327
rect -960 -1338 -928 -1334
rect -894 -1338 -865 -1334
rect -861 -1338 -780 -1334
rect -691 -1338 -614 -1334
rect -601 -1338 -570 -1334
rect -536 -1338 -507 -1334
rect -503 -1338 -422 -1334
rect -333 -1338 -263 -1334
rect -240 -1338 -212 -1334
rect -178 -1338 -149 -1334
rect -145 -1338 -64 -1334
rect 25 -1338 95 -1334
rect 111 -1338 146 -1334
rect 180 -1338 209 -1334
rect 213 -1338 294 -1334
rect 383 -1338 451 -1334
rect 474 -1338 502 -1334
rect 536 -1338 565 -1334
rect 569 -1338 650 -1334
rect 739 -1338 809 -1334
rect 825 -1338 860 -1334
rect 894 -1338 923 -1334
rect 927 -1338 1008 -1334
rect -618 -1342 -614 -1338
rect -267 -1342 -263 -1338
rect 91 -1342 95 -1338
rect 447 -1342 451 -1338
rect 805 -1342 809 -1338
rect -1226 -1347 -1169 -1343
rect -1130 -1346 -902 -1342
rect -887 -1346 -804 -1342
rect -783 -1346 -688 -1342
rect -618 -1346 -544 -1342
rect -529 -1346 -446 -1342
rect -425 -1346 -328 -1342
rect -267 -1346 -186 -1342
rect -171 -1346 -88 -1342
rect -67 -1346 29 -1342
rect 91 -1346 172 -1342
rect 187 -1346 270 -1342
rect 291 -1346 386 -1342
rect 447 -1346 528 -1342
rect 543 -1346 626 -1342
rect 647 -1346 742 -1342
rect 805 -1346 886 -1342
rect 901 -1346 984 -1342
rect 1005 -1346 1100 -1342
rect 1215 -1347 1272 -1343
rect -1247 -1354 -1219 -1350
rect -1215 -1354 -1179 -1350
rect -1175 -1354 -1159 -1350
rect -972 -1353 -924 -1349
rect -905 -1353 -776 -1349
rect -614 -1353 -566 -1349
rect -547 -1353 -418 -1349
rect -263 -1353 -208 -1349
rect -189 -1353 -60 -1349
rect 95 -1353 150 -1349
rect 169 -1353 298 -1349
rect 451 -1353 506 -1349
rect 525 -1353 654 -1349
rect 809 -1353 864 -1349
rect 883 -1353 1012 -1349
rect 1097 -1354 1222 -1350
rect 1226 -1354 1262 -1350
rect 1266 -1354 1282 -1350
rect -1279 -1361 -1223 -1357
rect -1219 -1361 -1193 -1357
rect -1189 -1361 -1145 -1357
rect -898 -1360 -794 -1356
rect -790 -1360 -760 -1356
rect -540 -1360 -436 -1356
rect -432 -1360 -402 -1356
rect -182 -1360 -78 -1356
rect -74 -1360 -44 -1356
rect 176 -1360 280 -1356
rect 284 -1360 314 -1356
rect 532 -1360 636 -1356
rect 640 -1360 670 -1356
rect 890 -1360 994 -1356
rect 998 -1360 1028 -1356
rect 1167 -1361 1218 -1357
rect 1222 -1361 1248 -1357
rect 1252 -1361 1296 -1357
rect -1182 -1368 -1124 -1364
rect -924 -1367 -872 -1363
rect -868 -1367 -838 -1363
rect -566 -1367 -514 -1363
rect -510 -1367 -480 -1363
rect -208 -1367 -156 -1363
rect -152 -1367 -122 -1363
rect 150 -1367 202 -1363
rect 206 -1367 236 -1363
rect 506 -1367 558 -1363
rect 562 -1367 592 -1363
rect 864 -1367 916 -1363
rect 920 -1367 950 -1363
rect 1259 -1368 1322 -1364
rect -1200 -1375 -1168 -1371
rect -879 -1375 -847 -1371
rect -801 -1375 -769 -1371
rect -521 -1375 -489 -1371
rect -443 -1375 -411 -1371
rect -163 -1375 -131 -1371
rect -167 -1378 -163 -1375
rect -131 -1378 -127 -1375
rect -85 -1375 -53 -1371
rect -89 -1378 -85 -1375
rect -53 -1378 -49 -1375
rect 195 -1375 227 -1371
rect 191 -1378 195 -1375
rect 227 -1378 231 -1375
rect 273 -1375 305 -1371
rect 269 -1378 273 -1375
rect 305 -1378 309 -1375
rect 551 -1375 583 -1371
rect 547 -1378 551 -1375
rect 583 -1378 587 -1375
rect 629 -1375 661 -1371
rect 625 -1378 629 -1375
rect 661 -1378 665 -1375
rect 909 -1375 941 -1371
rect 905 -1378 909 -1375
rect 941 -1378 945 -1375
rect 987 -1375 1019 -1371
rect 1241 -1375 1273 -1371
rect 983 -1378 987 -1375
rect 1019 -1378 1023 -1375
rect -210 -1386 -206 -1382
rect -184 -1386 -180 -1382
rect -141 -1386 -137 -1382
rect -106 -1386 -102 -1382
rect -62 -1386 -58 -1382
rect -45 -1386 -41 -1382
rect -9 -1386 -5 -1382
rect 12 -1386 16 -1382
rect 148 -1386 152 -1382
rect 174 -1386 178 -1382
rect 217 -1386 221 -1382
rect 252 -1386 256 -1382
rect 296 -1386 300 -1382
rect 313 -1386 317 -1382
rect 349 -1386 353 -1382
rect 370 -1386 374 -1382
rect 504 -1386 508 -1382
rect 530 -1386 534 -1382
rect 573 -1386 577 -1382
rect 608 -1386 612 -1382
rect 652 -1386 656 -1382
rect 669 -1386 673 -1382
rect 705 -1386 709 -1382
rect 726 -1386 730 -1382
rect 862 -1386 866 -1382
rect 888 -1386 892 -1382
rect 931 -1386 935 -1382
rect 966 -1386 970 -1382
rect 1010 -1386 1014 -1382
rect 1027 -1386 1031 -1382
rect 1063 -1386 1067 -1382
rect 1084 -1386 1088 -1382
rect 1804 -1386 1831 -1226
rect -1411 -1390 -1221 -1386
rect -1217 -1390 -1177 -1386
rect -1173 -1390 -1143 -1386
rect -1139 -1390 -926 -1386
rect -922 -1390 -900 -1386
rect -896 -1390 -857 -1386
rect -853 -1390 -822 -1386
rect -818 -1390 -778 -1386
rect -774 -1390 -761 -1386
rect -757 -1390 -725 -1386
rect -721 -1390 -704 -1386
rect -700 -1390 -568 -1386
rect -564 -1390 -542 -1386
rect -538 -1390 -499 -1386
rect -495 -1390 -464 -1386
rect -460 -1390 -420 -1386
rect -416 -1390 -403 -1386
rect -399 -1390 -367 -1386
rect -363 -1390 -346 -1386
rect -342 -1390 -210 -1386
rect -206 -1390 -184 -1386
rect -180 -1390 -141 -1386
rect -137 -1390 -106 -1386
rect -102 -1390 -62 -1386
rect -58 -1390 -45 -1386
rect -41 -1390 -9 -1386
rect -5 -1390 12 -1386
rect 16 -1390 148 -1386
rect 152 -1390 174 -1386
rect 178 -1390 217 -1386
rect 221 -1390 252 -1386
rect 256 -1390 296 -1386
rect 300 -1390 313 -1386
rect 317 -1390 349 -1386
rect 353 -1390 370 -1386
rect 374 -1390 504 -1386
rect 508 -1390 530 -1386
rect 534 -1390 573 -1386
rect 577 -1390 608 -1386
rect 612 -1390 652 -1386
rect 656 -1390 669 -1386
rect 673 -1390 705 -1386
rect 709 -1390 726 -1386
rect 730 -1390 862 -1386
rect 866 -1390 888 -1386
rect 892 -1390 931 -1386
rect 935 -1390 966 -1386
rect 970 -1390 1010 -1386
rect 1014 -1390 1027 -1386
rect 1031 -1390 1063 -1386
rect 1067 -1390 1084 -1386
rect 1088 -1390 1220 -1386
rect 1224 -1390 1264 -1386
rect 1268 -1390 1298 -1386
rect 1302 -1390 1831 -1386
rect -1253 -1397 -688 -1393
rect -1240 -1404 -1124 -1400
rect -972 -1404 -328 -1400
rect -240 -1404 386 -1400
rect 474 -1404 1100 -1400
rect 1188 -1404 1329 -1400
rect -601 -1411 29 -1407
rect 111 -1411 742 -1407
rect 827 -1411 1322 -1407
rect -2055 -1421 -1221 -1417
rect -1217 -1421 -1204 -1417
rect -1200 -1421 -1184 -1417
rect -1180 -1421 -1163 -1417
rect -1159 -1421 -1142 -1417
rect -1138 -1421 -1121 -1417
rect -1117 -1421 -1100 -1417
rect -1096 -1421 -1079 -1417
rect -1075 -1421 -1058 -1417
rect -1054 -1421 -1038 -1417
rect -1034 -1421 -926 -1417
rect -922 -1421 -909 -1417
rect -905 -1421 -889 -1417
rect -885 -1421 -868 -1417
rect -864 -1421 -847 -1417
rect -843 -1421 -826 -1417
rect -822 -1421 -805 -1417
rect -801 -1421 -784 -1417
rect -780 -1421 -763 -1417
rect -759 -1421 -743 -1417
rect -739 -1421 -568 -1417
rect -564 -1421 -551 -1417
rect -547 -1421 -531 -1417
rect -527 -1421 -510 -1417
rect -506 -1421 -489 -1417
rect -485 -1421 -468 -1417
rect -464 -1421 -447 -1417
rect -443 -1421 -426 -1417
rect -422 -1421 -405 -1417
rect -401 -1421 -385 -1417
rect -381 -1421 -210 -1417
rect -206 -1421 -193 -1417
rect -189 -1421 -173 -1417
rect -169 -1421 -152 -1417
rect -148 -1421 -131 -1417
rect -127 -1421 -110 -1417
rect -106 -1421 -89 -1417
rect -85 -1421 -68 -1417
rect -64 -1421 -47 -1417
rect -43 -1421 -27 -1417
rect -23 -1421 148 -1417
rect 152 -1421 165 -1417
rect 169 -1421 185 -1417
rect 189 -1421 206 -1417
rect 210 -1421 227 -1417
rect 231 -1421 248 -1417
rect 252 -1421 269 -1417
rect 273 -1421 290 -1417
rect 294 -1421 311 -1417
rect 315 -1421 331 -1417
rect 335 -1421 504 -1417
rect 508 -1421 521 -1417
rect 525 -1421 541 -1417
rect 545 -1421 562 -1417
rect 566 -1421 583 -1417
rect 587 -1421 604 -1417
rect 608 -1421 625 -1417
rect 629 -1421 646 -1417
rect 650 -1421 667 -1417
rect 671 -1421 687 -1417
rect 691 -1421 862 -1417
rect 866 -1421 879 -1417
rect 883 -1421 899 -1417
rect 903 -1421 920 -1417
rect 924 -1421 941 -1417
rect 945 -1421 962 -1417
rect 966 -1421 983 -1417
rect 987 -1421 1004 -1417
rect 1008 -1421 1025 -1417
rect 1029 -1421 1045 -1417
rect 1049 -1421 1364 -1417
rect -2054 -1588 -2027 -1421
rect -1199 -1469 -1165 -1465
rect -1101 -1469 -1081 -1465
rect -1066 -1469 -931 -1465
rect -904 -1469 -870 -1465
rect -806 -1469 -786 -1465
rect -771 -1469 -573 -1465
rect -546 -1469 -512 -1465
rect -448 -1469 -428 -1465
rect -413 -1469 -215 -1465
rect -188 -1469 -154 -1465
rect -90 -1469 -70 -1465
rect -55 -1469 143 -1465
rect 170 -1469 204 -1465
rect 268 -1469 288 -1465
rect 303 -1469 499 -1465
rect 526 -1469 560 -1465
rect 624 -1469 644 -1465
rect 659 -1469 857 -1465
rect 884 -1469 918 -1465
rect 982 -1469 1002 -1465
rect 1017 -1469 1053 -1465
rect -935 -1473 -931 -1469
rect -577 -1473 -573 -1469
rect -219 -1473 -215 -1469
rect 139 -1473 143 -1469
rect 495 -1473 499 -1469
rect 853 -1473 857 -1469
rect -1240 -1477 -1223 -1473
rect -1219 -1477 -1189 -1473
rect -1168 -1477 -1137 -1473
rect -1108 -1477 -1077 -1473
rect -1066 -1477 -1039 -1473
rect -935 -1477 -928 -1473
rect -924 -1477 -894 -1473
rect -873 -1477 -842 -1473
rect -813 -1477 -782 -1473
rect -771 -1477 -744 -1473
rect -577 -1477 -570 -1473
rect -566 -1477 -536 -1473
rect -515 -1477 -484 -1473
rect -455 -1477 -424 -1473
rect -413 -1477 -386 -1473
rect -219 -1477 -212 -1473
rect -208 -1477 -178 -1473
rect -157 -1477 -126 -1473
rect -97 -1477 -66 -1473
rect -55 -1477 -28 -1473
rect 139 -1477 146 -1473
rect 150 -1477 180 -1473
rect 201 -1477 232 -1473
rect 261 -1477 292 -1473
rect 303 -1477 330 -1473
rect 495 -1477 502 -1473
rect 506 -1477 536 -1473
rect 557 -1477 588 -1473
rect 617 -1477 648 -1473
rect 659 -1477 686 -1473
rect 853 -1477 860 -1473
rect 864 -1477 894 -1473
rect 915 -1477 946 -1473
rect 975 -1477 1006 -1473
rect 1017 -1477 1044 -1473
rect -1226 -1484 -1179 -1480
rect -1143 -1484 -1130 -1480
rect -1126 -1484 -1095 -1480
rect -1059 -1484 -1046 -1480
rect -1042 -1484 -1030 -1480
rect -931 -1484 -884 -1480
rect -848 -1484 -835 -1480
rect -831 -1484 -800 -1480
rect -764 -1484 -751 -1480
rect -747 -1484 -735 -1480
rect -573 -1484 -526 -1480
rect -490 -1484 -477 -1480
rect -473 -1484 -442 -1480
rect -406 -1484 -393 -1480
rect -389 -1484 -377 -1480
rect -215 -1484 -168 -1480
rect -132 -1484 -119 -1480
rect -115 -1484 -84 -1480
rect -48 -1484 -35 -1480
rect -31 -1484 -19 -1480
rect 143 -1484 190 -1480
rect 226 -1484 239 -1480
rect 243 -1484 274 -1480
rect 310 -1484 323 -1480
rect 327 -1484 339 -1480
rect 499 -1484 546 -1480
rect 582 -1484 595 -1480
rect 599 -1484 630 -1480
rect 666 -1484 679 -1480
rect 683 -1484 695 -1480
rect 857 -1484 904 -1480
rect 940 -1484 953 -1480
rect 957 -1484 988 -1480
rect 1024 -1484 1037 -1480
rect 1041 -1484 1053 -1480
rect -1234 -1491 -1219 -1487
rect -1215 -1491 -1105 -1487
rect -1084 -1491 -1053 -1487
rect -939 -1491 -924 -1487
rect -920 -1491 -810 -1487
rect -789 -1491 -758 -1487
rect -581 -1491 -566 -1487
rect -562 -1491 -452 -1487
rect -431 -1491 -400 -1487
rect -223 -1491 -208 -1487
rect -204 -1491 -94 -1487
rect -73 -1491 -42 -1487
rect 135 -1491 150 -1487
rect 154 -1491 264 -1487
rect 285 -1491 316 -1487
rect 491 -1491 506 -1487
rect 510 -1491 620 -1487
rect 641 -1491 672 -1487
rect 849 -1491 864 -1487
rect 868 -1491 978 -1487
rect 999 -1491 1030 -1487
rect -1184 -1498 -1161 -1494
rect -1142 -1498 -1123 -1494
rect -889 -1498 -866 -1494
rect -847 -1498 -828 -1494
rect -531 -1498 -508 -1494
rect -489 -1498 -470 -1494
rect -173 -1498 -150 -1494
rect -131 -1498 -112 -1494
rect 185 -1498 208 -1494
rect 227 -1498 246 -1494
rect 541 -1498 564 -1494
rect 583 -1498 602 -1494
rect 899 -1498 922 -1494
rect 941 -1498 960 -1494
rect 1804 -1509 1831 -1390
rect -1542 -1513 -1221 -1509
rect -1217 -1513 -1204 -1509
rect -1200 -1513 -1163 -1509
rect -1159 -1513 -1121 -1509
rect -1117 -1513 -1079 -1509
rect -1075 -1513 -1038 -1509
rect -1034 -1513 -926 -1509
rect -922 -1513 -909 -1509
rect -905 -1513 -868 -1509
rect -864 -1513 -826 -1509
rect -822 -1513 -784 -1509
rect -780 -1513 -743 -1509
rect -739 -1513 -568 -1509
rect -564 -1513 -551 -1509
rect -547 -1513 -510 -1509
rect -506 -1513 -468 -1509
rect -464 -1513 -426 -1509
rect -422 -1513 -385 -1509
rect -381 -1513 -210 -1509
rect -206 -1513 -193 -1509
rect -189 -1513 -152 -1509
rect -148 -1513 -110 -1509
rect -106 -1513 -68 -1509
rect -64 -1513 -27 -1509
rect -23 -1513 148 -1509
rect 152 -1513 165 -1509
rect 169 -1513 206 -1509
rect 210 -1513 248 -1509
rect 252 -1513 290 -1509
rect 294 -1513 331 -1509
rect 335 -1513 504 -1509
rect 508 -1513 521 -1509
rect 525 -1513 562 -1509
rect 566 -1513 604 -1509
rect 608 -1513 646 -1509
rect 650 -1513 687 -1509
rect 691 -1513 862 -1509
rect 866 -1513 879 -1509
rect 883 -1513 920 -1509
rect 924 -1513 962 -1509
rect 966 -1513 1004 -1509
rect 1008 -1513 1045 -1509
rect 1049 -1513 1831 -1509
rect -2054 -1592 -1221 -1588
rect -1217 -1592 -1204 -1588
rect -1200 -1592 -1184 -1588
rect -1180 -1592 -1163 -1588
rect -1159 -1592 -1142 -1588
rect -1138 -1592 -1121 -1588
rect -1117 -1592 -1100 -1588
rect -1096 -1592 -1079 -1588
rect -1075 -1592 -1058 -1588
rect -1054 -1592 -1038 -1588
rect -1034 -1592 -926 -1588
rect -922 -1592 -909 -1588
rect -905 -1592 -889 -1588
rect -885 -1592 -868 -1588
rect -864 -1592 -847 -1588
rect -843 -1592 -826 -1588
rect -822 -1592 -805 -1588
rect -801 -1592 -784 -1588
rect -780 -1592 -763 -1588
rect -759 -1592 -743 -1588
rect -739 -1592 -568 -1588
rect -564 -1592 -551 -1588
rect -547 -1592 -531 -1588
rect -527 -1592 -510 -1588
rect -506 -1592 -489 -1588
rect -485 -1592 -468 -1588
rect -464 -1592 -447 -1588
rect -443 -1592 -426 -1588
rect -422 -1592 -405 -1588
rect -401 -1592 -385 -1588
rect -381 -1592 -210 -1588
rect -206 -1592 -193 -1588
rect -189 -1592 -173 -1588
rect -169 -1592 -152 -1588
rect -148 -1592 -131 -1588
rect -127 -1592 -110 -1588
rect -106 -1592 -89 -1588
rect -85 -1592 -68 -1588
rect -64 -1592 -47 -1588
rect -43 -1592 -27 -1588
rect -23 -1592 148 -1588
rect 152 -1592 165 -1588
rect 169 -1592 185 -1588
rect 189 -1592 206 -1588
rect 210 -1592 227 -1588
rect 231 -1592 248 -1588
rect 252 -1592 269 -1588
rect 273 -1592 290 -1588
rect 294 -1592 311 -1588
rect 315 -1592 331 -1588
rect 335 -1592 504 -1588
rect 508 -1592 521 -1588
rect 525 -1592 541 -1588
rect 545 -1592 562 -1588
rect 566 -1592 583 -1588
rect 587 -1592 604 -1588
rect 608 -1592 625 -1588
rect 629 -1592 646 -1588
rect 650 -1592 667 -1588
rect 671 -1592 687 -1588
rect 691 -1592 862 -1588
rect 866 -1592 879 -1588
rect 883 -1592 899 -1588
rect 903 -1592 920 -1588
rect 924 -1592 941 -1588
rect 945 -1592 962 -1588
rect 966 -1592 983 -1588
rect 987 -1592 1004 -1588
rect 1008 -1592 1025 -1588
rect 1029 -1592 1045 -1588
rect 1049 -1592 1220 -1588
rect 1224 -1592 1237 -1588
rect 1241 -1592 1257 -1588
rect 1261 -1592 1278 -1588
rect 1282 -1592 1299 -1588
rect 1303 -1592 1320 -1588
rect 1324 -1592 1341 -1588
rect 1345 -1592 1362 -1588
rect 1366 -1592 1383 -1588
rect 1387 -1592 1403 -1588
rect 1407 -1592 1689 -1588
rect -2054 -1759 -2027 -1592
rect -1199 -1640 -1165 -1636
rect -1101 -1640 -1081 -1636
rect -1066 -1640 -1023 -1636
rect -904 -1640 -870 -1636
rect -806 -1640 -786 -1636
rect -771 -1640 -730 -1636
rect -546 -1640 -512 -1636
rect -448 -1640 -428 -1636
rect -413 -1640 -368 -1636
rect -188 -1640 -154 -1636
rect -90 -1640 -70 -1636
rect -55 -1640 -12 -1636
rect 170 -1640 204 -1636
rect 268 -1640 288 -1636
rect 303 -1640 346 -1636
rect 526 -1640 560 -1636
rect 624 -1640 644 -1636
rect 659 -1640 704 -1636
rect 884 -1640 918 -1636
rect 982 -1640 1002 -1636
rect 1017 -1640 1063 -1636
rect 1242 -1640 1276 -1636
rect 1340 -1640 1360 -1636
rect 1375 -1640 1424 -1636
rect -1253 -1648 -1223 -1644
rect -1219 -1648 -1189 -1644
rect -1168 -1648 -1137 -1644
rect -1108 -1648 -1077 -1644
rect -1066 -1648 -1039 -1644
rect -972 -1648 -928 -1644
rect -924 -1648 -894 -1644
rect -873 -1648 -842 -1644
rect -813 -1648 -782 -1644
rect -771 -1648 -744 -1644
rect -601 -1648 -570 -1644
rect -566 -1648 -536 -1644
rect -515 -1648 -484 -1644
rect -455 -1648 -424 -1644
rect -413 -1648 -386 -1644
rect -240 -1648 -212 -1644
rect -208 -1648 -178 -1644
rect -157 -1648 -126 -1644
rect -97 -1648 -66 -1644
rect -55 -1648 -28 -1644
rect 111 -1648 146 -1644
rect 150 -1648 180 -1644
rect 201 -1648 232 -1644
rect 261 -1648 292 -1644
rect 303 -1648 330 -1644
rect 474 -1648 502 -1644
rect 506 -1648 536 -1644
rect 557 -1648 588 -1644
rect 617 -1648 648 -1644
rect 659 -1648 686 -1644
rect 827 -1648 860 -1644
rect 864 -1648 894 -1644
rect 915 -1648 946 -1644
rect 975 -1648 1006 -1644
rect 1017 -1648 1044 -1644
rect 1188 -1648 1218 -1644
rect 1222 -1648 1252 -1644
rect 1273 -1648 1304 -1644
rect 1333 -1648 1364 -1644
rect 1375 -1648 1402 -1644
rect -1226 -1655 -1179 -1651
rect -1143 -1655 -1130 -1651
rect -1126 -1655 -1095 -1651
rect -1059 -1655 -1046 -1651
rect -1042 -1655 -1030 -1651
rect -931 -1655 -884 -1651
rect -848 -1655 -835 -1651
rect -831 -1655 -800 -1651
rect -764 -1655 -751 -1651
rect -747 -1655 -735 -1651
rect -573 -1655 -526 -1651
rect -490 -1655 -477 -1651
rect -473 -1655 -442 -1651
rect -406 -1655 -393 -1651
rect -389 -1655 -377 -1651
rect -215 -1655 -168 -1651
rect -132 -1655 -119 -1651
rect -115 -1655 -84 -1651
rect -48 -1655 -35 -1651
rect -31 -1655 -19 -1651
rect 143 -1655 190 -1651
rect 226 -1655 239 -1651
rect 243 -1655 274 -1651
rect 310 -1655 323 -1651
rect 327 -1655 339 -1651
rect 499 -1655 546 -1651
rect 582 -1655 595 -1651
rect 599 -1655 630 -1651
rect 666 -1655 679 -1651
rect 683 -1655 695 -1651
rect 857 -1655 904 -1651
rect 940 -1655 953 -1651
rect 957 -1655 988 -1651
rect 1024 -1655 1037 -1651
rect 1041 -1655 1053 -1651
rect 1215 -1655 1262 -1651
rect 1298 -1655 1311 -1651
rect 1315 -1655 1346 -1651
rect 1382 -1655 1395 -1651
rect 1399 -1655 1411 -1651
rect -1234 -1662 -1219 -1658
rect -1215 -1662 -1105 -1658
rect -1084 -1662 -1053 -1658
rect -939 -1662 -924 -1658
rect -920 -1662 -810 -1658
rect -789 -1662 -758 -1658
rect -581 -1662 -566 -1658
rect -562 -1662 -452 -1658
rect -431 -1662 -400 -1658
rect -223 -1662 -208 -1658
rect -204 -1662 -94 -1658
rect -73 -1662 -42 -1658
rect 135 -1662 150 -1658
rect 154 -1662 264 -1658
rect 285 -1662 316 -1658
rect 491 -1662 506 -1658
rect 510 -1662 620 -1658
rect 641 -1662 672 -1658
rect 849 -1662 864 -1658
rect 868 -1662 978 -1658
rect 999 -1662 1030 -1658
rect 1207 -1662 1222 -1658
rect 1226 -1662 1336 -1658
rect 1357 -1662 1388 -1658
rect -1184 -1669 -1161 -1665
rect -1142 -1669 -1123 -1665
rect -889 -1669 -866 -1665
rect -847 -1669 -828 -1665
rect -531 -1669 -508 -1665
rect -489 -1669 -470 -1665
rect -173 -1669 -150 -1665
rect -131 -1669 -112 -1665
rect 185 -1669 208 -1665
rect 227 -1669 246 -1665
rect 541 -1669 564 -1665
rect 583 -1669 602 -1665
rect 899 -1669 922 -1665
rect 941 -1669 960 -1665
rect 1257 -1669 1280 -1665
rect 1299 -1669 1318 -1665
rect 1804 -1680 1831 -1513
rect -1792 -1684 -1221 -1680
rect -1217 -1684 -1204 -1680
rect -1200 -1684 -1163 -1680
rect -1159 -1684 -1121 -1680
rect -1117 -1684 -1079 -1680
rect -1075 -1684 -1038 -1680
rect -1034 -1684 -926 -1680
rect -922 -1684 -909 -1680
rect -905 -1684 -868 -1680
rect -864 -1684 -826 -1680
rect -822 -1684 -784 -1680
rect -780 -1684 -743 -1680
rect -739 -1684 -568 -1680
rect -564 -1684 -551 -1680
rect -547 -1684 -510 -1680
rect -506 -1684 -468 -1680
rect -464 -1684 -426 -1680
rect -422 -1684 -385 -1680
rect -381 -1684 -210 -1680
rect -206 -1684 -193 -1680
rect -189 -1684 -152 -1680
rect -148 -1684 -110 -1680
rect -106 -1684 -68 -1680
rect -64 -1684 -27 -1680
rect -23 -1684 148 -1680
rect 152 -1684 165 -1680
rect 169 -1684 206 -1680
rect 210 -1684 248 -1680
rect 252 -1684 290 -1680
rect 294 -1684 331 -1680
rect 335 -1684 504 -1680
rect 508 -1684 521 -1680
rect 525 -1684 562 -1680
rect 566 -1684 604 -1680
rect 608 -1684 646 -1680
rect 650 -1684 687 -1680
rect 691 -1684 862 -1680
rect 866 -1684 879 -1680
rect 883 -1684 920 -1680
rect 924 -1684 962 -1680
rect 966 -1684 1004 -1680
rect 1008 -1684 1045 -1680
rect 1049 -1684 1220 -1680
rect 1224 -1684 1237 -1680
rect 1241 -1684 1278 -1680
rect 1282 -1684 1320 -1680
rect 1324 -1684 1362 -1680
rect 1366 -1684 1403 -1680
rect 1407 -1684 1831 -1680
rect -1253 -1691 -1023 -1687
rect -972 -1692 -730 -1688
rect -601 -1692 -368 -1688
rect -240 -1691 -12 -1687
rect 111 -1692 346 -1688
rect 474 -1691 704 -1687
rect 827 -1691 1063 -1687
rect 1188 -1692 1424 -1688
rect -2054 -1763 -1550 -1759
rect -1546 -1763 -1533 -1759
rect -1529 -1763 -1513 -1759
rect -1509 -1763 -1492 -1759
rect -1488 -1763 -1471 -1759
rect -1467 -1763 -1450 -1759
rect -1446 -1763 -1429 -1759
rect -1425 -1763 -1408 -1759
rect -1404 -1763 -1387 -1759
rect -1383 -1763 -1367 -1759
rect -1363 -1763 -1221 -1759
rect -1217 -1763 -1204 -1759
rect -1200 -1763 -1184 -1759
rect -1180 -1763 -1163 -1759
rect -1159 -1763 -1142 -1759
rect -1138 -1763 -1121 -1759
rect -1117 -1763 -1100 -1759
rect -1096 -1763 -1079 -1759
rect -1075 -1763 -1058 -1759
rect -1054 -1763 -1038 -1759
rect -1034 -1763 -926 -1759
rect -922 -1763 -909 -1759
rect -905 -1763 -889 -1759
rect -885 -1763 -868 -1759
rect -864 -1763 -847 -1759
rect -843 -1763 -826 -1759
rect -822 -1763 -805 -1759
rect -801 -1763 -784 -1759
rect -780 -1763 -763 -1759
rect -759 -1763 -743 -1759
rect -739 -1763 -568 -1759
rect -564 -1763 -551 -1759
rect -547 -1763 -531 -1759
rect -527 -1763 -510 -1759
rect -506 -1763 -489 -1759
rect -485 -1763 -468 -1759
rect -464 -1763 -447 -1759
rect -443 -1763 -426 -1759
rect -422 -1763 -405 -1759
rect -401 -1763 -385 -1759
rect -381 -1763 -210 -1759
rect -206 -1763 -193 -1759
rect -189 -1763 -173 -1759
rect -169 -1763 -152 -1759
rect -148 -1763 -131 -1759
rect -127 -1763 -110 -1759
rect -106 -1763 -89 -1759
rect -85 -1763 -68 -1759
rect -64 -1763 -47 -1759
rect -43 -1763 -27 -1759
rect -23 -1763 148 -1759
rect 152 -1763 165 -1759
rect 169 -1763 185 -1759
rect 189 -1763 206 -1759
rect 210 -1763 227 -1759
rect 231 -1763 248 -1759
rect 252 -1763 269 -1759
rect 273 -1763 290 -1759
rect 294 -1763 311 -1759
rect 315 -1763 331 -1759
rect 335 -1763 504 -1759
rect 508 -1763 521 -1759
rect 525 -1763 541 -1759
rect 545 -1763 562 -1759
rect 566 -1763 583 -1759
rect 587 -1763 604 -1759
rect 608 -1763 625 -1759
rect 629 -1763 646 -1759
rect 650 -1763 667 -1759
rect 671 -1763 687 -1759
rect 691 -1763 862 -1759
rect 866 -1763 879 -1759
rect 883 -1763 899 -1759
rect 903 -1763 920 -1759
rect 924 -1763 941 -1759
rect 945 -1763 962 -1759
rect 966 -1763 983 -1759
rect 987 -1763 1004 -1759
rect 1008 -1763 1025 -1759
rect 1029 -1763 1045 -1759
rect 1049 -1763 1220 -1759
rect 1224 -1763 1237 -1759
rect 1241 -1763 1257 -1759
rect 1261 -1763 1278 -1759
rect 1282 -1763 1299 -1759
rect 1303 -1763 1320 -1759
rect 1324 -1763 1341 -1759
rect 1345 -1763 1362 -1759
rect 1366 -1763 1383 -1759
rect 1387 -1763 1403 -1759
rect 1407 -1763 1682 -1759
rect -2054 -1866 -2027 -1763
rect -1395 -1803 -1351 -1799
rect -1528 -1811 -1494 -1807
rect -1430 -1811 -1410 -1807
rect -1199 -1811 -1165 -1807
rect -1101 -1811 -1081 -1807
rect -1066 -1811 -1016 -1807
rect -904 -1811 -870 -1807
rect -806 -1811 -786 -1807
rect -771 -1811 -723 -1807
rect -546 -1811 -512 -1807
rect -448 -1811 -428 -1807
rect -413 -1811 -366 -1807
rect -188 -1811 -154 -1807
rect -90 -1811 -70 -1807
rect -55 -1811 -9 -1807
rect 170 -1811 204 -1807
rect 268 -1811 288 -1807
rect 303 -1811 350 -1807
rect 526 -1811 560 -1807
rect 624 -1811 644 -1807
rect 659 -1811 703 -1807
rect 884 -1811 918 -1807
rect 982 -1811 1002 -1807
rect 1017 -1811 1060 -1807
rect 1242 -1811 1276 -1807
rect 1340 -1811 1360 -1807
rect 1375 -1811 1419 -1807
rect -1563 -1819 -1552 -1815
rect -1548 -1819 -1518 -1815
rect -1497 -1819 -1466 -1815
rect -1437 -1819 -1406 -1815
rect -1395 -1819 -1368 -1815
rect -1315 -1819 -1223 -1815
rect -1219 -1819 -1189 -1815
rect -1168 -1819 -1137 -1815
rect -1108 -1819 -1077 -1815
rect -1066 -1819 -1039 -1815
rect -945 -1819 -928 -1815
rect -924 -1819 -894 -1815
rect -873 -1819 -842 -1815
rect -813 -1819 -782 -1815
rect -771 -1819 -744 -1815
rect -587 -1819 -570 -1815
rect -566 -1819 -536 -1815
rect -515 -1819 -484 -1815
rect -455 -1819 -424 -1815
rect -413 -1819 -386 -1815
rect -229 -1819 -212 -1815
rect -208 -1819 -178 -1815
rect -157 -1819 -126 -1815
rect -97 -1819 -66 -1815
rect -55 -1819 -28 -1815
rect 129 -1819 146 -1815
rect 150 -1819 180 -1815
rect 201 -1819 232 -1815
rect 261 -1819 292 -1815
rect 303 -1819 330 -1815
rect 485 -1819 502 -1815
rect 506 -1819 536 -1815
rect 557 -1819 588 -1815
rect 617 -1819 648 -1815
rect 659 -1819 686 -1815
rect 843 -1819 860 -1815
rect 864 -1819 894 -1815
rect 915 -1819 946 -1815
rect 975 -1819 1006 -1815
rect 1017 -1819 1044 -1815
rect 1201 -1819 1218 -1815
rect 1222 -1819 1252 -1815
rect 1273 -1819 1304 -1815
rect 1333 -1819 1364 -1815
rect 1375 -1819 1402 -1815
rect -1555 -1826 -1508 -1822
rect -1472 -1826 -1459 -1822
rect -1455 -1826 -1424 -1822
rect -1388 -1826 -1375 -1822
rect -1371 -1826 -1359 -1822
rect -1226 -1826 -1179 -1822
rect -1143 -1826 -1130 -1822
rect -1126 -1826 -1095 -1822
rect -1059 -1826 -1046 -1822
rect -1042 -1826 -1030 -1822
rect -931 -1826 -884 -1822
rect -848 -1826 -835 -1822
rect -831 -1826 -800 -1822
rect -764 -1826 -751 -1822
rect -747 -1826 -735 -1822
rect -573 -1826 -526 -1822
rect -490 -1826 -477 -1822
rect -473 -1826 -442 -1822
rect -406 -1826 -393 -1822
rect -389 -1826 -377 -1822
rect -215 -1826 -168 -1822
rect -132 -1826 -119 -1822
rect -115 -1826 -84 -1822
rect -48 -1826 -35 -1822
rect -31 -1826 -19 -1822
rect 143 -1826 190 -1822
rect 226 -1826 239 -1822
rect 243 -1826 274 -1822
rect 310 -1826 323 -1822
rect 327 -1826 339 -1822
rect 499 -1826 546 -1822
rect 582 -1826 595 -1822
rect 599 -1826 630 -1822
rect 666 -1826 679 -1822
rect 683 -1826 695 -1822
rect 857 -1826 904 -1822
rect 940 -1826 953 -1822
rect 957 -1826 988 -1822
rect 1024 -1826 1037 -1822
rect 1041 -1826 1053 -1822
rect 1215 -1826 1262 -1822
rect 1298 -1826 1311 -1822
rect 1315 -1826 1346 -1822
rect 1382 -1826 1395 -1822
rect 1399 -1826 1411 -1822
rect -1563 -1833 -1548 -1829
rect -1544 -1833 -1434 -1829
rect -1413 -1833 -1382 -1829
rect -1234 -1833 -1219 -1829
rect -1215 -1833 -1105 -1829
rect -1084 -1833 -1053 -1829
rect -939 -1833 -924 -1829
rect -920 -1833 -810 -1829
rect -789 -1833 -758 -1829
rect -581 -1833 -566 -1829
rect -562 -1833 -452 -1829
rect -431 -1833 -400 -1829
rect -223 -1833 -208 -1829
rect -204 -1833 -94 -1829
rect -73 -1833 -42 -1829
rect 135 -1833 150 -1829
rect 154 -1833 264 -1829
rect 285 -1833 316 -1829
rect 491 -1833 506 -1829
rect 510 -1833 620 -1829
rect 641 -1833 672 -1829
rect 849 -1833 864 -1829
rect 868 -1833 978 -1829
rect 999 -1833 1030 -1829
rect 1207 -1833 1222 -1829
rect 1226 -1833 1336 -1829
rect 1357 -1833 1388 -1829
rect -1513 -1840 -1490 -1836
rect -1471 -1840 -1452 -1836
rect -1184 -1840 -1161 -1836
rect -1142 -1840 -1123 -1836
rect -889 -1840 -866 -1836
rect -847 -1840 -828 -1836
rect -531 -1840 -508 -1836
rect -489 -1840 -470 -1836
rect -173 -1840 -150 -1836
rect -131 -1840 -112 -1836
rect 185 -1840 208 -1836
rect 227 -1840 246 -1836
rect 541 -1840 564 -1836
rect 583 -1840 602 -1836
rect 899 -1840 922 -1836
rect 941 -1840 960 -1836
rect 1257 -1840 1280 -1836
rect 1299 -1840 1318 -1836
rect 1804 -1851 1831 -1684
rect -1789 -1855 -1550 -1851
rect -1546 -1855 -1533 -1851
rect -1529 -1855 -1492 -1851
rect -1488 -1855 -1450 -1851
rect -1446 -1855 -1408 -1851
rect -1404 -1855 -1367 -1851
rect -1363 -1855 -1221 -1851
rect -1217 -1855 -1204 -1851
rect -1200 -1855 -1163 -1851
rect -1159 -1855 -1121 -1851
rect -1117 -1855 -1079 -1851
rect -1075 -1855 -1038 -1851
rect -1034 -1855 -926 -1851
rect -922 -1855 -909 -1851
rect -905 -1855 -868 -1851
rect -864 -1855 -826 -1851
rect -822 -1855 -784 -1851
rect -780 -1855 -743 -1851
rect -739 -1855 -568 -1851
rect -564 -1855 -551 -1851
rect -547 -1855 -510 -1851
rect -506 -1855 -468 -1851
rect -464 -1855 -426 -1851
rect -422 -1855 -385 -1851
rect -381 -1855 -210 -1851
rect -206 -1855 -193 -1851
rect -189 -1855 -152 -1851
rect -148 -1855 -110 -1851
rect -106 -1855 -68 -1851
rect -64 -1855 -27 -1851
rect -23 -1855 148 -1851
rect 152 -1855 165 -1851
rect 169 -1855 206 -1851
rect 210 -1855 248 -1851
rect 252 -1855 290 -1851
rect 294 -1855 331 -1851
rect 335 -1855 504 -1851
rect 508 -1855 521 -1851
rect 525 -1855 562 -1851
rect 566 -1855 604 -1851
rect 608 -1855 646 -1851
rect 650 -1855 687 -1851
rect 691 -1855 862 -1851
rect 866 -1855 879 -1851
rect 883 -1855 920 -1851
rect 924 -1855 962 -1851
rect 966 -1855 1004 -1851
rect 1008 -1855 1045 -1851
rect 1049 -1855 1220 -1851
rect 1224 -1855 1237 -1851
rect 1241 -1855 1278 -1851
rect 1282 -1855 1320 -1851
rect 1324 -1855 1362 -1851
rect 1366 -1855 1403 -1851
rect 1407 -1855 1831 -1851
rect -2054 -1870 -1309 -1866
rect -1305 -1870 -1292 -1866
rect -1288 -1870 -935 -1866
rect -931 -1870 -918 -1866
rect -914 -1870 -577 -1866
rect -573 -1870 -560 -1866
rect -556 -1870 -219 -1866
rect -215 -1870 -202 -1866
rect -198 -1870 139 -1866
rect 143 -1870 156 -1866
rect 160 -1870 495 -1866
rect 499 -1870 512 -1866
rect 516 -1870 853 -1866
rect 857 -1870 870 -1866
rect 874 -1870 1211 -1866
rect 1215 -1870 1228 -1866
rect 1232 -1870 1589 -1866
rect -2054 -2025 -2027 -1870
rect -1304 -1902 -1016 -1898
rect -930 -1902 -723 -1898
rect -572 -1902 -366 -1898
rect -214 -1902 -9 -1898
rect 144 -1902 350 -1898
rect 500 -1902 703 -1898
rect 858 -1902 1060 -1898
rect 1216 -1902 1419 -1898
rect -1347 -1910 -1297 -1906
rect -1293 -1910 -923 -1906
rect -919 -1910 -565 -1906
rect -561 -1910 -207 -1906
rect -203 -1910 151 -1906
rect 155 -1910 507 -1906
rect 511 -1910 865 -1906
rect 869 -1910 1223 -1906
rect 1227 -1910 1589 -1906
rect -964 -1923 -909 -1919
rect -614 -1923 -551 -1919
rect -258 -1923 -193 -1919
rect 97 -1923 165 -1919
rect 455 -1923 521 -1919
rect 813 -1923 879 -1919
rect 1171 -1923 1237 -1919
rect 1804 -1958 1831 -1855
rect -1429 -1962 -1292 -1958
rect -1288 -1962 -918 -1958
rect -914 -1962 -560 -1958
rect -556 -1962 -202 -1958
rect -198 -1962 156 -1958
rect 160 -1962 512 -1958
rect 516 -1962 870 -1958
rect 874 -1962 1228 -1958
rect 1232 -1962 1831 -1958
rect -2054 -2029 -1225 -2025
rect -1221 -2029 -1208 -2025
rect -1204 -2029 -1168 -2025
rect -1164 -2029 -1147 -2025
rect -1143 -2029 -926 -2025
rect -922 -2029 -900 -2025
rect -896 -2029 -883 -2025
rect -879 -2029 -843 -2025
rect -839 -2029 -822 -2025
rect -818 -2029 -805 -2025
rect -801 -2029 -765 -2025
rect -761 -2029 -741 -2025
rect -737 -2029 -704 -2025
rect -700 -2029 -568 -2025
rect -564 -2029 -542 -2025
rect -538 -2029 -525 -2025
rect -521 -2029 -485 -2025
rect -481 -2029 -464 -2025
rect -460 -2029 -447 -2025
rect -443 -2029 -407 -2025
rect -403 -2029 -383 -2025
rect -379 -2029 -346 -2025
rect -342 -2029 -210 -2025
rect -206 -2029 -184 -2025
rect -180 -2029 -167 -2025
rect -163 -2029 -127 -2025
rect -123 -2029 -106 -2025
rect -102 -2029 -89 -2025
rect -85 -2029 -49 -2025
rect -45 -2029 -25 -2025
rect -21 -2029 12 -2025
rect 16 -2029 148 -2025
rect 152 -2029 174 -2025
rect 178 -2029 191 -2025
rect 195 -2029 231 -2025
rect 235 -2029 252 -2025
rect 256 -2029 269 -2025
rect 273 -2029 309 -2025
rect 313 -2029 333 -2025
rect 337 -2029 370 -2025
rect 374 -2029 504 -2025
rect 508 -2029 530 -2025
rect 534 -2029 547 -2025
rect 551 -2029 587 -2025
rect 591 -2029 608 -2025
rect 612 -2029 625 -2025
rect 629 -2029 665 -2025
rect 669 -2029 689 -2025
rect 693 -2029 726 -2025
rect 730 -2029 862 -2025
rect 866 -2029 888 -2025
rect 892 -2029 905 -2025
rect 909 -2029 945 -2025
rect 949 -2029 966 -2025
rect 970 -2029 983 -2025
rect 987 -2029 1023 -2025
rect 1027 -2029 1047 -2025
rect 1051 -2029 1084 -2025
rect 1088 -2029 1220 -2025
rect 1224 -2029 1246 -2025
rect 1250 -2029 1263 -2025
rect 1267 -2029 1303 -2025
rect 1307 -2029 1324 -2025
rect 1328 -2029 1341 -2025
rect 1345 -2029 1381 -2025
rect 1385 -2029 1405 -2025
rect 1409 -2029 1442 -2025
rect 1446 -2029 1589 -2025
rect -2054 -2169 -2027 -2029
rect -926 -2033 -922 -2029
rect -900 -2033 -896 -2029
rect -883 -2033 -879 -2029
rect -843 -2033 -839 -2029
rect -822 -2033 -818 -2029
rect -805 -2033 -801 -2029
rect -765 -2033 -761 -2029
rect -741 -2033 -737 -2029
rect -704 -2033 -700 -2029
rect -568 -2033 -564 -2029
rect -542 -2033 -538 -2029
rect -525 -2033 -521 -2029
rect -485 -2033 -481 -2029
rect -464 -2033 -460 -2029
rect -447 -2033 -443 -2029
rect -407 -2033 -403 -2029
rect -383 -2033 -379 -2029
rect -346 -2033 -342 -2029
rect -210 -2033 -206 -2029
rect -184 -2033 -180 -2029
rect -167 -2033 -163 -2029
rect -127 -2033 -123 -2029
rect -106 -2033 -102 -2029
rect -89 -2033 -85 -2029
rect -49 -2033 -45 -2029
rect -25 -2033 -21 -2029
rect 12 -2033 16 -2029
rect 148 -2033 152 -2029
rect 174 -2033 178 -2029
rect 191 -2033 195 -2029
rect 231 -2033 235 -2029
rect 252 -2033 256 -2029
rect 269 -2033 273 -2029
rect 309 -2033 313 -2029
rect 333 -2033 337 -2029
rect 370 -2033 374 -2029
rect 504 -2033 508 -2029
rect 530 -2033 534 -2029
rect 547 -2033 551 -2029
rect 587 -2033 591 -2029
rect 608 -2033 612 -2029
rect 625 -2033 629 -2029
rect 665 -2033 669 -2029
rect 689 -2033 693 -2029
rect 726 -2033 730 -2029
rect 862 -2033 866 -2029
rect 888 -2033 892 -2029
rect 905 -2033 909 -2029
rect 945 -2033 949 -2029
rect 966 -2033 970 -2029
rect 983 -2033 987 -2029
rect 1023 -2033 1027 -2029
rect 1047 -2033 1051 -2029
rect 1084 -2033 1088 -2029
rect 1220 -2033 1224 -2029
rect 1246 -2033 1250 -2029
rect 1263 -2033 1267 -2029
rect 1303 -2033 1307 -2029
rect 1324 -2033 1328 -2029
rect 1341 -2033 1345 -2029
rect 1381 -2033 1385 -2029
rect 1405 -2033 1409 -2029
rect 1442 -2033 1446 -2029
rect -920 -2048 -858 -2044
rect -854 -2048 -824 -2044
rect -776 -2048 -746 -2044
rect -562 -2048 -500 -2044
rect -496 -2048 -466 -2044
rect -418 -2048 -388 -2044
rect -204 -2048 -142 -2044
rect -138 -2048 -108 -2044
rect -60 -2048 -30 -2044
rect 154 -2048 216 -2044
rect 220 -2048 250 -2044
rect 298 -2048 328 -2044
rect 510 -2048 572 -2044
rect 576 -2048 606 -2044
rect 654 -2048 684 -2044
rect 868 -2048 930 -2044
rect 934 -2048 964 -2044
rect 1012 -2048 1042 -2044
rect 1226 -2048 1288 -2044
rect 1292 -2048 1322 -2044
rect 1370 -2048 1400 -2044
rect -913 -2055 -882 -2051
rect -555 -2055 -524 -2051
rect -197 -2055 -166 -2051
rect 161 -2055 192 -2051
rect 517 -2055 548 -2051
rect 875 -2055 906 -2051
rect 1233 -2055 1264 -2051
rect -931 -2062 -848 -2058
rect -809 -2062 -706 -2058
rect -573 -2062 -490 -2058
rect -451 -2062 -348 -2058
rect -215 -2062 -132 -2058
rect -93 -2062 10 -2058
rect 143 -2062 226 -2058
rect 265 -2062 368 -2058
rect 499 -2062 582 -2058
rect 621 -2062 724 -2058
rect 857 -2062 940 -2058
rect 979 -2062 1082 -2058
rect 1215 -2062 1298 -2058
rect 1337 -2062 1440 -2058
rect -972 -2069 -928 -2065
rect -894 -2069 -865 -2065
rect -861 -2069 -780 -2065
rect -691 -2069 -614 -2065
rect -601 -2069 -570 -2065
rect -536 -2069 -507 -2065
rect -503 -2069 -422 -2065
rect -333 -2066 -258 -2062
rect -618 -2073 -614 -2069
rect -262 -2073 -258 -2066
rect -240 -2069 -212 -2065
rect -178 -2069 -149 -2065
rect -145 -2069 -64 -2065
rect 25 -2069 97 -2065
rect 111 -2069 146 -2065
rect 180 -2069 209 -2065
rect 213 -2069 294 -2065
rect 383 -2069 455 -2065
rect 474 -2069 502 -2065
rect 536 -2069 565 -2065
rect 569 -2069 650 -2065
rect 739 -2069 813 -2065
rect 827 -2069 860 -2065
rect 894 -2069 923 -2065
rect 927 -2069 1008 -2065
rect 1097 -2067 1162 -2063
rect 93 -2073 97 -2069
rect 451 -2073 455 -2069
rect 809 -2073 813 -2069
rect 1158 -2073 1162 -2067
rect 1171 -2069 1218 -2065
rect 1252 -2069 1281 -2065
rect 1285 -2069 1366 -2065
rect -1230 -2078 -1173 -2074
rect -1134 -2077 -902 -2073
rect -887 -2077 -804 -2073
rect -783 -2077 -687 -2073
rect -618 -2077 -544 -2073
rect -529 -2077 -446 -2073
rect -425 -2077 -328 -2073
rect -262 -2077 -186 -2073
rect -171 -2077 -88 -2073
rect -67 -2077 29 -2073
rect 93 -2077 172 -2073
rect 187 -2077 270 -2073
rect 291 -2077 388 -2073
rect 451 -2077 528 -2073
rect 543 -2077 626 -2073
rect 647 -2077 743 -2073
rect 809 -2077 886 -2073
rect 901 -2077 984 -2073
rect 1005 -2077 1101 -2073
rect 1158 -2077 1244 -2073
rect 1259 -2077 1342 -2073
rect 1363 -2077 1466 -2073
rect -1253 -2085 -1223 -2081
rect -1219 -2085 -1183 -2081
rect -1179 -2085 -1163 -2081
rect -964 -2084 -924 -2080
rect -905 -2084 -776 -2080
rect -614 -2084 -566 -2080
rect -547 -2084 -418 -2080
rect -258 -2084 -208 -2080
rect -189 -2084 -60 -2080
rect 97 -2084 150 -2080
rect 169 -2084 298 -2080
rect 455 -2084 506 -2080
rect 525 -2084 654 -2080
rect 813 -2084 864 -2080
rect 883 -2084 1012 -2080
rect 1188 -2084 1222 -2080
rect 1241 -2084 1370 -2080
rect -1279 -2092 -1227 -2088
rect -1223 -2092 -1197 -2088
rect -1193 -2092 -1149 -2088
rect -898 -2091 -794 -2087
rect -790 -2091 -760 -2087
rect -540 -2091 -436 -2087
rect -432 -2091 -402 -2087
rect -182 -2091 -78 -2087
rect -74 -2091 -44 -2087
rect 176 -2091 280 -2087
rect 284 -2091 314 -2087
rect 532 -2091 636 -2087
rect 640 -2091 670 -2087
rect 890 -2091 994 -2087
rect 998 -2091 1028 -2087
rect 1248 -2091 1352 -2087
rect 1356 -2091 1386 -2087
rect -1186 -2099 -1115 -2095
rect -924 -2098 -872 -2094
rect -868 -2098 -838 -2094
rect -566 -2098 -514 -2094
rect -510 -2098 -480 -2094
rect -208 -2098 -156 -2094
rect -152 -2098 -122 -2094
rect 150 -2098 202 -2094
rect 206 -2098 236 -2094
rect 506 -2098 558 -2094
rect 562 -2098 592 -2094
rect 864 -2098 916 -2094
rect 920 -2098 950 -2094
rect 1222 -2098 1274 -2094
rect 1278 -2098 1308 -2094
rect -1204 -2106 -1172 -2102
rect -879 -2106 -847 -2102
rect -883 -2109 -879 -2106
rect -847 -2109 -843 -2106
rect -801 -2106 -769 -2102
rect -805 -2109 -801 -2106
rect -769 -2109 -765 -2106
rect -521 -2106 -489 -2102
rect -525 -2109 -521 -2106
rect -489 -2109 -485 -2106
rect -443 -2106 -411 -2102
rect -447 -2109 -443 -2106
rect -411 -2109 -407 -2106
rect -163 -2106 -131 -2102
rect -167 -2109 -163 -2106
rect -131 -2109 -127 -2106
rect -85 -2106 -53 -2102
rect -89 -2109 -85 -2106
rect -53 -2109 -49 -2106
rect 195 -2106 227 -2102
rect 191 -2109 195 -2106
rect 227 -2109 231 -2106
rect 273 -2106 305 -2102
rect 269 -2109 273 -2106
rect 305 -2109 309 -2106
rect 551 -2106 583 -2102
rect 547 -2109 551 -2106
rect 583 -2109 587 -2106
rect 629 -2106 661 -2102
rect 625 -2109 629 -2106
rect 661 -2109 665 -2106
rect 909 -2106 941 -2102
rect 905 -2109 909 -2106
rect 941 -2109 945 -2106
rect 987 -2106 1019 -2102
rect 983 -2109 987 -2106
rect 1019 -2109 1023 -2106
rect 1267 -2106 1299 -2102
rect 1263 -2109 1267 -2106
rect 1299 -2109 1303 -2106
rect 1345 -2106 1377 -2102
rect 1341 -2109 1345 -2106
rect 1377 -2109 1381 -2106
rect -926 -2117 -922 -2113
rect -900 -2117 -896 -2113
rect -857 -2117 -853 -2113
rect -822 -2117 -818 -2113
rect -778 -2117 -774 -2113
rect -761 -2117 -757 -2113
rect -725 -2117 -721 -2113
rect -704 -2117 -700 -2113
rect -568 -2117 -564 -2113
rect -542 -2117 -538 -2113
rect -499 -2117 -495 -2113
rect -464 -2117 -460 -2113
rect -420 -2117 -416 -2113
rect -403 -2117 -399 -2113
rect -367 -2117 -363 -2113
rect -346 -2117 -342 -2113
rect -210 -2117 -206 -2113
rect -184 -2117 -180 -2113
rect -141 -2117 -137 -2113
rect -106 -2117 -102 -2113
rect -62 -2117 -58 -2113
rect -45 -2117 -41 -2113
rect -9 -2117 -5 -2113
rect 12 -2117 16 -2113
rect 148 -2117 152 -2113
rect 174 -2117 178 -2113
rect 217 -2117 221 -2113
rect 252 -2117 256 -2113
rect 296 -2117 300 -2113
rect 313 -2117 317 -2113
rect 349 -2117 353 -2113
rect 370 -2117 374 -2113
rect 504 -2117 508 -2113
rect 530 -2117 534 -2113
rect 573 -2117 577 -2113
rect 608 -2117 612 -2113
rect 652 -2117 656 -2113
rect 669 -2117 673 -2113
rect 705 -2117 709 -2113
rect 726 -2117 730 -2113
rect 862 -2117 866 -2113
rect 888 -2117 892 -2113
rect 931 -2117 935 -2113
rect 966 -2117 970 -2113
rect 1010 -2117 1014 -2113
rect 1027 -2117 1031 -2113
rect 1063 -2117 1067 -2113
rect 1084 -2117 1088 -2113
rect 1220 -2117 1224 -2113
rect 1246 -2117 1250 -2113
rect 1289 -2117 1293 -2113
rect 1324 -2117 1328 -2113
rect 1368 -2117 1372 -2113
rect 1385 -2117 1389 -2113
rect 1421 -2117 1425 -2113
rect 1442 -2117 1446 -2113
rect 1804 -2117 1831 -1962
rect -1411 -2121 -1225 -2117
rect -1221 -2121 -1181 -2117
rect -1177 -2121 -1147 -2117
rect -1143 -2121 -926 -2117
rect -922 -2121 -900 -2117
rect -896 -2121 -857 -2117
rect -853 -2121 -822 -2117
rect -818 -2121 -778 -2117
rect -774 -2121 -761 -2117
rect -757 -2121 -725 -2117
rect -721 -2121 -704 -2117
rect -700 -2121 -568 -2117
rect -564 -2121 -542 -2117
rect -538 -2121 -499 -2117
rect -495 -2121 -464 -2117
rect -460 -2121 -420 -2117
rect -416 -2121 -403 -2117
rect -399 -2121 -367 -2117
rect -363 -2121 -346 -2117
rect -342 -2121 -210 -2117
rect -206 -2121 -184 -2117
rect -180 -2121 -141 -2117
rect -137 -2121 -106 -2117
rect -102 -2121 -62 -2117
rect -58 -2121 -45 -2117
rect -41 -2121 -9 -2117
rect -5 -2121 12 -2117
rect 16 -2121 148 -2117
rect 152 -2121 174 -2117
rect 178 -2121 217 -2117
rect 221 -2121 252 -2117
rect 256 -2121 296 -2117
rect 300 -2121 313 -2117
rect 317 -2121 349 -2117
rect 353 -2121 370 -2117
rect 374 -2121 504 -2117
rect 508 -2121 530 -2117
rect 534 -2121 573 -2117
rect 577 -2121 608 -2117
rect 612 -2121 652 -2117
rect 656 -2121 669 -2117
rect 673 -2121 705 -2117
rect 709 -2121 726 -2117
rect 730 -2121 862 -2117
rect 866 -2121 888 -2117
rect 892 -2121 931 -2117
rect 935 -2121 966 -2117
rect 970 -2121 1010 -2117
rect 1014 -2121 1027 -2117
rect 1031 -2121 1063 -2117
rect 1067 -2121 1084 -2117
rect 1088 -2121 1220 -2117
rect 1224 -2121 1246 -2117
rect 1250 -2121 1289 -2117
rect 1293 -2121 1324 -2117
rect 1328 -2121 1368 -2117
rect 1372 -2121 1385 -2117
rect 1389 -2121 1421 -2117
rect 1425 -2121 1442 -2117
rect 1446 -2121 1831 -2117
rect -1253 -2128 -687 -2124
rect -599 -2128 29 -2124
rect 115 -2128 743 -2124
rect 828 -2128 1466 -2124
rect -1241 -2135 -1115 -2131
rect -959 -2135 -328 -2131
rect -245 -2135 388 -2131
rect 469 -2135 1101 -2131
rect 1188 -2135 1451 -2131
rect -2054 -2173 -1225 -2169
rect -1221 -2173 -1208 -2169
rect -1204 -2173 -1188 -2169
rect -1184 -2173 -1167 -2169
rect -1163 -2173 -1146 -2169
rect -1142 -2173 -1125 -2169
rect -1121 -2173 -1104 -2169
rect -1100 -2173 -1083 -2169
rect -1079 -2173 -1062 -2169
rect -1058 -2173 -1042 -2169
rect -1038 -2173 -926 -2169
rect -922 -2173 -909 -2169
rect -905 -2173 -889 -2169
rect -885 -2173 -868 -2169
rect -864 -2173 -847 -2169
rect -843 -2173 -826 -2169
rect -822 -2173 -805 -2169
rect -801 -2173 -784 -2169
rect -780 -2173 -763 -2169
rect -759 -2173 -743 -2169
rect -739 -2173 -568 -2169
rect -564 -2173 -551 -2169
rect -547 -2173 -531 -2169
rect -527 -2173 -510 -2169
rect -506 -2173 -489 -2169
rect -485 -2173 -468 -2169
rect -464 -2173 -447 -2169
rect -443 -2173 -426 -2169
rect -422 -2173 -405 -2169
rect -401 -2173 -385 -2169
rect -381 -2173 -210 -2169
rect -206 -2173 -193 -2169
rect -189 -2173 -173 -2169
rect -169 -2173 -152 -2169
rect -148 -2173 -131 -2169
rect -127 -2173 -110 -2169
rect -106 -2173 -89 -2169
rect -85 -2173 -68 -2169
rect -64 -2173 -47 -2169
rect -43 -2173 -27 -2169
rect -23 -2173 148 -2169
rect 152 -2173 165 -2169
rect 169 -2173 185 -2169
rect 189 -2173 206 -2169
rect 210 -2173 227 -2169
rect 231 -2173 248 -2169
rect 252 -2173 269 -2169
rect 273 -2173 290 -2169
rect 294 -2173 311 -2169
rect 315 -2173 331 -2169
rect 335 -2173 504 -2169
rect 508 -2173 521 -2169
rect 525 -2173 541 -2169
rect 545 -2173 562 -2169
rect 566 -2173 583 -2169
rect 587 -2173 604 -2169
rect 608 -2173 625 -2169
rect 629 -2173 646 -2169
rect 650 -2173 667 -2169
rect 671 -2173 687 -2169
rect 691 -2173 1607 -2169
rect -2054 -2340 -2027 -2173
rect -1203 -2221 -1169 -2217
rect -1105 -2221 -1085 -2217
rect -1070 -2221 -931 -2217
rect -904 -2221 -870 -2217
rect -806 -2221 -786 -2217
rect -771 -2221 -573 -2217
rect -546 -2221 -512 -2217
rect -448 -2221 -428 -2217
rect -413 -2221 -215 -2217
rect -188 -2221 -154 -2217
rect -90 -2221 -70 -2217
rect -55 -2221 143 -2217
rect 170 -2221 204 -2217
rect 268 -2221 288 -2217
rect 303 -2221 499 -2217
rect 526 -2221 560 -2217
rect 624 -2221 644 -2217
rect 659 -2221 695 -2217
rect -935 -2225 -931 -2221
rect -577 -2225 -573 -2221
rect -219 -2225 -215 -2221
rect 139 -2225 143 -2221
rect 495 -2225 499 -2221
rect -1241 -2229 -1227 -2225
rect -1223 -2229 -1193 -2225
rect -1172 -2229 -1141 -2225
rect -1112 -2229 -1081 -2225
rect -1070 -2229 -1043 -2225
rect -935 -2229 -928 -2225
rect -924 -2229 -894 -2225
rect -873 -2229 -842 -2225
rect -813 -2229 -782 -2225
rect -771 -2229 -744 -2225
rect -577 -2229 -570 -2225
rect -566 -2229 -536 -2225
rect -515 -2229 -484 -2225
rect -455 -2229 -424 -2225
rect -413 -2229 -386 -2225
rect -219 -2229 -212 -2225
rect -208 -2229 -178 -2225
rect -157 -2229 -126 -2225
rect -97 -2229 -66 -2225
rect -55 -2229 -28 -2225
rect 139 -2229 146 -2225
rect 150 -2229 180 -2225
rect 201 -2229 232 -2225
rect 261 -2229 292 -2225
rect 303 -2229 330 -2225
rect 495 -2229 502 -2225
rect 506 -2229 536 -2225
rect 557 -2229 588 -2225
rect 617 -2229 648 -2225
rect 659 -2229 686 -2225
rect -1230 -2236 -1183 -2232
rect -1147 -2236 -1134 -2232
rect -1130 -2236 -1099 -2232
rect -1063 -2236 -1050 -2232
rect -1046 -2236 -1034 -2232
rect -931 -2236 -884 -2232
rect -848 -2236 -835 -2232
rect -831 -2236 -800 -2232
rect -764 -2236 -751 -2232
rect -747 -2236 -735 -2232
rect -573 -2236 -526 -2232
rect -490 -2236 -477 -2232
rect -473 -2236 -442 -2232
rect -406 -2236 -393 -2232
rect -389 -2236 -377 -2232
rect -215 -2236 -168 -2232
rect -132 -2236 -119 -2232
rect -115 -2236 -84 -2232
rect -48 -2236 -35 -2232
rect -31 -2236 -19 -2232
rect 143 -2236 190 -2232
rect 226 -2236 239 -2232
rect 243 -2236 274 -2232
rect 310 -2236 323 -2232
rect 327 -2236 339 -2232
rect 499 -2236 546 -2232
rect 582 -2236 595 -2232
rect 599 -2236 630 -2232
rect 666 -2236 679 -2232
rect 683 -2236 695 -2232
rect -1238 -2243 -1223 -2239
rect -1219 -2243 -1109 -2239
rect -1088 -2243 -1057 -2239
rect -939 -2243 -924 -2239
rect -920 -2243 -810 -2239
rect -789 -2243 -758 -2239
rect -581 -2243 -566 -2239
rect -562 -2243 -452 -2239
rect -431 -2243 -400 -2239
rect -223 -2243 -208 -2239
rect -204 -2243 -94 -2239
rect -73 -2243 -42 -2239
rect 135 -2243 150 -2239
rect 154 -2243 264 -2239
rect 285 -2243 316 -2239
rect 491 -2243 506 -2239
rect 510 -2243 620 -2239
rect 641 -2243 672 -2239
rect -1188 -2250 -1165 -2246
rect -1146 -2250 -1127 -2246
rect -889 -2250 -866 -2246
rect -847 -2250 -828 -2246
rect -531 -2250 -508 -2246
rect -489 -2250 -470 -2246
rect -173 -2250 -150 -2246
rect -131 -2250 -112 -2246
rect 185 -2250 208 -2246
rect 227 -2250 246 -2246
rect 541 -2250 564 -2246
rect 583 -2250 602 -2246
rect 1804 -2261 1831 -2121
rect -1857 -2265 -1225 -2261
rect -1221 -2265 -1208 -2261
rect -1204 -2265 -1167 -2261
rect -1163 -2265 -1125 -2261
rect -1121 -2265 -1083 -2261
rect -1079 -2265 -1042 -2261
rect -1038 -2265 -926 -2261
rect -922 -2265 -909 -2261
rect -905 -2265 -868 -2261
rect -864 -2265 -826 -2261
rect -822 -2265 -784 -2261
rect -780 -2265 -743 -2261
rect -739 -2265 -568 -2261
rect -564 -2265 -551 -2261
rect -547 -2265 -510 -2261
rect -506 -2265 -468 -2261
rect -464 -2265 -426 -2261
rect -422 -2265 -385 -2261
rect -381 -2265 -210 -2261
rect -206 -2265 -193 -2261
rect -189 -2265 -152 -2261
rect -148 -2265 -110 -2261
rect -106 -2265 -68 -2261
rect -64 -2265 -27 -2261
rect -23 -2265 148 -2261
rect 152 -2265 165 -2261
rect 169 -2265 206 -2261
rect 210 -2265 248 -2261
rect 252 -2265 290 -2261
rect 294 -2265 331 -2261
rect 335 -2265 504 -2261
rect 508 -2265 521 -2261
rect 525 -2265 562 -2261
rect 566 -2265 604 -2261
rect 608 -2265 646 -2261
rect 650 -2265 687 -2261
rect 691 -2265 1831 -2261
rect -2054 -2344 -1550 -2340
rect -1546 -2344 -1533 -2340
rect -1529 -2344 -1513 -2340
rect -1509 -2344 -1492 -2340
rect -1488 -2344 -1471 -2340
rect -1467 -2344 -1450 -2340
rect -1446 -2344 -1429 -2340
rect -1425 -2344 -1408 -2340
rect -1404 -2344 -1387 -2340
rect -1383 -2344 -1367 -2340
rect -1363 -2344 -1225 -2340
rect -1221 -2344 -1208 -2340
rect -1204 -2344 -1188 -2340
rect -1184 -2344 -1167 -2340
rect -1163 -2344 -1146 -2340
rect -1142 -2344 -1125 -2340
rect -1121 -2344 -1104 -2340
rect -1100 -2344 -1083 -2340
rect -1079 -2344 -1062 -2340
rect -1058 -2344 -1042 -2340
rect -1038 -2344 -926 -2340
rect -922 -2344 -909 -2340
rect -905 -2344 -889 -2340
rect -885 -2344 -868 -2340
rect -864 -2344 -847 -2340
rect -843 -2344 -826 -2340
rect -822 -2344 -805 -2340
rect -801 -2344 -784 -2340
rect -780 -2344 -763 -2340
rect -759 -2344 -743 -2340
rect -739 -2344 -568 -2340
rect -564 -2344 -551 -2340
rect -547 -2344 -531 -2340
rect -527 -2344 -510 -2340
rect -506 -2344 -489 -2340
rect -485 -2344 -468 -2340
rect -464 -2344 -447 -2340
rect -443 -2344 -426 -2340
rect -422 -2344 -405 -2340
rect -401 -2344 -385 -2340
rect -381 -2344 -210 -2340
rect -206 -2344 -193 -2340
rect -189 -2344 -173 -2340
rect -169 -2344 -152 -2340
rect -148 -2344 -131 -2340
rect -127 -2344 -110 -2340
rect -106 -2344 -89 -2340
rect -85 -2344 -68 -2340
rect -64 -2344 -47 -2340
rect -43 -2344 -27 -2340
rect -23 -2344 148 -2340
rect 152 -2344 165 -2340
rect 169 -2344 185 -2340
rect 189 -2344 206 -2340
rect 210 -2344 227 -2340
rect 231 -2344 248 -2340
rect 252 -2344 269 -2340
rect 273 -2344 290 -2340
rect 294 -2344 311 -2340
rect 315 -2344 331 -2340
rect 335 -2344 504 -2340
rect 508 -2344 521 -2340
rect 525 -2344 541 -2340
rect 545 -2344 562 -2340
rect 566 -2344 583 -2340
rect 587 -2344 604 -2340
rect 608 -2344 625 -2340
rect 629 -2344 646 -2340
rect 650 -2344 667 -2340
rect 671 -2344 687 -2340
rect 691 -2344 862 -2340
rect 866 -2344 879 -2340
rect 883 -2344 899 -2340
rect 903 -2344 920 -2340
rect 924 -2344 941 -2340
rect 945 -2344 962 -2340
rect 966 -2344 983 -2340
rect 987 -2344 1004 -2340
rect 1008 -2344 1025 -2340
rect 1029 -2344 1045 -2340
rect 1049 -2344 1220 -2340
rect 1224 -2344 1237 -2340
rect 1241 -2344 1257 -2340
rect 1261 -2344 1278 -2340
rect 1282 -2344 1299 -2340
rect 1303 -2344 1320 -2340
rect 1324 -2344 1341 -2340
rect 1345 -2344 1362 -2340
rect 1366 -2344 1383 -2340
rect 1387 -2344 1403 -2340
rect 1407 -2344 1616 -2340
rect -2054 -2511 -2027 -2344
rect -1528 -2392 -1494 -2388
rect -1430 -2392 -1410 -2388
rect -1395 -2392 -1350 -2388
rect -1203 -2392 -1169 -2388
rect -1105 -2392 -1085 -2388
rect -1070 -2392 -1024 -2388
rect -904 -2392 -870 -2388
rect -806 -2392 -786 -2388
rect -771 -2392 -723 -2388
rect -546 -2392 -512 -2388
rect -448 -2392 -428 -2388
rect -413 -2392 -366 -2388
rect -188 -2392 -154 -2388
rect -90 -2392 -70 -2388
rect -55 -2392 -8 -2388
rect 170 -2392 204 -2388
rect 268 -2392 288 -2388
rect 303 -2392 346 -2388
rect 526 -2392 560 -2388
rect 624 -2392 644 -2388
rect 659 -2392 705 -2388
rect 884 -2392 918 -2388
rect 982 -2392 1002 -2388
rect 1017 -2392 1062 -2388
rect 1242 -2392 1276 -2388
rect 1340 -2392 1360 -2388
rect 1375 -2392 1421 -2388
rect -1563 -2400 -1552 -2396
rect -1548 -2400 -1518 -2396
rect -1497 -2400 -1466 -2396
rect -1437 -2400 -1406 -2396
rect -1395 -2400 -1368 -2396
rect -1253 -2400 -1227 -2396
rect -1223 -2400 -1193 -2396
rect -1172 -2400 -1141 -2396
rect -1112 -2400 -1081 -2396
rect -1070 -2400 -1043 -2396
rect -959 -2400 -928 -2396
rect -924 -2400 -894 -2396
rect -873 -2400 -842 -2396
rect -813 -2400 -782 -2396
rect -771 -2400 -744 -2396
rect -599 -2400 -570 -2396
rect -566 -2400 -536 -2396
rect -515 -2400 -484 -2396
rect -455 -2400 -424 -2396
rect -413 -2400 -386 -2396
rect -245 -2400 -212 -2396
rect -208 -2400 -178 -2396
rect -157 -2400 -126 -2396
rect -97 -2400 -66 -2396
rect -55 -2400 -28 -2396
rect 115 -2400 146 -2396
rect 150 -2400 180 -2396
rect 201 -2400 232 -2396
rect 261 -2400 292 -2396
rect 303 -2400 330 -2396
rect 469 -2400 502 -2396
rect 506 -2400 536 -2396
rect 557 -2400 588 -2396
rect 617 -2400 648 -2396
rect 659 -2400 686 -2396
rect 828 -2400 860 -2396
rect 864 -2400 894 -2396
rect 915 -2400 946 -2396
rect 975 -2400 1006 -2396
rect 1017 -2400 1044 -2396
rect 1188 -2400 1218 -2396
rect 1222 -2400 1252 -2396
rect 1273 -2400 1304 -2396
rect 1333 -2400 1364 -2396
rect 1375 -2400 1402 -2396
rect -1555 -2407 -1508 -2403
rect -1472 -2407 -1459 -2403
rect -1455 -2407 -1424 -2403
rect -1388 -2407 -1375 -2403
rect -1371 -2407 -1359 -2403
rect -1230 -2407 -1183 -2403
rect -1147 -2407 -1134 -2403
rect -1130 -2407 -1099 -2403
rect -1063 -2407 -1050 -2403
rect -1046 -2407 -1034 -2403
rect -931 -2407 -884 -2403
rect -848 -2407 -835 -2403
rect -831 -2407 -800 -2403
rect -764 -2407 -751 -2403
rect -747 -2407 -735 -2403
rect -573 -2407 -526 -2403
rect -490 -2407 -477 -2403
rect -473 -2407 -442 -2403
rect -406 -2407 -393 -2403
rect -389 -2407 -377 -2403
rect -215 -2407 -168 -2403
rect -132 -2407 -119 -2403
rect -115 -2407 -84 -2403
rect -48 -2407 -35 -2403
rect -31 -2407 -19 -2403
rect 143 -2407 190 -2403
rect 226 -2407 239 -2403
rect 243 -2407 274 -2403
rect 310 -2407 323 -2403
rect 327 -2407 339 -2403
rect 499 -2407 546 -2403
rect 582 -2407 595 -2403
rect 599 -2407 630 -2403
rect 666 -2407 679 -2403
rect 683 -2407 695 -2403
rect 857 -2407 904 -2403
rect 940 -2407 953 -2403
rect 957 -2407 988 -2403
rect 1024 -2407 1037 -2403
rect 1041 -2407 1053 -2403
rect 1215 -2407 1262 -2403
rect 1298 -2407 1311 -2403
rect 1315 -2407 1346 -2403
rect 1382 -2407 1395 -2403
rect 1399 -2407 1411 -2403
rect -1563 -2414 -1548 -2410
rect -1544 -2414 -1434 -2410
rect -1413 -2414 -1382 -2410
rect -1238 -2414 -1223 -2410
rect -1219 -2414 -1109 -2410
rect -1088 -2414 -1057 -2410
rect -939 -2414 -924 -2410
rect -920 -2414 -810 -2410
rect -789 -2414 -758 -2410
rect -581 -2414 -566 -2410
rect -562 -2414 -452 -2410
rect -431 -2414 -400 -2410
rect -223 -2414 -208 -2410
rect -204 -2414 -94 -2410
rect -73 -2414 -42 -2410
rect 135 -2414 150 -2410
rect 154 -2414 264 -2410
rect 285 -2414 316 -2410
rect 491 -2414 506 -2410
rect 510 -2414 620 -2410
rect 641 -2414 672 -2410
rect 849 -2414 864 -2410
rect 868 -2414 978 -2410
rect 999 -2414 1030 -2410
rect 1207 -2414 1222 -2410
rect 1226 -2414 1336 -2410
rect 1357 -2414 1388 -2410
rect -1513 -2421 -1490 -2417
rect -1471 -2421 -1452 -2417
rect -1188 -2421 -1165 -2417
rect -1146 -2421 -1127 -2417
rect -889 -2421 -866 -2417
rect -847 -2421 -828 -2417
rect -531 -2421 -508 -2417
rect -489 -2421 -470 -2417
rect -173 -2421 -150 -2417
rect -131 -2421 -112 -2417
rect 185 -2421 208 -2417
rect 227 -2421 246 -2417
rect 541 -2421 564 -2417
rect 583 -2421 602 -2417
rect 899 -2421 922 -2417
rect 941 -2421 960 -2417
rect 1257 -2421 1280 -2417
rect 1299 -2421 1318 -2417
rect 1804 -2432 1831 -2265
rect -1851 -2436 -1550 -2432
rect -1546 -2436 -1533 -2432
rect -1529 -2436 -1492 -2432
rect -1488 -2436 -1450 -2432
rect -1446 -2436 -1408 -2432
rect -1404 -2436 -1367 -2432
rect -1363 -2436 -1225 -2432
rect -1221 -2436 -1208 -2432
rect -1204 -2436 -1167 -2432
rect -1163 -2436 -1125 -2432
rect -1121 -2436 -1083 -2432
rect -1079 -2436 -1042 -2432
rect -1038 -2436 -926 -2432
rect -922 -2436 -909 -2432
rect -905 -2436 -868 -2432
rect -864 -2436 -826 -2432
rect -822 -2436 -784 -2432
rect -780 -2436 -743 -2432
rect -739 -2436 -568 -2432
rect -564 -2436 -551 -2432
rect -547 -2436 -510 -2432
rect -506 -2436 -468 -2432
rect -464 -2436 -426 -2432
rect -422 -2436 -385 -2432
rect -381 -2436 -210 -2432
rect -206 -2436 -193 -2432
rect -189 -2436 -152 -2432
rect -148 -2436 -110 -2432
rect -106 -2436 -68 -2432
rect -64 -2436 -27 -2432
rect -23 -2436 148 -2432
rect 152 -2436 165 -2432
rect 169 -2436 206 -2432
rect 210 -2436 248 -2432
rect 252 -2436 290 -2432
rect 294 -2436 331 -2432
rect 335 -2436 504 -2432
rect 508 -2436 521 -2432
rect 525 -2436 562 -2432
rect 566 -2436 604 -2432
rect 608 -2436 646 -2432
rect 650 -2436 687 -2432
rect 691 -2436 862 -2432
rect 866 -2436 879 -2432
rect 883 -2436 920 -2432
rect 924 -2436 962 -2432
rect 966 -2436 1004 -2432
rect 1008 -2436 1045 -2432
rect 1049 -2436 1220 -2432
rect 1224 -2436 1237 -2432
rect 1241 -2436 1278 -2432
rect 1282 -2436 1320 -2432
rect 1324 -2436 1362 -2432
rect 1366 -2436 1403 -2432
rect 1407 -2436 1831 -2432
rect -1577 -2444 -1350 -2440
rect -1253 -2444 -1024 -2440
rect -959 -2443 -723 -2439
rect -599 -2444 -366 -2440
rect -245 -2444 -8 -2440
rect 115 -2443 346 -2439
rect 469 -2443 705 -2439
rect 828 -2444 1062 -2440
rect 1188 -2444 1421 -2440
rect -2054 -2515 -1550 -2511
rect -1546 -2515 -1533 -2511
rect -1529 -2515 -1513 -2511
rect -1509 -2515 -1492 -2511
rect -1488 -2515 -1471 -2511
rect -1467 -2515 -1450 -2511
rect -1446 -2515 -1429 -2511
rect -1425 -2515 -1408 -2511
rect -1404 -2515 -1387 -2511
rect -1383 -2515 -1367 -2511
rect -1363 -2515 -1225 -2511
rect -1221 -2515 -1208 -2511
rect -1204 -2515 -1188 -2511
rect -1184 -2515 -1167 -2511
rect -1163 -2515 -1146 -2511
rect -1142 -2515 -1125 -2511
rect -1121 -2515 -1104 -2511
rect -1100 -2515 -1083 -2511
rect -1079 -2515 -1062 -2511
rect -1058 -2515 -1042 -2511
rect -1038 -2515 -926 -2511
rect -922 -2515 -909 -2511
rect -905 -2515 -889 -2511
rect -885 -2515 -868 -2511
rect -864 -2515 -847 -2511
rect -843 -2515 -826 -2511
rect -822 -2515 -805 -2511
rect -801 -2515 -784 -2511
rect -780 -2515 -763 -2511
rect -759 -2515 -743 -2511
rect -739 -2515 -568 -2511
rect -564 -2515 -551 -2511
rect -547 -2515 -531 -2511
rect -527 -2515 -510 -2511
rect -506 -2515 -489 -2511
rect -485 -2515 -468 -2511
rect -464 -2515 -447 -2511
rect -443 -2515 -426 -2511
rect -422 -2515 -405 -2511
rect -401 -2515 -385 -2511
rect -381 -2515 -211 -2511
rect -207 -2515 -194 -2511
rect -190 -2515 -174 -2511
rect -170 -2515 -153 -2511
rect -149 -2515 -132 -2511
rect -128 -2515 -111 -2511
rect -107 -2515 -90 -2511
rect -86 -2515 -69 -2511
rect -65 -2515 -48 -2511
rect -44 -2515 -28 -2511
rect -24 -2515 148 -2511
rect 152 -2515 165 -2511
rect 169 -2515 185 -2511
rect 189 -2515 206 -2511
rect 210 -2515 227 -2511
rect 231 -2515 248 -2511
rect 252 -2515 269 -2511
rect 273 -2515 290 -2511
rect 294 -2515 311 -2511
rect 315 -2515 331 -2511
rect 335 -2515 504 -2511
rect 508 -2515 521 -2511
rect 525 -2515 541 -2511
rect 545 -2515 562 -2511
rect 566 -2515 583 -2511
rect 587 -2515 604 -2511
rect 608 -2515 625 -2511
rect 629 -2515 646 -2511
rect 650 -2515 667 -2511
rect 671 -2515 687 -2511
rect 691 -2515 862 -2511
rect 866 -2515 879 -2511
rect 883 -2515 899 -2511
rect 903 -2515 920 -2511
rect 924 -2515 941 -2511
rect 945 -2515 962 -2511
rect 966 -2515 983 -2511
rect 987 -2515 1004 -2511
rect 1008 -2515 1025 -2511
rect 1029 -2515 1045 -2511
rect 1049 -2515 1220 -2511
rect 1224 -2515 1237 -2511
rect 1241 -2515 1257 -2511
rect 1261 -2515 1278 -2511
rect 1282 -2515 1299 -2511
rect 1303 -2515 1320 -2511
rect 1324 -2515 1341 -2511
rect 1345 -2515 1362 -2511
rect 1366 -2515 1383 -2511
rect 1387 -2515 1403 -2511
rect 1407 -2515 1605 -2511
rect -2054 -2616 -2027 -2515
rect -1528 -2563 -1494 -2559
rect -1430 -2563 -1410 -2559
rect -1395 -2563 -1355 -2559
rect -1203 -2563 -1169 -2559
rect -1105 -2563 -1085 -2559
rect -1070 -2563 -1026 -2559
rect -904 -2563 -870 -2559
rect -806 -2563 -786 -2559
rect -771 -2563 -720 -2559
rect -546 -2563 -512 -2559
rect -448 -2563 -428 -2559
rect -413 -2563 -373 -2559
rect -189 -2563 -155 -2559
rect -91 -2563 -71 -2559
rect -56 -2563 -12 -2559
rect 170 -2563 204 -2559
rect 268 -2563 288 -2559
rect 303 -2563 347 -2559
rect 526 -2563 560 -2559
rect 624 -2563 644 -2559
rect 659 -2563 703 -2559
rect 884 -2563 918 -2559
rect 982 -2563 1002 -2559
rect 1017 -2563 1062 -2559
rect 1242 -2563 1276 -2559
rect 1340 -2563 1360 -2559
rect 1375 -2563 1419 -2559
rect -1577 -2571 -1552 -2567
rect -1548 -2571 -1518 -2567
rect -1497 -2571 -1466 -2567
rect -1437 -2571 -1406 -2567
rect -1395 -2571 -1368 -2567
rect -1315 -2571 -1227 -2567
rect -1223 -2571 -1193 -2567
rect -1172 -2571 -1141 -2567
rect -1112 -2571 -1081 -2567
rect -1070 -2571 -1043 -2567
rect -945 -2571 -928 -2567
rect -924 -2571 -894 -2567
rect -873 -2571 -842 -2567
rect -813 -2571 -782 -2567
rect -771 -2571 -744 -2567
rect -587 -2571 -570 -2567
rect -566 -2571 -536 -2567
rect -515 -2571 -484 -2567
rect -455 -2571 -424 -2567
rect -413 -2571 -386 -2567
rect -229 -2571 -213 -2567
rect -209 -2571 -179 -2567
rect -158 -2571 -127 -2567
rect -98 -2571 -67 -2567
rect -56 -2571 -29 -2567
rect 129 -2571 146 -2567
rect 150 -2571 180 -2567
rect 201 -2571 232 -2567
rect 261 -2571 292 -2567
rect 303 -2571 330 -2567
rect 485 -2571 502 -2567
rect 506 -2571 536 -2567
rect 557 -2571 588 -2567
rect 617 -2571 648 -2567
rect 659 -2571 686 -2567
rect 843 -2571 860 -2567
rect 864 -2571 894 -2567
rect 915 -2571 946 -2567
rect 975 -2571 1006 -2567
rect 1017 -2571 1044 -2567
rect 1201 -2571 1218 -2567
rect 1222 -2571 1252 -2567
rect 1273 -2571 1304 -2567
rect 1333 -2571 1364 -2567
rect 1375 -2571 1402 -2567
rect -1555 -2578 -1508 -2574
rect -1472 -2578 -1459 -2574
rect -1455 -2578 -1424 -2574
rect -1388 -2578 -1375 -2574
rect -1371 -2578 -1359 -2574
rect -1230 -2578 -1183 -2574
rect -1147 -2578 -1134 -2574
rect -1130 -2578 -1099 -2574
rect -1063 -2578 -1050 -2574
rect -1046 -2578 -1034 -2574
rect -931 -2578 -884 -2574
rect -848 -2578 -835 -2574
rect -831 -2578 -800 -2574
rect -764 -2578 -751 -2574
rect -747 -2578 -735 -2574
rect -573 -2578 -526 -2574
rect -490 -2578 -477 -2574
rect -473 -2578 -442 -2574
rect -406 -2578 -393 -2574
rect -389 -2578 -377 -2574
rect -216 -2578 -169 -2574
rect -133 -2578 -120 -2574
rect -116 -2578 -85 -2574
rect -49 -2578 -36 -2574
rect -32 -2578 -20 -2574
rect 143 -2578 190 -2574
rect 226 -2578 239 -2574
rect 243 -2578 274 -2574
rect 310 -2578 323 -2574
rect 327 -2578 339 -2574
rect 499 -2578 546 -2574
rect 582 -2578 595 -2574
rect 599 -2578 630 -2574
rect 666 -2578 679 -2574
rect 683 -2578 695 -2574
rect 857 -2578 904 -2574
rect 940 -2578 953 -2574
rect 957 -2578 988 -2574
rect 1024 -2578 1037 -2574
rect 1041 -2578 1053 -2574
rect 1215 -2578 1262 -2574
rect 1298 -2578 1311 -2574
rect 1315 -2578 1346 -2574
rect 1382 -2578 1395 -2574
rect 1399 -2578 1411 -2574
rect -1563 -2585 -1548 -2581
rect -1544 -2585 -1434 -2581
rect -1413 -2585 -1382 -2581
rect -1238 -2585 -1223 -2581
rect -1219 -2585 -1109 -2581
rect -1088 -2585 -1057 -2581
rect -939 -2585 -924 -2581
rect -920 -2585 -810 -2581
rect -789 -2585 -758 -2581
rect -581 -2585 -566 -2581
rect -562 -2585 -452 -2581
rect -431 -2585 -400 -2581
rect -224 -2585 -209 -2581
rect -205 -2585 -95 -2581
rect -74 -2585 -43 -2581
rect 135 -2585 150 -2581
rect 154 -2585 264 -2581
rect 285 -2585 316 -2581
rect 491 -2585 506 -2581
rect 510 -2585 620 -2581
rect 641 -2585 672 -2581
rect 849 -2585 864 -2581
rect 868 -2585 978 -2581
rect 999 -2585 1030 -2581
rect 1207 -2585 1222 -2581
rect 1226 -2585 1336 -2581
rect 1357 -2585 1388 -2581
rect -1513 -2592 -1490 -2588
rect -1471 -2592 -1452 -2588
rect -1188 -2592 -1165 -2588
rect -1146 -2592 -1127 -2588
rect -889 -2592 -866 -2588
rect -847 -2592 -828 -2588
rect -531 -2592 -508 -2588
rect -489 -2592 -470 -2588
rect -174 -2592 -151 -2588
rect -132 -2592 -113 -2588
rect 185 -2592 208 -2588
rect 227 -2592 246 -2588
rect 541 -2592 564 -2588
rect 583 -2592 602 -2588
rect 899 -2592 922 -2588
rect 941 -2592 960 -2588
rect 1257 -2592 1280 -2588
rect 1299 -2592 1318 -2588
rect 1804 -2603 1831 -2436
rect -1906 -2607 -1550 -2603
rect -1546 -2607 -1533 -2603
rect -1529 -2607 -1492 -2603
rect -1488 -2607 -1450 -2603
rect -1446 -2607 -1408 -2603
rect -1404 -2607 -1367 -2603
rect -1363 -2607 -1225 -2603
rect -1221 -2607 -1208 -2603
rect -1204 -2607 -1167 -2603
rect -1163 -2607 -1125 -2603
rect -1121 -2607 -1083 -2603
rect -1079 -2607 -1042 -2603
rect -1038 -2607 -926 -2603
rect -922 -2607 -909 -2603
rect -905 -2607 -868 -2603
rect -864 -2607 -826 -2603
rect -822 -2607 -784 -2603
rect -780 -2607 -743 -2603
rect -739 -2607 -568 -2603
rect -564 -2607 -551 -2603
rect -547 -2607 -510 -2603
rect -506 -2607 -468 -2603
rect -464 -2607 -426 -2603
rect -422 -2607 -385 -2603
rect -381 -2607 -211 -2603
rect -207 -2607 -194 -2603
rect -190 -2607 -153 -2603
rect -149 -2607 -111 -2603
rect -107 -2607 -69 -2603
rect -65 -2607 -28 -2603
rect -24 -2607 148 -2603
rect 152 -2607 165 -2603
rect 169 -2607 206 -2603
rect 210 -2607 248 -2603
rect 252 -2607 290 -2603
rect 294 -2607 331 -2603
rect 335 -2607 504 -2603
rect 508 -2607 521 -2603
rect 525 -2607 562 -2603
rect 566 -2607 604 -2603
rect 608 -2607 646 -2603
rect 650 -2607 687 -2603
rect 691 -2607 862 -2603
rect 866 -2607 879 -2603
rect 883 -2607 920 -2603
rect 924 -2607 962 -2603
rect 966 -2607 1004 -2603
rect 1008 -2607 1045 -2603
rect 1049 -2607 1220 -2603
rect 1224 -2607 1237 -2603
rect 1241 -2607 1278 -2603
rect 1282 -2607 1320 -2603
rect 1324 -2607 1362 -2603
rect 1366 -2607 1403 -2603
rect 1407 -2607 1831 -2603
rect -2054 -2620 -1309 -2616
rect -1305 -2620 -1292 -2616
rect -1288 -2620 -935 -2616
rect -931 -2620 -918 -2616
rect -914 -2620 -577 -2616
rect -573 -2620 -560 -2616
rect -556 -2620 -219 -2616
rect -215 -2620 -202 -2616
rect -198 -2620 139 -2616
rect 143 -2620 156 -2616
rect 160 -2620 495 -2616
rect 499 -2620 512 -2616
rect 516 -2620 853 -2616
rect 857 -2620 870 -2616
rect 874 -2620 1211 -2616
rect 1215 -2620 1228 -2616
rect 1232 -2620 1589 -2616
rect -2054 -2775 -2027 -2620
rect -1304 -2652 -1026 -2648
rect -930 -2652 -720 -2648
rect -572 -2652 -373 -2648
rect -214 -2652 -12 -2648
rect 144 -2652 347 -2648
rect 500 -2652 703 -2648
rect 858 -2652 1062 -2648
rect 1216 -2652 1419 -2648
rect -1351 -2660 -1297 -2656
rect -1293 -2660 -923 -2656
rect -919 -2660 -565 -2656
rect -561 -2660 -207 -2656
rect -203 -2660 151 -2656
rect 155 -2660 507 -2656
rect 511 -2660 865 -2656
rect 869 -2660 1223 -2656
rect 1227 -2660 1589 -2656
rect -975 -2673 -909 -2669
rect -612 -2673 -551 -2669
rect -259 -2673 -193 -2669
rect 101 -2673 165 -2669
rect 455 -2673 521 -2669
rect 814 -2673 879 -2669
rect 1171 -2673 1237 -2669
rect 1804 -2708 1831 -2607
rect -1411 -2712 -1292 -2708
rect -1288 -2712 -918 -2708
rect -914 -2712 -560 -2708
rect -556 -2712 -202 -2708
rect -198 -2712 156 -2708
rect 160 -2712 512 -2708
rect 516 -2712 870 -2708
rect 874 -2712 1228 -2708
rect 1232 -2712 1831 -2708
rect -2054 -2779 -1225 -2775
rect -1221 -2779 -1208 -2775
rect -1204 -2779 -1168 -2775
rect -1164 -2779 -1147 -2775
rect -1143 -2779 -926 -2775
rect -922 -2779 -900 -2775
rect -896 -2779 -883 -2775
rect -879 -2779 -843 -2775
rect -839 -2779 -822 -2775
rect -818 -2779 -805 -2775
rect -801 -2779 -765 -2775
rect -761 -2779 -741 -2775
rect -737 -2779 -704 -2775
rect -700 -2779 -568 -2775
rect -564 -2779 -542 -2775
rect -538 -2779 -525 -2775
rect -521 -2779 -485 -2775
rect -481 -2779 -464 -2775
rect -460 -2779 -447 -2775
rect -443 -2779 -407 -2775
rect -403 -2779 -383 -2775
rect -379 -2779 -346 -2775
rect -342 -2779 -210 -2775
rect -206 -2779 -184 -2775
rect -180 -2779 -167 -2775
rect -163 -2779 -127 -2775
rect -123 -2779 -106 -2775
rect -102 -2779 -89 -2775
rect -85 -2779 -49 -2775
rect -45 -2779 -25 -2775
rect -21 -2779 12 -2775
rect 16 -2779 148 -2775
rect 152 -2779 174 -2775
rect 178 -2779 191 -2775
rect 195 -2779 231 -2775
rect 235 -2779 252 -2775
rect 256 -2779 269 -2775
rect 273 -2779 309 -2775
rect 313 -2779 333 -2775
rect 337 -2779 370 -2775
rect 374 -2779 504 -2775
rect 508 -2779 530 -2775
rect 534 -2779 547 -2775
rect 551 -2779 587 -2775
rect 591 -2779 608 -2775
rect 612 -2779 625 -2775
rect 629 -2779 665 -2775
rect 669 -2779 689 -2775
rect 693 -2779 726 -2775
rect 730 -2779 862 -2775
rect 866 -2779 888 -2775
rect 892 -2779 905 -2775
rect 909 -2779 945 -2775
rect 949 -2779 966 -2775
rect 970 -2779 983 -2775
rect 987 -2779 1023 -2775
rect 1027 -2779 1047 -2775
rect 1051 -2779 1084 -2775
rect 1088 -2779 1220 -2775
rect 1224 -2779 1246 -2775
rect 1250 -2779 1263 -2775
rect 1267 -2779 1303 -2775
rect 1307 -2779 1324 -2775
rect 1328 -2779 1341 -2775
rect 1345 -2779 1381 -2775
rect 1385 -2779 1405 -2775
rect 1409 -2779 1442 -2775
rect 1446 -2779 1589 -2775
rect -2054 -2894 -2027 -2779
rect -926 -2783 -922 -2779
rect -900 -2783 -896 -2779
rect -883 -2783 -879 -2779
rect -843 -2783 -839 -2779
rect -822 -2783 -818 -2779
rect -805 -2783 -801 -2779
rect -765 -2783 -761 -2779
rect -741 -2783 -737 -2779
rect -704 -2783 -700 -2779
rect -568 -2783 -564 -2779
rect -542 -2783 -538 -2779
rect -525 -2783 -521 -2779
rect -485 -2783 -481 -2779
rect -464 -2783 -460 -2779
rect -447 -2783 -443 -2779
rect -407 -2783 -403 -2779
rect -383 -2783 -379 -2779
rect -346 -2783 -342 -2779
rect -210 -2783 -206 -2779
rect -184 -2783 -180 -2779
rect -167 -2783 -163 -2779
rect -127 -2783 -123 -2779
rect -106 -2783 -102 -2779
rect -89 -2783 -85 -2779
rect -49 -2783 -45 -2779
rect -25 -2783 -21 -2779
rect 12 -2783 16 -2779
rect 148 -2783 152 -2779
rect 174 -2783 178 -2779
rect 191 -2783 195 -2779
rect 231 -2783 235 -2779
rect 252 -2783 256 -2779
rect 269 -2783 273 -2779
rect 309 -2783 313 -2779
rect 333 -2783 337 -2779
rect 370 -2783 374 -2779
rect 504 -2783 508 -2779
rect 530 -2783 534 -2779
rect 547 -2783 551 -2779
rect 587 -2783 591 -2779
rect 608 -2783 612 -2779
rect 625 -2783 629 -2779
rect 665 -2783 669 -2779
rect 689 -2783 693 -2779
rect 726 -2783 730 -2779
rect 862 -2783 866 -2779
rect 888 -2783 892 -2779
rect 905 -2783 909 -2779
rect 945 -2783 949 -2779
rect 966 -2783 970 -2779
rect 983 -2783 987 -2779
rect 1023 -2783 1027 -2779
rect 1047 -2783 1051 -2779
rect 1084 -2783 1088 -2779
rect 1220 -2783 1224 -2779
rect 1246 -2783 1250 -2779
rect 1263 -2783 1267 -2779
rect 1303 -2783 1307 -2779
rect 1324 -2783 1328 -2779
rect 1341 -2783 1345 -2779
rect 1381 -2783 1385 -2779
rect 1405 -2783 1409 -2779
rect 1442 -2783 1446 -2779
rect -920 -2798 -858 -2794
rect -854 -2798 -824 -2794
rect -776 -2798 -746 -2794
rect -562 -2798 -500 -2794
rect -496 -2798 -466 -2794
rect -418 -2798 -388 -2794
rect -204 -2798 -142 -2794
rect -138 -2798 -108 -2794
rect -60 -2798 -30 -2794
rect 154 -2798 216 -2794
rect 220 -2798 250 -2794
rect 298 -2798 328 -2794
rect 510 -2798 572 -2794
rect 576 -2798 606 -2794
rect 654 -2798 684 -2794
rect 868 -2798 930 -2794
rect 934 -2798 964 -2794
rect 1012 -2798 1042 -2794
rect 1226 -2798 1288 -2794
rect 1292 -2798 1322 -2794
rect 1370 -2798 1400 -2794
rect -913 -2805 -882 -2801
rect -555 -2805 -524 -2801
rect -197 -2805 -166 -2801
rect 161 -2805 192 -2801
rect 517 -2805 548 -2801
rect 875 -2805 906 -2801
rect 1233 -2805 1264 -2801
rect -931 -2812 -848 -2808
rect -809 -2812 -706 -2808
rect -573 -2812 -490 -2808
rect -451 -2812 -348 -2808
rect -215 -2812 -132 -2808
rect -93 -2812 10 -2808
rect 143 -2812 226 -2808
rect 265 -2812 368 -2808
rect 499 -2812 582 -2808
rect 621 -2812 724 -2808
rect 857 -2812 940 -2808
rect 979 -2812 1082 -2808
rect 1215 -2812 1298 -2808
rect 1337 -2812 1440 -2808
rect -975 -2819 -928 -2815
rect -894 -2819 -865 -2815
rect -861 -2819 -780 -2815
rect -691 -2819 -612 -2815
rect -599 -2819 -570 -2815
rect -536 -2819 -507 -2815
rect -503 -2819 -422 -2815
rect -333 -2818 -259 -2814
rect -616 -2823 -612 -2819
rect -263 -2823 -259 -2818
rect -245 -2819 -212 -2815
rect -178 -2819 -149 -2815
rect -145 -2819 -64 -2815
rect 25 -2819 101 -2815
rect 115 -2819 146 -2815
rect 180 -2819 209 -2815
rect 213 -2819 294 -2815
rect 383 -2819 455 -2815
rect 469 -2819 502 -2815
rect 536 -2819 565 -2815
rect 569 -2819 650 -2815
rect 739 -2819 814 -2815
rect 828 -2819 860 -2815
rect 894 -2819 923 -2815
rect 927 -2819 1008 -2815
rect 1097 -2817 1164 -2813
rect 97 -2823 101 -2819
rect 451 -2823 455 -2819
rect 810 -2823 814 -2819
rect 1160 -2823 1164 -2817
rect 1171 -2819 1218 -2815
rect 1252 -2819 1281 -2815
rect 1285 -2819 1366 -2815
rect -1230 -2828 -1173 -2824
rect -1134 -2827 -902 -2823
rect -887 -2827 -804 -2823
rect -783 -2827 -688 -2823
rect -616 -2827 -544 -2823
rect -529 -2827 -446 -2823
rect -425 -2827 -329 -2823
rect -263 -2827 -186 -2823
rect -171 -2827 -88 -2823
rect -67 -2827 28 -2823
rect 97 -2827 172 -2823
rect 187 -2827 270 -2823
rect 291 -2827 389 -2823
rect 451 -2827 528 -2823
rect 543 -2827 626 -2823
rect 647 -2827 742 -2823
rect 810 -2827 886 -2823
rect 901 -2827 984 -2823
rect 1005 -2827 1103 -2823
rect 1160 -2827 1244 -2823
rect 1259 -2827 1342 -2823
rect 1363 -2827 1467 -2823
rect -1253 -2835 -1223 -2831
rect -1219 -2835 -1183 -2831
rect -1179 -2835 -1163 -2831
rect -959 -2834 -924 -2830
rect -905 -2834 -776 -2830
rect -612 -2834 -566 -2830
rect -547 -2834 -418 -2830
rect -259 -2834 -208 -2830
rect -189 -2834 -60 -2830
rect 101 -2834 150 -2830
rect 169 -2834 298 -2830
rect 455 -2834 506 -2830
rect 525 -2834 654 -2830
rect 814 -2834 864 -2830
rect 883 -2834 1012 -2830
rect 1188 -2834 1222 -2830
rect 1241 -2834 1370 -2830
rect -1279 -2842 -1227 -2838
rect -1223 -2842 -1197 -2838
rect -1193 -2842 -1149 -2838
rect -898 -2841 -794 -2837
rect -790 -2841 -760 -2837
rect -540 -2841 -436 -2837
rect -432 -2841 -402 -2837
rect -182 -2841 -78 -2837
rect -74 -2841 -44 -2837
rect 176 -2841 280 -2837
rect 284 -2841 314 -2837
rect 532 -2841 636 -2837
rect 640 -2841 670 -2837
rect 890 -2841 994 -2837
rect 998 -2841 1028 -2837
rect 1248 -2841 1352 -2837
rect 1356 -2841 1386 -2837
rect -1186 -2849 -1117 -2845
rect -924 -2848 -872 -2844
rect -868 -2848 -838 -2844
rect -566 -2848 -514 -2844
rect -510 -2848 -480 -2844
rect -208 -2848 -156 -2844
rect -152 -2848 -122 -2844
rect 150 -2848 202 -2844
rect 206 -2848 236 -2844
rect 506 -2848 558 -2844
rect 562 -2848 592 -2844
rect 864 -2848 916 -2844
rect 920 -2848 950 -2844
rect 1222 -2848 1274 -2844
rect 1278 -2848 1308 -2844
rect -1204 -2856 -1172 -2852
rect -879 -2856 -847 -2852
rect -883 -2859 -879 -2856
rect -847 -2859 -843 -2856
rect -801 -2856 -769 -2852
rect -805 -2859 -801 -2856
rect -769 -2859 -765 -2856
rect -521 -2856 -489 -2852
rect -525 -2859 -521 -2856
rect -489 -2859 -485 -2856
rect -443 -2856 -411 -2852
rect -447 -2859 -443 -2856
rect -411 -2859 -407 -2856
rect -163 -2856 -131 -2852
rect -167 -2859 -163 -2856
rect -131 -2859 -127 -2856
rect -85 -2856 -53 -2852
rect -89 -2859 -85 -2856
rect -53 -2859 -49 -2856
rect 195 -2856 227 -2852
rect 191 -2859 195 -2856
rect 227 -2859 231 -2856
rect 273 -2856 305 -2852
rect 269 -2859 273 -2856
rect 305 -2859 309 -2856
rect 551 -2856 583 -2852
rect 547 -2859 551 -2856
rect 583 -2859 587 -2856
rect 629 -2856 661 -2852
rect 625 -2859 629 -2856
rect 661 -2859 665 -2856
rect 909 -2856 941 -2852
rect 905 -2859 909 -2856
rect 941 -2859 945 -2856
rect 987 -2856 1019 -2852
rect 983 -2859 987 -2856
rect 1019 -2859 1023 -2856
rect 1267 -2856 1299 -2852
rect 1263 -2859 1267 -2856
rect 1299 -2859 1303 -2856
rect 1345 -2856 1377 -2852
rect 1341 -2859 1345 -2856
rect 1377 -2859 1381 -2856
rect -926 -2867 -922 -2863
rect -900 -2867 -896 -2863
rect -857 -2867 -853 -2863
rect -822 -2867 -818 -2863
rect -778 -2867 -774 -2863
rect -761 -2867 -757 -2863
rect -725 -2867 -721 -2863
rect -704 -2867 -700 -2863
rect -568 -2867 -564 -2863
rect -542 -2867 -538 -2863
rect -499 -2867 -495 -2863
rect -464 -2867 -460 -2863
rect -420 -2867 -416 -2863
rect -403 -2867 -399 -2863
rect -367 -2867 -363 -2863
rect -346 -2867 -342 -2863
rect -210 -2867 -206 -2863
rect -184 -2867 -180 -2863
rect -141 -2867 -137 -2863
rect -106 -2867 -102 -2863
rect -62 -2867 -58 -2863
rect -45 -2867 -41 -2863
rect -9 -2867 -5 -2863
rect 12 -2867 16 -2863
rect 148 -2867 152 -2863
rect 174 -2867 178 -2863
rect 217 -2867 221 -2863
rect 252 -2867 256 -2863
rect 296 -2867 300 -2863
rect 313 -2867 317 -2863
rect 349 -2867 353 -2863
rect 370 -2867 374 -2863
rect 504 -2867 508 -2863
rect 530 -2867 534 -2863
rect 573 -2867 577 -2863
rect 608 -2867 612 -2863
rect 652 -2867 656 -2863
rect 669 -2867 673 -2863
rect 705 -2867 709 -2863
rect 726 -2867 730 -2863
rect 862 -2867 866 -2863
rect 888 -2867 892 -2863
rect 931 -2867 935 -2863
rect 966 -2867 970 -2863
rect 1010 -2867 1014 -2863
rect 1027 -2867 1031 -2863
rect 1063 -2867 1067 -2863
rect 1084 -2867 1088 -2863
rect 1220 -2867 1224 -2863
rect 1246 -2867 1250 -2863
rect 1289 -2867 1293 -2863
rect 1324 -2867 1328 -2863
rect 1368 -2867 1372 -2863
rect 1385 -2867 1389 -2863
rect 1421 -2867 1425 -2863
rect 1442 -2867 1446 -2863
rect 1804 -2867 1831 -2712
rect -1411 -2871 -1225 -2867
rect -1221 -2871 -1181 -2867
rect -1177 -2871 -1147 -2867
rect -1143 -2871 -926 -2867
rect -922 -2871 -900 -2867
rect -896 -2871 -857 -2867
rect -853 -2871 -822 -2867
rect -818 -2871 -778 -2867
rect -774 -2871 -761 -2867
rect -757 -2871 -725 -2867
rect -721 -2871 -704 -2867
rect -700 -2871 -568 -2867
rect -564 -2871 -542 -2867
rect -538 -2871 -499 -2867
rect -495 -2871 -464 -2867
rect -460 -2871 -420 -2867
rect -416 -2871 -403 -2867
rect -399 -2871 -367 -2867
rect -363 -2871 -346 -2867
rect -342 -2871 -210 -2867
rect -206 -2871 -184 -2867
rect -180 -2871 -141 -2867
rect -137 -2871 -106 -2867
rect -102 -2871 -62 -2867
rect -58 -2871 -45 -2867
rect -41 -2871 -9 -2867
rect -5 -2871 12 -2867
rect 16 -2871 148 -2867
rect 152 -2871 174 -2867
rect 178 -2871 217 -2867
rect 221 -2871 252 -2867
rect 256 -2871 296 -2867
rect 300 -2871 313 -2867
rect 317 -2871 349 -2867
rect 353 -2871 370 -2867
rect 374 -2871 504 -2867
rect 508 -2871 530 -2867
rect 534 -2871 573 -2867
rect 577 -2871 608 -2867
rect 612 -2871 652 -2867
rect 656 -2871 669 -2867
rect 673 -2871 705 -2867
rect 709 -2871 726 -2867
rect 730 -2871 862 -2867
rect 866 -2871 888 -2867
rect 892 -2871 931 -2867
rect 935 -2871 966 -2867
rect 970 -2871 1010 -2867
rect 1014 -2871 1027 -2867
rect 1031 -2871 1063 -2867
rect 1067 -2871 1084 -2867
rect 1088 -2871 1220 -2867
rect 1224 -2871 1246 -2867
rect 1250 -2871 1289 -2867
rect 1293 -2871 1324 -2867
rect 1328 -2871 1368 -2867
rect 1372 -2871 1385 -2867
rect 1389 -2871 1421 -2867
rect 1425 -2871 1442 -2867
rect 1446 -2871 1831 -2867
rect -1253 -2878 -688 -2874
rect -599 -2878 28 -2874
rect 115 -2878 742 -2874
rect 827 -2878 1467 -2874
rect -1242 -2886 -1117 -2882
rect -959 -2885 -329 -2881
rect -245 -2885 389 -2881
rect 469 -2885 1103 -2881
rect 1188 -2885 1451 -2881
rect -2054 -2898 -1550 -2894
rect -1546 -2898 -1533 -2894
rect -1529 -2898 -1513 -2894
rect -1509 -2898 -1492 -2894
rect -1488 -2898 -1471 -2894
rect -1467 -2898 -1450 -2894
rect -1446 -2898 -1429 -2894
rect -1425 -2898 -1408 -2894
rect -1404 -2898 -1387 -2894
rect -1383 -2898 -1367 -2894
rect -1363 -2898 -1225 -2894
rect -1221 -2898 -1208 -2894
rect -1204 -2898 -1188 -2894
rect -1184 -2898 -1167 -2894
rect -1163 -2898 -1146 -2894
rect -1142 -2898 -1125 -2894
rect -1121 -2898 -1104 -2894
rect -1100 -2898 -1083 -2894
rect -1079 -2898 -1062 -2894
rect -1058 -2898 -1042 -2894
rect -1038 -2898 -926 -2894
rect -922 -2898 -909 -2894
rect -905 -2898 -889 -2894
rect -885 -2898 -868 -2894
rect -864 -2898 -847 -2894
rect -843 -2898 -826 -2894
rect -822 -2898 -805 -2894
rect -801 -2898 -784 -2894
rect -780 -2898 -763 -2894
rect -759 -2898 -743 -2894
rect -739 -2898 -568 -2894
rect -564 -2898 -551 -2894
rect -547 -2898 -531 -2894
rect -527 -2898 -510 -2894
rect -506 -2898 -489 -2894
rect -485 -2898 -468 -2894
rect -464 -2898 -447 -2894
rect -443 -2898 -426 -2894
rect -422 -2898 -405 -2894
rect -401 -2898 -385 -2894
rect -381 -2898 -210 -2894
rect -206 -2898 -193 -2894
rect -189 -2898 -173 -2894
rect -169 -2898 -152 -2894
rect -148 -2898 -131 -2894
rect -127 -2898 -110 -2894
rect -106 -2898 -89 -2894
rect -85 -2898 -68 -2894
rect -64 -2898 -47 -2894
rect -43 -2898 -27 -2894
rect -23 -2898 148 -2894
rect 152 -2898 165 -2894
rect 169 -2898 185 -2894
rect 189 -2898 206 -2894
rect 210 -2898 227 -2894
rect 231 -2898 248 -2894
rect 252 -2898 269 -2894
rect 273 -2898 290 -2894
rect 294 -2898 311 -2894
rect 315 -2898 331 -2894
rect 335 -2898 1604 -2894
rect -2054 -3065 -2027 -2898
rect -1528 -2946 -1494 -2942
rect -1430 -2946 -1410 -2942
rect -1395 -2946 -1352 -2942
rect -1203 -2946 -1169 -2942
rect -1105 -2946 -1085 -2942
rect -1070 -2946 -931 -2942
rect -904 -2946 -870 -2942
rect -806 -2946 -786 -2942
rect -771 -2946 -573 -2942
rect -546 -2946 -512 -2942
rect -448 -2946 -428 -2942
rect -413 -2946 -215 -2942
rect -188 -2946 -154 -2942
rect -90 -2946 -70 -2942
rect -55 -2946 143 -2942
rect 170 -2946 204 -2942
rect 268 -2946 288 -2942
rect 303 -2946 339 -2942
rect -935 -2950 -931 -2946
rect -577 -2950 -573 -2946
rect -219 -2950 -215 -2946
rect 139 -2950 143 -2946
rect -1563 -2954 -1552 -2950
rect -1548 -2954 -1518 -2950
rect -1497 -2954 -1466 -2950
rect -1437 -2954 -1406 -2950
rect -1395 -2954 -1368 -2950
rect -1242 -2954 -1227 -2950
rect -1223 -2954 -1193 -2950
rect -1172 -2954 -1141 -2950
rect -1112 -2954 -1081 -2950
rect -1070 -2954 -1043 -2950
rect -935 -2954 -928 -2950
rect -924 -2954 -894 -2950
rect -873 -2954 -842 -2950
rect -813 -2954 -782 -2950
rect -771 -2954 -744 -2950
rect -577 -2954 -570 -2950
rect -566 -2954 -536 -2950
rect -515 -2954 -484 -2950
rect -455 -2954 -424 -2950
rect -413 -2954 -386 -2950
rect -219 -2954 -212 -2950
rect -208 -2954 -178 -2950
rect -157 -2954 -126 -2950
rect -97 -2954 -66 -2950
rect -55 -2954 -28 -2950
rect 139 -2954 146 -2950
rect 150 -2954 180 -2950
rect 201 -2954 232 -2950
rect 261 -2954 292 -2950
rect 303 -2954 330 -2950
rect -1555 -2961 -1508 -2957
rect -1472 -2961 -1459 -2957
rect -1455 -2961 -1424 -2957
rect -1388 -2961 -1375 -2957
rect -1371 -2961 -1359 -2957
rect -1230 -2961 -1183 -2957
rect -1147 -2961 -1134 -2957
rect -1130 -2961 -1099 -2957
rect -1063 -2961 -1050 -2957
rect -1046 -2961 -1034 -2957
rect -931 -2961 -884 -2957
rect -848 -2961 -835 -2957
rect -831 -2961 -800 -2957
rect -764 -2961 -751 -2957
rect -747 -2961 -735 -2957
rect -573 -2961 -526 -2957
rect -490 -2961 -477 -2957
rect -473 -2961 -442 -2957
rect -406 -2961 -393 -2957
rect -389 -2961 -377 -2957
rect -215 -2961 -168 -2957
rect -132 -2961 -119 -2957
rect -115 -2961 -84 -2957
rect -48 -2961 -35 -2957
rect -31 -2961 -19 -2957
rect 143 -2961 190 -2957
rect 226 -2961 239 -2957
rect 243 -2961 274 -2957
rect 310 -2961 323 -2957
rect 327 -2961 339 -2957
rect -1563 -2968 -1548 -2964
rect -1544 -2968 -1434 -2964
rect -1413 -2968 -1382 -2964
rect -1238 -2968 -1223 -2964
rect -1219 -2968 -1109 -2964
rect -1088 -2968 -1057 -2964
rect -939 -2968 -924 -2964
rect -920 -2968 -810 -2964
rect -789 -2968 -758 -2964
rect -581 -2968 -566 -2964
rect -562 -2968 -452 -2964
rect -431 -2968 -400 -2964
rect -223 -2968 -208 -2964
rect -204 -2968 -94 -2964
rect -73 -2968 -42 -2964
rect 135 -2968 150 -2964
rect 154 -2968 264 -2964
rect 285 -2968 316 -2964
rect -1513 -2975 -1490 -2971
rect -1471 -2975 -1452 -2971
rect -1188 -2975 -1165 -2971
rect -1146 -2975 -1127 -2971
rect -889 -2975 -866 -2971
rect -847 -2975 -828 -2971
rect -531 -2975 -508 -2971
rect -489 -2975 -470 -2971
rect -173 -2975 -150 -2971
rect -131 -2975 -112 -2971
rect 185 -2975 208 -2971
rect 227 -2975 246 -2971
rect 1804 -2986 1831 -2871
rect -1735 -2990 -1550 -2986
rect -1546 -2990 -1533 -2986
rect -1529 -2990 -1492 -2986
rect -1488 -2990 -1450 -2986
rect -1446 -2990 -1408 -2986
rect -1404 -2990 -1367 -2986
rect -1363 -2990 -1225 -2986
rect -1221 -2990 -1208 -2986
rect -1204 -2990 -1167 -2986
rect -1163 -2990 -1125 -2986
rect -1121 -2990 -1083 -2986
rect -1079 -2990 -1042 -2986
rect -1038 -2990 -926 -2986
rect -922 -2990 -909 -2986
rect -905 -2990 -868 -2986
rect -864 -2990 -826 -2986
rect -822 -2990 -784 -2986
rect -780 -2990 -743 -2986
rect -739 -2990 -568 -2986
rect -564 -2990 -551 -2986
rect -547 -2990 -510 -2986
rect -506 -2990 -468 -2986
rect -464 -2990 -426 -2986
rect -422 -2990 -385 -2986
rect -381 -2990 -210 -2986
rect -206 -2990 -193 -2986
rect -189 -2990 -152 -2986
rect -148 -2990 -110 -2986
rect -106 -2990 -68 -2986
rect -64 -2990 -27 -2986
rect -23 -2990 148 -2986
rect 152 -2990 165 -2986
rect 169 -2990 206 -2986
rect 210 -2990 248 -2986
rect 252 -2990 290 -2986
rect 294 -2990 331 -2986
rect 335 -2990 1831 -2986
rect -1577 -2997 -1352 -2993
rect -2054 -3069 -1550 -3065
rect -1546 -3069 -1533 -3065
rect -1529 -3069 -1513 -3065
rect -1509 -3069 -1492 -3065
rect -1488 -3069 -1471 -3065
rect -1467 -3069 -1450 -3065
rect -1446 -3069 -1429 -3065
rect -1425 -3069 -1408 -3065
rect -1404 -3069 -1387 -3065
rect -1383 -3069 -1367 -3065
rect -1363 -3069 -1225 -3065
rect -1221 -3069 -1208 -3065
rect -1204 -3069 -1188 -3065
rect -1184 -3069 -1167 -3065
rect -1163 -3069 -1146 -3065
rect -1142 -3069 -1125 -3065
rect -1121 -3069 -1104 -3065
rect -1100 -3069 -1083 -3065
rect -1079 -3069 -1062 -3065
rect -1058 -3069 -1042 -3065
rect -1038 -3069 -926 -3065
rect -922 -3069 -909 -3065
rect -905 -3069 -889 -3065
rect -885 -3069 -868 -3065
rect -864 -3069 -847 -3065
rect -843 -3069 -826 -3065
rect -822 -3069 -805 -3065
rect -801 -3069 -784 -3065
rect -780 -3069 -763 -3065
rect -759 -3069 -743 -3065
rect -739 -3069 -568 -3065
rect -564 -3069 -551 -3065
rect -547 -3069 -531 -3065
rect -527 -3069 -510 -3065
rect -506 -3069 -489 -3065
rect -485 -3069 -468 -3065
rect -464 -3069 -447 -3065
rect -443 -3069 -426 -3065
rect -422 -3069 -405 -3065
rect -401 -3069 -385 -3065
rect -381 -3069 -210 -3065
rect -206 -3069 -193 -3065
rect -189 -3069 -173 -3065
rect -169 -3069 -152 -3065
rect -148 -3069 -131 -3065
rect -127 -3069 -110 -3065
rect -106 -3069 -89 -3065
rect -85 -3069 -68 -3065
rect -64 -3069 -47 -3065
rect -43 -3069 -27 -3065
rect -23 -3069 148 -3065
rect 152 -3069 165 -3065
rect 169 -3069 185 -3065
rect 189 -3069 206 -3065
rect 210 -3069 227 -3065
rect 231 -3069 248 -3065
rect 252 -3069 269 -3065
rect 273 -3069 290 -3065
rect 294 -3069 311 -3065
rect 315 -3069 331 -3065
rect 335 -3069 504 -3065
rect 508 -3069 521 -3065
rect 525 -3069 541 -3065
rect 545 -3069 562 -3065
rect 566 -3069 583 -3065
rect 587 -3069 604 -3065
rect 608 -3069 625 -3065
rect 629 -3069 646 -3065
rect 650 -3069 667 -3065
rect 671 -3069 687 -3065
rect 691 -3069 862 -3065
rect 866 -3069 879 -3065
rect 883 -3069 899 -3065
rect 903 -3069 920 -3065
rect 924 -3069 941 -3065
rect 945 -3069 962 -3065
rect 966 -3069 983 -3065
rect 987 -3069 1004 -3065
rect 1008 -3069 1025 -3065
rect 1029 -3069 1045 -3065
rect 1049 -3069 1220 -3065
rect 1224 -3069 1237 -3065
rect 1241 -3069 1257 -3065
rect 1261 -3069 1278 -3065
rect 1282 -3069 1299 -3065
rect 1303 -3069 1320 -3065
rect 1324 -3069 1341 -3065
rect 1345 -3069 1362 -3065
rect 1366 -3069 1383 -3065
rect 1387 -3069 1403 -3065
rect 1407 -3069 1618 -3065
rect -2054 -3236 -2027 -3069
rect -1528 -3117 -1494 -3113
rect -1430 -3117 -1410 -3113
rect -1395 -3117 -1355 -3113
rect -1203 -3117 -1169 -3113
rect -1105 -3117 -1085 -3113
rect -1070 -3117 -1026 -3113
rect -904 -3117 -870 -3113
rect -806 -3117 -786 -3113
rect -771 -3117 -725 -3113
rect -546 -3117 -512 -3113
rect -448 -3117 -428 -3113
rect -413 -3117 -367 -3113
rect -188 -3117 -154 -3113
rect -90 -3117 -70 -3113
rect -55 -3117 -13 -3113
rect 170 -3117 204 -3113
rect 268 -3117 288 -3113
rect 303 -3117 345 -3113
rect 526 -3117 560 -3113
rect 624 -3117 644 -3113
rect 659 -3117 701 -3113
rect 884 -3117 918 -3113
rect 982 -3117 1002 -3113
rect 1017 -3117 1060 -3113
rect 1242 -3117 1276 -3113
rect 1340 -3117 1360 -3113
rect 1375 -3117 1419 -3113
rect -1577 -3125 -1552 -3121
rect -1548 -3125 -1518 -3121
rect -1497 -3125 -1466 -3121
rect -1437 -3125 -1406 -3121
rect -1395 -3125 -1368 -3121
rect -1253 -3125 -1227 -3121
rect -1223 -3125 -1193 -3121
rect -1172 -3125 -1141 -3121
rect -1112 -3125 -1081 -3121
rect -1070 -3125 -1043 -3121
rect -959 -3125 -928 -3121
rect -924 -3125 -894 -3121
rect -873 -3125 -842 -3121
rect -813 -3125 -782 -3121
rect -771 -3125 -744 -3121
rect -599 -3125 -570 -3121
rect -566 -3125 -536 -3121
rect -515 -3125 -484 -3121
rect -455 -3125 -424 -3121
rect -413 -3125 -386 -3121
rect -245 -3125 -212 -3121
rect -208 -3125 -178 -3121
rect -157 -3125 -126 -3121
rect -97 -3125 -66 -3121
rect -55 -3125 -28 -3121
rect 115 -3125 146 -3121
rect 150 -3125 180 -3121
rect 201 -3125 232 -3121
rect 261 -3125 292 -3121
rect 303 -3125 330 -3121
rect 469 -3125 502 -3121
rect 506 -3125 536 -3121
rect 557 -3125 588 -3121
rect 617 -3125 648 -3121
rect 659 -3125 686 -3121
rect 827 -3125 860 -3121
rect 864 -3125 894 -3121
rect 915 -3125 946 -3121
rect 975 -3125 1006 -3121
rect 1017 -3125 1044 -3121
rect 1188 -3125 1218 -3121
rect 1222 -3125 1252 -3121
rect 1273 -3125 1304 -3121
rect 1333 -3125 1364 -3121
rect 1375 -3125 1402 -3121
rect -1555 -3132 -1508 -3128
rect -1472 -3132 -1459 -3128
rect -1455 -3132 -1424 -3128
rect -1388 -3132 -1375 -3128
rect -1371 -3132 -1359 -3128
rect -1230 -3132 -1183 -3128
rect -1147 -3132 -1134 -3128
rect -1130 -3132 -1099 -3128
rect -1063 -3132 -1050 -3128
rect -1046 -3132 -1034 -3128
rect -931 -3132 -884 -3128
rect -848 -3132 -835 -3128
rect -831 -3132 -800 -3128
rect -764 -3132 -751 -3128
rect -747 -3132 -735 -3128
rect -573 -3132 -526 -3128
rect -490 -3132 -477 -3128
rect -473 -3132 -442 -3128
rect -406 -3132 -393 -3128
rect -389 -3132 -377 -3128
rect -215 -3132 -168 -3128
rect -132 -3132 -119 -3128
rect -115 -3132 -84 -3128
rect -48 -3132 -35 -3128
rect -31 -3132 -19 -3128
rect 143 -3132 190 -3128
rect 226 -3132 239 -3128
rect 243 -3132 274 -3128
rect 310 -3132 323 -3128
rect 327 -3132 339 -3128
rect 499 -3132 546 -3128
rect 582 -3132 595 -3128
rect 599 -3132 630 -3128
rect 666 -3132 679 -3128
rect 683 -3132 695 -3128
rect 857 -3132 904 -3128
rect 940 -3132 953 -3128
rect 957 -3132 988 -3128
rect 1024 -3132 1037 -3128
rect 1041 -3132 1053 -3128
rect 1215 -3132 1262 -3128
rect 1298 -3132 1311 -3128
rect 1315 -3132 1346 -3128
rect 1382 -3132 1395 -3128
rect 1399 -3132 1411 -3128
rect -1563 -3139 -1548 -3135
rect -1544 -3139 -1434 -3135
rect -1413 -3139 -1382 -3135
rect -1238 -3139 -1223 -3135
rect -1219 -3139 -1109 -3135
rect -1088 -3139 -1057 -3135
rect -939 -3139 -924 -3135
rect -920 -3139 -810 -3135
rect -789 -3139 -758 -3135
rect -581 -3139 -566 -3135
rect -562 -3139 -452 -3135
rect -431 -3139 -400 -3135
rect -223 -3139 -208 -3135
rect -204 -3139 -94 -3135
rect -73 -3139 -42 -3135
rect 135 -3139 150 -3135
rect 154 -3139 264 -3135
rect 285 -3139 316 -3135
rect 491 -3139 506 -3135
rect 510 -3139 620 -3135
rect 641 -3139 672 -3135
rect 849 -3139 864 -3135
rect 868 -3139 978 -3135
rect 999 -3139 1030 -3135
rect 1207 -3139 1222 -3135
rect 1226 -3139 1336 -3135
rect 1357 -3139 1388 -3135
rect -1513 -3146 -1490 -3142
rect -1471 -3146 -1452 -3142
rect -1188 -3146 -1165 -3142
rect -1146 -3146 -1127 -3142
rect -889 -3146 -866 -3142
rect -847 -3146 -828 -3142
rect -531 -3146 -508 -3142
rect -489 -3146 -470 -3142
rect -173 -3146 -150 -3142
rect -131 -3146 -112 -3142
rect 185 -3146 208 -3142
rect 227 -3146 246 -3142
rect 541 -3146 564 -3142
rect 583 -3146 602 -3142
rect 899 -3146 922 -3142
rect 941 -3146 960 -3142
rect 1257 -3146 1280 -3142
rect 1299 -3146 1318 -3142
rect 1804 -3157 1831 -2990
rect -1765 -3161 -1550 -3157
rect -1546 -3161 -1533 -3157
rect -1529 -3161 -1492 -3157
rect -1488 -3161 -1450 -3157
rect -1446 -3161 -1408 -3157
rect -1404 -3161 -1367 -3157
rect -1363 -3161 -1225 -3157
rect -1221 -3161 -1208 -3157
rect -1204 -3161 -1167 -3157
rect -1163 -3161 -1125 -3157
rect -1121 -3161 -1083 -3157
rect -1079 -3161 -1042 -3157
rect -1038 -3161 -926 -3157
rect -922 -3161 -909 -3157
rect -905 -3161 -868 -3157
rect -864 -3161 -826 -3157
rect -822 -3161 -784 -3157
rect -780 -3161 -743 -3157
rect -739 -3161 -568 -3157
rect -564 -3161 -551 -3157
rect -547 -3161 -510 -3157
rect -506 -3161 -468 -3157
rect -464 -3161 -426 -3157
rect -422 -3161 -385 -3157
rect -381 -3161 -210 -3157
rect -206 -3161 -193 -3157
rect -189 -3161 -152 -3157
rect -148 -3161 -110 -3157
rect -106 -3161 -68 -3157
rect -64 -3161 -27 -3157
rect -23 -3161 148 -3157
rect 152 -3161 165 -3157
rect 169 -3161 206 -3157
rect 210 -3161 248 -3157
rect 252 -3161 290 -3157
rect 294 -3161 331 -3157
rect 335 -3161 504 -3157
rect 508 -3161 521 -3157
rect 525 -3161 562 -3157
rect 566 -3161 604 -3157
rect 608 -3161 646 -3157
rect 650 -3161 687 -3157
rect 691 -3161 862 -3157
rect 866 -3161 879 -3157
rect 883 -3161 920 -3157
rect 924 -3161 962 -3157
rect 966 -3161 1004 -3157
rect 1008 -3161 1045 -3157
rect 1049 -3161 1220 -3157
rect 1224 -3161 1237 -3157
rect 1241 -3161 1278 -3157
rect 1282 -3161 1320 -3157
rect 1324 -3161 1362 -3157
rect 1366 -3161 1403 -3157
rect 1407 -3161 1831 -3157
rect -1578 -3168 -1355 -3164
rect -1253 -3169 -1026 -3165
rect -959 -3169 -725 -3165
rect -599 -3168 -367 -3164
rect -245 -3169 -13 -3165
rect 115 -3168 345 -3164
rect 469 -3168 701 -3164
rect 827 -3168 1060 -3164
rect 1188 -3169 1419 -3165
rect -2054 -3240 -1550 -3236
rect -1546 -3240 -1533 -3236
rect -1529 -3240 -1513 -3236
rect -1509 -3240 -1492 -3236
rect -1488 -3240 -1471 -3236
rect -1467 -3240 -1450 -3236
rect -1446 -3240 -1429 -3236
rect -1425 -3240 -1408 -3236
rect -1404 -3240 -1387 -3236
rect -1383 -3240 -1367 -3236
rect -1363 -3240 -1225 -3236
rect -1221 -3240 -1208 -3236
rect -1204 -3240 -1188 -3236
rect -1184 -3240 -1167 -3236
rect -1163 -3240 -1146 -3236
rect -1142 -3240 -1125 -3236
rect -1121 -3240 -1104 -3236
rect -1100 -3240 -1083 -3236
rect -1079 -3240 -1062 -3236
rect -1058 -3240 -1042 -3236
rect -1038 -3240 -926 -3236
rect -922 -3240 -909 -3236
rect -905 -3240 -889 -3236
rect -885 -3240 -868 -3236
rect -864 -3240 -847 -3236
rect -843 -3240 -826 -3236
rect -822 -3240 -805 -3236
rect -801 -3240 -784 -3236
rect -780 -3240 -763 -3236
rect -759 -3240 -743 -3236
rect -739 -3240 -568 -3236
rect -564 -3240 -551 -3236
rect -547 -3240 -531 -3236
rect -527 -3240 -510 -3236
rect -506 -3240 -489 -3236
rect -485 -3240 -468 -3236
rect -464 -3240 -447 -3236
rect -443 -3240 -426 -3236
rect -422 -3240 -405 -3236
rect -401 -3240 -385 -3236
rect -381 -3240 -210 -3236
rect -206 -3240 -193 -3236
rect -189 -3240 -173 -3236
rect -169 -3240 -152 -3236
rect -148 -3240 -131 -3236
rect -127 -3240 -110 -3236
rect -106 -3240 -89 -3236
rect -85 -3240 -68 -3236
rect -64 -3240 -47 -3236
rect -43 -3240 -27 -3236
rect -23 -3240 148 -3236
rect 152 -3240 165 -3236
rect 169 -3240 185 -3236
rect 189 -3240 206 -3236
rect 210 -3240 227 -3236
rect 231 -3240 248 -3236
rect 252 -3240 269 -3236
rect 273 -3240 290 -3236
rect 294 -3240 311 -3236
rect 315 -3240 331 -3236
rect 335 -3240 504 -3236
rect 508 -3240 521 -3236
rect 525 -3240 541 -3236
rect 545 -3240 562 -3236
rect 566 -3240 583 -3236
rect 587 -3240 604 -3236
rect 608 -3240 625 -3236
rect 629 -3240 646 -3236
rect 650 -3240 667 -3236
rect 671 -3240 687 -3236
rect 691 -3240 862 -3236
rect 866 -3240 879 -3236
rect 883 -3240 899 -3236
rect 903 -3240 920 -3236
rect 924 -3240 941 -3236
rect 945 -3240 962 -3236
rect 966 -3240 983 -3236
rect 987 -3240 1004 -3236
rect 1008 -3240 1025 -3236
rect 1029 -3240 1045 -3236
rect 1049 -3240 1220 -3236
rect 1224 -3240 1237 -3236
rect 1241 -3240 1257 -3236
rect 1261 -3240 1278 -3236
rect 1282 -3240 1299 -3236
rect 1303 -3240 1320 -3236
rect 1324 -3240 1341 -3236
rect 1345 -3240 1362 -3236
rect 1366 -3240 1383 -3236
rect 1387 -3240 1403 -3236
rect 1407 -3240 1635 -3236
rect -2054 -3347 -2027 -3240
rect -1528 -3288 -1494 -3284
rect -1430 -3288 -1410 -3284
rect -1395 -3288 -1355 -3284
rect -1203 -3288 -1169 -3284
rect -1105 -3288 -1085 -3284
rect -1070 -3288 -1026 -3284
rect -904 -3288 -870 -3284
rect -806 -3288 -786 -3284
rect -771 -3288 -722 -3284
rect -546 -3288 -512 -3284
rect -448 -3288 -428 -3284
rect -413 -3288 -369 -3284
rect -188 -3288 -154 -3284
rect -90 -3288 -70 -3284
rect -55 -3288 -13 -3284
rect 170 -3288 204 -3284
rect 268 -3288 288 -3284
rect 303 -3288 347 -3284
rect 526 -3288 560 -3284
rect 624 -3288 644 -3284
rect 659 -3288 705 -3284
rect 884 -3288 918 -3284
rect 982 -3288 1002 -3284
rect 1017 -3288 1066 -3284
rect 1242 -3288 1276 -3284
rect 1340 -3288 1360 -3284
rect 1375 -3288 1422 -3284
rect -1578 -3296 -1552 -3292
rect -1548 -3296 -1518 -3292
rect -1497 -3296 -1466 -3292
rect -1437 -3296 -1406 -3292
rect -1395 -3296 -1368 -3292
rect -1315 -3296 -1227 -3292
rect -1223 -3296 -1193 -3292
rect -1172 -3296 -1141 -3292
rect -1112 -3296 -1081 -3292
rect -1070 -3296 -1043 -3292
rect -945 -3296 -928 -3292
rect -924 -3296 -894 -3292
rect -873 -3296 -842 -3292
rect -813 -3296 -782 -3292
rect -771 -3296 -744 -3292
rect -587 -3296 -570 -3292
rect -566 -3296 -536 -3292
rect -515 -3296 -484 -3292
rect -455 -3296 -424 -3292
rect -413 -3296 -386 -3292
rect -229 -3296 -212 -3292
rect -208 -3296 -178 -3292
rect -157 -3296 -126 -3292
rect -97 -3296 -66 -3292
rect -55 -3296 -28 -3292
rect 129 -3296 146 -3292
rect 150 -3296 180 -3292
rect 201 -3296 232 -3292
rect 261 -3296 292 -3292
rect 303 -3296 330 -3292
rect 485 -3296 502 -3292
rect 506 -3296 536 -3292
rect 557 -3296 588 -3292
rect 617 -3296 648 -3292
rect 659 -3296 686 -3292
rect 843 -3296 860 -3292
rect 864 -3296 894 -3292
rect 915 -3296 946 -3292
rect 975 -3296 1006 -3292
rect 1017 -3296 1044 -3292
rect 1201 -3296 1218 -3292
rect 1222 -3296 1252 -3292
rect 1273 -3296 1304 -3292
rect 1333 -3296 1364 -3292
rect 1375 -3296 1402 -3292
rect -1555 -3303 -1508 -3299
rect -1472 -3303 -1459 -3299
rect -1455 -3303 -1424 -3299
rect -1388 -3303 -1375 -3299
rect -1371 -3303 -1359 -3299
rect -1230 -3303 -1183 -3299
rect -1147 -3303 -1134 -3299
rect -1130 -3303 -1099 -3299
rect -1063 -3303 -1050 -3299
rect -1046 -3303 -1034 -3299
rect -931 -3303 -884 -3299
rect -848 -3303 -835 -3299
rect -831 -3303 -800 -3299
rect -764 -3303 -751 -3299
rect -747 -3303 -735 -3299
rect -573 -3303 -526 -3299
rect -490 -3303 -477 -3299
rect -473 -3303 -442 -3299
rect -406 -3303 -393 -3299
rect -389 -3303 -377 -3299
rect -215 -3303 -168 -3299
rect -132 -3303 -119 -3299
rect -115 -3303 -84 -3299
rect -48 -3303 -35 -3299
rect -31 -3303 -19 -3299
rect 143 -3303 190 -3299
rect 226 -3303 239 -3299
rect 243 -3303 274 -3299
rect 310 -3303 323 -3299
rect 327 -3303 339 -3299
rect 499 -3303 546 -3299
rect 582 -3303 595 -3299
rect 599 -3303 630 -3299
rect 666 -3303 679 -3299
rect 683 -3303 695 -3299
rect 857 -3303 904 -3299
rect 940 -3303 953 -3299
rect 957 -3303 988 -3299
rect 1024 -3303 1037 -3299
rect 1041 -3303 1053 -3299
rect 1215 -3303 1262 -3299
rect 1298 -3303 1311 -3299
rect 1315 -3303 1346 -3299
rect 1382 -3303 1395 -3299
rect 1399 -3303 1411 -3299
rect -1563 -3310 -1548 -3306
rect -1544 -3310 -1434 -3306
rect -1413 -3310 -1382 -3306
rect -1238 -3310 -1223 -3306
rect -1219 -3310 -1109 -3306
rect -1088 -3310 -1057 -3306
rect -939 -3310 -924 -3306
rect -920 -3310 -810 -3306
rect -789 -3310 -758 -3306
rect -581 -3310 -566 -3306
rect -562 -3310 -452 -3306
rect -431 -3310 -400 -3306
rect -223 -3310 -208 -3306
rect -204 -3310 -94 -3306
rect -73 -3310 -42 -3306
rect 135 -3310 150 -3306
rect 154 -3310 264 -3306
rect 285 -3310 316 -3306
rect 491 -3310 506 -3306
rect 510 -3310 620 -3306
rect 641 -3310 672 -3306
rect 849 -3310 864 -3306
rect 868 -3310 978 -3306
rect 999 -3310 1030 -3306
rect 1207 -3310 1222 -3306
rect 1226 -3310 1336 -3306
rect 1357 -3310 1388 -3306
rect -1513 -3317 -1490 -3313
rect -1471 -3317 -1452 -3313
rect -1188 -3317 -1165 -3313
rect -1146 -3317 -1127 -3313
rect -889 -3317 -866 -3313
rect -847 -3317 -828 -3313
rect -531 -3317 -508 -3313
rect -489 -3317 -470 -3313
rect -173 -3317 -150 -3313
rect -131 -3317 -112 -3313
rect 185 -3317 208 -3313
rect 227 -3317 246 -3313
rect 541 -3317 564 -3313
rect 583 -3317 602 -3313
rect 899 -3317 922 -3313
rect 941 -3317 960 -3313
rect 1257 -3317 1280 -3313
rect 1299 -3317 1318 -3313
rect 1804 -3328 1831 -3161
rect -1809 -3332 -1550 -3328
rect -1546 -3332 -1533 -3328
rect -1529 -3332 -1492 -3328
rect -1488 -3332 -1450 -3328
rect -1446 -3332 -1408 -3328
rect -1404 -3332 -1367 -3328
rect -1363 -3332 -1225 -3328
rect -1221 -3332 -1208 -3328
rect -1204 -3332 -1167 -3328
rect -1163 -3332 -1125 -3328
rect -1121 -3332 -1083 -3328
rect -1079 -3332 -1042 -3328
rect -1038 -3332 -926 -3328
rect -922 -3332 -909 -3328
rect -905 -3332 -868 -3328
rect -864 -3332 -826 -3328
rect -822 -3332 -784 -3328
rect -780 -3332 -743 -3328
rect -739 -3332 -568 -3328
rect -564 -3332 -551 -3328
rect -547 -3332 -510 -3328
rect -506 -3332 -468 -3328
rect -464 -3332 -426 -3328
rect -422 -3332 -385 -3328
rect -381 -3332 -210 -3328
rect -206 -3332 -193 -3328
rect -189 -3332 -152 -3328
rect -148 -3332 -110 -3328
rect -106 -3332 -68 -3328
rect -64 -3332 -27 -3328
rect -23 -3332 148 -3328
rect 152 -3332 165 -3328
rect 169 -3332 206 -3328
rect 210 -3332 248 -3328
rect 252 -3332 290 -3328
rect 294 -3332 331 -3328
rect 335 -3332 504 -3328
rect 508 -3332 521 -3328
rect 525 -3332 562 -3328
rect 566 -3332 604 -3328
rect 608 -3332 646 -3328
rect 650 -3332 687 -3328
rect 691 -3332 862 -3328
rect 866 -3332 879 -3328
rect 883 -3332 920 -3328
rect 924 -3332 962 -3328
rect 966 -3332 1004 -3328
rect 1008 -3332 1045 -3328
rect 1049 -3332 1220 -3328
rect 1224 -3332 1237 -3328
rect 1241 -3332 1278 -3328
rect 1282 -3332 1320 -3328
rect 1324 -3332 1362 -3328
rect 1366 -3332 1403 -3328
rect 1407 -3332 1831 -3328
rect -2054 -3351 -1309 -3347
rect -1305 -3351 -1292 -3347
rect -1288 -3351 -935 -3347
rect -931 -3351 -918 -3347
rect -914 -3351 -577 -3347
rect -573 -3351 -560 -3347
rect -556 -3351 -219 -3347
rect -215 -3351 -202 -3347
rect -198 -3351 139 -3347
rect 143 -3351 156 -3347
rect 160 -3351 495 -3347
rect 499 -3351 512 -3347
rect 516 -3351 853 -3347
rect 857 -3351 870 -3347
rect 874 -3351 1211 -3347
rect 1215 -3351 1228 -3347
rect 1232 -3351 1589 -3347
rect -2054 -3506 -2027 -3351
rect -1304 -3383 -1026 -3379
rect -930 -3383 -722 -3379
rect -572 -3383 -369 -3379
rect -214 -3383 -13 -3379
rect 144 -3383 347 -3379
rect 500 -3383 705 -3379
rect 858 -3383 1066 -3379
rect 1216 -3383 1422 -3379
rect -1351 -3391 -1297 -3387
rect -1293 -3391 -923 -3387
rect -919 -3391 -565 -3387
rect -561 -3391 -207 -3387
rect -203 -3391 151 -3387
rect 155 -3391 507 -3387
rect 511 -3391 865 -3387
rect 869 -3391 1223 -3387
rect 1227 -3391 1589 -3387
rect -975 -3404 -909 -3400
rect -612 -3404 -551 -3400
rect -259 -3404 -193 -3400
rect 101 -3404 165 -3400
rect 455 -3404 521 -3400
rect 813 -3404 879 -3400
rect 1171 -3404 1237 -3400
rect 1804 -3439 1831 -3332
rect -1411 -3443 -1292 -3439
rect -1288 -3443 -918 -3439
rect -914 -3443 -560 -3439
rect -556 -3443 -202 -3439
rect -198 -3443 156 -3439
rect 160 -3443 512 -3439
rect 516 -3443 870 -3439
rect 874 -3443 1228 -3439
rect 1232 -3443 1831 -3439
rect -2054 -3510 -1225 -3506
rect -1221 -3510 -1208 -3506
rect -1204 -3510 -1168 -3506
rect -1164 -3510 -1147 -3506
rect -1143 -3510 -926 -3506
rect -922 -3510 -900 -3506
rect -896 -3510 -883 -3506
rect -879 -3510 -843 -3506
rect -839 -3510 -822 -3506
rect -818 -3510 -805 -3506
rect -801 -3510 -765 -3506
rect -761 -3510 -741 -3506
rect -737 -3510 -704 -3506
rect -700 -3510 -568 -3506
rect -564 -3510 -542 -3506
rect -538 -3510 -525 -3506
rect -521 -3510 -485 -3506
rect -481 -3510 -464 -3506
rect -460 -3510 -447 -3506
rect -443 -3510 -407 -3506
rect -403 -3510 -383 -3506
rect -379 -3510 -346 -3506
rect -342 -3510 -210 -3506
rect -206 -3510 -184 -3506
rect -180 -3510 -167 -3506
rect -163 -3510 -127 -3506
rect -123 -3510 -106 -3506
rect -102 -3510 -89 -3506
rect -85 -3510 -49 -3506
rect -45 -3510 -25 -3506
rect -21 -3510 12 -3506
rect 16 -3510 148 -3506
rect 152 -3510 174 -3506
rect 178 -3510 191 -3506
rect 195 -3510 231 -3506
rect 235 -3510 252 -3506
rect 256 -3510 269 -3506
rect 273 -3510 309 -3506
rect 313 -3510 333 -3506
rect 337 -3510 370 -3506
rect 374 -3510 504 -3506
rect 508 -3510 530 -3506
rect 534 -3510 547 -3506
rect 551 -3510 587 -3506
rect 591 -3510 608 -3506
rect 612 -3510 625 -3506
rect 629 -3510 665 -3506
rect 669 -3510 689 -3506
rect 693 -3510 726 -3506
rect 730 -3510 862 -3506
rect 866 -3510 888 -3506
rect 892 -3510 905 -3506
rect 909 -3510 945 -3506
rect 949 -3510 966 -3506
rect 970 -3510 983 -3506
rect 987 -3510 1023 -3506
rect 1027 -3510 1047 -3506
rect 1051 -3510 1084 -3506
rect 1088 -3510 1220 -3506
rect 1224 -3510 1246 -3506
rect 1250 -3510 1263 -3506
rect 1267 -3510 1303 -3506
rect 1307 -3510 1324 -3506
rect 1328 -3510 1341 -3506
rect 1345 -3510 1381 -3506
rect 1385 -3510 1405 -3506
rect 1409 -3510 1442 -3506
rect 1446 -3510 1589 -3506
rect -2054 -3636 -2027 -3510
rect -926 -3514 -922 -3510
rect -900 -3514 -896 -3510
rect -883 -3514 -879 -3510
rect -843 -3514 -839 -3510
rect -822 -3514 -818 -3510
rect -805 -3514 -801 -3510
rect -765 -3514 -761 -3510
rect -741 -3514 -737 -3510
rect -704 -3514 -700 -3510
rect -568 -3514 -564 -3510
rect -542 -3514 -538 -3510
rect -525 -3514 -521 -3510
rect -485 -3514 -481 -3510
rect -464 -3514 -460 -3510
rect -447 -3514 -443 -3510
rect -407 -3514 -403 -3510
rect -383 -3514 -379 -3510
rect -346 -3514 -342 -3510
rect -210 -3514 -206 -3510
rect -184 -3514 -180 -3510
rect -167 -3514 -163 -3510
rect -127 -3514 -123 -3510
rect -106 -3514 -102 -3510
rect -89 -3514 -85 -3510
rect -49 -3514 -45 -3510
rect -25 -3514 -21 -3510
rect 12 -3514 16 -3510
rect 148 -3514 152 -3510
rect 174 -3514 178 -3510
rect 191 -3514 195 -3510
rect 231 -3514 235 -3510
rect 252 -3514 256 -3510
rect 269 -3514 273 -3510
rect 309 -3514 313 -3510
rect 333 -3514 337 -3510
rect 370 -3514 374 -3510
rect 504 -3514 508 -3510
rect 530 -3514 534 -3510
rect 547 -3514 551 -3510
rect 587 -3514 591 -3510
rect 608 -3514 612 -3510
rect 625 -3514 629 -3510
rect 665 -3514 669 -3510
rect 689 -3514 693 -3510
rect 726 -3514 730 -3510
rect 862 -3514 866 -3510
rect 888 -3514 892 -3510
rect 905 -3514 909 -3510
rect 945 -3514 949 -3510
rect 966 -3514 970 -3510
rect 983 -3514 987 -3510
rect 1023 -3514 1027 -3510
rect 1047 -3514 1051 -3510
rect 1084 -3514 1088 -3510
rect 1220 -3514 1224 -3510
rect 1246 -3514 1250 -3510
rect 1263 -3514 1267 -3510
rect 1303 -3514 1307 -3510
rect 1324 -3514 1328 -3510
rect 1341 -3514 1345 -3510
rect 1381 -3514 1385 -3510
rect 1405 -3514 1409 -3510
rect 1442 -3514 1446 -3510
rect -920 -3529 -858 -3525
rect -854 -3529 -824 -3525
rect -776 -3529 -746 -3525
rect -562 -3529 -500 -3525
rect -496 -3529 -466 -3525
rect -418 -3529 -388 -3525
rect -204 -3529 -142 -3525
rect -138 -3529 -108 -3525
rect -60 -3529 -30 -3525
rect 154 -3529 216 -3525
rect 220 -3529 250 -3525
rect 298 -3529 328 -3525
rect 510 -3529 572 -3525
rect 576 -3529 606 -3525
rect 654 -3529 684 -3525
rect 868 -3529 930 -3525
rect 934 -3529 964 -3525
rect 1012 -3529 1042 -3525
rect 1226 -3529 1288 -3525
rect 1292 -3529 1322 -3525
rect 1370 -3529 1400 -3525
rect -913 -3536 -882 -3532
rect -555 -3536 -524 -3532
rect -197 -3536 -166 -3532
rect 161 -3536 192 -3532
rect 517 -3536 548 -3532
rect 875 -3536 906 -3532
rect 1233 -3536 1264 -3532
rect -931 -3543 -848 -3539
rect -809 -3543 -706 -3539
rect -573 -3543 -490 -3539
rect -451 -3543 -348 -3539
rect -215 -3543 -132 -3539
rect -93 -3543 10 -3539
rect 143 -3543 226 -3539
rect 265 -3543 368 -3539
rect 499 -3543 582 -3539
rect 621 -3543 724 -3539
rect 857 -3543 940 -3539
rect 979 -3543 1082 -3539
rect 1215 -3543 1298 -3539
rect 1337 -3543 1440 -3539
rect -975 -3550 -928 -3546
rect -894 -3550 -865 -3546
rect -861 -3550 -780 -3546
rect -691 -3550 -612 -3546
rect -599 -3550 -570 -3546
rect -536 -3550 -507 -3546
rect -503 -3550 -422 -3546
rect -333 -3549 -259 -3545
rect -616 -3554 -612 -3550
rect -263 -3554 -259 -3549
rect -245 -3550 -212 -3546
rect -178 -3550 -149 -3546
rect -145 -3550 -64 -3546
rect 25 -3550 101 -3546
rect 115 -3550 146 -3546
rect 180 -3550 209 -3546
rect 213 -3550 294 -3546
rect 383 -3550 455 -3546
rect 469 -3550 502 -3546
rect 536 -3550 565 -3546
rect 569 -3550 650 -3546
rect 739 -3550 814 -3546
rect 828 -3550 860 -3546
rect 894 -3550 923 -3546
rect 927 -3550 1008 -3546
rect 1097 -3548 1164 -3544
rect 97 -3554 101 -3550
rect 451 -3554 455 -3550
rect 810 -3554 814 -3550
rect 1160 -3554 1164 -3548
rect 1171 -3550 1218 -3546
rect 1252 -3550 1281 -3546
rect 1285 -3550 1366 -3546
rect -1230 -3559 -1173 -3555
rect -1134 -3558 -902 -3554
rect -887 -3558 -804 -3554
rect -783 -3558 -687 -3554
rect -616 -3558 -544 -3554
rect -529 -3558 -446 -3554
rect -425 -3558 -328 -3554
rect -263 -3558 -186 -3554
rect -171 -3558 -88 -3554
rect -67 -3558 29 -3554
rect 97 -3558 172 -3554
rect 187 -3558 270 -3554
rect 291 -3558 388 -3554
rect 451 -3558 528 -3554
rect 543 -3558 626 -3554
rect 647 -3558 743 -3554
rect 810 -3558 886 -3554
rect 901 -3558 984 -3554
rect 1005 -3558 1101 -3554
rect 1160 -3558 1244 -3554
rect 1259 -3558 1342 -3554
rect 1363 -3558 1464 -3554
rect -1253 -3566 -1223 -3562
rect -1219 -3566 -1183 -3562
rect -1179 -3566 -1163 -3562
rect -959 -3565 -924 -3561
rect -905 -3565 -776 -3561
rect -612 -3565 -566 -3561
rect -547 -3565 -418 -3561
rect -259 -3565 -208 -3561
rect -189 -3565 -60 -3561
rect 101 -3565 150 -3561
rect 169 -3565 298 -3561
rect 455 -3565 506 -3561
rect 525 -3565 654 -3561
rect 814 -3565 864 -3561
rect 883 -3565 1012 -3561
rect 1188 -3565 1222 -3561
rect 1241 -3565 1370 -3561
rect -1279 -3573 -1227 -3569
rect -1223 -3573 -1197 -3569
rect -1193 -3573 -1149 -3569
rect -898 -3572 -794 -3568
rect -790 -3572 -760 -3568
rect -540 -3572 -436 -3568
rect -432 -3572 -402 -3568
rect -182 -3572 -78 -3568
rect -74 -3572 -44 -3568
rect 176 -3572 280 -3568
rect 284 -3572 314 -3568
rect 532 -3572 636 -3568
rect 640 -3572 670 -3568
rect 890 -3572 994 -3568
rect 998 -3572 1028 -3568
rect 1248 -3572 1352 -3568
rect 1356 -3572 1386 -3568
rect -1186 -3580 -1113 -3576
rect -924 -3579 -872 -3575
rect -868 -3579 -838 -3575
rect -566 -3579 -514 -3575
rect -510 -3579 -480 -3575
rect -208 -3579 -156 -3575
rect -152 -3579 -122 -3575
rect 150 -3579 202 -3575
rect 206 -3579 236 -3575
rect 506 -3579 558 -3575
rect 562 -3579 592 -3575
rect 864 -3579 916 -3575
rect 920 -3579 950 -3575
rect 1222 -3579 1274 -3575
rect 1278 -3579 1308 -3575
rect -1204 -3587 -1172 -3583
rect -879 -3587 -847 -3583
rect -883 -3590 -879 -3587
rect -847 -3590 -843 -3587
rect -801 -3587 -769 -3583
rect -805 -3590 -801 -3587
rect -769 -3590 -765 -3587
rect -521 -3587 -489 -3583
rect -525 -3590 -521 -3587
rect -489 -3590 -485 -3587
rect -443 -3587 -411 -3583
rect -447 -3590 -443 -3587
rect -411 -3590 -407 -3587
rect -163 -3587 -131 -3583
rect -167 -3590 -163 -3587
rect -131 -3590 -127 -3587
rect -85 -3587 -53 -3583
rect -89 -3590 -85 -3587
rect -53 -3590 -49 -3587
rect 195 -3587 227 -3583
rect 191 -3590 195 -3587
rect 227 -3590 231 -3587
rect 273 -3587 305 -3583
rect 269 -3590 273 -3587
rect 305 -3590 309 -3587
rect 551 -3587 583 -3583
rect 547 -3590 551 -3587
rect 583 -3590 587 -3587
rect 629 -3587 661 -3583
rect 625 -3590 629 -3587
rect 661 -3590 665 -3587
rect 909 -3587 941 -3583
rect 905 -3590 909 -3587
rect 941 -3590 945 -3587
rect 987 -3587 1019 -3583
rect 983 -3590 987 -3587
rect 1019 -3590 1023 -3587
rect 1267 -3587 1299 -3583
rect 1263 -3590 1267 -3587
rect 1299 -3590 1303 -3587
rect 1345 -3587 1377 -3583
rect 1341 -3590 1345 -3587
rect 1377 -3590 1381 -3587
rect -926 -3598 -922 -3594
rect -900 -3598 -896 -3594
rect -857 -3598 -853 -3594
rect -822 -3598 -818 -3594
rect -778 -3598 -774 -3594
rect -761 -3598 -757 -3594
rect -725 -3598 -721 -3594
rect -704 -3598 -700 -3594
rect -568 -3598 -564 -3594
rect -542 -3598 -538 -3594
rect -499 -3598 -495 -3594
rect -464 -3598 -460 -3594
rect -420 -3598 -416 -3594
rect -403 -3598 -399 -3594
rect -367 -3598 -363 -3594
rect -346 -3598 -342 -3594
rect -210 -3598 -206 -3594
rect -184 -3598 -180 -3594
rect -141 -3598 -137 -3594
rect -106 -3598 -102 -3594
rect -62 -3598 -58 -3594
rect -45 -3598 -41 -3594
rect -9 -3598 -5 -3594
rect 12 -3598 16 -3594
rect 148 -3598 152 -3594
rect 174 -3598 178 -3594
rect 217 -3598 221 -3594
rect 252 -3598 256 -3594
rect 296 -3598 300 -3594
rect 313 -3598 317 -3594
rect 349 -3598 353 -3594
rect 370 -3598 374 -3594
rect 504 -3598 508 -3594
rect 530 -3598 534 -3594
rect 573 -3598 577 -3594
rect 608 -3598 612 -3594
rect 652 -3598 656 -3594
rect 669 -3598 673 -3594
rect 705 -3598 709 -3594
rect 726 -3598 730 -3594
rect 862 -3598 866 -3594
rect 888 -3598 892 -3594
rect 931 -3598 935 -3594
rect 966 -3598 970 -3594
rect 1010 -3598 1014 -3594
rect 1027 -3598 1031 -3594
rect 1063 -3598 1067 -3594
rect 1084 -3598 1088 -3594
rect 1220 -3598 1224 -3594
rect 1246 -3598 1250 -3594
rect 1289 -3598 1293 -3594
rect 1324 -3598 1328 -3594
rect 1368 -3598 1372 -3594
rect 1385 -3598 1389 -3594
rect 1421 -3598 1425 -3594
rect 1442 -3598 1446 -3594
rect 1804 -3598 1831 -3443
rect -1411 -3602 -1225 -3598
rect -1221 -3602 -1181 -3598
rect -1177 -3602 -1147 -3598
rect -1143 -3602 -926 -3598
rect -922 -3602 -900 -3598
rect -896 -3602 -857 -3598
rect -853 -3602 -822 -3598
rect -818 -3602 -778 -3598
rect -774 -3602 -761 -3598
rect -757 -3602 -725 -3598
rect -721 -3602 -704 -3598
rect -700 -3602 -568 -3598
rect -564 -3602 -542 -3598
rect -538 -3602 -499 -3598
rect -495 -3602 -464 -3598
rect -460 -3602 -420 -3598
rect -416 -3602 -403 -3598
rect -399 -3602 -367 -3598
rect -363 -3602 -346 -3598
rect -342 -3602 -210 -3598
rect -206 -3602 -184 -3598
rect -180 -3602 -141 -3598
rect -137 -3602 -106 -3598
rect -102 -3602 -62 -3598
rect -58 -3602 -45 -3598
rect -41 -3602 -9 -3598
rect -5 -3602 12 -3598
rect 16 -3602 148 -3598
rect 152 -3602 174 -3598
rect 178 -3602 217 -3598
rect 221 -3602 252 -3598
rect 256 -3602 296 -3598
rect 300 -3602 313 -3598
rect 317 -3602 349 -3598
rect 353 -3602 370 -3598
rect 374 -3602 504 -3598
rect 508 -3602 530 -3598
rect 534 -3602 573 -3598
rect 577 -3602 608 -3598
rect 612 -3602 652 -3598
rect 656 -3602 669 -3598
rect 673 -3602 705 -3598
rect 709 -3602 726 -3598
rect 730 -3602 862 -3598
rect 866 -3602 888 -3598
rect 892 -3602 931 -3598
rect 935 -3602 966 -3598
rect 970 -3602 1010 -3598
rect 1014 -3602 1027 -3598
rect 1031 -3602 1063 -3598
rect 1067 -3602 1084 -3598
rect 1088 -3602 1220 -3598
rect 1224 -3602 1246 -3598
rect 1250 -3602 1289 -3598
rect 1293 -3602 1324 -3598
rect 1328 -3602 1368 -3598
rect 1372 -3602 1385 -3598
rect 1389 -3602 1421 -3598
rect 1425 -3602 1442 -3598
rect 1446 -3602 1831 -3598
rect -1253 -3609 -687 -3605
rect -599 -3609 29 -3605
rect 115 -3609 743 -3605
rect 828 -3609 1464 -3605
rect -1242 -3616 -1113 -3612
rect -959 -3616 -328 -3612
rect -245 -3616 388 -3612
rect 469 -3616 1101 -3612
rect 1188 -3616 1451 -3612
rect -2054 -3640 -1813 -3636
rect -1809 -3640 -1796 -3636
rect -1792 -3640 -1776 -3636
rect -1772 -3640 -1755 -3636
rect -1751 -3640 -1734 -3636
rect -1730 -3640 -1713 -3636
rect -1709 -3640 -1692 -3636
rect -1688 -3640 -1671 -3636
rect -1667 -3640 -1650 -3636
rect -1646 -3640 -1630 -3636
rect -1626 -3640 -1550 -3636
rect -1546 -3640 -1533 -3636
rect -1529 -3640 -1513 -3636
rect -1509 -3640 -1492 -3636
rect -1488 -3640 -1471 -3636
rect -1467 -3640 -1450 -3636
rect -1446 -3640 -1429 -3636
rect -1425 -3640 -1408 -3636
rect -1404 -3640 -1387 -3636
rect -1383 -3640 -1367 -3636
rect -1363 -3640 -1225 -3636
rect -1221 -3640 -1208 -3636
rect -1204 -3640 -1188 -3636
rect -1184 -3640 -1167 -3636
rect -1163 -3640 -1146 -3636
rect -1142 -3640 -1125 -3636
rect -1121 -3640 -1104 -3636
rect -1100 -3640 -1083 -3636
rect -1079 -3640 -1062 -3636
rect -1058 -3640 -1042 -3636
rect -1038 -3640 -925 -3636
rect -921 -3640 -908 -3636
rect -904 -3640 -888 -3636
rect -884 -3640 -867 -3636
rect -863 -3640 -846 -3636
rect -842 -3640 -825 -3636
rect -821 -3640 -804 -3636
rect -800 -3640 -783 -3636
rect -779 -3640 -762 -3636
rect -758 -3640 -742 -3636
rect -738 -3640 -568 -3636
rect -564 -3640 -551 -3636
rect -547 -3640 -531 -3636
rect -527 -3640 -510 -3636
rect -506 -3640 -489 -3636
rect -485 -3640 -468 -3636
rect -464 -3640 -447 -3636
rect -443 -3640 -426 -3636
rect -422 -3640 -405 -3636
rect -401 -3640 -385 -3636
rect -381 -3640 -210 -3636
rect -206 -3640 -193 -3636
rect -189 -3640 -173 -3636
rect -169 -3640 -152 -3636
rect -148 -3640 -131 -3636
rect -127 -3640 -110 -3636
rect -106 -3640 -89 -3636
rect -85 -3640 -68 -3636
rect -64 -3640 -47 -3636
rect -43 -3640 -27 -3636
rect -23 -3640 1751 -3636
rect -2054 -3807 -2027 -3640
rect -1791 -3688 -1757 -3684
rect -1693 -3688 -1673 -3684
rect -1658 -3688 -1555 -3684
rect -1528 -3688 -1494 -3684
rect -1430 -3688 -1410 -3684
rect -1395 -3688 -1353 -3684
rect -1203 -3688 -1169 -3684
rect -1105 -3688 -1085 -3684
rect -1070 -3688 -930 -3684
rect -903 -3688 -869 -3684
rect -805 -3688 -785 -3684
rect -770 -3688 -573 -3684
rect -546 -3688 -512 -3684
rect -448 -3688 -428 -3684
rect -413 -3688 -215 -3684
rect -188 -3688 -154 -3684
rect -90 -3688 -70 -3684
rect -55 -3688 -19 -3684
rect -1559 -3692 -1555 -3688
rect -934 -3692 -930 -3688
rect -577 -3692 -573 -3688
rect -219 -3692 -215 -3688
rect -1826 -3696 -1815 -3692
rect -1811 -3696 -1781 -3692
rect -1760 -3696 -1729 -3692
rect -1700 -3696 -1669 -3692
rect -1658 -3696 -1631 -3692
rect -1559 -3696 -1552 -3692
rect -1548 -3696 -1518 -3692
rect -1497 -3696 -1466 -3692
rect -1437 -3696 -1406 -3692
rect -1395 -3696 -1368 -3692
rect -1242 -3696 -1227 -3692
rect -1223 -3696 -1193 -3692
rect -1172 -3696 -1141 -3692
rect -1112 -3696 -1081 -3692
rect -1070 -3696 -1043 -3692
rect -934 -3696 -927 -3692
rect -923 -3696 -893 -3692
rect -872 -3696 -841 -3692
rect -812 -3696 -781 -3692
rect -770 -3696 -743 -3692
rect -577 -3696 -570 -3692
rect -566 -3696 -536 -3692
rect -515 -3696 -484 -3692
rect -455 -3696 -424 -3692
rect -413 -3696 -386 -3692
rect -219 -3696 -212 -3692
rect -208 -3696 -178 -3692
rect -157 -3696 -126 -3692
rect -97 -3696 -66 -3692
rect -55 -3696 -28 -3692
rect -1818 -3703 -1771 -3699
rect -1735 -3703 -1722 -3699
rect -1718 -3703 -1687 -3699
rect -1651 -3703 -1638 -3699
rect -1634 -3703 -1622 -3699
rect -1555 -3703 -1508 -3699
rect -1472 -3703 -1459 -3699
rect -1455 -3703 -1424 -3699
rect -1388 -3703 -1375 -3699
rect -1371 -3703 -1359 -3699
rect -1230 -3703 -1183 -3699
rect -1147 -3703 -1134 -3699
rect -1130 -3703 -1099 -3699
rect -1063 -3703 -1050 -3699
rect -1046 -3703 -1034 -3699
rect -930 -3703 -883 -3699
rect -847 -3703 -834 -3699
rect -830 -3703 -799 -3699
rect -763 -3703 -750 -3699
rect -746 -3703 -734 -3699
rect -573 -3703 -526 -3699
rect -490 -3703 -477 -3699
rect -473 -3703 -442 -3699
rect -406 -3703 -393 -3699
rect -389 -3703 -377 -3699
rect -215 -3703 -168 -3699
rect -132 -3703 -119 -3699
rect -115 -3703 -84 -3699
rect -48 -3703 -35 -3699
rect -31 -3703 -19 -3699
rect -1826 -3710 -1811 -3706
rect -1807 -3710 -1697 -3706
rect -1676 -3710 -1645 -3706
rect -1563 -3710 -1548 -3706
rect -1544 -3710 -1434 -3706
rect -1413 -3710 -1382 -3706
rect -1238 -3710 -1223 -3706
rect -1219 -3710 -1109 -3706
rect -1088 -3710 -1057 -3706
rect -938 -3710 -923 -3706
rect -919 -3710 -809 -3706
rect -788 -3710 -757 -3706
rect -581 -3710 -566 -3706
rect -562 -3710 -452 -3706
rect -431 -3710 -400 -3706
rect -223 -3710 -208 -3706
rect -204 -3710 -94 -3706
rect -73 -3710 -42 -3706
rect -1776 -3717 -1753 -3713
rect -1734 -3717 -1715 -3713
rect -1513 -3717 -1490 -3713
rect -1471 -3717 -1452 -3713
rect -1188 -3717 -1165 -3713
rect -1146 -3717 -1127 -3713
rect -888 -3717 -865 -3713
rect -846 -3717 -827 -3713
rect -531 -3717 -508 -3713
rect -489 -3717 -470 -3713
rect -173 -3717 -150 -3713
rect -131 -3717 -112 -3713
rect 1804 -3728 1831 -3602
rect -1918 -3732 -1813 -3728
rect -1809 -3732 -1796 -3728
rect -1792 -3732 -1755 -3728
rect -1751 -3732 -1713 -3728
rect -1709 -3732 -1671 -3728
rect -1667 -3732 -1630 -3728
rect -1626 -3732 -1550 -3728
rect -1546 -3732 -1533 -3728
rect -1529 -3732 -1492 -3728
rect -1488 -3732 -1450 -3728
rect -1446 -3732 -1408 -3728
rect -1404 -3732 -1367 -3728
rect -1363 -3732 -1225 -3728
rect -1221 -3732 -1208 -3728
rect -1204 -3732 -1167 -3728
rect -1163 -3732 -1125 -3728
rect -1121 -3732 -1083 -3728
rect -1079 -3732 -1042 -3728
rect -1038 -3732 -925 -3728
rect -921 -3732 -908 -3728
rect -904 -3732 -867 -3728
rect -863 -3732 -825 -3728
rect -821 -3732 -783 -3728
rect -779 -3732 -742 -3728
rect -738 -3732 -568 -3728
rect -564 -3732 -551 -3728
rect -547 -3732 -510 -3728
rect -506 -3732 -468 -3728
rect -464 -3732 -426 -3728
rect -422 -3732 -385 -3728
rect -381 -3732 -210 -3728
rect -206 -3732 -193 -3728
rect -189 -3732 -152 -3728
rect -148 -3732 -110 -3728
rect -106 -3732 -68 -3728
rect -64 -3732 -27 -3728
rect -23 -3732 1831 -3728
rect -1568 -3740 -1353 -3736
rect -2054 -3811 -1550 -3807
rect -1546 -3811 -1533 -3807
rect -1529 -3811 -1513 -3807
rect -1509 -3811 -1492 -3807
rect -1488 -3811 -1471 -3807
rect -1467 -3811 -1450 -3807
rect -1446 -3811 -1429 -3807
rect -1425 -3811 -1408 -3807
rect -1404 -3811 -1387 -3807
rect -1383 -3811 -1367 -3807
rect -1363 -3811 -1225 -3807
rect -1221 -3811 -1208 -3807
rect -1204 -3811 -1188 -3807
rect -1184 -3811 -1167 -3807
rect -1163 -3811 -1146 -3807
rect -1142 -3811 -1125 -3807
rect -1121 -3811 -1104 -3807
rect -1100 -3811 -1083 -3807
rect -1079 -3811 -1062 -3807
rect -1058 -3811 -1042 -3807
rect -1038 -3811 -925 -3807
rect -921 -3811 -908 -3807
rect -904 -3811 -888 -3807
rect -884 -3811 -867 -3807
rect -863 -3811 -846 -3807
rect -842 -3811 -825 -3807
rect -821 -3811 -804 -3807
rect -800 -3811 -783 -3807
rect -779 -3811 -762 -3807
rect -758 -3811 -742 -3807
rect -738 -3811 -568 -3807
rect -564 -3811 -551 -3807
rect -547 -3811 -531 -3807
rect -527 -3811 -510 -3807
rect -506 -3811 -489 -3807
rect -485 -3811 -468 -3807
rect -464 -3811 -447 -3807
rect -443 -3811 -426 -3807
rect -422 -3811 -405 -3807
rect -401 -3811 -385 -3807
rect -381 -3811 -210 -3807
rect -206 -3811 -193 -3807
rect -189 -3811 -173 -3807
rect -169 -3811 -152 -3807
rect -148 -3811 -131 -3807
rect -127 -3811 -110 -3807
rect -106 -3811 -89 -3807
rect -85 -3811 -68 -3807
rect -64 -3811 -47 -3807
rect -43 -3811 -27 -3807
rect -23 -3811 148 -3807
rect 152 -3811 165 -3807
rect 169 -3811 185 -3807
rect 189 -3811 206 -3807
rect 210 -3811 227 -3807
rect 231 -3811 248 -3807
rect 252 -3811 269 -3807
rect 273 -3811 290 -3807
rect 294 -3811 311 -3807
rect 315 -3811 331 -3807
rect 335 -3811 504 -3807
rect 508 -3811 521 -3807
rect 525 -3811 541 -3807
rect 545 -3811 562 -3807
rect 566 -3811 583 -3807
rect 587 -3811 604 -3807
rect 608 -3811 625 -3807
rect 629 -3811 646 -3807
rect 650 -3811 667 -3807
rect 671 -3811 687 -3807
rect 691 -3811 862 -3807
rect 866 -3811 879 -3807
rect 883 -3811 899 -3807
rect 903 -3811 920 -3807
rect 924 -3811 941 -3807
rect 945 -3811 962 -3807
rect 966 -3811 983 -3807
rect 987 -3811 1004 -3807
rect 1008 -3811 1025 -3807
rect 1029 -3811 1045 -3807
rect 1049 -3811 1220 -3807
rect 1224 -3811 1237 -3807
rect 1241 -3811 1257 -3807
rect 1261 -3811 1278 -3807
rect 1282 -3811 1299 -3807
rect 1303 -3811 1320 -3807
rect 1324 -3811 1341 -3807
rect 1345 -3811 1362 -3807
rect 1366 -3811 1383 -3807
rect 1387 -3811 1403 -3807
rect 1407 -3811 1745 -3807
rect -2054 -3982 -2027 -3811
rect -1528 -3859 -1494 -3855
rect -1430 -3859 -1410 -3855
rect -1395 -3859 -1355 -3855
rect -1203 -3859 -1169 -3855
rect -1105 -3859 -1085 -3855
rect -1070 -3859 -1028 -3855
rect -903 -3859 -869 -3855
rect -805 -3859 -785 -3855
rect -770 -3859 -723 -3855
rect -546 -3859 -512 -3855
rect -448 -3859 -428 -3855
rect -413 -3859 -369 -3855
rect -188 -3859 -154 -3855
rect -90 -3859 -70 -3855
rect -55 -3859 -9 -3855
rect 170 -3859 204 -3855
rect 268 -3859 288 -3855
rect 303 -3859 349 -3855
rect 526 -3859 560 -3855
rect 624 -3859 644 -3855
rect 659 -3859 702 -3855
rect 884 -3859 918 -3855
rect 982 -3859 1002 -3855
rect 1017 -3859 1060 -3855
rect 1242 -3859 1276 -3855
rect 1340 -3859 1360 -3855
rect 1375 -3859 1424 -3855
rect -1568 -3867 -1552 -3863
rect -1548 -3867 -1518 -3863
rect -1497 -3867 -1466 -3863
rect -1437 -3867 -1406 -3863
rect -1395 -3867 -1368 -3863
rect -1253 -3867 -1227 -3863
rect -1223 -3867 -1193 -3863
rect -1172 -3867 -1141 -3863
rect -1112 -3867 -1081 -3863
rect -1070 -3867 -1043 -3863
rect -959 -3867 -927 -3863
rect -923 -3867 -893 -3863
rect -872 -3867 -841 -3863
rect -812 -3867 -781 -3863
rect -770 -3867 -743 -3863
rect -599 -3867 -570 -3863
rect -566 -3867 -536 -3863
rect -515 -3867 -484 -3863
rect -455 -3867 -424 -3863
rect -413 -3867 -386 -3863
rect -245 -3867 -212 -3863
rect -208 -3867 -178 -3863
rect -157 -3867 -126 -3863
rect -97 -3867 -66 -3863
rect -55 -3867 -28 -3863
rect 115 -3867 146 -3863
rect 150 -3867 180 -3863
rect 201 -3867 232 -3863
rect 261 -3867 292 -3863
rect 303 -3867 330 -3863
rect 469 -3867 502 -3863
rect 506 -3867 536 -3863
rect 557 -3867 588 -3863
rect 617 -3867 648 -3863
rect 659 -3867 686 -3863
rect 828 -3867 860 -3863
rect 864 -3867 894 -3863
rect 915 -3867 946 -3863
rect 975 -3867 1006 -3863
rect 1017 -3867 1044 -3863
rect 1188 -3867 1218 -3863
rect 1222 -3867 1252 -3863
rect 1273 -3867 1304 -3863
rect 1333 -3867 1364 -3863
rect 1375 -3867 1402 -3863
rect -1555 -3874 -1508 -3870
rect -1472 -3874 -1459 -3870
rect -1455 -3874 -1424 -3870
rect -1388 -3874 -1375 -3870
rect -1371 -3874 -1359 -3870
rect -1230 -3874 -1183 -3870
rect -1147 -3874 -1134 -3870
rect -1130 -3874 -1099 -3870
rect -1063 -3874 -1050 -3870
rect -1046 -3874 -1034 -3870
rect -930 -3874 -883 -3870
rect -847 -3874 -834 -3870
rect -830 -3874 -799 -3870
rect -763 -3874 -750 -3870
rect -746 -3874 -734 -3870
rect -573 -3874 -526 -3870
rect -490 -3874 -477 -3870
rect -473 -3874 -442 -3870
rect -406 -3874 -393 -3870
rect -389 -3874 -377 -3870
rect -215 -3874 -168 -3870
rect -132 -3874 -119 -3870
rect -115 -3874 -84 -3870
rect -48 -3874 -35 -3870
rect -31 -3874 -19 -3870
rect 143 -3874 190 -3870
rect 226 -3874 239 -3870
rect 243 -3874 274 -3870
rect 310 -3874 323 -3870
rect 327 -3874 339 -3870
rect 499 -3874 546 -3870
rect 582 -3874 595 -3870
rect 599 -3874 630 -3870
rect 666 -3874 679 -3870
rect 683 -3874 695 -3870
rect 857 -3874 904 -3870
rect 940 -3874 953 -3870
rect 957 -3874 988 -3870
rect 1024 -3874 1037 -3870
rect 1041 -3874 1053 -3870
rect 1215 -3874 1262 -3870
rect 1298 -3874 1311 -3870
rect 1315 -3874 1346 -3870
rect 1382 -3874 1395 -3870
rect 1399 -3874 1411 -3870
rect -1563 -3881 -1548 -3877
rect -1544 -3881 -1434 -3877
rect -1413 -3881 -1382 -3877
rect -1238 -3881 -1223 -3877
rect -1219 -3881 -1109 -3877
rect -1088 -3881 -1057 -3877
rect -938 -3881 -923 -3877
rect -919 -3881 -809 -3877
rect -788 -3881 -757 -3877
rect -581 -3881 -566 -3877
rect -562 -3881 -452 -3877
rect -431 -3881 -400 -3877
rect -223 -3881 -208 -3877
rect -204 -3881 -94 -3877
rect -73 -3881 -42 -3877
rect 135 -3881 150 -3877
rect 154 -3881 264 -3877
rect 285 -3881 316 -3877
rect 491 -3881 506 -3877
rect 510 -3881 620 -3877
rect 641 -3881 672 -3877
rect 849 -3881 864 -3877
rect 868 -3881 978 -3877
rect 999 -3881 1030 -3877
rect 1207 -3881 1222 -3877
rect 1226 -3881 1336 -3877
rect 1357 -3881 1388 -3877
rect -1513 -3888 -1490 -3884
rect -1471 -3888 -1452 -3884
rect -1188 -3888 -1165 -3884
rect -1146 -3888 -1127 -3884
rect -888 -3888 -865 -3884
rect -846 -3888 -827 -3884
rect -531 -3888 -508 -3884
rect -489 -3888 -470 -3884
rect -173 -3888 -150 -3884
rect -131 -3888 -112 -3884
rect 185 -3888 208 -3884
rect 227 -3888 246 -3884
rect 541 -3888 564 -3884
rect 583 -3888 602 -3884
rect 899 -3888 922 -3884
rect 941 -3888 960 -3884
rect 1257 -3888 1280 -3884
rect 1299 -3888 1318 -3884
rect 1804 -3899 1831 -3732
rect -1591 -3903 -1550 -3899
rect -1546 -3903 -1533 -3899
rect -1529 -3903 -1492 -3899
rect -1488 -3903 -1450 -3899
rect -1446 -3903 -1408 -3899
rect -1404 -3903 -1367 -3899
rect -1363 -3903 -1225 -3899
rect -1221 -3903 -1208 -3899
rect -1204 -3903 -1167 -3899
rect -1163 -3903 -1125 -3899
rect -1121 -3903 -1083 -3899
rect -1079 -3903 -1042 -3899
rect -1038 -3903 -925 -3899
rect -921 -3903 -908 -3899
rect -904 -3903 -867 -3899
rect -863 -3903 -825 -3899
rect -821 -3903 -783 -3899
rect -779 -3903 -742 -3899
rect -738 -3903 -568 -3899
rect -564 -3903 -551 -3899
rect -547 -3903 -510 -3899
rect -506 -3903 -468 -3899
rect -464 -3903 -426 -3899
rect -422 -3903 -385 -3899
rect -381 -3903 -210 -3899
rect -206 -3903 -193 -3899
rect -189 -3903 -152 -3899
rect -148 -3903 -110 -3899
rect -106 -3903 -68 -3899
rect -64 -3903 -27 -3899
rect -23 -3903 148 -3899
rect 152 -3903 165 -3899
rect 169 -3903 206 -3899
rect 210 -3903 248 -3899
rect 252 -3903 290 -3899
rect 294 -3903 331 -3899
rect 335 -3903 504 -3899
rect 508 -3903 521 -3899
rect 525 -3903 562 -3899
rect 566 -3903 604 -3899
rect 608 -3903 646 -3899
rect 650 -3903 687 -3899
rect 691 -3903 862 -3899
rect 866 -3903 879 -3899
rect 883 -3903 920 -3899
rect 924 -3903 962 -3899
rect 966 -3903 1004 -3899
rect 1008 -3903 1045 -3899
rect 1049 -3903 1220 -3899
rect 1224 -3903 1237 -3899
rect 1241 -3903 1278 -3899
rect 1282 -3903 1320 -3899
rect 1324 -3903 1362 -3899
rect 1366 -3903 1403 -3899
rect 1407 -3903 1831 -3899
rect -1571 -3911 -1355 -3907
rect -1253 -3910 -1028 -3906
rect -959 -3911 -723 -3907
rect -599 -3910 -369 -3906
rect -245 -3910 -9 -3906
rect 115 -3910 349 -3906
rect 469 -3911 702 -3907
rect 828 -3910 1060 -3906
rect 1188 -3910 1424 -3906
rect -2054 -3986 -1550 -3982
rect -1546 -3986 -1533 -3982
rect -1529 -3986 -1513 -3982
rect -1509 -3986 -1492 -3982
rect -1488 -3986 -1471 -3982
rect -1467 -3986 -1450 -3982
rect -1446 -3986 -1429 -3982
rect -1425 -3986 -1408 -3982
rect -1404 -3986 -1387 -3982
rect -1383 -3986 -1367 -3982
rect -1363 -3986 -1225 -3982
rect -1221 -3986 -1208 -3982
rect -1204 -3986 -1188 -3982
rect -1184 -3986 -1167 -3982
rect -1163 -3986 -1146 -3982
rect -1142 -3986 -1125 -3982
rect -1121 -3986 -1104 -3982
rect -1100 -3986 -1083 -3982
rect -1079 -3986 -1062 -3982
rect -1058 -3986 -1042 -3982
rect -1038 -3986 -926 -3982
rect -922 -3986 -909 -3982
rect -905 -3986 -889 -3982
rect -885 -3986 -868 -3982
rect -864 -3986 -847 -3982
rect -843 -3986 -826 -3982
rect -822 -3986 -805 -3982
rect -801 -3986 -784 -3982
rect -780 -3986 -763 -3982
rect -759 -3986 -743 -3982
rect -739 -3986 -568 -3982
rect -564 -3986 -551 -3982
rect -547 -3986 -531 -3982
rect -527 -3986 -510 -3982
rect -506 -3986 -489 -3982
rect -485 -3986 -468 -3982
rect -464 -3986 -447 -3982
rect -443 -3986 -426 -3982
rect -422 -3986 -405 -3982
rect -401 -3986 -385 -3982
rect -381 -3986 -210 -3982
rect -206 -3986 -193 -3982
rect -189 -3986 -173 -3982
rect -169 -3986 -152 -3982
rect -148 -3986 -131 -3982
rect -127 -3986 -110 -3982
rect -106 -3986 -89 -3982
rect -85 -3986 -68 -3982
rect -64 -3986 -47 -3982
rect -43 -3986 -27 -3982
rect -23 -3986 148 -3982
rect 152 -3986 165 -3982
rect 169 -3986 185 -3982
rect 189 -3986 206 -3982
rect 210 -3986 227 -3982
rect 231 -3986 248 -3982
rect 252 -3986 269 -3982
rect 273 -3986 290 -3982
rect 294 -3986 311 -3982
rect 315 -3986 331 -3982
rect 335 -3986 504 -3982
rect 508 -3986 521 -3982
rect 525 -3986 541 -3982
rect 545 -3986 562 -3982
rect 566 -3986 583 -3982
rect 587 -3986 604 -3982
rect 608 -3986 625 -3982
rect 629 -3986 646 -3982
rect 650 -3986 667 -3982
rect 671 -3986 687 -3982
rect 691 -3986 862 -3982
rect 866 -3986 879 -3982
rect 883 -3986 899 -3982
rect 903 -3986 920 -3982
rect 924 -3986 941 -3982
rect 945 -3986 962 -3982
rect 966 -3986 983 -3982
rect 987 -3986 1004 -3982
rect 1008 -3986 1025 -3982
rect 1029 -3986 1045 -3982
rect 1049 -3986 1220 -3982
rect 1224 -3986 1237 -3982
rect 1241 -3986 1257 -3982
rect 1261 -3986 1278 -3982
rect 1282 -3986 1299 -3982
rect 1303 -3986 1320 -3982
rect 1324 -3986 1341 -3982
rect 1345 -3986 1362 -3982
rect 1366 -3986 1383 -3982
rect 1387 -3986 1403 -3982
rect 1407 -3986 1738 -3982
rect -2054 -4097 -2027 -3986
rect -1528 -4034 -1494 -4030
rect -1430 -4034 -1410 -4030
rect -1395 -4034 -1357 -4030
rect -1203 -4034 -1169 -4030
rect -1105 -4034 -1085 -4030
rect -1070 -4034 -1024 -4030
rect -904 -4034 -870 -4030
rect -806 -4034 -786 -4030
rect -771 -4034 -719 -4030
rect -546 -4034 -512 -4030
rect -448 -4034 -428 -4030
rect -413 -4034 -369 -4030
rect -188 -4034 -154 -4030
rect -90 -4034 -70 -4030
rect -55 -4034 -9 -4030
rect 170 -4034 204 -4030
rect 268 -4034 288 -4030
rect 303 -4034 348 -4030
rect 526 -4034 560 -4030
rect 624 -4034 644 -4030
rect 659 -4034 705 -4030
rect 884 -4034 918 -4030
rect 982 -4034 1002 -4030
rect 1017 -4034 1063 -4030
rect 1242 -4034 1276 -4030
rect 1340 -4034 1360 -4030
rect 1375 -4034 1418 -4030
rect -1571 -4042 -1552 -4038
rect -1548 -4042 -1518 -4038
rect -1497 -4042 -1466 -4038
rect -1437 -4042 -1406 -4038
rect -1395 -4042 -1368 -4038
rect -1315 -4042 -1227 -4038
rect -1223 -4042 -1193 -4038
rect -1172 -4042 -1141 -4038
rect -1112 -4042 -1081 -4038
rect -1070 -4042 -1043 -4038
rect -945 -4042 -928 -4038
rect -924 -4042 -894 -4038
rect -873 -4042 -842 -4038
rect -813 -4042 -782 -4038
rect -771 -4042 -744 -4038
rect -587 -4042 -570 -4038
rect -566 -4042 -536 -4038
rect -515 -4042 -484 -4038
rect -455 -4042 -424 -4038
rect -413 -4042 -386 -4038
rect -229 -4042 -212 -4038
rect -208 -4042 -178 -4038
rect -157 -4042 -126 -4038
rect -97 -4042 -66 -4038
rect -55 -4042 -28 -4038
rect 129 -4042 146 -4038
rect 150 -4042 180 -4038
rect 201 -4042 232 -4038
rect 261 -4042 292 -4038
rect 303 -4042 330 -4038
rect 485 -4042 502 -4038
rect 506 -4042 536 -4038
rect 557 -4042 588 -4038
rect 617 -4042 648 -4038
rect 659 -4042 686 -4038
rect 843 -4042 860 -4038
rect 864 -4042 894 -4038
rect 915 -4042 946 -4038
rect 975 -4042 1006 -4038
rect 1017 -4042 1044 -4038
rect 1201 -4042 1218 -4038
rect 1222 -4042 1252 -4038
rect 1273 -4042 1304 -4038
rect 1333 -4042 1364 -4038
rect 1375 -4042 1402 -4038
rect -1555 -4049 -1508 -4045
rect -1472 -4049 -1459 -4045
rect -1455 -4049 -1424 -4045
rect -1388 -4049 -1375 -4045
rect -1371 -4049 -1359 -4045
rect -1230 -4049 -1183 -4045
rect -1147 -4049 -1134 -4045
rect -1130 -4049 -1099 -4045
rect -1063 -4049 -1050 -4045
rect -1046 -4049 -1034 -4045
rect -931 -4049 -884 -4045
rect -848 -4049 -835 -4045
rect -831 -4049 -800 -4045
rect -764 -4049 -751 -4045
rect -747 -4049 -735 -4045
rect -573 -4049 -526 -4045
rect -490 -4049 -477 -4045
rect -473 -4049 -442 -4045
rect -406 -4049 -393 -4045
rect -389 -4049 -377 -4045
rect -215 -4049 -168 -4045
rect -132 -4049 -119 -4045
rect -115 -4049 -84 -4045
rect -48 -4049 -35 -4045
rect -31 -4049 -19 -4045
rect 143 -4049 190 -4045
rect 226 -4049 239 -4045
rect 243 -4049 274 -4045
rect 310 -4049 323 -4045
rect 327 -4049 339 -4045
rect 499 -4049 546 -4045
rect 582 -4049 595 -4045
rect 599 -4049 630 -4045
rect 666 -4049 679 -4045
rect 683 -4049 695 -4045
rect 857 -4049 904 -4045
rect 940 -4049 953 -4045
rect 957 -4049 988 -4045
rect 1024 -4049 1037 -4045
rect 1041 -4049 1053 -4045
rect 1215 -4049 1262 -4045
rect 1298 -4049 1311 -4045
rect 1315 -4049 1346 -4045
rect 1382 -4049 1395 -4045
rect 1399 -4049 1411 -4045
rect -1563 -4056 -1548 -4052
rect -1544 -4056 -1434 -4052
rect -1413 -4056 -1382 -4052
rect -1238 -4056 -1223 -4052
rect -1219 -4056 -1109 -4052
rect -1088 -4056 -1057 -4052
rect -939 -4056 -924 -4052
rect -920 -4056 -810 -4052
rect -789 -4056 -758 -4052
rect -581 -4056 -566 -4052
rect -562 -4056 -452 -4052
rect -431 -4056 -400 -4052
rect -223 -4056 -208 -4052
rect -204 -4056 -94 -4052
rect -73 -4056 -42 -4052
rect 135 -4056 150 -4052
rect 154 -4056 264 -4052
rect 285 -4056 316 -4052
rect 491 -4056 506 -4052
rect 510 -4056 620 -4052
rect 641 -4056 672 -4052
rect 849 -4056 864 -4052
rect 868 -4056 978 -4052
rect 999 -4056 1030 -4052
rect 1207 -4056 1222 -4052
rect 1226 -4056 1336 -4052
rect 1357 -4056 1388 -4052
rect -1513 -4063 -1490 -4059
rect -1471 -4063 -1452 -4059
rect -1188 -4063 -1165 -4059
rect -1146 -4063 -1127 -4059
rect -889 -4063 -866 -4059
rect -847 -4063 -828 -4059
rect -531 -4063 -508 -4059
rect -489 -4063 -470 -4059
rect -173 -4063 -150 -4059
rect -131 -4063 -112 -4059
rect 185 -4063 208 -4059
rect 227 -4063 246 -4059
rect 541 -4063 564 -4059
rect 583 -4063 602 -4059
rect 899 -4063 922 -4059
rect 941 -4063 960 -4059
rect 1257 -4063 1280 -4059
rect 1299 -4063 1318 -4059
rect 1804 -4074 1831 -3903
rect -1591 -4078 -1550 -4074
rect -1546 -4078 -1533 -4074
rect -1529 -4078 -1492 -4074
rect -1488 -4078 -1450 -4074
rect -1446 -4078 -1408 -4074
rect -1404 -4078 -1367 -4074
rect -1363 -4078 -1225 -4074
rect -1221 -4078 -1208 -4074
rect -1204 -4078 -1167 -4074
rect -1163 -4078 -1125 -4074
rect -1121 -4078 -1083 -4074
rect -1079 -4078 -1042 -4074
rect -1038 -4078 -926 -4074
rect -922 -4078 -909 -4074
rect -905 -4078 -868 -4074
rect -864 -4078 -826 -4074
rect -822 -4078 -784 -4074
rect -780 -4078 -743 -4074
rect -739 -4078 -568 -4074
rect -564 -4078 -551 -4074
rect -547 -4078 -510 -4074
rect -506 -4078 -468 -4074
rect -464 -4078 -426 -4074
rect -422 -4078 -385 -4074
rect -381 -4078 -210 -4074
rect -206 -4078 -193 -4074
rect -189 -4078 -152 -4074
rect -148 -4078 -110 -4074
rect -106 -4078 -68 -4074
rect -64 -4078 -27 -4074
rect -23 -4078 148 -4074
rect 152 -4078 165 -4074
rect 169 -4078 206 -4074
rect 210 -4078 248 -4074
rect 252 -4078 290 -4074
rect 294 -4078 331 -4074
rect 335 -4078 504 -4074
rect 508 -4078 521 -4074
rect 525 -4078 562 -4074
rect 566 -4078 604 -4074
rect 608 -4078 646 -4074
rect 650 -4078 687 -4074
rect 691 -4078 862 -4074
rect 866 -4078 879 -4074
rect 883 -4078 920 -4074
rect 924 -4078 962 -4074
rect 966 -4078 1004 -4074
rect 1008 -4078 1045 -4074
rect 1049 -4078 1220 -4074
rect 1224 -4078 1237 -4074
rect 1241 -4078 1278 -4074
rect 1282 -4078 1320 -4074
rect 1324 -4078 1362 -4074
rect 1366 -4078 1403 -4074
rect 1407 -4078 1831 -4074
rect -2054 -4101 -1309 -4097
rect -1305 -4101 -1292 -4097
rect -1288 -4101 -935 -4097
rect -931 -4101 -918 -4097
rect -914 -4101 -577 -4097
rect -573 -4101 -560 -4097
rect -556 -4101 -219 -4097
rect -215 -4101 -202 -4097
rect -198 -4101 139 -4097
rect 143 -4101 156 -4097
rect 160 -4101 495 -4097
rect 499 -4101 512 -4097
rect 516 -4101 853 -4097
rect 857 -4101 870 -4097
rect 874 -4101 1211 -4097
rect 1215 -4101 1228 -4097
rect 1232 -4101 1589 -4097
rect -2054 -4256 -2027 -4101
rect -1304 -4133 -1024 -4129
rect -930 -4133 -719 -4129
rect -572 -4133 -369 -4129
rect -214 -4133 -9 -4129
rect 144 -4133 348 -4129
rect 500 -4133 705 -4129
rect 858 -4133 1063 -4129
rect 1216 -4133 1418 -4129
rect -1353 -4141 -1297 -4137
rect -1293 -4141 -923 -4137
rect -919 -4141 -565 -4137
rect -561 -4141 -207 -4137
rect -203 -4141 151 -4137
rect 155 -4141 507 -4137
rect 511 -4141 865 -4137
rect 869 -4141 1223 -4137
rect 1227 -4141 1589 -4137
rect -975 -4154 -909 -4150
rect -612 -4154 -551 -4150
rect -259 -4154 -193 -4150
rect 101 -4154 165 -4150
rect 455 -4154 521 -4150
rect 814 -4154 879 -4150
rect 1171 -4154 1237 -4150
rect 1804 -4189 1831 -4078
rect -1411 -4193 -1292 -4189
rect -1288 -4193 -918 -4189
rect -914 -4193 -560 -4189
rect -556 -4193 -202 -4189
rect -198 -4193 156 -4189
rect 160 -4193 512 -4189
rect 516 -4193 870 -4189
rect 874 -4193 1228 -4189
rect 1232 -4193 1831 -4189
rect -2054 -4260 -1225 -4256
rect -1221 -4260 -1208 -4256
rect -1204 -4260 -1168 -4256
rect -1164 -4260 -1147 -4256
rect -1143 -4260 -926 -4256
rect -922 -4260 -900 -4256
rect -896 -4260 -883 -4256
rect -879 -4260 -843 -4256
rect -839 -4260 -822 -4256
rect -818 -4260 -805 -4256
rect -801 -4260 -765 -4256
rect -761 -4260 -741 -4256
rect -737 -4260 -704 -4256
rect -700 -4260 -568 -4256
rect -564 -4260 -542 -4256
rect -538 -4260 -525 -4256
rect -521 -4260 -485 -4256
rect -481 -4260 -464 -4256
rect -460 -4260 -447 -4256
rect -443 -4260 -407 -4256
rect -403 -4260 -383 -4256
rect -379 -4260 -346 -4256
rect -342 -4260 -210 -4256
rect -206 -4260 -184 -4256
rect -180 -4260 -167 -4256
rect -163 -4260 -127 -4256
rect -123 -4260 -106 -4256
rect -102 -4260 -89 -4256
rect -85 -4260 -49 -4256
rect -45 -4260 -25 -4256
rect -21 -4260 12 -4256
rect 16 -4260 148 -4256
rect 152 -4260 174 -4256
rect 178 -4260 191 -4256
rect 195 -4260 231 -4256
rect 235 -4260 252 -4256
rect 256 -4260 269 -4256
rect 273 -4260 309 -4256
rect 313 -4260 333 -4256
rect 337 -4260 370 -4256
rect 374 -4260 504 -4256
rect 508 -4260 530 -4256
rect 534 -4260 547 -4256
rect 551 -4260 587 -4256
rect 591 -4260 608 -4256
rect 612 -4260 625 -4256
rect 629 -4260 665 -4256
rect 669 -4260 689 -4256
rect 693 -4260 726 -4256
rect 730 -4260 862 -4256
rect 866 -4260 888 -4256
rect 892 -4260 905 -4256
rect 909 -4260 945 -4256
rect 949 -4260 966 -4256
rect 970 -4260 983 -4256
rect 987 -4260 1023 -4256
rect 1027 -4260 1047 -4256
rect 1051 -4260 1084 -4256
rect 1088 -4260 1220 -4256
rect 1224 -4260 1246 -4256
rect 1250 -4260 1263 -4256
rect 1267 -4260 1303 -4256
rect 1307 -4260 1324 -4256
rect 1328 -4260 1341 -4256
rect 1345 -4260 1381 -4256
rect 1385 -4260 1405 -4256
rect 1409 -4260 1442 -4256
rect 1446 -4260 1589 -4256
rect -2054 -4379 -2027 -4260
rect -926 -4264 -922 -4260
rect -900 -4264 -896 -4260
rect -883 -4264 -879 -4260
rect -843 -4264 -839 -4260
rect -822 -4264 -818 -4260
rect -805 -4264 -801 -4260
rect -765 -4264 -761 -4260
rect -741 -4264 -737 -4260
rect -704 -4264 -700 -4260
rect -568 -4264 -564 -4260
rect -542 -4264 -538 -4260
rect -525 -4264 -521 -4260
rect -485 -4264 -481 -4260
rect -464 -4264 -460 -4260
rect -447 -4264 -443 -4260
rect -407 -4264 -403 -4260
rect -383 -4264 -379 -4260
rect -346 -4264 -342 -4260
rect -210 -4264 -206 -4260
rect -184 -4264 -180 -4260
rect -167 -4264 -163 -4260
rect -127 -4264 -123 -4260
rect -106 -4264 -102 -4260
rect -89 -4264 -85 -4260
rect -49 -4264 -45 -4260
rect -25 -4264 -21 -4260
rect 12 -4264 16 -4260
rect 148 -4264 152 -4260
rect 174 -4264 178 -4260
rect 191 -4264 195 -4260
rect 231 -4264 235 -4260
rect 252 -4264 256 -4260
rect 269 -4264 273 -4260
rect 309 -4264 313 -4260
rect 333 -4264 337 -4260
rect 370 -4264 374 -4260
rect 504 -4264 508 -4260
rect 530 -4264 534 -4260
rect 547 -4264 551 -4260
rect 587 -4264 591 -4260
rect 608 -4264 612 -4260
rect 625 -4264 629 -4260
rect 665 -4264 669 -4260
rect 689 -4264 693 -4260
rect 726 -4264 730 -4260
rect 862 -4264 866 -4260
rect 888 -4264 892 -4260
rect 905 -4264 909 -4260
rect 945 -4264 949 -4260
rect 966 -4264 970 -4260
rect 983 -4264 987 -4260
rect 1023 -4264 1027 -4260
rect 1047 -4264 1051 -4260
rect 1084 -4264 1088 -4260
rect 1220 -4264 1224 -4260
rect 1246 -4264 1250 -4260
rect 1263 -4264 1267 -4260
rect 1303 -4264 1307 -4260
rect 1324 -4264 1328 -4260
rect 1341 -4264 1345 -4260
rect 1381 -4264 1385 -4260
rect 1405 -4264 1409 -4260
rect 1442 -4264 1446 -4260
rect -920 -4279 -858 -4275
rect -854 -4279 -824 -4275
rect -776 -4279 -746 -4275
rect -562 -4279 -500 -4275
rect -496 -4279 -466 -4275
rect -418 -4279 -388 -4275
rect -204 -4279 -142 -4275
rect -138 -4279 -108 -4275
rect -60 -4279 -30 -4275
rect 154 -4279 216 -4275
rect 220 -4279 250 -4275
rect 298 -4279 328 -4275
rect 510 -4279 572 -4275
rect 576 -4279 606 -4275
rect 654 -4279 684 -4275
rect 868 -4279 930 -4275
rect 934 -4279 964 -4275
rect 1012 -4279 1042 -4275
rect 1226 -4279 1288 -4275
rect 1292 -4279 1322 -4275
rect 1370 -4279 1400 -4275
rect -913 -4286 -882 -4282
rect -555 -4286 -524 -4282
rect -197 -4286 -166 -4282
rect 161 -4286 192 -4282
rect 517 -4286 548 -4282
rect 875 -4286 906 -4282
rect 1233 -4286 1264 -4282
rect -931 -4293 -848 -4289
rect -809 -4293 -706 -4289
rect -573 -4293 -490 -4289
rect -451 -4293 -348 -4289
rect -215 -4293 -132 -4289
rect -93 -4293 10 -4289
rect 143 -4293 226 -4289
rect 265 -4293 368 -4289
rect 499 -4293 582 -4289
rect 621 -4293 724 -4289
rect 857 -4293 940 -4289
rect 979 -4293 1082 -4289
rect 1215 -4293 1298 -4289
rect 1337 -4293 1440 -4289
rect -975 -4300 -928 -4296
rect -894 -4300 -865 -4296
rect -861 -4300 -780 -4296
rect -691 -4300 -612 -4296
rect -599 -4300 -570 -4296
rect -536 -4300 -507 -4296
rect -503 -4300 -422 -4296
rect -333 -4299 -259 -4295
rect -616 -4304 -612 -4300
rect -263 -4304 -259 -4299
rect -245 -4300 -212 -4296
rect -178 -4300 -149 -4296
rect -145 -4300 -64 -4296
rect 25 -4300 101 -4296
rect 115 -4300 146 -4296
rect 180 -4300 209 -4296
rect 213 -4300 294 -4296
rect 383 -4300 455 -4296
rect 469 -4300 502 -4296
rect 536 -4300 565 -4296
rect 569 -4300 650 -4296
rect 739 -4300 814 -4296
rect 828 -4300 860 -4296
rect 894 -4300 923 -4296
rect 927 -4300 1008 -4296
rect 1097 -4298 1164 -4294
rect 97 -4304 101 -4300
rect 451 -4304 455 -4300
rect 810 -4304 814 -4300
rect 1160 -4304 1164 -4298
rect 1171 -4300 1218 -4296
rect 1252 -4300 1281 -4296
rect 1285 -4300 1366 -4296
rect -1230 -4309 -1173 -4305
rect -1134 -4308 -902 -4304
rect -887 -4308 -804 -4304
rect -783 -4308 -687 -4304
rect -616 -4308 -544 -4304
rect -529 -4308 -446 -4304
rect -425 -4308 -328 -4304
rect -263 -4308 -186 -4304
rect -171 -4308 -88 -4304
rect -67 -4308 29 -4304
rect 97 -4308 172 -4304
rect 187 -4308 270 -4304
rect 291 -4308 388 -4304
rect 451 -4308 528 -4304
rect 543 -4308 626 -4304
rect 647 -4308 743 -4304
rect 810 -4308 886 -4304
rect 901 -4308 984 -4304
rect 1005 -4308 1101 -4304
rect 1160 -4308 1244 -4304
rect 1259 -4308 1342 -4304
rect 1363 -4308 1464 -4304
rect -1253 -4316 -1223 -4312
rect -1219 -4316 -1183 -4312
rect -1179 -4316 -1163 -4312
rect -959 -4315 -924 -4311
rect -905 -4315 -776 -4311
rect -612 -4315 -566 -4311
rect -547 -4315 -418 -4311
rect -259 -4315 -208 -4311
rect -189 -4315 -60 -4311
rect 101 -4315 150 -4311
rect 169 -4315 298 -4311
rect 455 -4315 506 -4311
rect 525 -4315 654 -4311
rect 814 -4315 864 -4311
rect 883 -4315 1012 -4311
rect 1188 -4315 1222 -4311
rect 1241 -4315 1370 -4311
rect -1279 -4323 -1227 -4319
rect -1223 -4323 -1197 -4319
rect -1193 -4323 -1149 -4319
rect -898 -4322 -794 -4318
rect -790 -4322 -760 -4318
rect -540 -4322 -436 -4318
rect -432 -4322 -402 -4318
rect -182 -4322 -78 -4318
rect -74 -4322 -44 -4318
rect 176 -4322 280 -4318
rect 284 -4322 314 -4318
rect 532 -4322 636 -4318
rect 640 -4322 670 -4318
rect 890 -4322 994 -4318
rect 998 -4322 1028 -4318
rect 1248 -4322 1352 -4318
rect 1356 -4322 1386 -4318
rect -1186 -4330 -1114 -4326
rect -924 -4329 -872 -4325
rect -868 -4329 -838 -4325
rect -566 -4329 -514 -4325
rect -510 -4329 -480 -4325
rect -208 -4329 -156 -4325
rect -152 -4329 -122 -4325
rect 150 -4329 202 -4325
rect 206 -4329 236 -4325
rect 506 -4329 558 -4325
rect 562 -4329 592 -4325
rect 864 -4329 916 -4325
rect 920 -4329 950 -4325
rect 1222 -4329 1274 -4325
rect 1278 -4329 1308 -4325
rect -1204 -4337 -1172 -4333
rect -879 -4337 -847 -4333
rect -883 -4340 -879 -4337
rect -847 -4340 -843 -4337
rect -801 -4337 -769 -4333
rect -805 -4340 -801 -4337
rect -769 -4340 -765 -4337
rect -521 -4337 -489 -4333
rect -525 -4340 -521 -4337
rect -489 -4340 -485 -4337
rect -443 -4337 -411 -4333
rect -447 -4340 -443 -4337
rect -411 -4340 -407 -4337
rect -163 -4337 -131 -4333
rect -167 -4340 -163 -4337
rect -131 -4340 -127 -4337
rect -85 -4337 -53 -4333
rect -89 -4340 -85 -4337
rect -53 -4340 -49 -4337
rect 195 -4337 227 -4333
rect 191 -4340 195 -4337
rect 227 -4340 231 -4337
rect 273 -4337 305 -4333
rect 269 -4340 273 -4337
rect 305 -4340 309 -4337
rect 551 -4337 583 -4333
rect 547 -4340 551 -4337
rect 583 -4340 587 -4337
rect 629 -4337 661 -4333
rect 625 -4340 629 -4337
rect 661 -4340 665 -4337
rect 909 -4337 941 -4333
rect 905 -4340 909 -4337
rect 941 -4340 945 -4337
rect 987 -4337 1019 -4333
rect 983 -4340 987 -4337
rect 1019 -4340 1023 -4337
rect 1267 -4337 1299 -4333
rect 1263 -4340 1267 -4337
rect 1299 -4340 1303 -4337
rect 1345 -4337 1377 -4333
rect 1341 -4340 1345 -4337
rect 1377 -4340 1381 -4337
rect -926 -4348 -922 -4344
rect -900 -4348 -896 -4344
rect -857 -4348 -853 -4344
rect -822 -4348 -818 -4344
rect -778 -4348 -774 -4344
rect -761 -4348 -757 -4344
rect -725 -4348 -721 -4344
rect -704 -4348 -700 -4344
rect -568 -4348 -564 -4344
rect -542 -4348 -538 -4344
rect -499 -4348 -495 -4344
rect -464 -4348 -460 -4344
rect -420 -4348 -416 -4344
rect -403 -4348 -399 -4344
rect -367 -4348 -363 -4344
rect -346 -4348 -342 -4344
rect -210 -4348 -206 -4344
rect -184 -4348 -180 -4344
rect -141 -4348 -137 -4344
rect -106 -4348 -102 -4344
rect -62 -4348 -58 -4344
rect -45 -4348 -41 -4344
rect -9 -4348 -5 -4344
rect 12 -4348 16 -4344
rect 148 -4348 152 -4344
rect 174 -4348 178 -4344
rect 217 -4348 221 -4344
rect 252 -4348 256 -4344
rect 296 -4348 300 -4344
rect 313 -4348 317 -4344
rect 349 -4348 353 -4344
rect 370 -4348 374 -4344
rect 504 -4348 508 -4344
rect 530 -4348 534 -4344
rect 573 -4348 577 -4344
rect 608 -4348 612 -4344
rect 652 -4348 656 -4344
rect 669 -4348 673 -4344
rect 705 -4348 709 -4344
rect 726 -4348 730 -4344
rect 862 -4348 866 -4344
rect 888 -4348 892 -4344
rect 931 -4348 935 -4344
rect 966 -4348 970 -4344
rect 1010 -4348 1014 -4344
rect 1027 -4348 1031 -4344
rect 1063 -4348 1067 -4344
rect 1084 -4348 1088 -4344
rect 1220 -4348 1224 -4344
rect 1246 -4348 1250 -4344
rect 1289 -4348 1293 -4344
rect 1324 -4348 1328 -4344
rect 1368 -4348 1372 -4344
rect 1385 -4348 1389 -4344
rect 1421 -4348 1425 -4344
rect 1442 -4348 1446 -4344
rect 1804 -4348 1831 -4193
rect -1411 -4352 -1225 -4348
rect -1221 -4352 -1181 -4348
rect -1177 -4352 -1147 -4348
rect -1143 -4352 -926 -4348
rect -922 -4352 -900 -4348
rect -896 -4352 -857 -4348
rect -853 -4352 -822 -4348
rect -818 -4352 -778 -4348
rect -774 -4352 -761 -4348
rect -757 -4352 -725 -4348
rect -721 -4352 -704 -4348
rect -700 -4352 -568 -4348
rect -564 -4352 -542 -4348
rect -538 -4352 -499 -4348
rect -495 -4352 -464 -4348
rect -460 -4352 -420 -4348
rect -416 -4352 -403 -4348
rect -399 -4352 -367 -4348
rect -363 -4352 -346 -4348
rect -342 -4352 -210 -4348
rect -206 -4352 -184 -4348
rect -180 -4352 -141 -4348
rect -137 -4352 -106 -4348
rect -102 -4352 -62 -4348
rect -58 -4352 -45 -4348
rect -41 -4352 -9 -4348
rect -5 -4352 12 -4348
rect 16 -4352 148 -4348
rect 152 -4352 174 -4348
rect 178 -4352 217 -4348
rect 221 -4352 252 -4348
rect 256 -4352 296 -4348
rect 300 -4352 313 -4348
rect 317 -4352 349 -4348
rect 353 -4352 370 -4348
rect 374 -4352 504 -4348
rect 508 -4352 530 -4348
rect 534 -4352 573 -4348
rect 577 -4352 608 -4348
rect 612 -4352 652 -4348
rect 656 -4352 669 -4348
rect 673 -4352 705 -4348
rect 709 -4352 726 -4348
rect 730 -4352 862 -4348
rect 866 -4352 888 -4348
rect 892 -4352 931 -4348
rect 935 -4352 966 -4348
rect 970 -4352 1010 -4348
rect 1014 -4352 1027 -4348
rect 1031 -4352 1063 -4348
rect 1067 -4352 1084 -4348
rect 1088 -4352 1220 -4348
rect 1224 -4352 1246 -4348
rect 1250 -4352 1289 -4348
rect 1293 -4352 1324 -4348
rect 1328 -4352 1368 -4348
rect 1372 -4352 1385 -4348
rect 1389 -4352 1421 -4348
rect 1425 -4352 1442 -4348
rect 1446 -4352 1831 -4348
rect -1253 -4359 -687 -4355
rect -599 -4359 29 -4355
rect 115 -4359 743 -4355
rect 828 -4359 1464 -4355
rect -1242 -4366 -1114 -4362
rect -959 -4366 -328 -4362
rect -245 -4366 388 -4362
rect 469 -4366 1101 -4362
rect 1188 -4366 1451 -4362
rect -2056 -4383 -1805 -4379
rect -1801 -4383 -1788 -4379
rect -1784 -4383 -1768 -4379
rect -1764 -4383 -1747 -4379
rect -1743 -4383 -1726 -4379
rect -1722 -4383 -1705 -4379
rect -1701 -4383 -1684 -4379
rect -1680 -4383 -1663 -4379
rect -1659 -4383 -1642 -4379
rect -1638 -4383 -1622 -4379
rect -1618 -4383 -1542 -4379
rect -1538 -4383 -1525 -4379
rect -1521 -4383 -1505 -4379
rect -1501 -4383 -1484 -4379
rect -1480 -4383 -1463 -4379
rect -1459 -4383 -1442 -4379
rect -1438 -4383 -1421 -4379
rect -1417 -4383 -1400 -4379
rect -1396 -4383 -1379 -4379
rect -1375 -4383 -1359 -4379
rect -1355 -4383 -1225 -4379
rect -1221 -4383 -1208 -4379
rect -1204 -4383 -1188 -4379
rect -1184 -4383 -1167 -4379
rect -1163 -4383 -1146 -4379
rect -1142 -4383 -1125 -4379
rect -1121 -4383 -1104 -4379
rect -1100 -4383 -1083 -4379
rect -1079 -4383 -1062 -4379
rect -1058 -4383 -1042 -4379
rect -1038 -4383 -926 -4379
rect -922 -4383 -909 -4379
rect -905 -4383 -889 -4379
rect -885 -4383 -868 -4379
rect -864 -4383 -847 -4379
rect -843 -4383 -826 -4379
rect -822 -4383 -805 -4379
rect -801 -4383 -784 -4379
rect -780 -4383 -763 -4379
rect -759 -4383 -743 -4379
rect -739 -4383 -568 -4379
rect -564 -4383 -551 -4379
rect -547 -4383 -531 -4379
rect -527 -4383 -510 -4379
rect -506 -4383 -489 -4379
rect -485 -4383 -468 -4379
rect -464 -4383 -447 -4379
rect -443 -4383 -426 -4379
rect -422 -4383 -405 -4379
rect -401 -4383 -385 -4379
rect -381 -4383 1612 -4379
rect -2054 -4550 -2027 -4383
rect -1783 -4431 -1749 -4427
rect -1685 -4431 -1665 -4427
rect -1650 -4431 -1547 -4427
rect -1520 -4431 -1486 -4427
rect -1422 -4431 -1402 -4427
rect -1387 -4431 -1346 -4427
rect -1203 -4431 -1169 -4427
rect -1105 -4431 -1085 -4427
rect -1070 -4431 -931 -4427
rect -904 -4431 -870 -4427
rect -806 -4431 -786 -4427
rect -771 -4431 -573 -4427
rect -546 -4431 -512 -4427
rect -448 -4431 -428 -4427
rect -413 -4431 -377 -4427
rect -1551 -4435 -1547 -4431
rect -935 -4435 -931 -4431
rect -577 -4435 -573 -4431
rect -1818 -4439 -1807 -4435
rect -1803 -4439 -1773 -4435
rect -1752 -4439 -1721 -4435
rect -1692 -4439 -1661 -4435
rect -1650 -4439 -1623 -4435
rect -1551 -4439 -1544 -4435
rect -1540 -4439 -1510 -4435
rect -1489 -4439 -1458 -4435
rect -1429 -4439 -1398 -4435
rect -1387 -4439 -1360 -4435
rect -1242 -4439 -1227 -4435
rect -1223 -4439 -1193 -4435
rect -1172 -4439 -1141 -4435
rect -1112 -4439 -1081 -4435
rect -1070 -4439 -1043 -4435
rect -935 -4439 -928 -4435
rect -924 -4439 -894 -4435
rect -873 -4439 -842 -4435
rect -813 -4439 -782 -4435
rect -771 -4439 -744 -4435
rect -577 -4439 -570 -4435
rect -566 -4439 -536 -4435
rect -515 -4439 -484 -4435
rect -455 -4439 -424 -4435
rect -413 -4439 -386 -4435
rect -1810 -4446 -1763 -4442
rect -1727 -4446 -1714 -4442
rect -1710 -4446 -1679 -4442
rect -1643 -4446 -1630 -4442
rect -1626 -4446 -1614 -4442
rect -1547 -4446 -1500 -4442
rect -1464 -4446 -1451 -4442
rect -1447 -4446 -1416 -4442
rect -1380 -4446 -1367 -4442
rect -1363 -4446 -1351 -4442
rect -1230 -4446 -1183 -4442
rect -1147 -4446 -1134 -4442
rect -1130 -4446 -1099 -4442
rect -1063 -4446 -1050 -4442
rect -1046 -4446 -1034 -4442
rect -931 -4446 -884 -4442
rect -848 -4446 -835 -4442
rect -831 -4446 -800 -4442
rect -764 -4446 -751 -4442
rect -747 -4446 -735 -4442
rect -573 -4446 -526 -4442
rect -490 -4446 -477 -4442
rect -473 -4446 -442 -4442
rect -406 -4446 -393 -4442
rect -389 -4446 -377 -4442
rect -1818 -4453 -1803 -4449
rect -1799 -4453 -1689 -4449
rect -1668 -4453 -1637 -4449
rect -1555 -4453 -1540 -4449
rect -1536 -4453 -1426 -4449
rect -1405 -4453 -1374 -4449
rect -1238 -4453 -1223 -4449
rect -1219 -4453 -1109 -4449
rect -1088 -4453 -1057 -4449
rect -939 -4453 -924 -4449
rect -920 -4453 -810 -4449
rect -789 -4453 -758 -4449
rect -581 -4453 -566 -4449
rect -562 -4453 -452 -4449
rect -431 -4453 -400 -4449
rect -1768 -4460 -1745 -4456
rect -1726 -4460 -1707 -4456
rect -1505 -4460 -1482 -4456
rect -1463 -4460 -1444 -4456
rect -1188 -4460 -1165 -4456
rect -1146 -4460 -1127 -4456
rect -889 -4460 -866 -4456
rect -847 -4460 -828 -4456
rect -531 -4460 -508 -4456
rect -489 -4460 -470 -4456
rect 1804 -4471 1831 -4352
rect -1954 -4475 -1805 -4471
rect -1801 -4475 -1788 -4471
rect -1784 -4475 -1747 -4471
rect -1743 -4475 -1705 -4471
rect -1701 -4475 -1663 -4471
rect -1659 -4475 -1622 -4471
rect -1618 -4475 -1542 -4471
rect -1538 -4475 -1525 -4471
rect -1521 -4475 -1484 -4471
rect -1480 -4475 -1442 -4471
rect -1438 -4475 -1400 -4471
rect -1396 -4475 -1359 -4471
rect -1355 -4475 -1225 -4471
rect -1221 -4475 -1208 -4471
rect -1204 -4475 -1167 -4471
rect -1163 -4475 -1125 -4471
rect -1121 -4475 -1083 -4471
rect -1079 -4475 -1042 -4471
rect -1038 -4475 -926 -4471
rect -922 -4475 -909 -4471
rect -905 -4475 -868 -4471
rect -864 -4475 -826 -4471
rect -822 -4475 -784 -4471
rect -780 -4475 -743 -4471
rect -739 -4475 -568 -4471
rect -564 -4475 -551 -4471
rect -547 -4475 -510 -4471
rect -506 -4475 -468 -4471
rect -464 -4475 -426 -4471
rect -422 -4475 -385 -4471
rect -381 -4475 1831 -4471
rect -1827 -4482 -1346 -4478
rect -2054 -4554 -1805 -4550
rect -1801 -4554 -1788 -4550
rect -1784 -4554 -1768 -4550
rect -1764 -4554 -1747 -4550
rect -1743 -4554 -1726 -4550
rect -1722 -4554 -1705 -4550
rect -1701 -4554 -1684 -4550
rect -1680 -4554 -1663 -4550
rect -1659 -4554 -1642 -4550
rect -1638 -4554 -1622 -4550
rect -1618 -4554 -1542 -4550
rect -1538 -4554 -1525 -4550
rect -1521 -4554 -1505 -4550
rect -1501 -4554 -1484 -4550
rect -1480 -4554 -1463 -4550
rect -1459 -4554 -1442 -4550
rect -1438 -4554 -1421 -4550
rect -1417 -4554 -1400 -4550
rect -1396 -4554 -1379 -4550
rect -1375 -4554 -1359 -4550
rect -1355 -4554 -1225 -4550
rect -1221 -4554 -1208 -4550
rect -1204 -4554 -1188 -4550
rect -1184 -4554 -1167 -4550
rect -1163 -4554 -1146 -4550
rect -1142 -4554 -1125 -4550
rect -1121 -4554 -1104 -4550
rect -1100 -4554 -1083 -4550
rect -1079 -4554 -1062 -4550
rect -1058 -4554 -1042 -4550
rect -1038 -4554 -926 -4550
rect -922 -4554 -909 -4550
rect -905 -4554 -889 -4550
rect -885 -4554 -868 -4550
rect -864 -4554 -847 -4550
rect -843 -4554 -826 -4550
rect -822 -4554 -805 -4550
rect -801 -4554 -784 -4550
rect -780 -4554 -763 -4550
rect -759 -4554 -743 -4550
rect -739 -4554 -568 -4550
rect -564 -4554 -551 -4550
rect -547 -4554 -531 -4550
rect -527 -4554 -510 -4550
rect -506 -4554 -489 -4550
rect -485 -4554 -468 -4550
rect -464 -4554 -447 -4550
rect -443 -4554 -426 -4550
rect -422 -4554 -405 -4550
rect -401 -4554 -385 -4550
rect -381 -4554 -210 -4550
rect -206 -4554 -193 -4550
rect -189 -4554 -173 -4550
rect -169 -4554 -152 -4550
rect -148 -4554 -131 -4550
rect -127 -4554 -110 -4550
rect -106 -4554 -89 -4550
rect -85 -4554 -68 -4550
rect -64 -4554 -47 -4550
rect -43 -4554 -27 -4550
rect -23 -4554 148 -4550
rect 152 -4554 165 -4550
rect 169 -4554 185 -4550
rect 189 -4554 206 -4550
rect 210 -4554 227 -4550
rect 231 -4554 248 -4550
rect 252 -4554 269 -4550
rect 273 -4554 290 -4550
rect 294 -4554 311 -4550
rect 315 -4554 331 -4550
rect 335 -4554 504 -4550
rect 508 -4554 521 -4550
rect 525 -4554 541 -4550
rect 545 -4554 562 -4550
rect 566 -4554 583 -4550
rect 587 -4554 604 -4550
rect 608 -4554 625 -4550
rect 629 -4554 646 -4550
rect 650 -4554 667 -4550
rect 671 -4554 687 -4550
rect 691 -4554 862 -4550
rect 866 -4554 879 -4550
rect 883 -4554 899 -4550
rect 903 -4554 920 -4550
rect 924 -4554 941 -4550
rect 945 -4554 962 -4550
rect 966 -4554 983 -4550
rect 987 -4554 1004 -4550
rect 1008 -4554 1025 -4550
rect 1029 -4554 1045 -4550
rect 1049 -4554 1220 -4550
rect 1224 -4554 1237 -4550
rect 1241 -4554 1257 -4550
rect 1261 -4554 1278 -4550
rect 1282 -4554 1299 -4550
rect 1303 -4554 1320 -4550
rect 1324 -4554 1341 -4550
rect 1345 -4554 1362 -4550
rect 1366 -4554 1383 -4550
rect 1387 -4554 1403 -4550
rect 1407 -4554 1613 -4550
rect -2054 -4721 -2027 -4554
rect -1783 -4602 -1749 -4598
rect -1685 -4602 -1665 -4598
rect -1650 -4602 -1547 -4598
rect -1520 -4602 -1486 -4598
rect -1422 -4602 -1402 -4598
rect -1387 -4602 -1347 -4598
rect -1203 -4602 -1169 -4598
rect -1105 -4602 -1085 -4598
rect -1070 -4602 -1023 -4598
rect -904 -4602 -870 -4598
rect -806 -4602 -786 -4598
rect -771 -4602 -729 -4598
rect -546 -4602 -512 -4598
rect -448 -4602 -428 -4598
rect -413 -4602 -370 -4598
rect -188 -4602 -154 -4598
rect -90 -4602 -70 -4598
rect -55 -4602 -9 -4598
rect 170 -4602 204 -4598
rect 268 -4602 288 -4598
rect 303 -4602 348 -4598
rect 526 -4602 560 -4598
rect 624 -4602 644 -4598
rect 659 -4602 700 -4598
rect 884 -4602 918 -4598
rect 982 -4602 1002 -4598
rect 1017 -4602 1059 -4598
rect 1242 -4602 1276 -4598
rect 1340 -4602 1360 -4598
rect 1375 -4602 1419 -4598
rect -1551 -4606 -1547 -4602
rect -1827 -4610 -1807 -4606
rect -1803 -4610 -1773 -4606
rect -1752 -4610 -1721 -4606
rect -1692 -4610 -1661 -4606
rect -1650 -4610 -1623 -4606
rect -1551 -4610 -1544 -4606
rect -1540 -4610 -1510 -4606
rect -1489 -4610 -1458 -4606
rect -1429 -4610 -1398 -4606
rect -1387 -4610 -1360 -4606
rect -1253 -4610 -1227 -4606
rect -1223 -4610 -1193 -4606
rect -1172 -4610 -1141 -4606
rect -1112 -4610 -1081 -4606
rect -1070 -4610 -1043 -4606
rect -959 -4610 -928 -4606
rect -924 -4610 -894 -4606
rect -873 -4610 -842 -4606
rect -813 -4610 -782 -4606
rect -771 -4610 -744 -4606
rect -599 -4610 -570 -4606
rect -566 -4610 -536 -4606
rect -515 -4610 -484 -4606
rect -455 -4610 -424 -4606
rect -413 -4610 -386 -4606
rect -245 -4610 -212 -4606
rect -208 -4610 -178 -4606
rect -157 -4610 -126 -4606
rect -97 -4610 -66 -4606
rect -55 -4610 -28 -4606
rect 115 -4610 146 -4606
rect 150 -4610 180 -4606
rect 201 -4610 232 -4606
rect 261 -4610 292 -4606
rect 303 -4610 330 -4606
rect 469 -4610 502 -4606
rect 506 -4610 536 -4606
rect 557 -4610 588 -4606
rect 617 -4610 648 -4606
rect 659 -4610 686 -4606
rect 828 -4610 860 -4606
rect 864 -4610 894 -4606
rect 915 -4610 946 -4606
rect 975 -4610 1006 -4606
rect 1017 -4610 1044 -4606
rect 1188 -4610 1218 -4606
rect 1222 -4610 1252 -4606
rect 1273 -4610 1304 -4606
rect 1333 -4610 1364 -4606
rect 1375 -4610 1402 -4606
rect -1810 -4617 -1763 -4613
rect -1727 -4617 -1714 -4613
rect -1710 -4617 -1679 -4613
rect -1643 -4617 -1630 -4613
rect -1626 -4617 -1614 -4613
rect -1547 -4617 -1500 -4613
rect -1464 -4617 -1451 -4613
rect -1447 -4617 -1416 -4613
rect -1380 -4617 -1367 -4613
rect -1363 -4617 -1351 -4613
rect -1230 -4617 -1183 -4613
rect -1147 -4617 -1134 -4613
rect -1130 -4617 -1099 -4613
rect -1063 -4617 -1050 -4613
rect -1046 -4617 -1034 -4613
rect -931 -4617 -884 -4613
rect -848 -4617 -835 -4613
rect -831 -4617 -800 -4613
rect -764 -4617 -751 -4613
rect -747 -4617 -735 -4613
rect -573 -4617 -526 -4613
rect -490 -4617 -477 -4613
rect -473 -4617 -442 -4613
rect -406 -4617 -393 -4613
rect -389 -4617 -377 -4613
rect -215 -4617 -168 -4613
rect -132 -4617 -119 -4613
rect -115 -4617 -84 -4613
rect -48 -4617 -35 -4613
rect -31 -4617 -19 -4613
rect 143 -4617 190 -4613
rect 226 -4617 239 -4613
rect 243 -4617 274 -4613
rect 310 -4617 323 -4613
rect 327 -4617 339 -4613
rect 499 -4617 546 -4613
rect 582 -4617 595 -4613
rect 599 -4617 630 -4613
rect 666 -4617 679 -4613
rect 683 -4617 695 -4613
rect 857 -4617 904 -4613
rect 940 -4617 953 -4613
rect 957 -4617 988 -4613
rect 1024 -4617 1037 -4613
rect 1041 -4617 1053 -4613
rect 1215 -4617 1262 -4613
rect 1298 -4617 1311 -4613
rect 1315 -4617 1346 -4613
rect 1382 -4617 1395 -4613
rect 1399 -4617 1411 -4613
rect -1818 -4624 -1803 -4620
rect -1799 -4624 -1689 -4620
rect -1668 -4624 -1637 -4620
rect -1555 -4624 -1540 -4620
rect -1536 -4624 -1426 -4620
rect -1405 -4624 -1374 -4620
rect -1238 -4624 -1223 -4620
rect -1219 -4624 -1109 -4620
rect -1088 -4624 -1057 -4620
rect -939 -4624 -924 -4620
rect -920 -4624 -810 -4620
rect -789 -4624 -758 -4620
rect -581 -4624 -566 -4620
rect -562 -4624 -452 -4620
rect -431 -4624 -400 -4620
rect -223 -4624 -208 -4620
rect -204 -4624 -94 -4620
rect -73 -4624 -42 -4620
rect 135 -4624 150 -4620
rect 154 -4624 264 -4620
rect 285 -4624 316 -4620
rect 491 -4624 506 -4620
rect 510 -4624 620 -4620
rect 641 -4624 672 -4620
rect 849 -4624 864 -4620
rect 868 -4624 978 -4620
rect 999 -4624 1030 -4620
rect 1207 -4624 1222 -4620
rect 1226 -4624 1336 -4620
rect 1357 -4624 1388 -4620
rect -1768 -4631 -1745 -4627
rect -1726 -4631 -1707 -4627
rect -1505 -4631 -1482 -4627
rect -1463 -4631 -1444 -4627
rect -1188 -4631 -1165 -4627
rect -1146 -4631 -1127 -4627
rect -889 -4631 -866 -4627
rect -847 -4631 -828 -4627
rect -531 -4631 -508 -4627
rect -489 -4631 -470 -4627
rect -173 -4631 -150 -4627
rect -131 -4631 -112 -4627
rect 185 -4631 208 -4627
rect 227 -4631 246 -4627
rect 541 -4631 564 -4627
rect 583 -4631 602 -4627
rect 899 -4631 922 -4627
rect 941 -4631 960 -4627
rect 1257 -4631 1280 -4627
rect 1299 -4631 1318 -4627
rect 1804 -4642 1831 -4475
rect -1972 -4646 -1805 -4642
rect -1801 -4646 -1788 -4642
rect -1784 -4646 -1747 -4642
rect -1743 -4646 -1705 -4642
rect -1701 -4646 -1663 -4642
rect -1659 -4646 -1622 -4642
rect -1618 -4646 -1542 -4642
rect -1538 -4646 -1525 -4642
rect -1521 -4646 -1484 -4642
rect -1480 -4646 -1442 -4642
rect -1438 -4646 -1400 -4642
rect -1396 -4646 -1359 -4642
rect -1355 -4646 -1225 -4642
rect -1221 -4646 -1208 -4642
rect -1204 -4646 -1167 -4642
rect -1163 -4646 -1125 -4642
rect -1121 -4646 -1083 -4642
rect -1079 -4646 -1042 -4642
rect -1038 -4646 -926 -4642
rect -922 -4646 -909 -4642
rect -905 -4646 -868 -4642
rect -864 -4646 -826 -4642
rect -822 -4646 -784 -4642
rect -780 -4646 -743 -4642
rect -739 -4646 -568 -4642
rect -564 -4646 -551 -4642
rect -547 -4646 -510 -4642
rect -506 -4646 -468 -4642
rect -464 -4646 -426 -4642
rect -422 -4646 -385 -4642
rect -381 -4646 -210 -4642
rect -206 -4646 -193 -4642
rect -189 -4646 -152 -4642
rect -148 -4646 -110 -4642
rect -106 -4646 -68 -4642
rect -64 -4646 -27 -4642
rect -23 -4646 148 -4642
rect 152 -4646 165 -4642
rect 169 -4646 206 -4642
rect 210 -4646 248 -4642
rect 252 -4646 290 -4642
rect 294 -4646 331 -4642
rect 335 -4646 504 -4642
rect 508 -4646 521 -4642
rect 525 -4646 562 -4642
rect 566 -4646 604 -4642
rect 608 -4646 646 -4642
rect 650 -4646 687 -4642
rect 691 -4646 862 -4642
rect 866 -4646 879 -4642
rect 883 -4646 920 -4642
rect 924 -4646 962 -4642
rect 966 -4646 1004 -4642
rect 1008 -4646 1045 -4642
rect 1049 -4646 1220 -4642
rect 1224 -4646 1237 -4642
rect 1241 -4646 1278 -4642
rect 1282 -4646 1320 -4642
rect 1324 -4646 1362 -4642
rect 1366 -4646 1403 -4642
rect 1407 -4646 1831 -4642
rect -1562 -4654 -1347 -4650
rect -1253 -4654 -1023 -4650
rect -959 -4653 -729 -4649
rect -599 -4653 -370 -4649
rect -245 -4653 -9 -4649
rect 115 -4655 348 -4651
rect 469 -4654 700 -4650
rect 828 -4653 1059 -4649
rect 1188 -4653 1419 -4649
rect -2054 -4725 -1542 -4721
rect -1538 -4725 -1525 -4721
rect -1521 -4725 -1505 -4721
rect -1501 -4725 -1484 -4721
rect -1480 -4725 -1463 -4721
rect -1459 -4725 -1442 -4721
rect -1438 -4725 -1421 -4721
rect -1417 -4725 -1400 -4721
rect -1396 -4725 -1379 -4721
rect -1375 -4725 -1359 -4721
rect -1355 -4725 -1225 -4721
rect -1221 -4725 -1208 -4721
rect -1204 -4725 -1188 -4721
rect -1184 -4725 -1167 -4721
rect -1163 -4725 -1146 -4721
rect -1142 -4725 -1125 -4721
rect -1121 -4725 -1104 -4721
rect -1100 -4725 -1083 -4721
rect -1079 -4725 -1062 -4721
rect -1058 -4725 -1042 -4721
rect -1038 -4725 -926 -4721
rect -922 -4725 -909 -4721
rect -905 -4725 -889 -4721
rect -885 -4725 -868 -4721
rect -864 -4725 -847 -4721
rect -843 -4725 -826 -4721
rect -822 -4725 -805 -4721
rect -801 -4725 -784 -4721
rect -780 -4725 -763 -4721
rect -759 -4725 -743 -4721
rect -739 -4725 -568 -4721
rect -564 -4725 -551 -4721
rect -547 -4725 -531 -4721
rect -527 -4725 -510 -4721
rect -506 -4725 -489 -4721
rect -485 -4725 -468 -4721
rect -464 -4725 -447 -4721
rect -443 -4725 -426 -4721
rect -422 -4725 -405 -4721
rect -401 -4725 -385 -4721
rect -381 -4725 -210 -4721
rect -206 -4725 -193 -4721
rect -189 -4725 -173 -4721
rect -169 -4725 -152 -4721
rect -148 -4725 -131 -4721
rect -127 -4725 -110 -4721
rect -106 -4725 -89 -4721
rect -85 -4725 -68 -4721
rect -64 -4725 -47 -4721
rect -43 -4725 -27 -4721
rect -23 -4725 148 -4721
rect 152 -4725 165 -4721
rect 169 -4725 185 -4721
rect 189 -4725 206 -4721
rect 210 -4725 227 -4721
rect 231 -4725 248 -4721
rect 252 -4725 269 -4721
rect 273 -4725 290 -4721
rect 294 -4725 311 -4721
rect 315 -4725 331 -4721
rect 335 -4725 504 -4721
rect 508 -4725 521 -4721
rect 525 -4725 541 -4721
rect 545 -4725 562 -4721
rect 566 -4725 583 -4721
rect 587 -4725 604 -4721
rect 608 -4725 625 -4721
rect 629 -4725 646 -4721
rect 650 -4725 667 -4721
rect 671 -4725 687 -4721
rect 691 -4725 862 -4721
rect 866 -4725 879 -4721
rect 883 -4725 899 -4721
rect 903 -4725 920 -4721
rect 924 -4725 941 -4721
rect 945 -4725 962 -4721
rect 966 -4725 983 -4721
rect 987 -4725 1004 -4721
rect 1008 -4725 1025 -4721
rect 1029 -4725 1045 -4721
rect 1049 -4725 1220 -4721
rect 1224 -4725 1237 -4721
rect 1241 -4725 1257 -4721
rect 1261 -4725 1278 -4721
rect 1282 -4725 1299 -4721
rect 1303 -4725 1320 -4721
rect 1324 -4725 1341 -4721
rect 1345 -4725 1362 -4721
rect 1366 -4725 1383 -4721
rect 1387 -4725 1403 -4721
rect 1407 -4725 1649 -4721
rect -2054 -4836 -2027 -4725
rect -1520 -4773 -1486 -4769
rect -1422 -4773 -1402 -4769
rect -1387 -4773 -1346 -4769
rect -1203 -4773 -1169 -4769
rect -1105 -4773 -1085 -4769
rect -1070 -4773 -1022 -4769
rect -904 -4773 -870 -4769
rect -806 -4773 -786 -4769
rect -771 -4773 -722 -4769
rect -546 -4773 -512 -4769
rect -448 -4773 -428 -4769
rect -413 -4773 -369 -4769
rect -188 -4773 -154 -4769
rect -90 -4773 -70 -4769
rect -55 -4773 -11 -4769
rect 170 -4773 204 -4769
rect 268 -4773 288 -4769
rect 303 -4773 347 -4769
rect 526 -4773 560 -4769
rect 624 -4773 644 -4769
rect 659 -4773 706 -4769
rect 884 -4773 918 -4769
rect 982 -4773 1002 -4769
rect 1017 -4773 1062 -4769
rect 1242 -4773 1276 -4769
rect 1340 -4773 1360 -4769
rect 1375 -4773 1420 -4769
rect -1562 -4781 -1544 -4777
rect -1540 -4781 -1510 -4777
rect -1489 -4781 -1458 -4777
rect -1429 -4781 -1398 -4777
rect -1387 -4781 -1360 -4777
rect -1315 -4781 -1227 -4777
rect -1223 -4781 -1193 -4777
rect -1172 -4781 -1141 -4777
rect -1112 -4781 -1081 -4777
rect -1070 -4781 -1043 -4777
rect -945 -4781 -928 -4777
rect -924 -4781 -894 -4777
rect -873 -4781 -842 -4777
rect -813 -4781 -782 -4777
rect -771 -4781 -744 -4777
rect -587 -4781 -570 -4777
rect -566 -4781 -536 -4777
rect -515 -4781 -484 -4777
rect -455 -4781 -424 -4777
rect -413 -4781 -386 -4777
rect -229 -4781 -212 -4777
rect -208 -4781 -178 -4777
rect -157 -4781 -126 -4777
rect -97 -4781 -66 -4777
rect -55 -4781 -28 -4777
rect 129 -4781 146 -4777
rect 150 -4781 180 -4777
rect 201 -4781 232 -4777
rect 261 -4781 292 -4777
rect 303 -4781 330 -4777
rect 485 -4781 502 -4777
rect 506 -4781 536 -4777
rect 557 -4781 588 -4777
rect 617 -4781 648 -4777
rect 659 -4781 686 -4777
rect 843 -4781 860 -4777
rect 864 -4781 894 -4777
rect 915 -4781 946 -4777
rect 975 -4781 1006 -4777
rect 1017 -4781 1044 -4777
rect 1201 -4781 1218 -4777
rect 1222 -4781 1252 -4777
rect 1273 -4781 1304 -4777
rect 1333 -4781 1364 -4777
rect 1375 -4781 1402 -4777
rect -1547 -4788 -1500 -4784
rect -1464 -4788 -1451 -4784
rect -1447 -4788 -1416 -4784
rect -1380 -4788 -1367 -4784
rect -1363 -4788 -1351 -4784
rect -1230 -4788 -1183 -4784
rect -1147 -4788 -1134 -4784
rect -1130 -4788 -1099 -4784
rect -1063 -4788 -1050 -4784
rect -1046 -4788 -1034 -4784
rect -931 -4788 -884 -4784
rect -848 -4788 -835 -4784
rect -831 -4788 -800 -4784
rect -764 -4788 -751 -4784
rect -747 -4788 -735 -4784
rect -573 -4788 -526 -4784
rect -490 -4788 -477 -4784
rect -473 -4788 -442 -4784
rect -406 -4788 -393 -4784
rect -389 -4788 -377 -4784
rect -215 -4788 -168 -4784
rect -132 -4788 -119 -4784
rect -115 -4788 -84 -4784
rect -48 -4788 -35 -4784
rect -31 -4788 -19 -4784
rect 143 -4788 190 -4784
rect 226 -4788 239 -4784
rect 243 -4788 274 -4784
rect 310 -4788 323 -4784
rect 327 -4788 339 -4784
rect 499 -4788 546 -4784
rect 582 -4788 595 -4784
rect 599 -4788 630 -4784
rect 666 -4788 679 -4784
rect 683 -4788 695 -4784
rect 857 -4788 904 -4784
rect 940 -4788 953 -4784
rect 957 -4788 988 -4784
rect 1024 -4788 1037 -4784
rect 1041 -4788 1053 -4784
rect 1215 -4788 1262 -4784
rect 1298 -4788 1311 -4784
rect 1315 -4788 1346 -4784
rect 1382 -4788 1395 -4784
rect 1399 -4788 1411 -4784
rect -1555 -4795 -1540 -4791
rect -1536 -4795 -1426 -4791
rect -1405 -4795 -1374 -4791
rect -1238 -4795 -1223 -4791
rect -1219 -4795 -1109 -4791
rect -1088 -4795 -1057 -4791
rect -939 -4795 -924 -4791
rect -920 -4795 -810 -4791
rect -789 -4795 -758 -4791
rect -581 -4795 -566 -4791
rect -562 -4795 -452 -4791
rect -431 -4795 -400 -4791
rect -223 -4795 -208 -4791
rect -204 -4795 -94 -4791
rect -73 -4795 -42 -4791
rect 135 -4795 150 -4791
rect 154 -4795 264 -4791
rect 285 -4795 316 -4791
rect 491 -4795 506 -4791
rect 510 -4795 620 -4791
rect 641 -4795 672 -4791
rect 849 -4795 864 -4791
rect 868 -4795 978 -4791
rect 999 -4795 1030 -4791
rect 1207 -4795 1222 -4791
rect 1226 -4795 1336 -4791
rect 1357 -4795 1388 -4791
rect -1505 -4802 -1482 -4798
rect -1463 -4802 -1444 -4798
rect -1188 -4802 -1165 -4798
rect -1146 -4802 -1127 -4798
rect -889 -4802 -866 -4798
rect -847 -4802 -828 -4798
rect -531 -4802 -508 -4798
rect -489 -4802 -470 -4798
rect -173 -4802 -150 -4798
rect -131 -4802 -112 -4798
rect 185 -4802 208 -4798
rect 227 -4802 246 -4798
rect 541 -4802 564 -4798
rect 583 -4802 602 -4798
rect 899 -4802 922 -4798
rect 941 -4802 960 -4798
rect 1257 -4802 1280 -4798
rect 1299 -4802 1318 -4798
rect 1804 -4813 1831 -4646
rect -1642 -4817 -1542 -4813
rect -1538 -4817 -1525 -4813
rect -1521 -4817 -1484 -4813
rect -1480 -4817 -1442 -4813
rect -1438 -4817 -1400 -4813
rect -1396 -4817 -1359 -4813
rect -1355 -4817 -1225 -4813
rect -1221 -4817 -1208 -4813
rect -1204 -4817 -1167 -4813
rect -1163 -4817 -1125 -4813
rect -1121 -4817 -1083 -4813
rect -1079 -4817 -1042 -4813
rect -1038 -4817 -926 -4813
rect -922 -4817 -909 -4813
rect -905 -4817 -868 -4813
rect -864 -4817 -826 -4813
rect -822 -4817 -784 -4813
rect -780 -4817 -743 -4813
rect -739 -4817 -568 -4813
rect -564 -4817 -551 -4813
rect -547 -4817 -510 -4813
rect -506 -4817 -468 -4813
rect -464 -4817 -426 -4813
rect -422 -4817 -385 -4813
rect -381 -4817 -210 -4813
rect -206 -4817 -193 -4813
rect -189 -4817 -152 -4813
rect -148 -4817 -110 -4813
rect -106 -4817 -68 -4813
rect -64 -4817 -27 -4813
rect -23 -4817 148 -4813
rect 152 -4817 165 -4813
rect 169 -4817 206 -4813
rect 210 -4817 248 -4813
rect 252 -4817 290 -4813
rect 294 -4817 331 -4813
rect 335 -4817 504 -4813
rect 508 -4817 521 -4813
rect 525 -4817 562 -4813
rect 566 -4817 604 -4813
rect 608 -4817 646 -4813
rect 650 -4817 687 -4813
rect 691 -4817 862 -4813
rect 866 -4817 879 -4813
rect 883 -4817 920 -4813
rect 924 -4817 962 -4813
rect 966 -4817 1004 -4813
rect 1008 -4817 1045 -4813
rect 1049 -4817 1220 -4813
rect 1224 -4817 1237 -4813
rect 1241 -4817 1278 -4813
rect 1282 -4817 1320 -4813
rect 1324 -4817 1362 -4813
rect 1366 -4817 1403 -4813
rect 1407 -4817 1831 -4813
rect -2054 -4840 -1309 -4836
rect -1305 -4840 -1292 -4836
rect -1288 -4840 -935 -4836
rect -931 -4840 -918 -4836
rect -914 -4840 -577 -4836
rect -573 -4840 -560 -4836
rect -556 -4840 -219 -4836
rect -215 -4840 -202 -4836
rect -198 -4840 139 -4836
rect 143 -4840 156 -4836
rect 160 -4840 495 -4836
rect 499 -4840 512 -4836
rect 516 -4840 853 -4836
rect 857 -4840 870 -4836
rect 874 -4840 1211 -4836
rect 1215 -4840 1228 -4836
rect 1232 -4840 1589 -4836
rect -2054 -4995 -2027 -4840
rect -1304 -4872 -1022 -4868
rect -930 -4872 -722 -4868
rect -572 -4872 -369 -4868
rect -214 -4872 -11 -4868
rect 144 -4872 347 -4868
rect 496 -4872 706 -4868
rect 858 -4872 1062 -4868
rect 1216 -4872 1420 -4868
rect -1342 -4880 -1297 -4876
rect -1293 -4880 -923 -4876
rect -919 -4880 -565 -4876
rect -561 -4880 -207 -4876
rect -203 -4880 151 -4876
rect 155 -4880 507 -4876
rect 511 -4880 865 -4876
rect 869 -4880 1223 -4876
rect 1227 -4880 1589 -4876
rect -975 -4893 -909 -4889
rect -612 -4893 -551 -4889
rect -259 -4893 -193 -4889
rect 101 -4893 165 -4889
rect 455 -4893 521 -4889
rect 814 -4893 879 -4889
rect 1171 -4893 1237 -4889
rect 1804 -4928 1831 -4817
rect -1411 -4932 -1292 -4928
rect -1288 -4932 -918 -4928
rect -914 -4932 -560 -4928
rect -556 -4932 -202 -4928
rect -198 -4932 156 -4928
rect 160 -4932 512 -4928
rect 516 -4932 870 -4928
rect 874 -4932 1228 -4928
rect 1232 -4932 1831 -4928
rect -2054 -4999 -1225 -4995
rect -1221 -4999 -1208 -4995
rect -1204 -4999 -1168 -4995
rect -1164 -4999 -1147 -4995
rect -1143 -4999 -926 -4995
rect -922 -4999 -900 -4995
rect -896 -4999 -883 -4995
rect -879 -4999 -843 -4995
rect -839 -4999 -822 -4995
rect -818 -4999 -805 -4995
rect -801 -4999 -765 -4995
rect -761 -4999 -741 -4995
rect -737 -4999 -704 -4995
rect -700 -4999 -568 -4995
rect -564 -4999 -542 -4995
rect -538 -4999 -525 -4995
rect -521 -4999 -485 -4995
rect -481 -4999 -464 -4995
rect -460 -4999 -447 -4995
rect -443 -4999 -407 -4995
rect -403 -4999 -383 -4995
rect -379 -4999 -346 -4995
rect -342 -4999 -210 -4995
rect -206 -4999 -184 -4995
rect -180 -4999 -167 -4995
rect -163 -4999 -127 -4995
rect -123 -4999 -106 -4995
rect -102 -4999 -89 -4995
rect -85 -4999 -49 -4995
rect -45 -4999 -25 -4995
rect -21 -4999 12 -4995
rect 16 -4999 148 -4995
rect 152 -4999 174 -4995
rect 178 -4999 191 -4995
rect 195 -4999 231 -4995
rect 235 -4999 252 -4995
rect 256 -4999 269 -4995
rect 273 -4999 309 -4995
rect 313 -4999 333 -4995
rect 337 -4999 370 -4995
rect 374 -4999 504 -4995
rect 508 -4999 530 -4995
rect 534 -4999 547 -4995
rect 551 -4999 587 -4995
rect 591 -4999 608 -4995
rect 612 -4999 625 -4995
rect 629 -4999 665 -4995
rect 669 -4999 689 -4995
rect 693 -4999 726 -4995
rect 730 -4999 862 -4995
rect 866 -4999 888 -4995
rect 892 -4999 905 -4995
rect 909 -4999 945 -4995
rect 949 -4999 966 -4995
rect 970 -4999 983 -4995
rect 987 -4999 1023 -4995
rect 1027 -4999 1047 -4995
rect 1051 -4999 1084 -4995
rect 1088 -4999 1220 -4995
rect 1224 -4999 1246 -4995
rect 1250 -4999 1263 -4995
rect 1267 -4999 1303 -4995
rect 1307 -4999 1324 -4995
rect 1328 -4999 1341 -4995
rect 1345 -4999 1381 -4995
rect 1385 -4999 1405 -4995
rect 1409 -4999 1442 -4995
rect 1446 -4999 1589 -4995
rect -2054 -5114 -2027 -4999
rect -926 -5003 -922 -4999
rect -900 -5003 -896 -4999
rect -883 -5003 -879 -4999
rect -843 -5003 -839 -4999
rect -822 -5003 -818 -4999
rect -805 -5003 -801 -4999
rect -765 -5003 -761 -4999
rect -741 -5003 -737 -4999
rect -704 -5003 -700 -4999
rect -568 -5003 -564 -4999
rect -542 -5003 -538 -4999
rect -525 -5003 -521 -4999
rect -485 -5003 -481 -4999
rect -464 -5003 -460 -4999
rect -447 -5003 -443 -4999
rect -407 -5003 -403 -4999
rect -383 -5003 -379 -4999
rect -346 -5003 -342 -4999
rect -210 -5003 -206 -4999
rect -184 -5003 -180 -4999
rect -167 -5003 -163 -4999
rect -127 -5003 -123 -4999
rect -106 -5003 -102 -4999
rect -89 -5003 -85 -4999
rect -49 -5003 -45 -4999
rect -25 -5003 -21 -4999
rect 12 -5003 16 -4999
rect 148 -5003 152 -4999
rect 174 -5003 178 -4999
rect 191 -5003 195 -4999
rect 231 -5003 235 -4999
rect 252 -5003 256 -4999
rect 269 -5003 273 -4999
rect 309 -5003 313 -4999
rect 333 -5003 337 -4999
rect 370 -5003 374 -4999
rect 504 -5003 508 -4999
rect 530 -5003 534 -4999
rect 547 -5003 551 -4999
rect 587 -5003 591 -4999
rect 608 -5003 612 -4999
rect 625 -5003 629 -4999
rect 665 -5003 669 -4999
rect 689 -5003 693 -4999
rect 726 -5003 730 -4999
rect 862 -5003 866 -4999
rect 888 -5003 892 -4999
rect 905 -5003 909 -4999
rect 945 -5003 949 -4999
rect 966 -5003 970 -4999
rect 983 -5003 987 -4999
rect 1023 -5003 1027 -4999
rect 1047 -5003 1051 -4999
rect 1084 -5003 1088 -4999
rect 1220 -5003 1224 -4999
rect 1246 -5003 1250 -4999
rect 1263 -5003 1267 -4999
rect 1303 -5003 1307 -4999
rect 1324 -5003 1328 -4999
rect 1341 -5003 1345 -4999
rect 1381 -5003 1385 -4999
rect 1405 -5003 1409 -4999
rect 1442 -5003 1446 -4999
rect -920 -5018 -858 -5014
rect -854 -5018 -824 -5014
rect -776 -5018 -746 -5014
rect -562 -5018 -500 -5014
rect -496 -5018 -466 -5014
rect -418 -5018 -388 -5014
rect -204 -5018 -142 -5014
rect -138 -5018 -108 -5014
rect -60 -5018 -30 -5014
rect 154 -5018 216 -5014
rect 220 -5018 250 -5014
rect 298 -5018 328 -5014
rect 510 -5018 572 -5014
rect 576 -5018 606 -5014
rect 654 -5018 684 -5014
rect 868 -5018 930 -5014
rect 934 -5018 964 -5014
rect 1012 -5018 1042 -5014
rect 1226 -5018 1288 -5014
rect 1292 -5018 1322 -5014
rect 1370 -5018 1400 -5014
rect -913 -5025 -882 -5021
rect -555 -5025 -524 -5021
rect -197 -5025 -166 -5021
rect 161 -5025 192 -5021
rect 517 -5025 548 -5021
rect 875 -5025 906 -5021
rect 1233 -5025 1264 -5021
rect -931 -5032 -848 -5028
rect -809 -5032 -706 -5028
rect -573 -5032 -490 -5028
rect -451 -5032 -348 -5028
rect -215 -5032 -132 -5028
rect -93 -5032 10 -5028
rect 143 -5032 226 -5028
rect 265 -5032 368 -5028
rect 499 -5032 582 -5028
rect 621 -5032 724 -5028
rect 857 -5032 940 -5028
rect 979 -5032 1082 -5028
rect 1215 -5032 1298 -5028
rect 1337 -5032 1440 -5028
rect -975 -5039 -928 -5035
rect -894 -5039 -865 -5035
rect -861 -5039 -780 -5035
rect -691 -5039 -612 -5035
rect -599 -5039 -570 -5035
rect -536 -5039 -507 -5035
rect -503 -5039 -422 -5035
rect -333 -5038 -259 -5034
rect -616 -5043 -612 -5039
rect -263 -5043 -259 -5038
rect -245 -5039 -212 -5035
rect -178 -5039 -149 -5035
rect -145 -5039 -64 -5035
rect 25 -5039 101 -5035
rect 115 -5039 146 -5035
rect 180 -5039 209 -5035
rect 213 -5039 294 -5035
rect 383 -5039 455 -5035
rect 469 -5039 502 -5035
rect 536 -5039 565 -5035
rect 569 -5039 650 -5035
rect 739 -5039 814 -5035
rect 828 -5039 860 -5035
rect 894 -5039 923 -5035
rect 927 -5039 1008 -5035
rect 1097 -5037 1164 -5033
rect 97 -5043 101 -5039
rect 451 -5043 455 -5039
rect 810 -5043 814 -5039
rect 1160 -5043 1164 -5037
rect 1171 -5039 1218 -5035
rect 1252 -5039 1281 -5035
rect 1285 -5039 1366 -5035
rect -1230 -5048 -1173 -5044
rect -1134 -5047 -902 -5043
rect -887 -5047 -804 -5043
rect -783 -5047 -687 -5043
rect -616 -5047 -544 -5043
rect -529 -5047 -446 -5043
rect -425 -5047 -328 -5043
rect -263 -5047 -186 -5043
rect -171 -5047 -88 -5043
rect -67 -5047 29 -5043
rect 97 -5047 172 -5043
rect 187 -5047 270 -5043
rect 291 -5047 388 -5043
rect 451 -5047 528 -5043
rect 543 -5047 626 -5043
rect 647 -5047 743 -5043
rect 810 -5047 886 -5043
rect 901 -5047 984 -5043
rect 1005 -5047 1101 -5043
rect 1160 -5047 1244 -5043
rect 1259 -5047 1342 -5043
rect 1363 -5047 1464 -5043
rect -1253 -5055 -1223 -5051
rect -1219 -5055 -1183 -5051
rect -1179 -5055 -1163 -5051
rect -959 -5054 -924 -5050
rect -905 -5054 -776 -5050
rect -612 -5054 -566 -5050
rect -547 -5054 -418 -5050
rect -259 -5054 -208 -5050
rect -189 -5054 -60 -5050
rect 101 -5054 150 -5050
rect 169 -5054 298 -5050
rect 455 -5054 506 -5050
rect 525 -5054 654 -5050
rect 814 -5054 864 -5050
rect 883 -5054 1012 -5050
rect 1188 -5054 1222 -5050
rect 1241 -5054 1370 -5050
rect -1279 -5062 -1227 -5058
rect -1223 -5062 -1197 -5058
rect -1193 -5062 -1149 -5058
rect -898 -5061 -794 -5057
rect -790 -5061 -760 -5057
rect -540 -5061 -436 -5057
rect -432 -5061 -402 -5057
rect -182 -5061 -78 -5057
rect -74 -5061 -44 -5057
rect 176 -5061 280 -5057
rect 284 -5061 314 -5057
rect 532 -5061 636 -5057
rect 640 -5061 670 -5057
rect 890 -5061 994 -5057
rect 998 -5061 1028 -5057
rect 1248 -5061 1352 -5057
rect 1356 -5061 1386 -5057
rect -1186 -5069 -1102 -5065
rect -924 -5068 -872 -5064
rect -868 -5068 -838 -5064
rect -566 -5068 -514 -5064
rect -510 -5068 -480 -5064
rect -208 -5068 -156 -5064
rect -152 -5068 -122 -5064
rect 150 -5068 202 -5064
rect 206 -5068 236 -5064
rect 506 -5068 558 -5064
rect 562 -5068 592 -5064
rect 864 -5068 916 -5064
rect 920 -5068 950 -5064
rect 1222 -5068 1274 -5064
rect 1278 -5068 1308 -5064
rect -1204 -5076 -1172 -5072
rect -879 -5076 -847 -5072
rect -883 -5079 -879 -5076
rect -847 -5079 -843 -5076
rect -801 -5076 -769 -5072
rect -805 -5079 -801 -5076
rect -769 -5079 -765 -5076
rect -521 -5076 -489 -5072
rect -525 -5079 -521 -5076
rect -489 -5079 -485 -5076
rect -443 -5076 -411 -5072
rect -447 -5079 -443 -5076
rect -411 -5079 -407 -5076
rect -163 -5076 -131 -5072
rect -167 -5079 -163 -5076
rect -131 -5079 -127 -5076
rect -85 -5076 -53 -5072
rect -89 -5079 -85 -5076
rect -53 -5079 -49 -5076
rect 195 -5076 227 -5072
rect 191 -5079 195 -5076
rect 227 -5079 231 -5076
rect 273 -5076 305 -5072
rect 269 -5079 273 -5076
rect 305 -5079 309 -5076
rect 551 -5076 583 -5072
rect 547 -5079 551 -5076
rect 583 -5079 587 -5076
rect 629 -5076 661 -5072
rect 625 -5079 629 -5076
rect 661 -5079 665 -5076
rect 909 -5076 941 -5072
rect 905 -5079 909 -5076
rect 941 -5079 945 -5076
rect 987 -5076 1019 -5072
rect 983 -5079 987 -5076
rect 1019 -5079 1023 -5076
rect 1267 -5076 1299 -5072
rect 1263 -5079 1267 -5076
rect 1299 -5079 1303 -5076
rect 1345 -5076 1377 -5072
rect 1341 -5079 1345 -5076
rect 1377 -5079 1381 -5076
rect -926 -5087 -922 -5083
rect -900 -5087 -896 -5083
rect -857 -5087 -853 -5083
rect -822 -5087 -818 -5083
rect -778 -5087 -774 -5083
rect -761 -5087 -757 -5083
rect -725 -5087 -721 -5083
rect -704 -5087 -700 -5083
rect -568 -5087 -564 -5083
rect -542 -5087 -538 -5083
rect -499 -5087 -495 -5083
rect -464 -5087 -460 -5083
rect -420 -5087 -416 -5083
rect -403 -5087 -399 -5083
rect -367 -5087 -363 -5083
rect -346 -5087 -342 -5083
rect -210 -5087 -206 -5083
rect -184 -5087 -180 -5083
rect -141 -5087 -137 -5083
rect -106 -5087 -102 -5083
rect -62 -5087 -58 -5083
rect -45 -5087 -41 -5083
rect -9 -5087 -5 -5083
rect 12 -5087 16 -5083
rect 148 -5087 152 -5083
rect 174 -5087 178 -5083
rect 217 -5087 221 -5083
rect 252 -5087 256 -5083
rect 296 -5087 300 -5083
rect 313 -5087 317 -5083
rect 349 -5087 353 -5083
rect 370 -5087 374 -5083
rect 504 -5087 508 -5083
rect 530 -5087 534 -5083
rect 573 -5087 577 -5083
rect 608 -5087 612 -5083
rect 652 -5087 656 -5083
rect 669 -5087 673 -5083
rect 705 -5087 709 -5083
rect 726 -5087 730 -5083
rect 862 -5087 866 -5083
rect 888 -5087 892 -5083
rect 931 -5087 935 -5083
rect 966 -5087 970 -5083
rect 1010 -5087 1014 -5083
rect 1027 -5087 1031 -5083
rect 1063 -5087 1067 -5083
rect 1084 -5087 1088 -5083
rect 1220 -5087 1224 -5083
rect 1246 -5087 1250 -5083
rect 1289 -5087 1293 -5083
rect 1324 -5087 1328 -5083
rect 1368 -5087 1372 -5083
rect 1385 -5087 1389 -5083
rect 1421 -5087 1425 -5083
rect 1442 -5087 1446 -5083
rect 1804 -5087 1831 -4932
rect -1411 -5091 -1225 -5087
rect -1221 -5091 -1181 -5087
rect -1177 -5091 -1147 -5087
rect -1143 -5091 -926 -5087
rect -922 -5091 -900 -5087
rect -896 -5091 -857 -5087
rect -853 -5091 -822 -5087
rect -818 -5091 -778 -5087
rect -774 -5091 -761 -5087
rect -757 -5091 -725 -5087
rect -721 -5091 -704 -5087
rect -700 -5091 -568 -5087
rect -564 -5091 -542 -5087
rect -538 -5091 -499 -5087
rect -495 -5091 -464 -5087
rect -460 -5091 -420 -5087
rect -416 -5091 -403 -5087
rect -399 -5091 -367 -5087
rect -363 -5091 -346 -5087
rect -342 -5091 -210 -5087
rect -206 -5091 -184 -5087
rect -180 -5091 -141 -5087
rect -137 -5091 -106 -5087
rect -102 -5091 -62 -5087
rect -58 -5091 -45 -5087
rect -41 -5091 -9 -5087
rect -5 -5091 12 -5087
rect 16 -5091 148 -5087
rect 152 -5091 174 -5087
rect 178 -5091 217 -5087
rect 221 -5091 252 -5087
rect 256 -5091 296 -5087
rect 300 -5091 313 -5087
rect 317 -5091 349 -5087
rect 353 -5091 370 -5087
rect 374 -5091 504 -5087
rect 508 -5091 530 -5087
rect 534 -5091 573 -5087
rect 577 -5091 608 -5087
rect 612 -5091 652 -5087
rect 656 -5091 669 -5087
rect 673 -5091 705 -5087
rect 709 -5091 726 -5087
rect 730 -5091 862 -5087
rect 866 -5091 888 -5087
rect 892 -5091 931 -5087
rect 935 -5091 966 -5087
rect 970 -5091 1010 -5087
rect 1014 -5091 1027 -5087
rect 1031 -5091 1063 -5087
rect 1067 -5091 1084 -5087
rect 1088 -5091 1220 -5087
rect 1224 -5091 1246 -5087
rect 1250 -5091 1289 -5087
rect 1293 -5091 1324 -5087
rect 1328 -5091 1368 -5087
rect 1372 -5091 1385 -5087
rect 1389 -5091 1421 -5087
rect 1425 -5091 1442 -5087
rect 1446 -5091 1831 -5087
rect -1253 -5098 -687 -5094
rect -599 -5098 29 -5094
rect 112 -5098 743 -5094
rect 826 -5098 1464 -5094
rect -1242 -5106 -1102 -5102
rect -959 -5105 -328 -5101
rect -245 -5105 388 -5101
rect 468 -5105 1101 -5101
rect 1181 -5105 1451 -5101
rect -2054 -5118 -1801 -5114
rect -1797 -5118 -1784 -5114
rect -1780 -5118 -1764 -5114
rect -1760 -5118 -1743 -5114
rect -1739 -5118 -1722 -5114
rect -1718 -5118 -1701 -5114
rect -1697 -5118 -1680 -5114
rect -1676 -5118 -1659 -5114
rect -1655 -5118 -1638 -5114
rect -1634 -5118 -1618 -5114
rect -1614 -5118 -1538 -5114
rect -1534 -5118 -1521 -5114
rect -1517 -5118 -1501 -5114
rect -1497 -5118 -1480 -5114
rect -1476 -5118 -1459 -5114
rect -1455 -5118 -1438 -5114
rect -1434 -5118 -1417 -5114
rect -1413 -5118 -1396 -5114
rect -1392 -5118 -1375 -5114
rect -1371 -5118 -1355 -5114
rect -1351 -5118 -1225 -5114
rect -1221 -5118 -1208 -5114
rect -1204 -5118 -1188 -5114
rect -1184 -5118 -1167 -5114
rect -1163 -5118 -1146 -5114
rect -1142 -5118 -1125 -5114
rect -1121 -5118 -1104 -5114
rect -1100 -5118 -1083 -5114
rect -1079 -5118 -1062 -5114
rect -1058 -5118 -1042 -5114
rect -1038 -5118 -926 -5114
rect -922 -5118 -909 -5114
rect -905 -5118 -889 -5114
rect -885 -5118 -868 -5114
rect -864 -5118 -847 -5114
rect -843 -5118 -826 -5114
rect -822 -5118 -805 -5114
rect -801 -5118 -784 -5114
rect -780 -5118 -763 -5114
rect -759 -5118 -743 -5114
rect -739 -5118 -714 -5114
rect -2054 -5285 -2027 -5118
rect -1779 -5166 -1745 -5162
rect -1681 -5166 -1661 -5162
rect -1646 -5166 -1543 -5162
rect -1516 -5166 -1482 -5162
rect -1418 -5166 -1398 -5162
rect -1383 -5166 -1340 -5162
rect -1203 -5166 -1169 -5162
rect -1105 -5166 -1085 -5162
rect -1070 -5166 -931 -5162
rect -904 -5166 -870 -5162
rect -806 -5166 -786 -5162
rect -771 -5166 -735 -5162
rect -1547 -5170 -1543 -5166
rect -935 -5170 -931 -5166
rect -1814 -5174 -1803 -5170
rect -1799 -5174 -1769 -5170
rect -1748 -5174 -1717 -5170
rect -1688 -5174 -1657 -5170
rect -1646 -5174 -1619 -5170
rect -1547 -5174 -1540 -5170
rect -1536 -5174 -1506 -5170
rect -1485 -5174 -1454 -5170
rect -1425 -5174 -1394 -5170
rect -1383 -5174 -1356 -5170
rect -1242 -5174 -1227 -5170
rect -1223 -5174 -1193 -5170
rect -1172 -5174 -1141 -5170
rect -1112 -5174 -1081 -5170
rect -1070 -5174 -1043 -5170
rect -935 -5174 -928 -5170
rect -924 -5174 -894 -5170
rect -873 -5174 -842 -5170
rect -813 -5174 -782 -5170
rect -771 -5174 -744 -5170
rect -1806 -5181 -1759 -5177
rect -1723 -5181 -1710 -5177
rect -1706 -5181 -1675 -5177
rect -1639 -5181 -1626 -5177
rect -1622 -5181 -1610 -5177
rect -1543 -5181 -1496 -5177
rect -1460 -5181 -1447 -5177
rect -1443 -5181 -1412 -5177
rect -1376 -5181 -1363 -5177
rect -1359 -5181 -1347 -5177
rect -1230 -5181 -1183 -5177
rect -1147 -5181 -1134 -5177
rect -1130 -5181 -1099 -5177
rect -1063 -5181 -1050 -5177
rect -1046 -5181 -1034 -5177
rect -931 -5181 -884 -5177
rect -848 -5181 -835 -5177
rect -831 -5181 -800 -5177
rect -764 -5181 -751 -5177
rect -747 -5181 -735 -5177
rect -1814 -5188 -1799 -5184
rect -1795 -5188 -1685 -5184
rect -1664 -5188 -1633 -5184
rect -1551 -5188 -1536 -5184
rect -1532 -5188 -1422 -5184
rect -1401 -5188 -1370 -5184
rect -1238 -5188 -1223 -5184
rect -1219 -5188 -1109 -5184
rect -1088 -5188 -1057 -5184
rect -939 -5188 -924 -5184
rect -920 -5188 -810 -5184
rect -789 -5188 -758 -5184
rect -1764 -5195 -1741 -5191
rect -1722 -5195 -1703 -5191
rect -1501 -5195 -1478 -5191
rect -1459 -5195 -1440 -5191
rect -1188 -5195 -1165 -5191
rect -1146 -5195 -1127 -5191
rect -889 -5195 -866 -5191
rect -847 -5195 -828 -5191
rect 1804 -5206 1831 -5091
rect -1932 -5210 -1801 -5206
rect -1797 -5210 -1784 -5206
rect -1780 -5210 -1743 -5206
rect -1739 -5210 -1701 -5206
rect -1697 -5210 -1659 -5206
rect -1655 -5210 -1618 -5206
rect -1614 -5210 -1538 -5206
rect -1534 -5210 -1521 -5206
rect -1517 -5210 -1480 -5206
rect -1476 -5210 -1438 -5206
rect -1434 -5210 -1396 -5206
rect -1392 -5210 -1355 -5206
rect -1351 -5210 -1225 -5206
rect -1221 -5210 -1208 -5206
rect -1204 -5210 -1167 -5206
rect -1163 -5210 -1125 -5206
rect -1121 -5210 -1083 -5206
rect -1079 -5210 -1042 -5206
rect -1038 -5210 -926 -5206
rect -922 -5210 -909 -5206
rect -905 -5210 -868 -5206
rect -864 -5210 -826 -5206
rect -822 -5210 -784 -5206
rect -780 -5210 -743 -5206
rect -739 -5210 1831 -5206
rect -1821 -5218 -1340 -5214
rect -2054 -5289 -1801 -5285
rect -1797 -5289 -1784 -5285
rect -1780 -5289 -1764 -5285
rect -1760 -5289 -1743 -5285
rect -1739 -5289 -1722 -5285
rect -1718 -5289 -1701 -5285
rect -1697 -5289 -1680 -5285
rect -1676 -5289 -1659 -5285
rect -1655 -5289 -1638 -5285
rect -1634 -5289 -1618 -5285
rect -1614 -5289 -1538 -5285
rect -1534 -5289 -1521 -5285
rect -1517 -5289 -1501 -5285
rect -1497 -5289 -1480 -5285
rect -1476 -5289 -1459 -5285
rect -1455 -5289 -1438 -5285
rect -1434 -5289 -1417 -5285
rect -1413 -5289 -1396 -5285
rect -1392 -5289 -1375 -5285
rect -1371 -5289 -1355 -5285
rect -1351 -5289 -1225 -5285
rect -1221 -5289 -1208 -5285
rect -1204 -5289 -1188 -5285
rect -1184 -5289 -1167 -5285
rect -1163 -5289 -1146 -5285
rect -1142 -5289 -1125 -5285
rect -1121 -5289 -1104 -5285
rect -1100 -5289 -1083 -5285
rect -1079 -5289 -1062 -5285
rect -1058 -5289 -1042 -5285
rect -1038 -5289 -926 -5285
rect -922 -5289 -909 -5285
rect -905 -5289 -889 -5285
rect -885 -5289 -868 -5285
rect -864 -5289 -847 -5285
rect -843 -5289 -826 -5285
rect -822 -5289 -805 -5285
rect -801 -5289 -784 -5285
rect -780 -5289 -763 -5285
rect -759 -5289 -743 -5285
rect -739 -5289 -568 -5285
rect -564 -5289 -551 -5285
rect -547 -5289 -531 -5285
rect -527 -5289 -510 -5285
rect -506 -5289 -489 -5285
rect -485 -5289 -468 -5285
rect -464 -5289 -447 -5285
rect -443 -5289 -426 -5285
rect -422 -5289 -405 -5285
rect -401 -5289 -385 -5285
rect -381 -5289 -210 -5285
rect -206 -5289 -193 -5285
rect -189 -5289 -173 -5285
rect -169 -5289 -152 -5285
rect -148 -5289 -131 -5285
rect -127 -5289 -110 -5285
rect -106 -5289 -89 -5285
rect -85 -5289 -68 -5285
rect -64 -5289 -47 -5285
rect -43 -5289 -27 -5285
rect -23 -5289 148 -5285
rect 152 -5289 165 -5285
rect 169 -5289 185 -5285
rect 189 -5289 206 -5285
rect 210 -5289 227 -5285
rect 231 -5289 248 -5285
rect 252 -5289 269 -5285
rect 273 -5289 290 -5285
rect 294 -5289 311 -5285
rect 315 -5289 331 -5285
rect 335 -5289 504 -5285
rect 508 -5289 521 -5285
rect 525 -5289 541 -5285
rect 545 -5289 562 -5285
rect 566 -5289 583 -5285
rect 587 -5289 604 -5285
rect 608 -5289 625 -5285
rect 629 -5289 646 -5285
rect 650 -5289 667 -5285
rect 671 -5289 687 -5285
rect 691 -5289 862 -5285
rect 866 -5289 879 -5285
rect 883 -5289 899 -5285
rect 903 -5289 920 -5285
rect 924 -5289 941 -5285
rect 945 -5289 962 -5285
rect 966 -5289 983 -5285
rect 987 -5289 1004 -5285
rect 1008 -5289 1025 -5285
rect 1029 -5289 1045 -5285
rect 1049 -5289 1220 -5285
rect 1224 -5289 1237 -5285
rect 1241 -5289 1257 -5285
rect 1261 -5289 1278 -5285
rect 1282 -5289 1299 -5285
rect 1303 -5289 1320 -5285
rect 1324 -5289 1341 -5285
rect 1345 -5289 1362 -5285
rect 1366 -5289 1383 -5285
rect 1387 -5289 1403 -5285
rect 1407 -5289 1622 -5285
rect -2054 -5445 -2027 -5289
rect -1779 -5337 -1745 -5333
rect -1681 -5337 -1661 -5333
rect -1646 -5337 -1543 -5333
rect -1516 -5337 -1482 -5333
rect -1418 -5337 -1398 -5333
rect -1383 -5337 -1340 -5333
rect -1203 -5337 -1169 -5333
rect -1105 -5337 -1085 -5333
rect -1070 -5337 -1024 -5333
rect -904 -5337 -870 -5333
rect -806 -5337 -786 -5333
rect -771 -5337 -725 -5333
rect -546 -5337 -512 -5333
rect -448 -5337 -428 -5333
rect -413 -5337 -369 -5333
rect -188 -5337 -154 -5333
rect -90 -5337 -70 -5333
rect -55 -5337 -7 -5333
rect 170 -5337 204 -5333
rect 268 -5337 288 -5333
rect 303 -5337 349 -5333
rect 526 -5337 560 -5333
rect 624 -5337 644 -5333
rect 659 -5337 705 -5333
rect 884 -5337 918 -5333
rect 982 -5337 1002 -5333
rect 1017 -5337 1061 -5333
rect 1242 -5337 1276 -5333
rect 1340 -5337 1360 -5333
rect 1375 -5337 1423 -5333
rect -1547 -5341 -1543 -5337
rect -1821 -5345 -1803 -5341
rect -1799 -5345 -1769 -5341
rect -1748 -5345 -1717 -5341
rect -1688 -5345 -1657 -5341
rect -1646 -5345 -1619 -5341
rect -1547 -5345 -1540 -5341
rect -1536 -5345 -1506 -5341
rect -1485 -5345 -1454 -5341
rect -1425 -5345 -1394 -5341
rect -1383 -5345 -1356 -5341
rect -1253 -5345 -1227 -5341
rect -1223 -5345 -1193 -5341
rect -1172 -5345 -1141 -5341
rect -1112 -5345 -1081 -5341
rect -1070 -5345 -1043 -5341
rect -959 -5345 -928 -5341
rect -924 -5345 -894 -5341
rect -873 -5345 -842 -5341
rect -813 -5345 -782 -5341
rect -771 -5345 -744 -5341
rect -599 -5345 -570 -5341
rect -566 -5345 -536 -5341
rect -515 -5345 -484 -5341
rect -455 -5345 -424 -5341
rect -413 -5345 -386 -5341
rect -245 -5345 -212 -5341
rect -208 -5345 -178 -5341
rect -157 -5345 -126 -5341
rect -97 -5345 -66 -5341
rect -55 -5345 -28 -5341
rect 112 -5345 146 -5341
rect 150 -5345 180 -5341
rect 201 -5345 232 -5341
rect 261 -5345 292 -5341
rect 303 -5345 330 -5341
rect 468 -5345 502 -5341
rect 506 -5345 536 -5341
rect 557 -5345 588 -5341
rect 617 -5345 648 -5341
rect 659 -5345 686 -5341
rect 826 -5345 860 -5341
rect 864 -5345 894 -5341
rect 915 -5345 946 -5341
rect 975 -5345 1006 -5341
rect 1017 -5345 1044 -5341
rect 1181 -5345 1218 -5341
rect 1222 -5345 1252 -5341
rect 1273 -5345 1304 -5341
rect 1333 -5345 1364 -5341
rect 1375 -5345 1402 -5341
rect -1806 -5352 -1759 -5348
rect -1723 -5352 -1710 -5348
rect -1706 -5352 -1675 -5348
rect -1639 -5352 -1626 -5348
rect -1622 -5352 -1610 -5348
rect -1543 -5352 -1496 -5348
rect -1460 -5352 -1447 -5348
rect -1443 -5352 -1412 -5348
rect -1376 -5352 -1363 -5348
rect -1359 -5352 -1347 -5348
rect -1230 -5352 -1183 -5348
rect -1147 -5352 -1134 -5348
rect -1130 -5352 -1099 -5348
rect -1063 -5352 -1050 -5348
rect -1046 -5352 -1034 -5348
rect -931 -5352 -884 -5348
rect -848 -5352 -835 -5348
rect -831 -5352 -800 -5348
rect -764 -5352 -751 -5348
rect -747 -5352 -735 -5348
rect -573 -5352 -526 -5348
rect -490 -5352 -477 -5348
rect -473 -5352 -442 -5348
rect -406 -5352 -393 -5348
rect -389 -5352 -377 -5348
rect -215 -5352 -168 -5348
rect -132 -5352 -119 -5348
rect -115 -5352 -84 -5348
rect -48 -5352 -35 -5348
rect -31 -5352 -19 -5348
rect 143 -5352 190 -5348
rect 226 -5352 239 -5348
rect 243 -5352 274 -5348
rect 310 -5352 323 -5348
rect 327 -5352 339 -5348
rect 499 -5352 546 -5348
rect 582 -5352 595 -5348
rect 599 -5352 630 -5348
rect 666 -5352 679 -5348
rect 683 -5352 695 -5348
rect 857 -5352 904 -5348
rect 940 -5352 953 -5348
rect 957 -5352 988 -5348
rect 1024 -5352 1037 -5348
rect 1041 -5352 1053 -5348
rect 1215 -5352 1262 -5348
rect 1298 -5352 1311 -5348
rect 1315 -5352 1346 -5348
rect 1382 -5352 1395 -5348
rect 1399 -5352 1411 -5348
rect -1814 -5359 -1799 -5355
rect -1795 -5359 -1685 -5355
rect -1664 -5359 -1633 -5355
rect -1551 -5359 -1536 -5355
rect -1532 -5359 -1422 -5355
rect -1401 -5359 -1370 -5355
rect -1238 -5359 -1223 -5355
rect -1219 -5359 -1109 -5355
rect -1088 -5359 -1057 -5355
rect -939 -5359 -924 -5355
rect -920 -5359 -810 -5355
rect -789 -5359 -758 -5355
rect -581 -5359 -566 -5355
rect -562 -5359 -452 -5355
rect -431 -5359 -400 -5355
rect -223 -5359 -208 -5355
rect -204 -5359 -94 -5355
rect -73 -5359 -42 -5355
rect 135 -5359 150 -5355
rect 154 -5359 264 -5355
rect 285 -5359 316 -5355
rect 491 -5359 506 -5355
rect 510 -5359 620 -5355
rect 641 -5359 672 -5355
rect 849 -5359 864 -5355
rect 868 -5359 978 -5355
rect 999 -5359 1030 -5355
rect 1207 -5359 1222 -5355
rect 1226 -5359 1336 -5355
rect 1357 -5359 1388 -5355
rect -1764 -5366 -1741 -5362
rect -1722 -5366 -1703 -5362
rect -1501 -5366 -1478 -5362
rect -1459 -5366 -1440 -5362
rect -1188 -5366 -1165 -5362
rect -1146 -5366 -1127 -5362
rect -889 -5366 -866 -5362
rect -847 -5366 -828 -5362
rect -531 -5366 -508 -5362
rect -489 -5366 -470 -5362
rect -173 -5366 -150 -5362
rect -131 -5366 -112 -5362
rect 185 -5366 208 -5362
rect 227 -5366 246 -5362
rect 541 -5366 564 -5362
rect 583 -5366 602 -5362
rect 899 -5366 922 -5362
rect 941 -5366 960 -5362
rect 1257 -5366 1280 -5362
rect 1299 -5366 1318 -5362
rect 1804 -5377 1831 -5210
rect -1930 -5381 -1801 -5377
rect -1797 -5381 -1784 -5377
rect -1780 -5381 -1743 -5377
rect -1739 -5381 -1701 -5377
rect -1697 -5381 -1659 -5377
rect -1655 -5381 -1618 -5377
rect -1614 -5381 -1538 -5377
rect -1534 -5381 -1521 -5377
rect -1517 -5381 -1480 -5377
rect -1476 -5381 -1438 -5377
rect -1434 -5381 -1396 -5377
rect -1392 -5381 -1355 -5377
rect -1351 -5381 -1225 -5377
rect -1221 -5381 -1208 -5377
rect -1204 -5381 -1167 -5377
rect -1163 -5381 -1125 -5377
rect -1121 -5381 -1083 -5377
rect -1079 -5381 -1042 -5377
rect -1038 -5381 -926 -5377
rect -922 -5381 -909 -5377
rect -905 -5381 -868 -5377
rect -864 -5381 -826 -5377
rect -822 -5381 -784 -5377
rect -780 -5381 -743 -5377
rect -739 -5381 -568 -5377
rect -564 -5381 -551 -5377
rect -547 -5381 -510 -5377
rect -506 -5381 -468 -5377
rect -464 -5381 -426 -5377
rect -422 -5381 -385 -5377
rect -381 -5381 -210 -5377
rect -206 -5381 -193 -5377
rect -189 -5381 -152 -5377
rect -148 -5381 -110 -5377
rect -106 -5381 -68 -5377
rect -64 -5381 -27 -5377
rect -23 -5381 148 -5377
rect 152 -5381 165 -5377
rect 169 -5381 206 -5377
rect 210 -5381 248 -5377
rect 252 -5381 290 -5377
rect 294 -5381 331 -5377
rect 335 -5381 504 -5377
rect 508 -5381 521 -5377
rect 525 -5381 562 -5377
rect 566 -5381 604 -5377
rect 608 -5381 646 -5377
rect 650 -5381 687 -5377
rect 691 -5381 862 -5377
rect 866 -5381 879 -5377
rect 883 -5381 920 -5377
rect 924 -5381 962 -5377
rect 966 -5381 1004 -5377
rect 1008 -5381 1045 -5377
rect 1049 -5381 1220 -5377
rect 1224 -5381 1237 -5377
rect 1241 -5381 1278 -5377
rect 1282 -5381 1320 -5377
rect 1324 -5381 1362 -5377
rect 1366 -5381 1403 -5377
rect 1407 -5381 1831 -5377
rect -1822 -5389 -1340 -5385
rect -1253 -5388 -1024 -5384
rect -959 -5388 -725 -5384
rect -599 -5389 -369 -5385
rect -245 -5388 -7 -5384
rect 112 -5388 349 -5384
rect 468 -5390 705 -5386
rect 826 -5389 1061 -5385
rect 1181 -5388 1423 -5384
rect -2054 -5449 -1801 -5445
rect -1797 -5449 -1784 -5445
rect -1780 -5449 -1764 -5445
rect -1760 -5449 -1743 -5445
rect -1739 -5449 -1722 -5445
rect -1718 -5449 -1701 -5445
rect -1697 -5449 -1680 -5445
rect -1676 -5449 -1659 -5445
rect -1655 -5449 -1638 -5445
rect -1634 -5449 -1618 -5445
rect -1614 -5449 -1538 -5445
rect -1534 -5449 -1521 -5445
rect -1517 -5449 -1501 -5445
rect -1497 -5449 -1480 -5445
rect -1476 -5449 -1459 -5445
rect -1455 -5449 -1438 -5445
rect -1434 -5449 -1417 -5445
rect -1413 -5449 -1396 -5445
rect -1392 -5449 -1375 -5445
rect -1371 -5449 -1355 -5445
rect -1351 -5449 -1225 -5445
rect -1221 -5449 -1208 -5445
rect -1204 -5449 -1188 -5445
rect -1184 -5449 -1167 -5445
rect -1163 -5449 -1146 -5445
rect -1142 -5449 -1125 -5445
rect -1121 -5449 -1104 -5445
rect -1100 -5449 -1083 -5445
rect -1079 -5449 -1062 -5445
rect -1058 -5449 -1042 -5445
rect -1038 -5449 -926 -5445
rect -922 -5449 -909 -5445
rect -905 -5449 -889 -5445
rect -885 -5449 -868 -5445
rect -864 -5449 -847 -5445
rect -843 -5449 -826 -5445
rect -822 -5449 -805 -5445
rect -801 -5449 -784 -5445
rect -780 -5449 -763 -5445
rect -759 -5449 -743 -5445
rect -739 -5449 -568 -5445
rect -564 -5449 -551 -5445
rect -547 -5449 -531 -5445
rect -527 -5449 -510 -5445
rect -506 -5449 -489 -5445
rect -485 -5449 -468 -5445
rect -464 -5449 -447 -5445
rect -443 -5449 -426 -5445
rect -422 -5449 -405 -5445
rect -401 -5449 -385 -5445
rect -381 -5449 -210 -5445
rect -206 -5449 -193 -5445
rect -189 -5449 -173 -5445
rect -169 -5449 -152 -5445
rect -148 -5449 -131 -5445
rect -127 -5449 -110 -5445
rect -106 -5449 -89 -5445
rect -85 -5449 -68 -5445
rect -64 -5449 -47 -5445
rect -43 -5449 -27 -5445
rect -23 -5449 148 -5445
rect 152 -5449 165 -5445
rect 169 -5449 185 -5445
rect 189 -5449 206 -5445
rect 210 -5449 227 -5445
rect 231 -5449 248 -5445
rect 252 -5449 269 -5445
rect 273 -5449 290 -5445
rect 294 -5449 311 -5445
rect 315 -5449 331 -5445
rect 335 -5449 504 -5445
rect 508 -5449 521 -5445
rect 525 -5449 541 -5445
rect 545 -5449 562 -5445
rect 566 -5449 583 -5445
rect 587 -5449 604 -5445
rect 608 -5449 625 -5445
rect 629 -5449 646 -5445
rect 650 -5449 667 -5445
rect 671 -5449 687 -5445
rect 691 -5449 862 -5445
rect 866 -5449 879 -5445
rect 883 -5449 899 -5445
rect 903 -5449 920 -5445
rect 924 -5449 941 -5445
rect 945 -5449 962 -5445
rect 966 -5449 983 -5445
rect 987 -5449 1004 -5445
rect 1008 -5449 1025 -5445
rect 1029 -5449 1045 -5445
rect 1049 -5449 1220 -5445
rect 1224 -5449 1237 -5445
rect 1241 -5449 1257 -5445
rect 1261 -5449 1278 -5445
rect 1282 -5449 1299 -5445
rect 1303 -5449 1320 -5445
rect 1324 -5449 1341 -5445
rect 1345 -5449 1362 -5445
rect 1366 -5449 1383 -5445
rect 1387 -5449 1403 -5445
rect 1407 -5449 1609 -5445
rect -2054 -5559 -2027 -5449
rect -1779 -5497 -1745 -5493
rect -1681 -5497 -1661 -5493
rect -1646 -5497 -1543 -5493
rect -1516 -5497 -1482 -5493
rect -1418 -5497 -1398 -5493
rect -1383 -5497 -1342 -5493
rect -1203 -5497 -1169 -5493
rect -1105 -5497 -1085 -5493
rect -1070 -5497 -1020 -5493
rect -904 -5497 -870 -5493
rect -806 -5497 -786 -5493
rect -771 -5497 -725 -5493
rect -546 -5497 -512 -5493
rect -448 -5497 -428 -5493
rect -413 -5497 -368 -5493
rect -188 -5497 -154 -5493
rect -90 -5497 -70 -5493
rect -55 -5497 -12 -5493
rect 170 -5497 204 -5493
rect 268 -5497 288 -5493
rect 303 -5497 348 -5493
rect 526 -5497 560 -5493
rect 624 -5497 644 -5493
rect 659 -5497 705 -5493
rect 884 -5497 918 -5493
rect 982 -5497 1002 -5493
rect 1017 -5497 1062 -5493
rect 1242 -5497 1276 -5493
rect 1340 -5497 1360 -5493
rect 1375 -5497 1423 -5493
rect -1547 -5501 -1543 -5497
rect -1822 -5505 -1803 -5501
rect -1799 -5505 -1769 -5501
rect -1748 -5505 -1717 -5501
rect -1688 -5505 -1657 -5501
rect -1646 -5505 -1619 -5501
rect -1547 -5505 -1540 -5501
rect -1536 -5505 -1506 -5501
rect -1485 -5505 -1454 -5501
rect -1425 -5505 -1394 -5501
rect -1383 -5505 -1356 -5501
rect -1315 -5505 -1227 -5501
rect -1223 -5505 -1193 -5501
rect -1172 -5505 -1141 -5501
rect -1112 -5505 -1081 -5501
rect -1070 -5505 -1043 -5501
rect -945 -5505 -928 -5501
rect -924 -5505 -894 -5501
rect -873 -5505 -842 -5501
rect -813 -5505 -782 -5501
rect -771 -5505 -744 -5501
rect -587 -5505 -570 -5501
rect -566 -5505 -536 -5501
rect -515 -5505 -484 -5501
rect -455 -5505 -424 -5501
rect -413 -5505 -386 -5501
rect -229 -5505 -212 -5501
rect -208 -5505 -178 -5501
rect -157 -5505 -126 -5501
rect -97 -5505 -66 -5501
rect -55 -5505 -28 -5501
rect 129 -5505 146 -5501
rect 150 -5505 180 -5501
rect 201 -5505 232 -5501
rect 261 -5505 292 -5501
rect 303 -5505 330 -5501
rect 485 -5505 502 -5501
rect 506 -5505 536 -5501
rect 557 -5505 588 -5501
rect 617 -5505 648 -5501
rect 659 -5505 686 -5501
rect 843 -5505 860 -5501
rect 864 -5505 894 -5501
rect 915 -5505 946 -5501
rect 975 -5505 1006 -5501
rect 1017 -5505 1044 -5501
rect 1201 -5505 1218 -5501
rect 1222 -5505 1252 -5501
rect 1273 -5505 1304 -5501
rect 1333 -5505 1364 -5501
rect 1375 -5505 1402 -5501
rect -1806 -5512 -1759 -5508
rect -1723 -5512 -1710 -5508
rect -1706 -5512 -1675 -5508
rect -1639 -5512 -1626 -5508
rect -1622 -5512 -1610 -5508
rect -1543 -5512 -1496 -5508
rect -1460 -5512 -1447 -5508
rect -1443 -5512 -1412 -5508
rect -1376 -5512 -1363 -5508
rect -1359 -5512 -1347 -5508
rect -1230 -5512 -1183 -5508
rect -1147 -5512 -1134 -5508
rect -1130 -5512 -1099 -5508
rect -1063 -5512 -1050 -5508
rect -1046 -5512 -1034 -5508
rect -931 -5512 -884 -5508
rect -848 -5512 -835 -5508
rect -831 -5512 -800 -5508
rect -764 -5512 -751 -5508
rect -747 -5512 -735 -5508
rect -573 -5512 -526 -5508
rect -490 -5512 -477 -5508
rect -473 -5512 -442 -5508
rect -406 -5512 -393 -5508
rect -389 -5512 -377 -5508
rect -215 -5512 -168 -5508
rect -132 -5512 -119 -5508
rect -115 -5512 -84 -5508
rect -48 -5512 -35 -5508
rect -31 -5512 -19 -5508
rect 143 -5512 190 -5508
rect 226 -5512 239 -5508
rect 243 -5512 274 -5508
rect 310 -5512 323 -5508
rect 327 -5512 339 -5508
rect 499 -5512 546 -5508
rect 582 -5512 595 -5508
rect 599 -5512 630 -5508
rect 666 -5512 679 -5508
rect 683 -5512 695 -5508
rect 857 -5512 904 -5508
rect 940 -5512 953 -5508
rect 957 -5512 988 -5508
rect 1024 -5512 1037 -5508
rect 1041 -5512 1053 -5508
rect 1215 -5512 1262 -5508
rect 1298 -5512 1311 -5508
rect 1315 -5512 1346 -5508
rect 1382 -5512 1395 -5508
rect 1399 -5512 1411 -5508
rect -1814 -5519 -1799 -5515
rect -1795 -5519 -1685 -5515
rect -1664 -5519 -1633 -5515
rect -1551 -5519 -1536 -5515
rect -1532 -5519 -1422 -5515
rect -1401 -5519 -1370 -5515
rect -1238 -5519 -1223 -5515
rect -1219 -5519 -1109 -5515
rect -1088 -5519 -1057 -5515
rect -939 -5519 -924 -5515
rect -920 -5519 -810 -5515
rect -789 -5519 -758 -5515
rect -581 -5519 -566 -5515
rect -562 -5519 -452 -5515
rect -431 -5519 -400 -5515
rect -223 -5519 -208 -5515
rect -204 -5519 -94 -5515
rect -73 -5519 -42 -5515
rect 135 -5519 150 -5515
rect 154 -5519 264 -5515
rect 285 -5519 316 -5515
rect 491 -5519 506 -5515
rect 510 -5519 620 -5515
rect 641 -5519 672 -5515
rect 849 -5519 864 -5515
rect 868 -5519 978 -5515
rect 999 -5519 1030 -5515
rect 1207 -5519 1222 -5515
rect 1226 -5519 1336 -5515
rect 1357 -5519 1388 -5515
rect -1764 -5526 -1741 -5522
rect -1722 -5526 -1703 -5522
rect -1501 -5526 -1478 -5522
rect -1459 -5526 -1440 -5522
rect -1188 -5526 -1165 -5522
rect -1146 -5526 -1127 -5522
rect -889 -5526 -866 -5522
rect -847 -5526 -828 -5522
rect -531 -5526 -508 -5522
rect -489 -5526 -470 -5522
rect -173 -5526 -150 -5522
rect -131 -5526 -112 -5522
rect 185 -5526 208 -5522
rect 227 -5526 246 -5522
rect 541 -5526 564 -5522
rect 583 -5526 602 -5522
rect 899 -5526 922 -5522
rect 941 -5526 960 -5522
rect 1257 -5526 1280 -5522
rect 1299 -5526 1318 -5522
rect 1804 -5537 1831 -5381
rect -1945 -5541 -1801 -5537
rect -1797 -5541 -1784 -5537
rect -1780 -5541 -1743 -5537
rect -1739 -5541 -1701 -5537
rect -1697 -5541 -1659 -5537
rect -1655 -5541 -1618 -5537
rect -1614 -5541 -1538 -5537
rect -1534 -5541 -1521 -5537
rect -1517 -5541 -1480 -5537
rect -1476 -5541 -1438 -5537
rect -1434 -5541 -1396 -5537
rect -1392 -5541 -1355 -5537
rect -1351 -5541 -1225 -5537
rect -1221 -5541 -1208 -5537
rect -1204 -5541 -1167 -5537
rect -1163 -5541 -1125 -5537
rect -1121 -5541 -1083 -5537
rect -1079 -5541 -1042 -5537
rect -1038 -5541 -926 -5537
rect -922 -5541 -909 -5537
rect -905 -5541 -868 -5537
rect -864 -5541 -826 -5537
rect -822 -5541 -784 -5537
rect -780 -5541 -743 -5537
rect -739 -5541 -568 -5537
rect -564 -5541 -551 -5537
rect -547 -5541 -510 -5537
rect -506 -5541 -468 -5537
rect -464 -5541 -426 -5537
rect -422 -5541 -385 -5537
rect -381 -5541 -210 -5537
rect -206 -5541 -193 -5537
rect -189 -5541 -152 -5537
rect -148 -5541 -110 -5537
rect -106 -5541 -68 -5537
rect -64 -5541 -27 -5537
rect -23 -5541 148 -5537
rect 152 -5541 165 -5537
rect 169 -5541 206 -5537
rect 210 -5541 248 -5537
rect 252 -5541 290 -5537
rect 294 -5541 331 -5537
rect 335 -5541 504 -5537
rect 508 -5541 521 -5537
rect 525 -5541 562 -5537
rect 566 -5541 604 -5537
rect 608 -5541 646 -5537
rect 650 -5541 687 -5537
rect 691 -5541 862 -5537
rect 866 -5541 879 -5537
rect 883 -5541 920 -5537
rect 924 -5541 962 -5537
rect 966 -5541 1004 -5537
rect 1008 -5541 1045 -5537
rect 1049 -5541 1220 -5537
rect 1224 -5541 1237 -5537
rect 1241 -5541 1278 -5537
rect 1282 -5541 1320 -5537
rect 1324 -5541 1362 -5537
rect 1366 -5541 1403 -5537
rect 1407 -5541 1831 -5537
rect -2054 -5563 -1309 -5559
rect -1305 -5563 -1292 -5559
rect -1288 -5563 -935 -5559
rect -931 -5563 -918 -5559
rect -914 -5563 -577 -5559
rect -573 -5563 -560 -5559
rect -556 -5563 -219 -5559
rect -215 -5563 -202 -5559
rect -198 -5563 139 -5559
rect 143 -5563 156 -5559
rect 160 -5563 495 -5559
rect 499 -5563 512 -5559
rect 516 -5563 853 -5559
rect 857 -5563 870 -5559
rect 874 -5563 1211 -5559
rect 1215 -5563 1228 -5559
rect 1232 -5563 1589 -5559
rect -2054 -5718 -2027 -5563
rect -1304 -5595 -1020 -5591
rect -930 -5595 -725 -5591
rect -572 -5595 -368 -5591
rect -214 -5595 -12 -5591
rect 144 -5595 348 -5591
rect 500 -5595 705 -5591
rect 858 -5595 1062 -5591
rect 1216 -5595 1423 -5591
rect -1338 -5603 -1297 -5599
rect -1293 -5603 -923 -5599
rect -919 -5603 -565 -5599
rect -561 -5603 -207 -5599
rect -203 -5603 151 -5599
rect 155 -5603 507 -5599
rect 511 -5603 865 -5599
rect 869 -5603 1223 -5599
rect 1227 -5603 1589 -5599
rect -975 -5616 -909 -5612
rect -612 -5616 -551 -5612
rect -259 -5616 -193 -5612
rect 101 -5616 165 -5612
rect 455 -5616 521 -5612
rect 814 -5616 879 -5612
rect 1171 -5616 1237 -5612
rect 1804 -5651 1831 -5541
rect -1411 -5655 -1292 -5651
rect -1288 -5655 -918 -5651
rect -914 -5655 -560 -5651
rect -556 -5655 -202 -5651
rect -198 -5655 156 -5651
rect 160 -5655 512 -5651
rect 516 -5655 870 -5651
rect 874 -5655 1228 -5651
rect 1232 -5655 1831 -5651
rect -2054 -5722 -1225 -5718
rect -1221 -5722 -1208 -5718
rect -1204 -5722 -1168 -5718
rect -1164 -5722 -1147 -5718
rect -1143 -5722 -926 -5718
rect -922 -5722 -900 -5718
rect -896 -5722 -883 -5718
rect -879 -5722 -843 -5718
rect -839 -5722 -822 -5718
rect -818 -5722 -805 -5718
rect -801 -5722 -765 -5718
rect -761 -5722 -741 -5718
rect -737 -5722 -704 -5718
rect -700 -5722 -568 -5718
rect -564 -5722 -542 -5718
rect -538 -5722 -525 -5718
rect -521 -5722 -485 -5718
rect -481 -5722 -464 -5718
rect -460 -5722 -447 -5718
rect -443 -5722 -407 -5718
rect -403 -5722 -383 -5718
rect -379 -5722 -346 -5718
rect -342 -5722 -210 -5718
rect -206 -5722 -184 -5718
rect -180 -5722 -167 -5718
rect -163 -5722 -127 -5718
rect -123 -5722 -106 -5718
rect -102 -5722 -89 -5718
rect -85 -5722 -49 -5718
rect -45 -5722 -25 -5718
rect -21 -5722 12 -5718
rect 16 -5722 148 -5718
rect 152 -5722 174 -5718
rect 178 -5722 191 -5718
rect 195 -5722 231 -5718
rect 235 -5722 252 -5718
rect 256 -5722 269 -5718
rect 273 -5722 309 -5718
rect 313 -5722 333 -5718
rect 337 -5722 370 -5718
rect 374 -5722 504 -5718
rect 508 -5722 530 -5718
rect 534 -5722 547 -5718
rect 551 -5722 587 -5718
rect 591 -5722 608 -5718
rect 612 -5722 625 -5718
rect 629 -5722 665 -5718
rect 669 -5722 689 -5718
rect 693 -5722 726 -5718
rect 730 -5722 862 -5718
rect 866 -5722 888 -5718
rect 892 -5722 905 -5718
rect 909 -5722 945 -5718
rect 949 -5722 966 -5718
rect 970 -5722 983 -5718
rect 987 -5722 1023 -5718
rect 1027 -5722 1047 -5718
rect 1051 -5722 1084 -5718
rect 1088 -5722 1220 -5718
rect 1224 -5722 1246 -5718
rect 1250 -5722 1263 -5718
rect 1267 -5722 1303 -5718
rect 1307 -5722 1324 -5718
rect 1328 -5722 1341 -5718
rect 1345 -5722 1381 -5718
rect 1385 -5722 1405 -5718
rect 1409 -5722 1442 -5718
rect 1446 -5722 1589 -5718
rect -2054 -5841 -2027 -5722
rect -926 -5726 -922 -5722
rect -900 -5726 -896 -5722
rect -883 -5726 -879 -5722
rect -843 -5726 -839 -5722
rect -822 -5726 -818 -5722
rect -805 -5726 -801 -5722
rect -765 -5726 -761 -5722
rect -741 -5726 -737 -5722
rect -704 -5726 -700 -5722
rect -568 -5726 -564 -5722
rect -542 -5726 -538 -5722
rect -525 -5726 -521 -5722
rect -485 -5726 -481 -5722
rect -464 -5726 -460 -5722
rect -447 -5726 -443 -5722
rect -407 -5726 -403 -5722
rect -383 -5726 -379 -5722
rect -346 -5726 -342 -5722
rect -210 -5726 -206 -5722
rect -184 -5726 -180 -5722
rect -167 -5726 -163 -5722
rect -127 -5726 -123 -5722
rect -106 -5726 -102 -5722
rect -89 -5726 -85 -5722
rect -49 -5726 -45 -5722
rect -25 -5726 -21 -5722
rect 12 -5726 16 -5722
rect 148 -5726 152 -5722
rect 174 -5726 178 -5722
rect 191 -5726 195 -5722
rect 231 -5726 235 -5722
rect 252 -5726 256 -5722
rect 269 -5726 273 -5722
rect 309 -5726 313 -5722
rect 333 -5726 337 -5722
rect 370 -5726 374 -5722
rect 504 -5726 508 -5722
rect 530 -5726 534 -5722
rect 547 -5726 551 -5722
rect 587 -5726 591 -5722
rect 608 -5726 612 -5722
rect 625 -5726 629 -5722
rect 665 -5726 669 -5722
rect 689 -5726 693 -5722
rect 726 -5726 730 -5722
rect 862 -5726 866 -5722
rect 888 -5726 892 -5722
rect 905 -5726 909 -5722
rect 945 -5726 949 -5722
rect 966 -5726 970 -5722
rect 983 -5726 987 -5722
rect 1023 -5726 1027 -5722
rect 1047 -5726 1051 -5722
rect 1084 -5726 1088 -5722
rect 1220 -5726 1224 -5722
rect 1246 -5726 1250 -5722
rect 1263 -5726 1267 -5722
rect 1303 -5726 1307 -5722
rect 1324 -5726 1328 -5722
rect 1341 -5726 1345 -5722
rect 1381 -5726 1385 -5722
rect 1405 -5726 1409 -5722
rect 1442 -5726 1446 -5722
rect -920 -5741 -858 -5737
rect -854 -5741 -824 -5737
rect -776 -5741 -746 -5737
rect -562 -5741 -500 -5737
rect -496 -5741 -466 -5737
rect -418 -5741 -388 -5737
rect -204 -5741 -142 -5737
rect -138 -5741 -108 -5737
rect -60 -5741 -30 -5737
rect 154 -5741 216 -5737
rect 220 -5741 250 -5737
rect 298 -5741 328 -5737
rect 510 -5741 572 -5737
rect 576 -5741 606 -5737
rect 654 -5741 684 -5737
rect 868 -5741 930 -5737
rect 934 -5741 964 -5737
rect 1012 -5741 1042 -5737
rect 1226 -5741 1288 -5737
rect 1292 -5741 1322 -5737
rect 1370 -5741 1400 -5737
rect -913 -5748 -882 -5744
rect -555 -5748 -524 -5744
rect -197 -5748 -166 -5744
rect 161 -5748 192 -5744
rect 517 -5748 548 -5744
rect 875 -5748 906 -5744
rect 1233 -5748 1264 -5744
rect -931 -5755 -848 -5751
rect -809 -5755 -706 -5751
rect -573 -5755 -490 -5751
rect -451 -5755 -348 -5751
rect -215 -5755 -132 -5751
rect -93 -5755 10 -5751
rect 143 -5755 226 -5751
rect 265 -5755 368 -5751
rect 499 -5755 582 -5751
rect 621 -5755 724 -5751
rect 857 -5755 940 -5751
rect 979 -5755 1082 -5751
rect 1215 -5755 1298 -5751
rect 1337 -5755 1440 -5751
rect -975 -5762 -928 -5758
rect -894 -5762 -865 -5758
rect -861 -5762 -780 -5758
rect -691 -5762 -612 -5758
rect -599 -5762 -570 -5758
rect -536 -5762 -507 -5758
rect -503 -5762 -422 -5758
rect -333 -5761 -259 -5757
rect -616 -5766 -612 -5762
rect -263 -5766 -259 -5761
rect -245 -5762 -212 -5758
rect -178 -5762 -149 -5758
rect -145 -5762 -64 -5758
rect 25 -5762 101 -5758
rect 112 -5762 146 -5758
rect 180 -5762 209 -5758
rect 213 -5762 294 -5758
rect 383 -5762 455 -5758
rect 468 -5762 502 -5758
rect 536 -5762 565 -5758
rect 569 -5762 650 -5758
rect 739 -5762 814 -5758
rect 826 -5762 860 -5758
rect 894 -5762 923 -5758
rect 927 -5762 1008 -5758
rect 1097 -5760 1164 -5756
rect 97 -5766 101 -5762
rect 451 -5766 455 -5762
rect 810 -5766 814 -5762
rect 1160 -5766 1164 -5760
rect 1171 -5762 1218 -5758
rect 1252 -5762 1281 -5758
rect 1285 -5762 1366 -5758
rect -1230 -5771 -1173 -5767
rect -1134 -5770 -902 -5766
rect -887 -5770 -804 -5766
rect -783 -5770 -683 -5766
rect -616 -5770 -544 -5766
rect -529 -5770 -446 -5766
rect -425 -5770 -326 -5766
rect -263 -5770 -186 -5766
rect -171 -5770 -88 -5766
rect -67 -5770 33 -5766
rect 97 -5770 172 -5766
rect 187 -5770 270 -5766
rect 291 -5770 392 -5766
rect 451 -5770 528 -5766
rect 543 -5770 626 -5766
rect 647 -5770 748 -5766
rect 810 -5770 886 -5766
rect 901 -5770 984 -5766
rect 1005 -5770 1106 -5766
rect 1160 -5770 1244 -5766
rect 1259 -5770 1342 -5766
rect 1363 -5770 1466 -5766
rect -1253 -5778 -1223 -5774
rect -1219 -5778 -1183 -5774
rect -1179 -5778 -1163 -5774
rect -959 -5777 -924 -5773
rect -905 -5777 -776 -5773
rect -612 -5777 -566 -5773
rect -547 -5777 -418 -5773
rect -259 -5777 -208 -5773
rect -189 -5777 -60 -5773
rect 101 -5777 150 -5773
rect 169 -5777 298 -5773
rect 455 -5777 506 -5773
rect 525 -5777 654 -5773
rect 814 -5777 864 -5773
rect 883 -5777 1012 -5773
rect 1181 -5777 1222 -5773
rect 1241 -5777 1370 -5773
rect -1279 -5785 -1227 -5781
rect -1223 -5785 -1197 -5781
rect -1193 -5785 -1149 -5781
rect -898 -5784 -794 -5780
rect -790 -5784 -760 -5780
rect -540 -5784 -436 -5780
rect -432 -5784 -402 -5780
rect -182 -5784 -78 -5780
rect -74 -5784 -44 -5780
rect 176 -5784 280 -5780
rect 284 -5784 314 -5780
rect 532 -5784 636 -5780
rect 640 -5784 670 -5780
rect 890 -5784 994 -5780
rect 998 -5784 1028 -5780
rect 1248 -5784 1352 -5780
rect 1356 -5784 1386 -5780
rect -1186 -5792 -1103 -5788
rect -924 -5791 -872 -5787
rect -868 -5791 -838 -5787
rect -566 -5791 -514 -5787
rect -510 -5791 -480 -5787
rect -208 -5791 -156 -5787
rect -152 -5791 -122 -5787
rect 150 -5791 202 -5787
rect 206 -5791 236 -5787
rect 506 -5791 558 -5787
rect 562 -5791 592 -5787
rect 864 -5791 916 -5787
rect 920 -5791 950 -5787
rect 1222 -5791 1274 -5787
rect 1278 -5791 1308 -5787
rect -1204 -5799 -1172 -5795
rect -879 -5799 -847 -5795
rect -883 -5802 -879 -5799
rect -847 -5802 -843 -5799
rect -801 -5799 -769 -5795
rect -805 -5802 -801 -5799
rect -769 -5802 -765 -5799
rect -521 -5799 -489 -5795
rect -525 -5802 -521 -5799
rect -489 -5802 -485 -5799
rect -443 -5799 -411 -5795
rect -447 -5802 -443 -5799
rect -411 -5802 -407 -5799
rect -163 -5799 -131 -5795
rect -167 -5802 -163 -5799
rect -131 -5802 -127 -5799
rect -85 -5799 -53 -5795
rect -89 -5802 -85 -5799
rect -53 -5802 -49 -5799
rect 195 -5799 227 -5795
rect 191 -5802 195 -5799
rect 227 -5802 231 -5799
rect 273 -5799 305 -5795
rect 269 -5802 273 -5799
rect 305 -5802 309 -5799
rect 551 -5799 583 -5795
rect 547 -5802 551 -5799
rect 583 -5802 587 -5799
rect 629 -5799 661 -5795
rect 625 -5802 629 -5799
rect 661 -5802 665 -5799
rect 909 -5799 941 -5795
rect 905 -5802 909 -5799
rect 941 -5802 945 -5799
rect 987 -5799 1019 -5795
rect 983 -5802 987 -5799
rect 1019 -5802 1023 -5799
rect 1267 -5799 1299 -5795
rect 1263 -5802 1267 -5799
rect 1299 -5802 1303 -5799
rect 1345 -5799 1377 -5795
rect 1341 -5802 1345 -5799
rect 1377 -5802 1381 -5799
rect -926 -5810 -922 -5806
rect -900 -5810 -896 -5806
rect -857 -5810 -853 -5806
rect -822 -5810 -818 -5806
rect -778 -5810 -774 -5806
rect -761 -5810 -757 -5806
rect -725 -5810 -721 -5806
rect -704 -5810 -700 -5806
rect -568 -5810 -564 -5806
rect -542 -5810 -538 -5806
rect -499 -5810 -495 -5806
rect -464 -5810 -460 -5806
rect -420 -5810 -416 -5806
rect -403 -5810 -399 -5806
rect -367 -5810 -363 -5806
rect -346 -5810 -342 -5806
rect -210 -5810 -206 -5806
rect -184 -5810 -180 -5806
rect -141 -5810 -137 -5806
rect -106 -5810 -102 -5806
rect -62 -5810 -58 -5806
rect -45 -5810 -41 -5806
rect -9 -5810 -5 -5806
rect 12 -5810 16 -5806
rect 148 -5810 152 -5806
rect 174 -5810 178 -5806
rect 217 -5810 221 -5806
rect 252 -5810 256 -5806
rect 296 -5810 300 -5806
rect 313 -5810 317 -5806
rect 349 -5810 353 -5806
rect 370 -5810 374 -5806
rect 504 -5810 508 -5806
rect 530 -5810 534 -5806
rect 573 -5810 577 -5806
rect 608 -5810 612 -5806
rect 652 -5810 656 -5806
rect 669 -5810 673 -5806
rect 705 -5810 709 -5806
rect 726 -5810 730 -5806
rect 862 -5810 866 -5806
rect 888 -5810 892 -5806
rect 931 -5810 935 -5806
rect 966 -5810 970 -5806
rect 1010 -5810 1014 -5806
rect 1027 -5810 1031 -5806
rect 1063 -5810 1067 -5806
rect 1084 -5810 1088 -5806
rect 1220 -5810 1224 -5806
rect 1246 -5810 1250 -5806
rect 1289 -5810 1293 -5806
rect 1324 -5810 1328 -5806
rect 1368 -5810 1372 -5806
rect 1385 -5810 1389 -5806
rect 1421 -5810 1425 -5806
rect 1442 -5810 1446 -5806
rect 1804 -5810 1831 -5655
rect -1965 -5814 -1225 -5810
rect -1221 -5814 -1181 -5810
rect -1177 -5814 -1147 -5810
rect -1143 -5814 -926 -5810
rect -922 -5814 -900 -5810
rect -896 -5814 -857 -5810
rect -853 -5814 -822 -5810
rect -818 -5814 -778 -5810
rect -774 -5814 -761 -5810
rect -757 -5814 -725 -5810
rect -721 -5814 -704 -5810
rect -700 -5814 -568 -5810
rect -564 -5814 -542 -5810
rect -538 -5814 -499 -5810
rect -495 -5814 -464 -5810
rect -460 -5814 -420 -5810
rect -416 -5814 -403 -5810
rect -399 -5814 -367 -5810
rect -363 -5814 -346 -5810
rect -342 -5814 -210 -5810
rect -206 -5814 -184 -5810
rect -180 -5814 -141 -5810
rect -137 -5814 -106 -5810
rect -102 -5814 -62 -5810
rect -58 -5814 -45 -5810
rect -41 -5814 -9 -5810
rect -5 -5814 12 -5810
rect 16 -5814 148 -5810
rect 152 -5814 174 -5810
rect 178 -5814 217 -5810
rect 221 -5814 252 -5810
rect 256 -5814 296 -5810
rect 300 -5814 313 -5810
rect 317 -5814 349 -5810
rect 353 -5814 370 -5810
rect 374 -5814 504 -5810
rect 508 -5814 530 -5810
rect 534 -5814 573 -5810
rect 577 -5814 608 -5810
rect 612 -5814 652 -5810
rect 656 -5814 669 -5810
rect 673 -5814 705 -5810
rect 709 -5814 726 -5810
rect 730 -5814 862 -5810
rect 866 -5814 888 -5810
rect 892 -5814 931 -5810
rect 935 -5814 966 -5810
rect 970 -5814 1010 -5810
rect 1014 -5814 1027 -5810
rect 1031 -5814 1063 -5810
rect 1067 -5814 1084 -5810
rect 1088 -5814 1220 -5810
rect 1224 -5814 1246 -5810
rect 1250 -5814 1289 -5810
rect 1293 -5814 1324 -5810
rect 1328 -5814 1368 -5810
rect 1372 -5814 1385 -5810
rect 1389 -5814 1421 -5810
rect 1425 -5814 1442 -5810
rect 1446 -5814 1831 -5810
rect -1242 -5824 -1103 -5820
rect -945 -5821 -683 -5817
rect -582 -5821 -326 -5817
rect -229 -5821 33 -5817
rect 133 -5822 392 -5818
rect 488 -5821 748 -5817
rect 846 -5821 1106 -5817
rect 1203 -5821 1466 -5817
rect -2054 -5845 -1225 -5841
rect -1221 -5845 -1208 -5841
rect -1204 -5845 -1188 -5841
rect -1184 -5845 -1167 -5841
rect -1163 -5845 -1146 -5841
rect -1142 -5845 -1125 -5841
rect -1121 -5845 -1104 -5841
rect -1100 -5845 -1083 -5841
rect -1079 -5845 -1062 -5841
rect -1058 -5845 -1042 -5841
rect -1038 -5845 -926 -5841
rect -922 -5845 -909 -5841
rect -905 -5845 -889 -5841
rect -885 -5845 -868 -5841
rect -864 -5845 -847 -5841
rect -843 -5845 -826 -5841
rect -822 -5845 -805 -5841
rect -801 -5845 -784 -5841
rect -780 -5845 -763 -5841
rect -759 -5845 -743 -5841
rect -739 -5845 -568 -5841
rect -564 -5845 -551 -5841
rect -547 -5845 -531 -5841
rect -527 -5845 -510 -5841
rect -506 -5845 -489 -5841
rect -485 -5845 -468 -5841
rect -464 -5845 -447 -5841
rect -443 -5845 -426 -5841
rect -422 -5845 -405 -5841
rect -401 -5845 -385 -5841
rect -381 -5845 -210 -5841
rect -206 -5845 -193 -5841
rect -189 -5845 -173 -5841
rect -169 -5845 -152 -5841
rect -148 -5845 -131 -5841
rect -127 -5845 -110 -5841
rect -106 -5845 -89 -5841
rect -85 -5845 -68 -5841
rect -64 -5845 -47 -5841
rect -43 -5845 -27 -5841
rect -23 -5845 148 -5841
rect 152 -5845 165 -5841
rect 169 -5845 185 -5841
rect 189 -5845 206 -5841
rect 210 -5845 227 -5841
rect 231 -5845 248 -5841
rect 252 -5845 269 -5841
rect 273 -5845 290 -5841
rect 294 -5845 311 -5841
rect 315 -5845 331 -5841
rect 335 -5845 504 -5841
rect 508 -5845 521 -5841
rect 525 -5845 541 -5841
rect 545 -5845 562 -5841
rect 566 -5845 583 -5841
rect 587 -5845 604 -5841
rect 608 -5845 625 -5841
rect 629 -5845 646 -5841
rect 650 -5845 667 -5841
rect 671 -5845 687 -5841
rect 691 -5845 862 -5841
rect 866 -5845 879 -5841
rect 883 -5845 899 -5841
rect 903 -5845 920 -5841
rect 924 -5845 941 -5841
rect 945 -5845 962 -5841
rect 966 -5845 983 -5841
rect 987 -5845 1004 -5841
rect 1008 -5845 1025 -5841
rect 1029 -5845 1045 -5841
rect 1049 -5845 1220 -5841
rect 1224 -5845 1237 -5841
rect 1241 -5845 1257 -5841
rect 1261 -5845 1278 -5841
rect 1282 -5845 1299 -5841
rect 1303 -5845 1320 -5841
rect 1324 -5845 1341 -5841
rect 1345 -5845 1362 -5841
rect 1366 -5845 1383 -5841
rect 1387 -5845 1403 -5841
rect 1407 -5845 1564 -5841
rect 1568 -5845 1581 -5841
rect 1585 -5845 1601 -5841
rect 1605 -5845 1622 -5841
rect 1626 -5845 1643 -5841
rect 1647 -5845 1664 -5841
rect 1668 -5845 1685 -5841
rect 1689 -5845 1706 -5841
rect 1710 -5845 1727 -5841
rect 1731 -5845 1747 -5841
rect 1751 -5845 1755 -5841
rect -2054 -5997 -2027 -5845
rect -1203 -5893 -1169 -5889
rect -1105 -5893 -1085 -5889
rect -1070 -5893 -1034 -5889
rect -904 -5893 -870 -5889
rect -806 -5893 -786 -5889
rect -771 -5893 -735 -5889
rect -546 -5893 -512 -5889
rect -448 -5893 -428 -5889
rect -413 -5893 -377 -5889
rect -188 -5893 -154 -5889
rect -90 -5893 -70 -5889
rect -55 -5893 -19 -5889
rect 170 -5893 204 -5889
rect 268 -5893 288 -5889
rect 303 -5893 339 -5889
rect 526 -5893 560 -5889
rect 624 -5893 644 -5889
rect 659 -5893 695 -5889
rect 884 -5893 918 -5889
rect 982 -5893 1002 -5889
rect 1017 -5893 1053 -5889
rect 1242 -5893 1276 -5889
rect 1340 -5893 1360 -5889
rect 1375 -5893 1411 -5889
rect 1586 -5893 1620 -5889
rect 1684 -5893 1704 -5889
rect 1719 -5893 1755 -5889
rect -1242 -5901 -1227 -5897
rect -1223 -5901 -1193 -5897
rect -1172 -5901 -1141 -5897
rect -1112 -5901 -1081 -5897
rect -1070 -5901 -1043 -5897
rect -945 -5901 -928 -5897
rect -924 -5901 -894 -5897
rect -873 -5901 -842 -5897
rect -813 -5901 -782 -5897
rect -771 -5901 -744 -5897
rect -582 -5901 -570 -5897
rect -566 -5901 -536 -5897
rect -515 -5901 -484 -5897
rect -455 -5901 -424 -5897
rect -413 -5901 -386 -5897
rect -229 -5901 -212 -5897
rect -208 -5901 -178 -5897
rect -157 -5901 -126 -5897
rect -97 -5901 -66 -5897
rect -55 -5901 -28 -5897
rect 133 -5901 146 -5897
rect 150 -5901 180 -5897
rect 201 -5901 232 -5897
rect 261 -5901 292 -5897
rect 303 -5901 330 -5897
rect 488 -5901 502 -5897
rect 506 -5901 536 -5897
rect 557 -5901 588 -5897
rect 617 -5901 648 -5897
rect 659 -5901 686 -5897
rect 846 -5901 860 -5897
rect 864 -5901 894 -5897
rect 915 -5901 946 -5897
rect 975 -5901 1006 -5897
rect 1017 -5901 1044 -5897
rect 1203 -5901 1218 -5897
rect 1222 -5901 1252 -5897
rect 1273 -5901 1304 -5897
rect 1333 -5901 1364 -5897
rect 1375 -5901 1402 -5897
rect 1455 -5901 1562 -5897
rect 1566 -5901 1596 -5897
rect 1617 -5901 1648 -5897
rect 1677 -5901 1708 -5897
rect 1719 -5901 1746 -5897
rect -1230 -5908 -1183 -5904
rect -1147 -5908 -1134 -5904
rect -1130 -5908 -1099 -5904
rect -1063 -5908 -1050 -5904
rect -1046 -5908 -1034 -5904
rect -931 -5908 -884 -5904
rect -848 -5908 -835 -5904
rect -831 -5908 -800 -5904
rect -764 -5908 -751 -5904
rect -747 -5908 -735 -5904
rect -573 -5908 -526 -5904
rect -490 -5908 -477 -5904
rect -473 -5908 -442 -5904
rect -406 -5908 -393 -5904
rect -389 -5908 -377 -5904
rect -215 -5908 -168 -5904
rect -132 -5908 -119 -5904
rect -115 -5908 -84 -5904
rect -48 -5908 -35 -5904
rect -31 -5908 -19 -5904
rect 143 -5908 190 -5904
rect 226 -5908 239 -5904
rect 243 -5908 274 -5904
rect 310 -5908 323 -5904
rect 327 -5908 339 -5904
rect 499 -5908 546 -5904
rect 582 -5908 595 -5904
rect 599 -5908 630 -5904
rect 666 -5908 679 -5904
rect 683 -5908 695 -5904
rect 857 -5908 904 -5904
rect 940 -5908 953 -5904
rect 957 -5908 988 -5904
rect 1024 -5908 1037 -5904
rect 1041 -5908 1053 -5904
rect 1215 -5908 1262 -5904
rect 1298 -5908 1311 -5904
rect 1315 -5908 1346 -5904
rect 1382 -5908 1395 -5904
rect 1399 -5908 1411 -5904
rect 1559 -5908 1606 -5904
rect 1642 -5908 1655 -5904
rect 1659 -5908 1690 -5904
rect 1726 -5908 1739 -5904
rect 1743 -5908 1755 -5904
rect -1238 -5915 -1223 -5911
rect -1219 -5915 -1109 -5911
rect -1088 -5915 -1057 -5911
rect -939 -5915 -924 -5911
rect -920 -5915 -810 -5911
rect -789 -5915 -758 -5911
rect -581 -5915 -566 -5911
rect -562 -5915 -452 -5911
rect -431 -5915 -400 -5911
rect -223 -5915 -208 -5911
rect -204 -5915 -94 -5911
rect -73 -5915 -42 -5911
rect 135 -5915 150 -5911
rect 154 -5915 264 -5911
rect 285 -5915 316 -5911
rect 491 -5915 506 -5911
rect 510 -5915 620 -5911
rect 641 -5915 672 -5911
rect 849 -5915 864 -5911
rect 868 -5915 978 -5911
rect 999 -5915 1030 -5911
rect 1207 -5915 1222 -5911
rect 1226 -5915 1336 -5911
rect 1357 -5915 1388 -5911
rect 1551 -5915 1566 -5911
rect 1570 -5915 1680 -5911
rect 1701 -5915 1732 -5911
rect -1188 -5922 -1165 -5918
rect -1146 -5922 -1127 -5918
rect -889 -5922 -866 -5918
rect -847 -5922 -828 -5918
rect -531 -5922 -508 -5918
rect -489 -5922 -470 -5918
rect -173 -5922 -150 -5918
rect -131 -5922 -112 -5918
rect 185 -5922 208 -5918
rect 227 -5922 246 -5918
rect 541 -5922 564 -5918
rect 583 -5922 602 -5918
rect 899 -5922 922 -5918
rect 941 -5922 960 -5918
rect 1257 -5922 1280 -5918
rect 1299 -5922 1318 -5918
rect 1601 -5922 1624 -5918
rect 1643 -5922 1662 -5918
rect 1804 -5933 1831 -5814
rect -1968 -5937 -1225 -5933
rect -1221 -5937 -1208 -5933
rect -1204 -5937 -1167 -5933
rect -1163 -5937 -1125 -5933
rect -1121 -5937 -1083 -5933
rect -1079 -5937 -1042 -5933
rect -1038 -5937 -926 -5933
rect -922 -5937 -909 -5933
rect -905 -5937 -868 -5933
rect -864 -5937 -826 -5933
rect -822 -5937 -784 -5933
rect -780 -5937 -743 -5933
rect -739 -5937 -568 -5933
rect -564 -5937 -551 -5933
rect -547 -5937 -510 -5933
rect -506 -5937 -468 -5933
rect -464 -5937 -426 -5933
rect -422 -5937 -385 -5933
rect -381 -5937 -210 -5933
rect -206 -5937 -193 -5933
rect -189 -5937 -152 -5933
rect -148 -5937 -110 -5933
rect -106 -5937 -68 -5933
rect -64 -5937 -27 -5933
rect -23 -5937 148 -5933
rect 152 -5937 165 -5933
rect 169 -5937 206 -5933
rect 210 -5937 248 -5933
rect 252 -5937 290 -5933
rect 294 -5937 331 -5933
rect 335 -5937 504 -5933
rect 508 -5937 521 -5933
rect 525 -5937 562 -5933
rect 566 -5937 604 -5933
rect 608 -5937 646 -5933
rect 650 -5937 687 -5933
rect 691 -5937 862 -5933
rect 866 -5937 879 -5933
rect 883 -5937 920 -5933
rect 924 -5937 962 -5933
rect 966 -5937 1004 -5933
rect 1008 -5937 1045 -5933
rect 1049 -5937 1220 -5933
rect 1224 -5937 1237 -5933
rect 1241 -5937 1278 -5933
rect 1282 -5937 1320 -5933
rect 1324 -5937 1362 -5933
rect 1366 -5937 1403 -5933
rect 1407 -5937 1564 -5933
rect 1568 -5937 1581 -5933
rect 1585 -5937 1622 -5933
rect 1626 -5937 1664 -5933
rect 1668 -5937 1706 -5933
rect 1710 -5937 1747 -5933
rect 1751 -5937 1831 -5933
rect 1804 -5989 1831 -5937
<< ntransistor >>
rect -1302 -868 -1300 -864
rect -1294 -868 -1292 -864
rect -1284 -868 -1282 -864
rect -931 -868 -929 -864
rect -923 -868 -921 -864
rect -913 -868 -911 -864
rect -572 -868 -570 -864
rect -564 -868 -562 -864
rect -554 -868 -552 -864
rect -214 -868 -212 -864
rect -206 -868 -204 -864
rect -196 -868 -194 -864
rect 143 -868 145 -864
rect 151 -868 153 -864
rect 161 -868 163 -864
rect 500 -868 502 -864
rect 508 -868 510 -864
rect 518 -868 520 -864
rect 858 -868 860 -864
rect 866 -868 868 -864
rect 876 -868 878 -864
rect 1216 -868 1218 -864
rect 1224 -868 1226 -864
rect 1234 -868 1236 -864
rect -1225 -1102 -1223 -1098
rect -1215 -1102 -1213 -1098
rect -1199 -1102 -1197 -1098
rect -1191 -1102 -1189 -1098
rect -1175 -1102 -1173 -1098
rect -1167 -1102 -1165 -1098
rect -1157 -1102 -1155 -1098
rect -1149 -1102 -1147 -1098
rect -1133 -1102 -1131 -1098
rect -1125 -1102 -1123 -1098
rect -1115 -1102 -1113 -1098
rect -1107 -1102 -1105 -1098
rect -1091 -1102 -1089 -1098
rect -1083 -1102 -1081 -1098
rect -1073 -1102 -1071 -1098
rect -1065 -1102 -1063 -1098
rect -1049 -1102 -1047 -1098
rect -1041 -1102 -1039 -1098
rect -930 -1102 -928 -1098
rect -920 -1102 -918 -1098
rect -904 -1102 -902 -1098
rect -896 -1102 -894 -1098
rect -880 -1102 -878 -1098
rect -872 -1102 -870 -1098
rect -862 -1102 -860 -1098
rect -854 -1102 -852 -1098
rect -838 -1102 -836 -1098
rect -830 -1102 -828 -1098
rect -820 -1102 -818 -1098
rect -812 -1102 -810 -1098
rect -796 -1102 -794 -1098
rect -788 -1102 -786 -1098
rect -778 -1102 -776 -1098
rect -770 -1102 -768 -1098
rect -754 -1102 -752 -1098
rect -746 -1102 -744 -1098
rect -572 -1102 -570 -1098
rect -562 -1102 -560 -1098
rect -546 -1102 -544 -1098
rect -538 -1102 -536 -1098
rect -522 -1102 -520 -1098
rect -514 -1102 -512 -1098
rect -504 -1102 -502 -1098
rect -496 -1102 -494 -1098
rect -480 -1102 -478 -1098
rect -472 -1102 -470 -1098
rect -462 -1102 -460 -1098
rect -454 -1102 -452 -1098
rect -438 -1102 -436 -1098
rect -430 -1102 -428 -1098
rect -420 -1102 -418 -1098
rect -412 -1102 -410 -1098
rect -396 -1102 -394 -1098
rect -388 -1102 -386 -1098
rect -214 -1102 -212 -1098
rect -204 -1102 -202 -1098
rect -188 -1102 -186 -1098
rect -180 -1102 -178 -1098
rect -164 -1102 -162 -1098
rect -156 -1102 -154 -1098
rect -146 -1102 -144 -1098
rect -138 -1102 -136 -1098
rect -122 -1102 -120 -1098
rect -114 -1102 -112 -1098
rect -104 -1102 -102 -1098
rect -96 -1102 -94 -1098
rect -80 -1102 -78 -1098
rect -72 -1102 -70 -1098
rect -62 -1102 -60 -1098
rect -54 -1102 -52 -1098
rect -38 -1102 -36 -1098
rect -30 -1102 -28 -1098
rect 144 -1102 146 -1098
rect 154 -1102 156 -1098
rect 170 -1102 172 -1098
rect 178 -1102 180 -1098
rect 194 -1102 196 -1098
rect 202 -1102 204 -1098
rect 212 -1102 214 -1098
rect 220 -1102 222 -1098
rect 236 -1102 238 -1098
rect 244 -1102 246 -1098
rect 254 -1102 256 -1098
rect 262 -1102 264 -1098
rect 278 -1102 280 -1098
rect 286 -1102 288 -1098
rect 296 -1102 298 -1098
rect 304 -1102 306 -1098
rect 320 -1102 322 -1098
rect 328 -1102 330 -1098
rect 500 -1102 502 -1098
rect 510 -1102 512 -1098
rect 526 -1102 528 -1098
rect 534 -1102 536 -1098
rect 550 -1102 552 -1098
rect 558 -1102 560 -1098
rect 568 -1102 570 -1098
rect 576 -1102 578 -1098
rect 592 -1102 594 -1098
rect 600 -1102 602 -1098
rect 610 -1102 612 -1098
rect 618 -1102 620 -1098
rect 634 -1102 636 -1098
rect 642 -1102 644 -1098
rect 652 -1102 654 -1098
rect 660 -1102 662 -1098
rect 676 -1102 678 -1098
rect 684 -1102 686 -1098
rect 858 -1102 860 -1098
rect 868 -1102 870 -1098
rect 884 -1102 886 -1098
rect 892 -1102 894 -1098
rect 908 -1102 910 -1098
rect 916 -1102 918 -1098
rect 926 -1102 928 -1098
rect 934 -1102 936 -1098
rect 950 -1102 952 -1098
rect 958 -1102 960 -1098
rect 968 -1102 970 -1098
rect 976 -1102 978 -1098
rect 992 -1102 994 -1098
rect 1000 -1102 1002 -1098
rect 1010 -1102 1012 -1098
rect 1018 -1102 1020 -1098
rect 1034 -1102 1036 -1098
rect 1042 -1102 1044 -1098
rect -1304 -1218 -1302 -1214
rect -1296 -1218 -1294 -1214
rect -1286 -1218 -1284 -1214
rect -930 -1218 -928 -1214
rect -922 -1218 -920 -1214
rect -912 -1218 -910 -1214
rect -572 -1218 -570 -1214
rect -564 -1218 -562 -1214
rect -554 -1218 -552 -1214
rect -214 -1218 -212 -1214
rect -206 -1218 -204 -1214
rect -196 -1218 -194 -1214
rect 144 -1218 146 -1214
rect 152 -1218 154 -1214
rect 162 -1218 164 -1214
rect 500 -1218 502 -1214
rect 508 -1218 510 -1214
rect 518 -1218 520 -1214
rect 858 -1218 860 -1214
rect 866 -1218 868 -1214
rect 876 -1218 878 -1214
rect 1216 -1218 1218 -1214
rect 1224 -1218 1226 -1214
rect 1234 -1218 1236 -1214
rect -1225 -1382 -1223 -1378
rect -1215 -1382 -1213 -1378
rect -1199 -1382 -1197 -1378
rect -1189 -1382 -1187 -1378
rect -1181 -1382 -1179 -1378
rect -1171 -1382 -1169 -1378
rect -1155 -1382 -1153 -1378
rect -1147 -1382 -1145 -1378
rect -1137 -1382 -1135 -1378
rect -930 -1382 -928 -1378
rect -920 -1382 -918 -1378
rect -904 -1382 -902 -1378
rect -894 -1382 -892 -1378
rect -878 -1382 -876 -1378
rect -868 -1382 -866 -1378
rect -860 -1382 -858 -1378
rect -850 -1382 -848 -1378
rect -834 -1382 -832 -1378
rect -826 -1382 -824 -1378
rect -816 -1382 -814 -1378
rect -800 -1382 -798 -1378
rect -790 -1382 -788 -1378
rect -782 -1382 -780 -1378
rect -772 -1382 -770 -1378
rect -756 -1382 -754 -1378
rect -748 -1382 -746 -1378
rect -732 -1382 -730 -1378
rect -716 -1382 -714 -1378
rect -708 -1382 -706 -1378
rect -698 -1382 -696 -1378
rect -572 -1382 -570 -1378
rect -562 -1382 -560 -1378
rect -546 -1382 -544 -1378
rect -536 -1382 -534 -1378
rect -520 -1382 -518 -1378
rect -510 -1382 -508 -1378
rect -502 -1382 -500 -1378
rect -492 -1382 -490 -1378
rect -476 -1382 -474 -1378
rect -468 -1382 -466 -1378
rect -458 -1382 -456 -1378
rect -442 -1382 -440 -1378
rect -432 -1382 -430 -1378
rect -424 -1382 -422 -1378
rect -414 -1382 -412 -1378
rect -398 -1382 -396 -1378
rect -390 -1382 -388 -1378
rect -374 -1382 -372 -1378
rect -358 -1382 -356 -1378
rect -350 -1382 -348 -1378
rect -340 -1382 -338 -1378
rect -214 -1382 -212 -1378
rect -204 -1382 -202 -1378
rect -188 -1382 -186 -1378
rect -178 -1382 -176 -1378
rect -162 -1382 -160 -1378
rect -152 -1382 -150 -1378
rect -144 -1382 -142 -1378
rect -134 -1382 -132 -1378
rect -118 -1382 -116 -1378
rect -110 -1382 -108 -1378
rect -100 -1382 -98 -1378
rect -84 -1382 -82 -1378
rect -74 -1382 -72 -1378
rect -66 -1382 -64 -1378
rect -56 -1382 -54 -1378
rect -40 -1382 -38 -1378
rect -32 -1382 -30 -1378
rect -16 -1382 -14 -1378
rect 0 -1382 2 -1378
rect 8 -1382 10 -1378
rect 18 -1382 20 -1378
rect 144 -1382 146 -1378
rect 154 -1382 156 -1378
rect 170 -1382 172 -1378
rect 180 -1382 182 -1378
rect 196 -1382 198 -1378
rect 206 -1382 208 -1378
rect 214 -1382 216 -1378
rect 224 -1382 226 -1378
rect 240 -1382 242 -1378
rect 248 -1382 250 -1378
rect 258 -1382 260 -1378
rect 274 -1382 276 -1378
rect 284 -1382 286 -1378
rect 292 -1382 294 -1378
rect 302 -1382 304 -1378
rect 318 -1382 320 -1378
rect 326 -1382 328 -1378
rect 342 -1382 344 -1378
rect 358 -1382 360 -1378
rect 366 -1382 368 -1378
rect 376 -1382 378 -1378
rect 500 -1382 502 -1378
rect 510 -1382 512 -1378
rect 526 -1382 528 -1378
rect 536 -1382 538 -1378
rect 552 -1382 554 -1378
rect 562 -1382 564 -1378
rect 570 -1382 572 -1378
rect 580 -1382 582 -1378
rect 596 -1382 598 -1378
rect 604 -1382 606 -1378
rect 614 -1382 616 -1378
rect 630 -1382 632 -1378
rect 640 -1382 642 -1378
rect 648 -1382 650 -1378
rect 658 -1382 660 -1378
rect 674 -1382 676 -1378
rect 682 -1382 684 -1378
rect 698 -1382 700 -1378
rect 714 -1382 716 -1378
rect 722 -1382 724 -1378
rect 732 -1382 734 -1378
rect 858 -1382 860 -1378
rect 868 -1382 870 -1378
rect 884 -1382 886 -1378
rect 894 -1382 896 -1378
rect 910 -1382 912 -1378
rect 920 -1382 922 -1378
rect 928 -1382 930 -1378
rect 938 -1382 940 -1378
rect 954 -1382 956 -1378
rect 962 -1382 964 -1378
rect 972 -1382 974 -1378
rect 988 -1382 990 -1378
rect 998 -1382 1000 -1378
rect 1006 -1382 1008 -1378
rect 1016 -1382 1018 -1378
rect 1032 -1382 1034 -1378
rect 1040 -1382 1042 -1378
rect 1056 -1382 1058 -1378
rect 1072 -1382 1074 -1378
rect 1080 -1382 1082 -1378
rect 1090 -1382 1092 -1378
rect 1216 -1382 1218 -1378
rect 1226 -1382 1228 -1378
rect 1242 -1382 1244 -1378
rect 1252 -1382 1254 -1378
rect 1260 -1382 1262 -1378
rect 1270 -1382 1272 -1378
rect 1286 -1382 1288 -1378
rect 1294 -1382 1296 -1378
rect 1304 -1382 1306 -1378
rect -1225 -1505 -1223 -1501
rect -1215 -1505 -1213 -1501
rect -1199 -1505 -1197 -1501
rect -1191 -1505 -1189 -1501
rect -1175 -1505 -1173 -1501
rect -1167 -1505 -1165 -1501
rect -1157 -1505 -1155 -1501
rect -1149 -1505 -1147 -1501
rect -1133 -1505 -1131 -1501
rect -1125 -1505 -1123 -1501
rect -1115 -1505 -1113 -1501
rect -1107 -1505 -1105 -1501
rect -1091 -1505 -1089 -1501
rect -1083 -1505 -1081 -1501
rect -1073 -1505 -1071 -1501
rect -1065 -1505 -1063 -1501
rect -1049 -1505 -1047 -1501
rect -1041 -1505 -1039 -1501
rect -930 -1505 -928 -1501
rect -920 -1505 -918 -1501
rect -904 -1505 -902 -1501
rect -896 -1505 -894 -1501
rect -880 -1505 -878 -1501
rect -872 -1505 -870 -1501
rect -862 -1505 -860 -1501
rect -854 -1505 -852 -1501
rect -838 -1505 -836 -1501
rect -830 -1505 -828 -1501
rect -820 -1505 -818 -1501
rect -812 -1505 -810 -1501
rect -796 -1505 -794 -1501
rect -788 -1505 -786 -1501
rect -778 -1505 -776 -1501
rect -770 -1505 -768 -1501
rect -754 -1505 -752 -1501
rect -746 -1505 -744 -1501
rect -572 -1505 -570 -1501
rect -562 -1505 -560 -1501
rect -546 -1505 -544 -1501
rect -538 -1505 -536 -1501
rect -522 -1505 -520 -1501
rect -514 -1505 -512 -1501
rect -504 -1505 -502 -1501
rect -496 -1505 -494 -1501
rect -480 -1505 -478 -1501
rect -472 -1505 -470 -1501
rect -462 -1505 -460 -1501
rect -454 -1505 -452 -1501
rect -438 -1505 -436 -1501
rect -430 -1505 -428 -1501
rect -420 -1505 -418 -1501
rect -412 -1505 -410 -1501
rect -396 -1505 -394 -1501
rect -388 -1505 -386 -1501
rect -214 -1505 -212 -1501
rect -204 -1505 -202 -1501
rect -188 -1505 -186 -1501
rect -180 -1505 -178 -1501
rect -164 -1505 -162 -1501
rect -156 -1505 -154 -1501
rect -146 -1505 -144 -1501
rect -138 -1505 -136 -1501
rect -122 -1505 -120 -1501
rect -114 -1505 -112 -1501
rect -104 -1505 -102 -1501
rect -96 -1505 -94 -1501
rect -80 -1505 -78 -1501
rect -72 -1505 -70 -1501
rect -62 -1505 -60 -1501
rect -54 -1505 -52 -1501
rect -38 -1505 -36 -1501
rect -30 -1505 -28 -1501
rect 144 -1505 146 -1501
rect 154 -1505 156 -1501
rect 170 -1505 172 -1501
rect 178 -1505 180 -1501
rect 194 -1505 196 -1501
rect 202 -1505 204 -1501
rect 212 -1505 214 -1501
rect 220 -1505 222 -1501
rect 236 -1505 238 -1501
rect 244 -1505 246 -1501
rect 254 -1505 256 -1501
rect 262 -1505 264 -1501
rect 278 -1505 280 -1501
rect 286 -1505 288 -1501
rect 296 -1505 298 -1501
rect 304 -1505 306 -1501
rect 320 -1505 322 -1501
rect 328 -1505 330 -1501
rect 500 -1505 502 -1501
rect 510 -1505 512 -1501
rect 526 -1505 528 -1501
rect 534 -1505 536 -1501
rect 550 -1505 552 -1501
rect 558 -1505 560 -1501
rect 568 -1505 570 -1501
rect 576 -1505 578 -1501
rect 592 -1505 594 -1501
rect 600 -1505 602 -1501
rect 610 -1505 612 -1501
rect 618 -1505 620 -1501
rect 634 -1505 636 -1501
rect 642 -1505 644 -1501
rect 652 -1505 654 -1501
rect 660 -1505 662 -1501
rect 676 -1505 678 -1501
rect 684 -1505 686 -1501
rect 858 -1505 860 -1501
rect 868 -1505 870 -1501
rect 884 -1505 886 -1501
rect 892 -1505 894 -1501
rect 908 -1505 910 -1501
rect 916 -1505 918 -1501
rect 926 -1505 928 -1501
rect 934 -1505 936 -1501
rect 950 -1505 952 -1501
rect 958 -1505 960 -1501
rect 968 -1505 970 -1501
rect 976 -1505 978 -1501
rect 992 -1505 994 -1501
rect 1000 -1505 1002 -1501
rect 1010 -1505 1012 -1501
rect 1018 -1505 1020 -1501
rect 1034 -1505 1036 -1501
rect 1042 -1505 1044 -1501
rect -1225 -1676 -1223 -1672
rect -1215 -1676 -1213 -1672
rect -1199 -1676 -1197 -1672
rect -1191 -1676 -1189 -1672
rect -1175 -1676 -1173 -1672
rect -1167 -1676 -1165 -1672
rect -1157 -1676 -1155 -1672
rect -1149 -1676 -1147 -1672
rect -1133 -1676 -1131 -1672
rect -1125 -1676 -1123 -1672
rect -1115 -1676 -1113 -1672
rect -1107 -1676 -1105 -1672
rect -1091 -1676 -1089 -1672
rect -1083 -1676 -1081 -1672
rect -1073 -1676 -1071 -1672
rect -1065 -1676 -1063 -1672
rect -1049 -1676 -1047 -1672
rect -1041 -1676 -1039 -1672
rect -930 -1676 -928 -1672
rect -920 -1676 -918 -1672
rect -904 -1676 -902 -1672
rect -896 -1676 -894 -1672
rect -880 -1676 -878 -1672
rect -872 -1676 -870 -1672
rect -862 -1676 -860 -1672
rect -854 -1676 -852 -1672
rect -838 -1676 -836 -1672
rect -830 -1676 -828 -1672
rect -820 -1676 -818 -1672
rect -812 -1676 -810 -1672
rect -796 -1676 -794 -1672
rect -788 -1676 -786 -1672
rect -778 -1676 -776 -1672
rect -770 -1676 -768 -1672
rect -754 -1676 -752 -1672
rect -746 -1676 -744 -1672
rect -572 -1676 -570 -1672
rect -562 -1676 -560 -1672
rect -546 -1676 -544 -1672
rect -538 -1676 -536 -1672
rect -522 -1676 -520 -1672
rect -514 -1676 -512 -1672
rect -504 -1676 -502 -1672
rect -496 -1676 -494 -1672
rect -480 -1676 -478 -1672
rect -472 -1676 -470 -1672
rect -462 -1676 -460 -1672
rect -454 -1676 -452 -1672
rect -438 -1676 -436 -1672
rect -430 -1676 -428 -1672
rect -420 -1676 -418 -1672
rect -412 -1676 -410 -1672
rect -396 -1676 -394 -1672
rect -388 -1676 -386 -1672
rect -214 -1676 -212 -1672
rect -204 -1676 -202 -1672
rect -188 -1676 -186 -1672
rect -180 -1676 -178 -1672
rect -164 -1676 -162 -1672
rect -156 -1676 -154 -1672
rect -146 -1676 -144 -1672
rect -138 -1676 -136 -1672
rect -122 -1676 -120 -1672
rect -114 -1676 -112 -1672
rect -104 -1676 -102 -1672
rect -96 -1676 -94 -1672
rect -80 -1676 -78 -1672
rect -72 -1676 -70 -1672
rect -62 -1676 -60 -1672
rect -54 -1676 -52 -1672
rect -38 -1676 -36 -1672
rect -30 -1676 -28 -1672
rect 144 -1676 146 -1672
rect 154 -1676 156 -1672
rect 170 -1676 172 -1672
rect 178 -1676 180 -1672
rect 194 -1676 196 -1672
rect 202 -1676 204 -1672
rect 212 -1676 214 -1672
rect 220 -1676 222 -1672
rect 236 -1676 238 -1672
rect 244 -1676 246 -1672
rect 254 -1676 256 -1672
rect 262 -1676 264 -1672
rect 278 -1676 280 -1672
rect 286 -1676 288 -1672
rect 296 -1676 298 -1672
rect 304 -1676 306 -1672
rect 320 -1676 322 -1672
rect 328 -1676 330 -1672
rect 500 -1676 502 -1672
rect 510 -1676 512 -1672
rect 526 -1676 528 -1672
rect 534 -1676 536 -1672
rect 550 -1676 552 -1672
rect 558 -1676 560 -1672
rect 568 -1676 570 -1672
rect 576 -1676 578 -1672
rect 592 -1676 594 -1672
rect 600 -1676 602 -1672
rect 610 -1676 612 -1672
rect 618 -1676 620 -1672
rect 634 -1676 636 -1672
rect 642 -1676 644 -1672
rect 652 -1676 654 -1672
rect 660 -1676 662 -1672
rect 676 -1676 678 -1672
rect 684 -1676 686 -1672
rect 858 -1676 860 -1672
rect 868 -1676 870 -1672
rect 884 -1676 886 -1672
rect 892 -1676 894 -1672
rect 908 -1676 910 -1672
rect 916 -1676 918 -1672
rect 926 -1676 928 -1672
rect 934 -1676 936 -1672
rect 950 -1676 952 -1672
rect 958 -1676 960 -1672
rect 968 -1676 970 -1672
rect 976 -1676 978 -1672
rect 992 -1676 994 -1672
rect 1000 -1676 1002 -1672
rect 1010 -1676 1012 -1672
rect 1018 -1676 1020 -1672
rect 1034 -1676 1036 -1672
rect 1042 -1676 1044 -1672
rect 1216 -1676 1218 -1672
rect 1226 -1676 1228 -1672
rect 1242 -1676 1244 -1672
rect 1250 -1676 1252 -1672
rect 1266 -1676 1268 -1672
rect 1274 -1676 1276 -1672
rect 1284 -1676 1286 -1672
rect 1292 -1676 1294 -1672
rect 1308 -1676 1310 -1672
rect 1316 -1676 1318 -1672
rect 1326 -1676 1328 -1672
rect 1334 -1676 1336 -1672
rect 1350 -1676 1352 -1672
rect 1358 -1676 1360 -1672
rect 1368 -1676 1370 -1672
rect 1376 -1676 1378 -1672
rect 1392 -1676 1394 -1672
rect 1400 -1676 1402 -1672
rect -1554 -1847 -1552 -1843
rect -1544 -1847 -1542 -1843
rect -1528 -1847 -1526 -1843
rect -1520 -1847 -1518 -1843
rect -1504 -1847 -1502 -1843
rect -1496 -1847 -1494 -1843
rect -1486 -1847 -1484 -1843
rect -1478 -1847 -1476 -1843
rect -1462 -1847 -1460 -1843
rect -1454 -1847 -1452 -1843
rect -1444 -1847 -1442 -1843
rect -1436 -1847 -1434 -1843
rect -1420 -1847 -1418 -1843
rect -1412 -1847 -1410 -1843
rect -1402 -1847 -1400 -1843
rect -1394 -1847 -1392 -1843
rect -1378 -1847 -1376 -1843
rect -1370 -1847 -1368 -1843
rect -1225 -1847 -1223 -1843
rect -1215 -1847 -1213 -1843
rect -1199 -1847 -1197 -1843
rect -1191 -1847 -1189 -1843
rect -1175 -1847 -1173 -1843
rect -1167 -1847 -1165 -1843
rect -1157 -1847 -1155 -1843
rect -1149 -1847 -1147 -1843
rect -1133 -1847 -1131 -1843
rect -1125 -1847 -1123 -1843
rect -1115 -1847 -1113 -1843
rect -1107 -1847 -1105 -1843
rect -1091 -1847 -1089 -1843
rect -1083 -1847 -1081 -1843
rect -1073 -1847 -1071 -1843
rect -1065 -1847 -1063 -1843
rect -1049 -1847 -1047 -1843
rect -1041 -1847 -1039 -1843
rect -930 -1847 -928 -1843
rect -920 -1847 -918 -1843
rect -904 -1847 -902 -1843
rect -896 -1847 -894 -1843
rect -880 -1847 -878 -1843
rect -872 -1847 -870 -1843
rect -862 -1847 -860 -1843
rect -854 -1847 -852 -1843
rect -838 -1847 -836 -1843
rect -830 -1847 -828 -1843
rect -820 -1847 -818 -1843
rect -812 -1847 -810 -1843
rect -796 -1847 -794 -1843
rect -788 -1847 -786 -1843
rect -778 -1847 -776 -1843
rect -770 -1847 -768 -1843
rect -754 -1847 -752 -1843
rect -746 -1847 -744 -1843
rect -572 -1847 -570 -1843
rect -562 -1847 -560 -1843
rect -546 -1847 -544 -1843
rect -538 -1847 -536 -1843
rect -522 -1847 -520 -1843
rect -514 -1847 -512 -1843
rect -504 -1847 -502 -1843
rect -496 -1847 -494 -1843
rect -480 -1847 -478 -1843
rect -472 -1847 -470 -1843
rect -462 -1847 -460 -1843
rect -454 -1847 -452 -1843
rect -438 -1847 -436 -1843
rect -430 -1847 -428 -1843
rect -420 -1847 -418 -1843
rect -412 -1847 -410 -1843
rect -396 -1847 -394 -1843
rect -388 -1847 -386 -1843
rect -214 -1847 -212 -1843
rect -204 -1847 -202 -1843
rect -188 -1847 -186 -1843
rect -180 -1847 -178 -1843
rect -164 -1847 -162 -1843
rect -156 -1847 -154 -1843
rect -146 -1847 -144 -1843
rect -138 -1847 -136 -1843
rect -122 -1847 -120 -1843
rect -114 -1847 -112 -1843
rect -104 -1847 -102 -1843
rect -96 -1847 -94 -1843
rect -80 -1847 -78 -1843
rect -72 -1847 -70 -1843
rect -62 -1847 -60 -1843
rect -54 -1847 -52 -1843
rect -38 -1847 -36 -1843
rect -30 -1847 -28 -1843
rect 144 -1847 146 -1843
rect 154 -1847 156 -1843
rect 170 -1847 172 -1843
rect 178 -1847 180 -1843
rect 194 -1847 196 -1843
rect 202 -1847 204 -1843
rect 212 -1847 214 -1843
rect 220 -1847 222 -1843
rect 236 -1847 238 -1843
rect 244 -1847 246 -1843
rect 254 -1847 256 -1843
rect 262 -1847 264 -1843
rect 278 -1847 280 -1843
rect 286 -1847 288 -1843
rect 296 -1847 298 -1843
rect 304 -1847 306 -1843
rect 320 -1847 322 -1843
rect 328 -1847 330 -1843
rect 500 -1847 502 -1843
rect 510 -1847 512 -1843
rect 526 -1847 528 -1843
rect 534 -1847 536 -1843
rect 550 -1847 552 -1843
rect 558 -1847 560 -1843
rect 568 -1847 570 -1843
rect 576 -1847 578 -1843
rect 592 -1847 594 -1843
rect 600 -1847 602 -1843
rect 610 -1847 612 -1843
rect 618 -1847 620 -1843
rect 634 -1847 636 -1843
rect 642 -1847 644 -1843
rect 652 -1847 654 -1843
rect 660 -1847 662 -1843
rect 676 -1847 678 -1843
rect 684 -1847 686 -1843
rect 858 -1847 860 -1843
rect 868 -1847 870 -1843
rect 884 -1847 886 -1843
rect 892 -1847 894 -1843
rect 908 -1847 910 -1843
rect 916 -1847 918 -1843
rect 926 -1847 928 -1843
rect 934 -1847 936 -1843
rect 950 -1847 952 -1843
rect 958 -1847 960 -1843
rect 968 -1847 970 -1843
rect 976 -1847 978 -1843
rect 992 -1847 994 -1843
rect 1000 -1847 1002 -1843
rect 1010 -1847 1012 -1843
rect 1018 -1847 1020 -1843
rect 1034 -1847 1036 -1843
rect 1042 -1847 1044 -1843
rect 1216 -1847 1218 -1843
rect 1226 -1847 1228 -1843
rect 1242 -1847 1244 -1843
rect 1250 -1847 1252 -1843
rect 1266 -1847 1268 -1843
rect 1274 -1847 1276 -1843
rect 1284 -1847 1286 -1843
rect 1292 -1847 1294 -1843
rect 1308 -1847 1310 -1843
rect 1316 -1847 1318 -1843
rect 1326 -1847 1328 -1843
rect 1334 -1847 1336 -1843
rect 1350 -1847 1352 -1843
rect 1358 -1847 1360 -1843
rect 1368 -1847 1370 -1843
rect 1376 -1847 1378 -1843
rect 1392 -1847 1394 -1843
rect 1400 -1847 1402 -1843
rect -1304 -1954 -1302 -1950
rect -1296 -1954 -1294 -1950
rect -1286 -1954 -1284 -1950
rect -930 -1954 -928 -1950
rect -922 -1954 -920 -1950
rect -912 -1954 -910 -1950
rect -572 -1954 -570 -1950
rect -564 -1954 -562 -1950
rect -554 -1954 -552 -1950
rect -214 -1954 -212 -1950
rect -206 -1954 -204 -1950
rect -196 -1954 -194 -1950
rect 144 -1954 146 -1950
rect 152 -1954 154 -1950
rect 162 -1954 164 -1950
rect 500 -1954 502 -1950
rect 508 -1954 510 -1950
rect 518 -1954 520 -1950
rect 858 -1954 860 -1950
rect 866 -1954 868 -1950
rect 876 -1954 878 -1950
rect 1216 -1954 1218 -1950
rect 1224 -1954 1226 -1950
rect 1234 -1954 1236 -1950
rect -1229 -2113 -1227 -2109
rect -1219 -2113 -1217 -2109
rect -1203 -2113 -1201 -2109
rect -1193 -2113 -1191 -2109
rect -1185 -2113 -1183 -2109
rect -1175 -2113 -1173 -2109
rect -1159 -2113 -1157 -2109
rect -1151 -2113 -1149 -2109
rect -1141 -2113 -1139 -2109
rect -930 -2113 -928 -2109
rect -920 -2113 -918 -2109
rect -904 -2113 -902 -2109
rect -894 -2113 -892 -2109
rect -878 -2113 -876 -2109
rect -868 -2113 -866 -2109
rect -860 -2113 -858 -2109
rect -850 -2113 -848 -2109
rect -834 -2113 -832 -2109
rect -826 -2113 -824 -2109
rect -816 -2113 -814 -2109
rect -800 -2113 -798 -2109
rect -790 -2113 -788 -2109
rect -782 -2113 -780 -2109
rect -772 -2113 -770 -2109
rect -756 -2113 -754 -2109
rect -748 -2113 -746 -2109
rect -732 -2113 -730 -2109
rect -716 -2113 -714 -2109
rect -708 -2113 -706 -2109
rect -698 -2113 -696 -2109
rect -572 -2113 -570 -2109
rect -562 -2113 -560 -2109
rect -546 -2113 -544 -2109
rect -536 -2113 -534 -2109
rect -520 -2113 -518 -2109
rect -510 -2113 -508 -2109
rect -502 -2113 -500 -2109
rect -492 -2113 -490 -2109
rect -476 -2113 -474 -2109
rect -468 -2113 -466 -2109
rect -458 -2113 -456 -2109
rect -442 -2113 -440 -2109
rect -432 -2113 -430 -2109
rect -424 -2113 -422 -2109
rect -414 -2113 -412 -2109
rect -398 -2113 -396 -2109
rect -390 -2113 -388 -2109
rect -374 -2113 -372 -2109
rect -358 -2113 -356 -2109
rect -350 -2113 -348 -2109
rect -340 -2113 -338 -2109
rect -214 -2113 -212 -2109
rect -204 -2113 -202 -2109
rect -188 -2113 -186 -2109
rect -178 -2113 -176 -2109
rect -162 -2113 -160 -2109
rect -152 -2113 -150 -2109
rect -144 -2113 -142 -2109
rect -134 -2113 -132 -2109
rect -118 -2113 -116 -2109
rect -110 -2113 -108 -2109
rect -100 -2113 -98 -2109
rect -84 -2113 -82 -2109
rect -74 -2113 -72 -2109
rect -66 -2113 -64 -2109
rect -56 -2113 -54 -2109
rect -40 -2113 -38 -2109
rect -32 -2113 -30 -2109
rect -16 -2113 -14 -2109
rect 0 -2113 2 -2109
rect 8 -2113 10 -2109
rect 18 -2113 20 -2109
rect 144 -2113 146 -2109
rect 154 -2113 156 -2109
rect 170 -2113 172 -2109
rect 180 -2113 182 -2109
rect 196 -2113 198 -2109
rect 206 -2113 208 -2109
rect 214 -2113 216 -2109
rect 224 -2113 226 -2109
rect 240 -2113 242 -2109
rect 248 -2113 250 -2109
rect 258 -2113 260 -2109
rect 274 -2113 276 -2109
rect 284 -2113 286 -2109
rect 292 -2113 294 -2109
rect 302 -2113 304 -2109
rect 318 -2113 320 -2109
rect 326 -2113 328 -2109
rect 342 -2113 344 -2109
rect 358 -2113 360 -2109
rect 366 -2113 368 -2109
rect 376 -2113 378 -2109
rect 500 -2113 502 -2109
rect 510 -2113 512 -2109
rect 526 -2113 528 -2109
rect 536 -2113 538 -2109
rect 552 -2113 554 -2109
rect 562 -2113 564 -2109
rect 570 -2113 572 -2109
rect 580 -2113 582 -2109
rect 596 -2113 598 -2109
rect 604 -2113 606 -2109
rect 614 -2113 616 -2109
rect 630 -2113 632 -2109
rect 640 -2113 642 -2109
rect 648 -2113 650 -2109
rect 658 -2113 660 -2109
rect 674 -2113 676 -2109
rect 682 -2113 684 -2109
rect 698 -2113 700 -2109
rect 714 -2113 716 -2109
rect 722 -2113 724 -2109
rect 732 -2113 734 -2109
rect 858 -2113 860 -2109
rect 868 -2113 870 -2109
rect 884 -2113 886 -2109
rect 894 -2113 896 -2109
rect 910 -2113 912 -2109
rect 920 -2113 922 -2109
rect 928 -2113 930 -2109
rect 938 -2113 940 -2109
rect 954 -2113 956 -2109
rect 962 -2113 964 -2109
rect 972 -2113 974 -2109
rect 988 -2113 990 -2109
rect 998 -2113 1000 -2109
rect 1006 -2113 1008 -2109
rect 1016 -2113 1018 -2109
rect 1032 -2113 1034 -2109
rect 1040 -2113 1042 -2109
rect 1056 -2113 1058 -2109
rect 1072 -2113 1074 -2109
rect 1080 -2113 1082 -2109
rect 1090 -2113 1092 -2109
rect 1216 -2113 1218 -2109
rect 1226 -2113 1228 -2109
rect 1242 -2113 1244 -2109
rect 1252 -2113 1254 -2109
rect 1268 -2113 1270 -2109
rect 1278 -2113 1280 -2109
rect 1286 -2113 1288 -2109
rect 1296 -2113 1298 -2109
rect 1312 -2113 1314 -2109
rect 1320 -2113 1322 -2109
rect 1330 -2113 1332 -2109
rect 1346 -2113 1348 -2109
rect 1356 -2113 1358 -2109
rect 1364 -2113 1366 -2109
rect 1374 -2113 1376 -2109
rect 1390 -2113 1392 -2109
rect 1398 -2113 1400 -2109
rect 1414 -2113 1416 -2109
rect 1430 -2113 1432 -2109
rect 1438 -2113 1440 -2109
rect 1448 -2113 1450 -2109
rect -1229 -2257 -1227 -2253
rect -1219 -2257 -1217 -2253
rect -1203 -2257 -1201 -2253
rect -1195 -2257 -1193 -2253
rect -1179 -2257 -1177 -2253
rect -1171 -2257 -1169 -2253
rect -1161 -2257 -1159 -2253
rect -1153 -2257 -1151 -2253
rect -1137 -2257 -1135 -2253
rect -1129 -2257 -1127 -2253
rect -1119 -2257 -1117 -2253
rect -1111 -2257 -1109 -2253
rect -1095 -2257 -1093 -2253
rect -1087 -2257 -1085 -2253
rect -1077 -2257 -1075 -2253
rect -1069 -2257 -1067 -2253
rect -1053 -2257 -1051 -2253
rect -1045 -2257 -1043 -2253
rect -930 -2257 -928 -2253
rect -920 -2257 -918 -2253
rect -904 -2257 -902 -2253
rect -896 -2257 -894 -2253
rect -880 -2257 -878 -2253
rect -872 -2257 -870 -2253
rect -862 -2257 -860 -2253
rect -854 -2257 -852 -2253
rect -838 -2257 -836 -2253
rect -830 -2257 -828 -2253
rect -820 -2257 -818 -2253
rect -812 -2257 -810 -2253
rect -796 -2257 -794 -2253
rect -788 -2257 -786 -2253
rect -778 -2257 -776 -2253
rect -770 -2257 -768 -2253
rect -754 -2257 -752 -2253
rect -746 -2257 -744 -2253
rect -572 -2257 -570 -2253
rect -562 -2257 -560 -2253
rect -546 -2257 -544 -2253
rect -538 -2257 -536 -2253
rect -522 -2257 -520 -2253
rect -514 -2257 -512 -2253
rect -504 -2257 -502 -2253
rect -496 -2257 -494 -2253
rect -480 -2257 -478 -2253
rect -472 -2257 -470 -2253
rect -462 -2257 -460 -2253
rect -454 -2257 -452 -2253
rect -438 -2257 -436 -2253
rect -430 -2257 -428 -2253
rect -420 -2257 -418 -2253
rect -412 -2257 -410 -2253
rect -396 -2257 -394 -2253
rect -388 -2257 -386 -2253
rect -214 -2257 -212 -2253
rect -204 -2257 -202 -2253
rect -188 -2257 -186 -2253
rect -180 -2257 -178 -2253
rect -164 -2257 -162 -2253
rect -156 -2257 -154 -2253
rect -146 -2257 -144 -2253
rect -138 -2257 -136 -2253
rect -122 -2257 -120 -2253
rect -114 -2257 -112 -2253
rect -104 -2257 -102 -2253
rect -96 -2257 -94 -2253
rect -80 -2257 -78 -2253
rect -72 -2257 -70 -2253
rect -62 -2257 -60 -2253
rect -54 -2257 -52 -2253
rect -38 -2257 -36 -2253
rect -30 -2257 -28 -2253
rect 144 -2257 146 -2253
rect 154 -2257 156 -2253
rect 170 -2257 172 -2253
rect 178 -2257 180 -2253
rect 194 -2257 196 -2253
rect 202 -2257 204 -2253
rect 212 -2257 214 -2253
rect 220 -2257 222 -2253
rect 236 -2257 238 -2253
rect 244 -2257 246 -2253
rect 254 -2257 256 -2253
rect 262 -2257 264 -2253
rect 278 -2257 280 -2253
rect 286 -2257 288 -2253
rect 296 -2257 298 -2253
rect 304 -2257 306 -2253
rect 320 -2257 322 -2253
rect 328 -2257 330 -2253
rect 500 -2257 502 -2253
rect 510 -2257 512 -2253
rect 526 -2257 528 -2253
rect 534 -2257 536 -2253
rect 550 -2257 552 -2253
rect 558 -2257 560 -2253
rect 568 -2257 570 -2253
rect 576 -2257 578 -2253
rect 592 -2257 594 -2253
rect 600 -2257 602 -2253
rect 610 -2257 612 -2253
rect 618 -2257 620 -2253
rect 634 -2257 636 -2253
rect 642 -2257 644 -2253
rect 652 -2257 654 -2253
rect 660 -2257 662 -2253
rect 676 -2257 678 -2253
rect 684 -2257 686 -2253
rect -1554 -2428 -1552 -2424
rect -1544 -2428 -1542 -2424
rect -1528 -2428 -1526 -2424
rect -1520 -2428 -1518 -2424
rect -1504 -2428 -1502 -2424
rect -1496 -2428 -1494 -2424
rect -1486 -2428 -1484 -2424
rect -1478 -2428 -1476 -2424
rect -1462 -2428 -1460 -2424
rect -1454 -2428 -1452 -2424
rect -1444 -2428 -1442 -2424
rect -1436 -2428 -1434 -2424
rect -1420 -2428 -1418 -2424
rect -1412 -2428 -1410 -2424
rect -1402 -2428 -1400 -2424
rect -1394 -2428 -1392 -2424
rect -1378 -2428 -1376 -2424
rect -1370 -2428 -1368 -2424
rect -1229 -2428 -1227 -2424
rect -1219 -2428 -1217 -2424
rect -1203 -2428 -1201 -2424
rect -1195 -2428 -1193 -2424
rect -1179 -2428 -1177 -2424
rect -1171 -2428 -1169 -2424
rect -1161 -2428 -1159 -2424
rect -1153 -2428 -1151 -2424
rect -1137 -2428 -1135 -2424
rect -1129 -2428 -1127 -2424
rect -1119 -2428 -1117 -2424
rect -1111 -2428 -1109 -2424
rect -1095 -2428 -1093 -2424
rect -1087 -2428 -1085 -2424
rect -1077 -2428 -1075 -2424
rect -1069 -2428 -1067 -2424
rect -1053 -2428 -1051 -2424
rect -1045 -2428 -1043 -2424
rect -930 -2428 -928 -2424
rect -920 -2428 -918 -2424
rect -904 -2428 -902 -2424
rect -896 -2428 -894 -2424
rect -880 -2428 -878 -2424
rect -872 -2428 -870 -2424
rect -862 -2428 -860 -2424
rect -854 -2428 -852 -2424
rect -838 -2428 -836 -2424
rect -830 -2428 -828 -2424
rect -820 -2428 -818 -2424
rect -812 -2428 -810 -2424
rect -796 -2428 -794 -2424
rect -788 -2428 -786 -2424
rect -778 -2428 -776 -2424
rect -770 -2428 -768 -2424
rect -754 -2428 -752 -2424
rect -746 -2428 -744 -2424
rect -572 -2428 -570 -2424
rect -562 -2428 -560 -2424
rect -546 -2428 -544 -2424
rect -538 -2428 -536 -2424
rect -522 -2428 -520 -2424
rect -514 -2428 -512 -2424
rect -504 -2428 -502 -2424
rect -496 -2428 -494 -2424
rect -480 -2428 -478 -2424
rect -472 -2428 -470 -2424
rect -462 -2428 -460 -2424
rect -454 -2428 -452 -2424
rect -438 -2428 -436 -2424
rect -430 -2428 -428 -2424
rect -420 -2428 -418 -2424
rect -412 -2428 -410 -2424
rect -396 -2428 -394 -2424
rect -388 -2428 -386 -2424
rect -214 -2428 -212 -2424
rect -204 -2428 -202 -2424
rect -188 -2428 -186 -2424
rect -180 -2428 -178 -2424
rect -164 -2428 -162 -2424
rect -156 -2428 -154 -2424
rect -146 -2428 -144 -2424
rect -138 -2428 -136 -2424
rect -122 -2428 -120 -2424
rect -114 -2428 -112 -2424
rect -104 -2428 -102 -2424
rect -96 -2428 -94 -2424
rect -80 -2428 -78 -2424
rect -72 -2428 -70 -2424
rect -62 -2428 -60 -2424
rect -54 -2428 -52 -2424
rect -38 -2428 -36 -2424
rect -30 -2428 -28 -2424
rect 144 -2428 146 -2424
rect 154 -2428 156 -2424
rect 170 -2428 172 -2424
rect 178 -2428 180 -2424
rect 194 -2428 196 -2424
rect 202 -2428 204 -2424
rect 212 -2428 214 -2424
rect 220 -2428 222 -2424
rect 236 -2428 238 -2424
rect 244 -2428 246 -2424
rect 254 -2428 256 -2424
rect 262 -2428 264 -2424
rect 278 -2428 280 -2424
rect 286 -2428 288 -2424
rect 296 -2428 298 -2424
rect 304 -2428 306 -2424
rect 320 -2428 322 -2424
rect 328 -2428 330 -2424
rect 500 -2428 502 -2424
rect 510 -2428 512 -2424
rect 526 -2428 528 -2424
rect 534 -2428 536 -2424
rect 550 -2428 552 -2424
rect 558 -2428 560 -2424
rect 568 -2428 570 -2424
rect 576 -2428 578 -2424
rect 592 -2428 594 -2424
rect 600 -2428 602 -2424
rect 610 -2428 612 -2424
rect 618 -2428 620 -2424
rect 634 -2428 636 -2424
rect 642 -2428 644 -2424
rect 652 -2428 654 -2424
rect 660 -2428 662 -2424
rect 676 -2428 678 -2424
rect 684 -2428 686 -2424
rect 858 -2428 860 -2424
rect 868 -2428 870 -2424
rect 884 -2428 886 -2424
rect 892 -2428 894 -2424
rect 908 -2428 910 -2424
rect 916 -2428 918 -2424
rect 926 -2428 928 -2424
rect 934 -2428 936 -2424
rect 950 -2428 952 -2424
rect 958 -2428 960 -2424
rect 968 -2428 970 -2424
rect 976 -2428 978 -2424
rect 992 -2428 994 -2424
rect 1000 -2428 1002 -2424
rect 1010 -2428 1012 -2424
rect 1018 -2428 1020 -2424
rect 1034 -2428 1036 -2424
rect 1042 -2428 1044 -2424
rect 1216 -2428 1218 -2424
rect 1226 -2428 1228 -2424
rect 1242 -2428 1244 -2424
rect 1250 -2428 1252 -2424
rect 1266 -2428 1268 -2424
rect 1274 -2428 1276 -2424
rect 1284 -2428 1286 -2424
rect 1292 -2428 1294 -2424
rect 1308 -2428 1310 -2424
rect 1316 -2428 1318 -2424
rect 1326 -2428 1328 -2424
rect 1334 -2428 1336 -2424
rect 1350 -2428 1352 -2424
rect 1358 -2428 1360 -2424
rect 1368 -2428 1370 -2424
rect 1376 -2428 1378 -2424
rect 1392 -2428 1394 -2424
rect 1400 -2428 1402 -2424
rect -1554 -2599 -1552 -2595
rect -1544 -2599 -1542 -2595
rect -1528 -2599 -1526 -2595
rect -1520 -2599 -1518 -2595
rect -1504 -2599 -1502 -2595
rect -1496 -2599 -1494 -2595
rect -1486 -2599 -1484 -2595
rect -1478 -2599 -1476 -2595
rect -1462 -2599 -1460 -2595
rect -1454 -2599 -1452 -2595
rect -1444 -2599 -1442 -2595
rect -1436 -2599 -1434 -2595
rect -1420 -2599 -1418 -2595
rect -1412 -2599 -1410 -2595
rect -1402 -2599 -1400 -2595
rect -1394 -2599 -1392 -2595
rect -1378 -2599 -1376 -2595
rect -1370 -2599 -1368 -2595
rect -1229 -2599 -1227 -2595
rect -1219 -2599 -1217 -2595
rect -1203 -2599 -1201 -2595
rect -1195 -2599 -1193 -2595
rect -1179 -2599 -1177 -2595
rect -1171 -2599 -1169 -2595
rect -1161 -2599 -1159 -2595
rect -1153 -2599 -1151 -2595
rect -1137 -2599 -1135 -2595
rect -1129 -2599 -1127 -2595
rect -1119 -2599 -1117 -2595
rect -1111 -2599 -1109 -2595
rect -1095 -2599 -1093 -2595
rect -1087 -2599 -1085 -2595
rect -1077 -2599 -1075 -2595
rect -1069 -2599 -1067 -2595
rect -1053 -2599 -1051 -2595
rect -1045 -2599 -1043 -2595
rect -930 -2599 -928 -2595
rect -920 -2599 -918 -2595
rect -904 -2599 -902 -2595
rect -896 -2599 -894 -2595
rect -880 -2599 -878 -2595
rect -872 -2599 -870 -2595
rect -862 -2599 -860 -2595
rect -854 -2599 -852 -2595
rect -838 -2599 -836 -2595
rect -830 -2599 -828 -2595
rect -820 -2599 -818 -2595
rect -812 -2599 -810 -2595
rect -796 -2599 -794 -2595
rect -788 -2599 -786 -2595
rect -778 -2599 -776 -2595
rect -770 -2599 -768 -2595
rect -754 -2599 -752 -2595
rect -746 -2599 -744 -2595
rect -572 -2599 -570 -2595
rect -562 -2599 -560 -2595
rect -546 -2599 -544 -2595
rect -538 -2599 -536 -2595
rect -522 -2599 -520 -2595
rect -514 -2599 -512 -2595
rect -504 -2599 -502 -2595
rect -496 -2599 -494 -2595
rect -480 -2599 -478 -2595
rect -472 -2599 -470 -2595
rect -462 -2599 -460 -2595
rect -454 -2599 -452 -2595
rect -438 -2599 -436 -2595
rect -430 -2599 -428 -2595
rect -420 -2599 -418 -2595
rect -412 -2599 -410 -2595
rect -396 -2599 -394 -2595
rect -388 -2599 -386 -2595
rect -215 -2599 -213 -2595
rect -205 -2599 -203 -2595
rect -189 -2599 -187 -2595
rect -181 -2599 -179 -2595
rect -165 -2599 -163 -2595
rect -157 -2599 -155 -2595
rect -147 -2599 -145 -2595
rect -139 -2599 -137 -2595
rect -123 -2599 -121 -2595
rect -115 -2599 -113 -2595
rect -105 -2599 -103 -2595
rect -97 -2599 -95 -2595
rect -81 -2599 -79 -2595
rect -73 -2599 -71 -2595
rect -63 -2599 -61 -2595
rect -55 -2599 -53 -2595
rect -39 -2599 -37 -2595
rect -31 -2599 -29 -2595
rect 144 -2599 146 -2595
rect 154 -2599 156 -2595
rect 170 -2599 172 -2595
rect 178 -2599 180 -2595
rect 194 -2599 196 -2595
rect 202 -2599 204 -2595
rect 212 -2599 214 -2595
rect 220 -2599 222 -2595
rect 236 -2599 238 -2595
rect 244 -2599 246 -2595
rect 254 -2599 256 -2595
rect 262 -2599 264 -2595
rect 278 -2599 280 -2595
rect 286 -2599 288 -2595
rect 296 -2599 298 -2595
rect 304 -2599 306 -2595
rect 320 -2599 322 -2595
rect 328 -2599 330 -2595
rect 500 -2599 502 -2595
rect 510 -2599 512 -2595
rect 526 -2599 528 -2595
rect 534 -2599 536 -2595
rect 550 -2599 552 -2595
rect 558 -2599 560 -2595
rect 568 -2599 570 -2595
rect 576 -2599 578 -2595
rect 592 -2599 594 -2595
rect 600 -2599 602 -2595
rect 610 -2599 612 -2595
rect 618 -2599 620 -2595
rect 634 -2599 636 -2595
rect 642 -2599 644 -2595
rect 652 -2599 654 -2595
rect 660 -2599 662 -2595
rect 676 -2599 678 -2595
rect 684 -2599 686 -2595
rect 858 -2599 860 -2595
rect 868 -2599 870 -2595
rect 884 -2599 886 -2595
rect 892 -2599 894 -2595
rect 908 -2599 910 -2595
rect 916 -2599 918 -2595
rect 926 -2599 928 -2595
rect 934 -2599 936 -2595
rect 950 -2599 952 -2595
rect 958 -2599 960 -2595
rect 968 -2599 970 -2595
rect 976 -2599 978 -2595
rect 992 -2599 994 -2595
rect 1000 -2599 1002 -2595
rect 1010 -2599 1012 -2595
rect 1018 -2599 1020 -2595
rect 1034 -2599 1036 -2595
rect 1042 -2599 1044 -2595
rect 1216 -2599 1218 -2595
rect 1226 -2599 1228 -2595
rect 1242 -2599 1244 -2595
rect 1250 -2599 1252 -2595
rect 1266 -2599 1268 -2595
rect 1274 -2599 1276 -2595
rect 1284 -2599 1286 -2595
rect 1292 -2599 1294 -2595
rect 1308 -2599 1310 -2595
rect 1316 -2599 1318 -2595
rect 1326 -2599 1328 -2595
rect 1334 -2599 1336 -2595
rect 1350 -2599 1352 -2595
rect 1358 -2599 1360 -2595
rect 1368 -2599 1370 -2595
rect 1376 -2599 1378 -2595
rect 1392 -2599 1394 -2595
rect 1400 -2599 1402 -2595
rect -1304 -2704 -1302 -2700
rect -1296 -2704 -1294 -2700
rect -1286 -2704 -1284 -2700
rect -930 -2704 -928 -2700
rect -922 -2704 -920 -2700
rect -912 -2704 -910 -2700
rect -572 -2704 -570 -2700
rect -564 -2704 -562 -2700
rect -554 -2704 -552 -2700
rect -214 -2704 -212 -2700
rect -206 -2704 -204 -2700
rect -196 -2704 -194 -2700
rect 144 -2704 146 -2700
rect 152 -2704 154 -2700
rect 162 -2704 164 -2700
rect 500 -2704 502 -2700
rect 508 -2704 510 -2700
rect 518 -2704 520 -2700
rect 858 -2704 860 -2700
rect 866 -2704 868 -2700
rect 876 -2704 878 -2700
rect 1216 -2704 1218 -2700
rect 1224 -2704 1226 -2700
rect 1234 -2704 1236 -2700
rect -1229 -2863 -1227 -2859
rect -1219 -2863 -1217 -2859
rect -1203 -2863 -1201 -2859
rect -1193 -2863 -1191 -2859
rect -1185 -2863 -1183 -2859
rect -1175 -2863 -1173 -2859
rect -1159 -2863 -1157 -2859
rect -1151 -2863 -1149 -2859
rect -1141 -2863 -1139 -2859
rect -930 -2863 -928 -2859
rect -920 -2863 -918 -2859
rect -904 -2863 -902 -2859
rect -894 -2863 -892 -2859
rect -878 -2863 -876 -2859
rect -868 -2863 -866 -2859
rect -860 -2863 -858 -2859
rect -850 -2863 -848 -2859
rect -834 -2863 -832 -2859
rect -826 -2863 -824 -2859
rect -816 -2863 -814 -2859
rect -800 -2863 -798 -2859
rect -790 -2863 -788 -2859
rect -782 -2863 -780 -2859
rect -772 -2863 -770 -2859
rect -756 -2863 -754 -2859
rect -748 -2863 -746 -2859
rect -732 -2863 -730 -2859
rect -716 -2863 -714 -2859
rect -708 -2863 -706 -2859
rect -698 -2863 -696 -2859
rect -572 -2863 -570 -2859
rect -562 -2863 -560 -2859
rect -546 -2863 -544 -2859
rect -536 -2863 -534 -2859
rect -520 -2863 -518 -2859
rect -510 -2863 -508 -2859
rect -502 -2863 -500 -2859
rect -492 -2863 -490 -2859
rect -476 -2863 -474 -2859
rect -468 -2863 -466 -2859
rect -458 -2863 -456 -2859
rect -442 -2863 -440 -2859
rect -432 -2863 -430 -2859
rect -424 -2863 -422 -2859
rect -414 -2863 -412 -2859
rect -398 -2863 -396 -2859
rect -390 -2863 -388 -2859
rect -374 -2863 -372 -2859
rect -358 -2863 -356 -2859
rect -350 -2863 -348 -2859
rect -340 -2863 -338 -2859
rect -214 -2863 -212 -2859
rect -204 -2863 -202 -2859
rect -188 -2863 -186 -2859
rect -178 -2863 -176 -2859
rect -162 -2863 -160 -2859
rect -152 -2863 -150 -2859
rect -144 -2863 -142 -2859
rect -134 -2863 -132 -2859
rect -118 -2863 -116 -2859
rect -110 -2863 -108 -2859
rect -100 -2863 -98 -2859
rect -84 -2863 -82 -2859
rect -74 -2863 -72 -2859
rect -66 -2863 -64 -2859
rect -56 -2863 -54 -2859
rect -40 -2863 -38 -2859
rect -32 -2863 -30 -2859
rect -16 -2863 -14 -2859
rect 0 -2863 2 -2859
rect 8 -2863 10 -2859
rect 18 -2863 20 -2859
rect 144 -2863 146 -2859
rect 154 -2863 156 -2859
rect 170 -2863 172 -2859
rect 180 -2863 182 -2859
rect 196 -2863 198 -2859
rect 206 -2863 208 -2859
rect 214 -2863 216 -2859
rect 224 -2863 226 -2859
rect 240 -2863 242 -2859
rect 248 -2863 250 -2859
rect 258 -2863 260 -2859
rect 274 -2863 276 -2859
rect 284 -2863 286 -2859
rect 292 -2863 294 -2859
rect 302 -2863 304 -2859
rect 318 -2863 320 -2859
rect 326 -2863 328 -2859
rect 342 -2863 344 -2859
rect 358 -2863 360 -2859
rect 366 -2863 368 -2859
rect 376 -2863 378 -2859
rect 500 -2863 502 -2859
rect 510 -2863 512 -2859
rect 526 -2863 528 -2859
rect 536 -2863 538 -2859
rect 552 -2863 554 -2859
rect 562 -2863 564 -2859
rect 570 -2863 572 -2859
rect 580 -2863 582 -2859
rect 596 -2863 598 -2859
rect 604 -2863 606 -2859
rect 614 -2863 616 -2859
rect 630 -2863 632 -2859
rect 640 -2863 642 -2859
rect 648 -2863 650 -2859
rect 658 -2863 660 -2859
rect 674 -2863 676 -2859
rect 682 -2863 684 -2859
rect 698 -2863 700 -2859
rect 714 -2863 716 -2859
rect 722 -2863 724 -2859
rect 732 -2863 734 -2859
rect 858 -2863 860 -2859
rect 868 -2863 870 -2859
rect 884 -2863 886 -2859
rect 894 -2863 896 -2859
rect 910 -2863 912 -2859
rect 920 -2863 922 -2859
rect 928 -2863 930 -2859
rect 938 -2863 940 -2859
rect 954 -2863 956 -2859
rect 962 -2863 964 -2859
rect 972 -2863 974 -2859
rect 988 -2863 990 -2859
rect 998 -2863 1000 -2859
rect 1006 -2863 1008 -2859
rect 1016 -2863 1018 -2859
rect 1032 -2863 1034 -2859
rect 1040 -2863 1042 -2859
rect 1056 -2863 1058 -2859
rect 1072 -2863 1074 -2859
rect 1080 -2863 1082 -2859
rect 1090 -2863 1092 -2859
rect 1216 -2863 1218 -2859
rect 1226 -2863 1228 -2859
rect 1242 -2863 1244 -2859
rect 1252 -2863 1254 -2859
rect 1268 -2863 1270 -2859
rect 1278 -2863 1280 -2859
rect 1286 -2863 1288 -2859
rect 1296 -2863 1298 -2859
rect 1312 -2863 1314 -2859
rect 1320 -2863 1322 -2859
rect 1330 -2863 1332 -2859
rect 1346 -2863 1348 -2859
rect 1356 -2863 1358 -2859
rect 1364 -2863 1366 -2859
rect 1374 -2863 1376 -2859
rect 1390 -2863 1392 -2859
rect 1398 -2863 1400 -2859
rect 1414 -2863 1416 -2859
rect 1430 -2863 1432 -2859
rect 1438 -2863 1440 -2859
rect 1448 -2863 1450 -2859
rect -1554 -2982 -1552 -2978
rect -1544 -2982 -1542 -2978
rect -1528 -2982 -1526 -2978
rect -1520 -2982 -1518 -2978
rect -1504 -2982 -1502 -2978
rect -1496 -2982 -1494 -2978
rect -1486 -2982 -1484 -2978
rect -1478 -2982 -1476 -2978
rect -1462 -2982 -1460 -2978
rect -1454 -2982 -1452 -2978
rect -1444 -2982 -1442 -2978
rect -1436 -2982 -1434 -2978
rect -1420 -2982 -1418 -2978
rect -1412 -2982 -1410 -2978
rect -1402 -2982 -1400 -2978
rect -1394 -2982 -1392 -2978
rect -1378 -2982 -1376 -2978
rect -1370 -2982 -1368 -2978
rect -1229 -2982 -1227 -2978
rect -1219 -2982 -1217 -2978
rect -1203 -2982 -1201 -2978
rect -1195 -2982 -1193 -2978
rect -1179 -2982 -1177 -2978
rect -1171 -2982 -1169 -2978
rect -1161 -2982 -1159 -2978
rect -1153 -2982 -1151 -2978
rect -1137 -2982 -1135 -2978
rect -1129 -2982 -1127 -2978
rect -1119 -2982 -1117 -2978
rect -1111 -2982 -1109 -2978
rect -1095 -2982 -1093 -2978
rect -1087 -2982 -1085 -2978
rect -1077 -2982 -1075 -2978
rect -1069 -2982 -1067 -2978
rect -1053 -2982 -1051 -2978
rect -1045 -2982 -1043 -2978
rect -930 -2982 -928 -2978
rect -920 -2982 -918 -2978
rect -904 -2982 -902 -2978
rect -896 -2982 -894 -2978
rect -880 -2982 -878 -2978
rect -872 -2982 -870 -2978
rect -862 -2982 -860 -2978
rect -854 -2982 -852 -2978
rect -838 -2982 -836 -2978
rect -830 -2982 -828 -2978
rect -820 -2982 -818 -2978
rect -812 -2982 -810 -2978
rect -796 -2982 -794 -2978
rect -788 -2982 -786 -2978
rect -778 -2982 -776 -2978
rect -770 -2982 -768 -2978
rect -754 -2982 -752 -2978
rect -746 -2982 -744 -2978
rect -572 -2982 -570 -2978
rect -562 -2982 -560 -2978
rect -546 -2982 -544 -2978
rect -538 -2982 -536 -2978
rect -522 -2982 -520 -2978
rect -514 -2982 -512 -2978
rect -504 -2982 -502 -2978
rect -496 -2982 -494 -2978
rect -480 -2982 -478 -2978
rect -472 -2982 -470 -2978
rect -462 -2982 -460 -2978
rect -454 -2982 -452 -2978
rect -438 -2982 -436 -2978
rect -430 -2982 -428 -2978
rect -420 -2982 -418 -2978
rect -412 -2982 -410 -2978
rect -396 -2982 -394 -2978
rect -388 -2982 -386 -2978
rect -214 -2982 -212 -2978
rect -204 -2982 -202 -2978
rect -188 -2982 -186 -2978
rect -180 -2982 -178 -2978
rect -164 -2982 -162 -2978
rect -156 -2982 -154 -2978
rect -146 -2982 -144 -2978
rect -138 -2982 -136 -2978
rect -122 -2982 -120 -2978
rect -114 -2982 -112 -2978
rect -104 -2982 -102 -2978
rect -96 -2982 -94 -2978
rect -80 -2982 -78 -2978
rect -72 -2982 -70 -2978
rect -62 -2982 -60 -2978
rect -54 -2982 -52 -2978
rect -38 -2982 -36 -2978
rect -30 -2982 -28 -2978
rect 144 -2982 146 -2978
rect 154 -2982 156 -2978
rect 170 -2982 172 -2978
rect 178 -2982 180 -2978
rect 194 -2982 196 -2978
rect 202 -2982 204 -2978
rect 212 -2982 214 -2978
rect 220 -2982 222 -2978
rect 236 -2982 238 -2978
rect 244 -2982 246 -2978
rect 254 -2982 256 -2978
rect 262 -2982 264 -2978
rect 278 -2982 280 -2978
rect 286 -2982 288 -2978
rect 296 -2982 298 -2978
rect 304 -2982 306 -2978
rect 320 -2982 322 -2978
rect 328 -2982 330 -2978
rect -1554 -3153 -1552 -3149
rect -1544 -3153 -1542 -3149
rect -1528 -3153 -1526 -3149
rect -1520 -3153 -1518 -3149
rect -1504 -3153 -1502 -3149
rect -1496 -3153 -1494 -3149
rect -1486 -3153 -1484 -3149
rect -1478 -3153 -1476 -3149
rect -1462 -3153 -1460 -3149
rect -1454 -3153 -1452 -3149
rect -1444 -3153 -1442 -3149
rect -1436 -3153 -1434 -3149
rect -1420 -3153 -1418 -3149
rect -1412 -3153 -1410 -3149
rect -1402 -3153 -1400 -3149
rect -1394 -3153 -1392 -3149
rect -1378 -3153 -1376 -3149
rect -1370 -3153 -1368 -3149
rect -1229 -3153 -1227 -3149
rect -1219 -3153 -1217 -3149
rect -1203 -3153 -1201 -3149
rect -1195 -3153 -1193 -3149
rect -1179 -3153 -1177 -3149
rect -1171 -3153 -1169 -3149
rect -1161 -3153 -1159 -3149
rect -1153 -3153 -1151 -3149
rect -1137 -3153 -1135 -3149
rect -1129 -3153 -1127 -3149
rect -1119 -3153 -1117 -3149
rect -1111 -3153 -1109 -3149
rect -1095 -3153 -1093 -3149
rect -1087 -3153 -1085 -3149
rect -1077 -3153 -1075 -3149
rect -1069 -3153 -1067 -3149
rect -1053 -3153 -1051 -3149
rect -1045 -3153 -1043 -3149
rect -930 -3153 -928 -3149
rect -920 -3153 -918 -3149
rect -904 -3153 -902 -3149
rect -896 -3153 -894 -3149
rect -880 -3153 -878 -3149
rect -872 -3153 -870 -3149
rect -862 -3153 -860 -3149
rect -854 -3153 -852 -3149
rect -838 -3153 -836 -3149
rect -830 -3153 -828 -3149
rect -820 -3153 -818 -3149
rect -812 -3153 -810 -3149
rect -796 -3153 -794 -3149
rect -788 -3153 -786 -3149
rect -778 -3153 -776 -3149
rect -770 -3153 -768 -3149
rect -754 -3153 -752 -3149
rect -746 -3153 -744 -3149
rect -572 -3153 -570 -3149
rect -562 -3153 -560 -3149
rect -546 -3153 -544 -3149
rect -538 -3153 -536 -3149
rect -522 -3153 -520 -3149
rect -514 -3153 -512 -3149
rect -504 -3153 -502 -3149
rect -496 -3153 -494 -3149
rect -480 -3153 -478 -3149
rect -472 -3153 -470 -3149
rect -462 -3153 -460 -3149
rect -454 -3153 -452 -3149
rect -438 -3153 -436 -3149
rect -430 -3153 -428 -3149
rect -420 -3153 -418 -3149
rect -412 -3153 -410 -3149
rect -396 -3153 -394 -3149
rect -388 -3153 -386 -3149
rect -214 -3153 -212 -3149
rect -204 -3153 -202 -3149
rect -188 -3153 -186 -3149
rect -180 -3153 -178 -3149
rect -164 -3153 -162 -3149
rect -156 -3153 -154 -3149
rect -146 -3153 -144 -3149
rect -138 -3153 -136 -3149
rect -122 -3153 -120 -3149
rect -114 -3153 -112 -3149
rect -104 -3153 -102 -3149
rect -96 -3153 -94 -3149
rect -80 -3153 -78 -3149
rect -72 -3153 -70 -3149
rect -62 -3153 -60 -3149
rect -54 -3153 -52 -3149
rect -38 -3153 -36 -3149
rect -30 -3153 -28 -3149
rect 144 -3153 146 -3149
rect 154 -3153 156 -3149
rect 170 -3153 172 -3149
rect 178 -3153 180 -3149
rect 194 -3153 196 -3149
rect 202 -3153 204 -3149
rect 212 -3153 214 -3149
rect 220 -3153 222 -3149
rect 236 -3153 238 -3149
rect 244 -3153 246 -3149
rect 254 -3153 256 -3149
rect 262 -3153 264 -3149
rect 278 -3153 280 -3149
rect 286 -3153 288 -3149
rect 296 -3153 298 -3149
rect 304 -3153 306 -3149
rect 320 -3153 322 -3149
rect 328 -3153 330 -3149
rect 500 -3153 502 -3149
rect 510 -3153 512 -3149
rect 526 -3153 528 -3149
rect 534 -3153 536 -3149
rect 550 -3153 552 -3149
rect 558 -3153 560 -3149
rect 568 -3153 570 -3149
rect 576 -3153 578 -3149
rect 592 -3153 594 -3149
rect 600 -3153 602 -3149
rect 610 -3153 612 -3149
rect 618 -3153 620 -3149
rect 634 -3153 636 -3149
rect 642 -3153 644 -3149
rect 652 -3153 654 -3149
rect 660 -3153 662 -3149
rect 676 -3153 678 -3149
rect 684 -3153 686 -3149
rect 858 -3153 860 -3149
rect 868 -3153 870 -3149
rect 884 -3153 886 -3149
rect 892 -3153 894 -3149
rect 908 -3153 910 -3149
rect 916 -3153 918 -3149
rect 926 -3153 928 -3149
rect 934 -3153 936 -3149
rect 950 -3153 952 -3149
rect 958 -3153 960 -3149
rect 968 -3153 970 -3149
rect 976 -3153 978 -3149
rect 992 -3153 994 -3149
rect 1000 -3153 1002 -3149
rect 1010 -3153 1012 -3149
rect 1018 -3153 1020 -3149
rect 1034 -3153 1036 -3149
rect 1042 -3153 1044 -3149
rect 1216 -3153 1218 -3149
rect 1226 -3153 1228 -3149
rect 1242 -3153 1244 -3149
rect 1250 -3153 1252 -3149
rect 1266 -3153 1268 -3149
rect 1274 -3153 1276 -3149
rect 1284 -3153 1286 -3149
rect 1292 -3153 1294 -3149
rect 1308 -3153 1310 -3149
rect 1316 -3153 1318 -3149
rect 1326 -3153 1328 -3149
rect 1334 -3153 1336 -3149
rect 1350 -3153 1352 -3149
rect 1358 -3153 1360 -3149
rect 1368 -3153 1370 -3149
rect 1376 -3153 1378 -3149
rect 1392 -3153 1394 -3149
rect 1400 -3153 1402 -3149
rect -1554 -3324 -1552 -3320
rect -1544 -3324 -1542 -3320
rect -1528 -3324 -1526 -3320
rect -1520 -3324 -1518 -3320
rect -1504 -3324 -1502 -3320
rect -1496 -3324 -1494 -3320
rect -1486 -3324 -1484 -3320
rect -1478 -3324 -1476 -3320
rect -1462 -3324 -1460 -3320
rect -1454 -3324 -1452 -3320
rect -1444 -3324 -1442 -3320
rect -1436 -3324 -1434 -3320
rect -1420 -3324 -1418 -3320
rect -1412 -3324 -1410 -3320
rect -1402 -3324 -1400 -3320
rect -1394 -3324 -1392 -3320
rect -1378 -3324 -1376 -3320
rect -1370 -3324 -1368 -3320
rect -1229 -3324 -1227 -3320
rect -1219 -3324 -1217 -3320
rect -1203 -3324 -1201 -3320
rect -1195 -3324 -1193 -3320
rect -1179 -3324 -1177 -3320
rect -1171 -3324 -1169 -3320
rect -1161 -3324 -1159 -3320
rect -1153 -3324 -1151 -3320
rect -1137 -3324 -1135 -3320
rect -1129 -3324 -1127 -3320
rect -1119 -3324 -1117 -3320
rect -1111 -3324 -1109 -3320
rect -1095 -3324 -1093 -3320
rect -1087 -3324 -1085 -3320
rect -1077 -3324 -1075 -3320
rect -1069 -3324 -1067 -3320
rect -1053 -3324 -1051 -3320
rect -1045 -3324 -1043 -3320
rect -930 -3324 -928 -3320
rect -920 -3324 -918 -3320
rect -904 -3324 -902 -3320
rect -896 -3324 -894 -3320
rect -880 -3324 -878 -3320
rect -872 -3324 -870 -3320
rect -862 -3324 -860 -3320
rect -854 -3324 -852 -3320
rect -838 -3324 -836 -3320
rect -830 -3324 -828 -3320
rect -820 -3324 -818 -3320
rect -812 -3324 -810 -3320
rect -796 -3324 -794 -3320
rect -788 -3324 -786 -3320
rect -778 -3324 -776 -3320
rect -770 -3324 -768 -3320
rect -754 -3324 -752 -3320
rect -746 -3324 -744 -3320
rect -572 -3324 -570 -3320
rect -562 -3324 -560 -3320
rect -546 -3324 -544 -3320
rect -538 -3324 -536 -3320
rect -522 -3324 -520 -3320
rect -514 -3324 -512 -3320
rect -504 -3324 -502 -3320
rect -496 -3324 -494 -3320
rect -480 -3324 -478 -3320
rect -472 -3324 -470 -3320
rect -462 -3324 -460 -3320
rect -454 -3324 -452 -3320
rect -438 -3324 -436 -3320
rect -430 -3324 -428 -3320
rect -420 -3324 -418 -3320
rect -412 -3324 -410 -3320
rect -396 -3324 -394 -3320
rect -388 -3324 -386 -3320
rect -214 -3324 -212 -3320
rect -204 -3324 -202 -3320
rect -188 -3324 -186 -3320
rect -180 -3324 -178 -3320
rect -164 -3324 -162 -3320
rect -156 -3324 -154 -3320
rect -146 -3324 -144 -3320
rect -138 -3324 -136 -3320
rect -122 -3324 -120 -3320
rect -114 -3324 -112 -3320
rect -104 -3324 -102 -3320
rect -96 -3324 -94 -3320
rect -80 -3324 -78 -3320
rect -72 -3324 -70 -3320
rect -62 -3324 -60 -3320
rect -54 -3324 -52 -3320
rect -38 -3324 -36 -3320
rect -30 -3324 -28 -3320
rect 144 -3324 146 -3320
rect 154 -3324 156 -3320
rect 170 -3324 172 -3320
rect 178 -3324 180 -3320
rect 194 -3324 196 -3320
rect 202 -3324 204 -3320
rect 212 -3324 214 -3320
rect 220 -3324 222 -3320
rect 236 -3324 238 -3320
rect 244 -3324 246 -3320
rect 254 -3324 256 -3320
rect 262 -3324 264 -3320
rect 278 -3324 280 -3320
rect 286 -3324 288 -3320
rect 296 -3324 298 -3320
rect 304 -3324 306 -3320
rect 320 -3324 322 -3320
rect 328 -3324 330 -3320
rect 500 -3324 502 -3320
rect 510 -3324 512 -3320
rect 526 -3324 528 -3320
rect 534 -3324 536 -3320
rect 550 -3324 552 -3320
rect 558 -3324 560 -3320
rect 568 -3324 570 -3320
rect 576 -3324 578 -3320
rect 592 -3324 594 -3320
rect 600 -3324 602 -3320
rect 610 -3324 612 -3320
rect 618 -3324 620 -3320
rect 634 -3324 636 -3320
rect 642 -3324 644 -3320
rect 652 -3324 654 -3320
rect 660 -3324 662 -3320
rect 676 -3324 678 -3320
rect 684 -3324 686 -3320
rect 858 -3324 860 -3320
rect 868 -3324 870 -3320
rect 884 -3324 886 -3320
rect 892 -3324 894 -3320
rect 908 -3324 910 -3320
rect 916 -3324 918 -3320
rect 926 -3324 928 -3320
rect 934 -3324 936 -3320
rect 950 -3324 952 -3320
rect 958 -3324 960 -3320
rect 968 -3324 970 -3320
rect 976 -3324 978 -3320
rect 992 -3324 994 -3320
rect 1000 -3324 1002 -3320
rect 1010 -3324 1012 -3320
rect 1018 -3324 1020 -3320
rect 1034 -3324 1036 -3320
rect 1042 -3324 1044 -3320
rect 1216 -3324 1218 -3320
rect 1226 -3324 1228 -3320
rect 1242 -3324 1244 -3320
rect 1250 -3324 1252 -3320
rect 1266 -3324 1268 -3320
rect 1274 -3324 1276 -3320
rect 1284 -3324 1286 -3320
rect 1292 -3324 1294 -3320
rect 1308 -3324 1310 -3320
rect 1316 -3324 1318 -3320
rect 1326 -3324 1328 -3320
rect 1334 -3324 1336 -3320
rect 1350 -3324 1352 -3320
rect 1358 -3324 1360 -3320
rect 1368 -3324 1370 -3320
rect 1376 -3324 1378 -3320
rect 1392 -3324 1394 -3320
rect 1400 -3324 1402 -3320
rect -1304 -3435 -1302 -3431
rect -1296 -3435 -1294 -3431
rect -1286 -3435 -1284 -3431
rect -930 -3435 -928 -3431
rect -922 -3435 -920 -3431
rect -912 -3435 -910 -3431
rect -572 -3435 -570 -3431
rect -564 -3435 -562 -3431
rect -554 -3435 -552 -3431
rect -214 -3435 -212 -3431
rect -206 -3435 -204 -3431
rect -196 -3435 -194 -3431
rect 144 -3435 146 -3431
rect 152 -3435 154 -3431
rect 162 -3435 164 -3431
rect 500 -3435 502 -3431
rect 508 -3435 510 -3431
rect 518 -3435 520 -3431
rect 858 -3435 860 -3431
rect 866 -3435 868 -3431
rect 876 -3435 878 -3431
rect 1216 -3435 1218 -3431
rect 1224 -3435 1226 -3431
rect 1234 -3435 1236 -3431
rect -1229 -3594 -1227 -3590
rect -1219 -3594 -1217 -3590
rect -1203 -3594 -1201 -3590
rect -1193 -3594 -1191 -3590
rect -1185 -3594 -1183 -3590
rect -1175 -3594 -1173 -3590
rect -1159 -3594 -1157 -3590
rect -1151 -3594 -1149 -3590
rect -1141 -3594 -1139 -3590
rect -930 -3594 -928 -3590
rect -920 -3594 -918 -3590
rect -904 -3594 -902 -3590
rect -894 -3594 -892 -3590
rect -878 -3594 -876 -3590
rect -868 -3594 -866 -3590
rect -860 -3594 -858 -3590
rect -850 -3594 -848 -3590
rect -834 -3594 -832 -3590
rect -826 -3594 -824 -3590
rect -816 -3594 -814 -3590
rect -800 -3594 -798 -3590
rect -790 -3594 -788 -3590
rect -782 -3594 -780 -3590
rect -772 -3594 -770 -3590
rect -756 -3594 -754 -3590
rect -748 -3594 -746 -3590
rect -732 -3594 -730 -3590
rect -716 -3594 -714 -3590
rect -708 -3594 -706 -3590
rect -698 -3594 -696 -3590
rect -572 -3594 -570 -3590
rect -562 -3594 -560 -3590
rect -546 -3594 -544 -3590
rect -536 -3594 -534 -3590
rect -520 -3594 -518 -3590
rect -510 -3594 -508 -3590
rect -502 -3594 -500 -3590
rect -492 -3594 -490 -3590
rect -476 -3594 -474 -3590
rect -468 -3594 -466 -3590
rect -458 -3594 -456 -3590
rect -442 -3594 -440 -3590
rect -432 -3594 -430 -3590
rect -424 -3594 -422 -3590
rect -414 -3594 -412 -3590
rect -398 -3594 -396 -3590
rect -390 -3594 -388 -3590
rect -374 -3594 -372 -3590
rect -358 -3594 -356 -3590
rect -350 -3594 -348 -3590
rect -340 -3594 -338 -3590
rect -214 -3594 -212 -3590
rect -204 -3594 -202 -3590
rect -188 -3594 -186 -3590
rect -178 -3594 -176 -3590
rect -162 -3594 -160 -3590
rect -152 -3594 -150 -3590
rect -144 -3594 -142 -3590
rect -134 -3594 -132 -3590
rect -118 -3594 -116 -3590
rect -110 -3594 -108 -3590
rect -100 -3594 -98 -3590
rect -84 -3594 -82 -3590
rect -74 -3594 -72 -3590
rect -66 -3594 -64 -3590
rect -56 -3594 -54 -3590
rect -40 -3594 -38 -3590
rect -32 -3594 -30 -3590
rect -16 -3594 -14 -3590
rect 0 -3594 2 -3590
rect 8 -3594 10 -3590
rect 18 -3594 20 -3590
rect 144 -3594 146 -3590
rect 154 -3594 156 -3590
rect 170 -3594 172 -3590
rect 180 -3594 182 -3590
rect 196 -3594 198 -3590
rect 206 -3594 208 -3590
rect 214 -3594 216 -3590
rect 224 -3594 226 -3590
rect 240 -3594 242 -3590
rect 248 -3594 250 -3590
rect 258 -3594 260 -3590
rect 274 -3594 276 -3590
rect 284 -3594 286 -3590
rect 292 -3594 294 -3590
rect 302 -3594 304 -3590
rect 318 -3594 320 -3590
rect 326 -3594 328 -3590
rect 342 -3594 344 -3590
rect 358 -3594 360 -3590
rect 366 -3594 368 -3590
rect 376 -3594 378 -3590
rect 500 -3594 502 -3590
rect 510 -3594 512 -3590
rect 526 -3594 528 -3590
rect 536 -3594 538 -3590
rect 552 -3594 554 -3590
rect 562 -3594 564 -3590
rect 570 -3594 572 -3590
rect 580 -3594 582 -3590
rect 596 -3594 598 -3590
rect 604 -3594 606 -3590
rect 614 -3594 616 -3590
rect 630 -3594 632 -3590
rect 640 -3594 642 -3590
rect 648 -3594 650 -3590
rect 658 -3594 660 -3590
rect 674 -3594 676 -3590
rect 682 -3594 684 -3590
rect 698 -3594 700 -3590
rect 714 -3594 716 -3590
rect 722 -3594 724 -3590
rect 732 -3594 734 -3590
rect 858 -3594 860 -3590
rect 868 -3594 870 -3590
rect 884 -3594 886 -3590
rect 894 -3594 896 -3590
rect 910 -3594 912 -3590
rect 920 -3594 922 -3590
rect 928 -3594 930 -3590
rect 938 -3594 940 -3590
rect 954 -3594 956 -3590
rect 962 -3594 964 -3590
rect 972 -3594 974 -3590
rect 988 -3594 990 -3590
rect 998 -3594 1000 -3590
rect 1006 -3594 1008 -3590
rect 1016 -3594 1018 -3590
rect 1032 -3594 1034 -3590
rect 1040 -3594 1042 -3590
rect 1056 -3594 1058 -3590
rect 1072 -3594 1074 -3590
rect 1080 -3594 1082 -3590
rect 1090 -3594 1092 -3590
rect 1216 -3594 1218 -3590
rect 1226 -3594 1228 -3590
rect 1242 -3594 1244 -3590
rect 1252 -3594 1254 -3590
rect 1268 -3594 1270 -3590
rect 1278 -3594 1280 -3590
rect 1286 -3594 1288 -3590
rect 1296 -3594 1298 -3590
rect 1312 -3594 1314 -3590
rect 1320 -3594 1322 -3590
rect 1330 -3594 1332 -3590
rect 1346 -3594 1348 -3590
rect 1356 -3594 1358 -3590
rect 1364 -3594 1366 -3590
rect 1374 -3594 1376 -3590
rect 1390 -3594 1392 -3590
rect 1398 -3594 1400 -3590
rect 1414 -3594 1416 -3590
rect 1430 -3594 1432 -3590
rect 1438 -3594 1440 -3590
rect 1448 -3594 1450 -3590
rect -1817 -3724 -1815 -3720
rect -1807 -3724 -1805 -3720
rect -1791 -3724 -1789 -3720
rect -1783 -3724 -1781 -3720
rect -1767 -3724 -1765 -3720
rect -1759 -3724 -1757 -3720
rect -1749 -3724 -1747 -3720
rect -1741 -3724 -1739 -3720
rect -1725 -3724 -1723 -3720
rect -1717 -3724 -1715 -3720
rect -1707 -3724 -1705 -3720
rect -1699 -3724 -1697 -3720
rect -1683 -3724 -1681 -3720
rect -1675 -3724 -1673 -3720
rect -1665 -3724 -1663 -3720
rect -1657 -3724 -1655 -3720
rect -1641 -3724 -1639 -3720
rect -1633 -3724 -1631 -3720
rect -1554 -3724 -1552 -3720
rect -1544 -3724 -1542 -3720
rect -1528 -3724 -1526 -3720
rect -1520 -3724 -1518 -3720
rect -1504 -3724 -1502 -3720
rect -1496 -3724 -1494 -3720
rect -1486 -3724 -1484 -3720
rect -1478 -3724 -1476 -3720
rect -1462 -3724 -1460 -3720
rect -1454 -3724 -1452 -3720
rect -1444 -3724 -1442 -3720
rect -1436 -3724 -1434 -3720
rect -1420 -3724 -1418 -3720
rect -1412 -3724 -1410 -3720
rect -1402 -3724 -1400 -3720
rect -1394 -3724 -1392 -3720
rect -1378 -3724 -1376 -3720
rect -1370 -3724 -1368 -3720
rect -1229 -3724 -1227 -3720
rect -1219 -3724 -1217 -3720
rect -1203 -3724 -1201 -3720
rect -1195 -3724 -1193 -3720
rect -1179 -3724 -1177 -3720
rect -1171 -3724 -1169 -3720
rect -1161 -3724 -1159 -3720
rect -1153 -3724 -1151 -3720
rect -1137 -3724 -1135 -3720
rect -1129 -3724 -1127 -3720
rect -1119 -3724 -1117 -3720
rect -1111 -3724 -1109 -3720
rect -1095 -3724 -1093 -3720
rect -1087 -3724 -1085 -3720
rect -1077 -3724 -1075 -3720
rect -1069 -3724 -1067 -3720
rect -1053 -3724 -1051 -3720
rect -1045 -3724 -1043 -3720
rect -929 -3724 -927 -3720
rect -919 -3724 -917 -3720
rect -903 -3724 -901 -3720
rect -895 -3724 -893 -3720
rect -879 -3724 -877 -3720
rect -871 -3724 -869 -3720
rect -861 -3724 -859 -3720
rect -853 -3724 -851 -3720
rect -837 -3724 -835 -3720
rect -829 -3724 -827 -3720
rect -819 -3724 -817 -3720
rect -811 -3724 -809 -3720
rect -795 -3724 -793 -3720
rect -787 -3724 -785 -3720
rect -777 -3724 -775 -3720
rect -769 -3724 -767 -3720
rect -753 -3724 -751 -3720
rect -745 -3724 -743 -3720
rect -572 -3724 -570 -3720
rect -562 -3724 -560 -3720
rect -546 -3724 -544 -3720
rect -538 -3724 -536 -3720
rect -522 -3724 -520 -3720
rect -514 -3724 -512 -3720
rect -504 -3724 -502 -3720
rect -496 -3724 -494 -3720
rect -480 -3724 -478 -3720
rect -472 -3724 -470 -3720
rect -462 -3724 -460 -3720
rect -454 -3724 -452 -3720
rect -438 -3724 -436 -3720
rect -430 -3724 -428 -3720
rect -420 -3724 -418 -3720
rect -412 -3724 -410 -3720
rect -396 -3724 -394 -3720
rect -388 -3724 -386 -3720
rect -214 -3724 -212 -3720
rect -204 -3724 -202 -3720
rect -188 -3724 -186 -3720
rect -180 -3724 -178 -3720
rect -164 -3724 -162 -3720
rect -156 -3724 -154 -3720
rect -146 -3724 -144 -3720
rect -138 -3724 -136 -3720
rect -122 -3724 -120 -3720
rect -114 -3724 -112 -3720
rect -104 -3724 -102 -3720
rect -96 -3724 -94 -3720
rect -80 -3724 -78 -3720
rect -72 -3724 -70 -3720
rect -62 -3724 -60 -3720
rect -54 -3724 -52 -3720
rect -38 -3724 -36 -3720
rect -30 -3724 -28 -3720
rect -1554 -3895 -1552 -3891
rect -1544 -3895 -1542 -3891
rect -1528 -3895 -1526 -3891
rect -1520 -3895 -1518 -3891
rect -1504 -3895 -1502 -3891
rect -1496 -3895 -1494 -3891
rect -1486 -3895 -1484 -3891
rect -1478 -3895 -1476 -3891
rect -1462 -3895 -1460 -3891
rect -1454 -3895 -1452 -3891
rect -1444 -3895 -1442 -3891
rect -1436 -3895 -1434 -3891
rect -1420 -3895 -1418 -3891
rect -1412 -3895 -1410 -3891
rect -1402 -3895 -1400 -3891
rect -1394 -3895 -1392 -3891
rect -1378 -3895 -1376 -3891
rect -1370 -3895 -1368 -3891
rect -1229 -3895 -1227 -3891
rect -1219 -3895 -1217 -3891
rect -1203 -3895 -1201 -3891
rect -1195 -3895 -1193 -3891
rect -1179 -3895 -1177 -3891
rect -1171 -3895 -1169 -3891
rect -1161 -3895 -1159 -3891
rect -1153 -3895 -1151 -3891
rect -1137 -3895 -1135 -3891
rect -1129 -3895 -1127 -3891
rect -1119 -3895 -1117 -3891
rect -1111 -3895 -1109 -3891
rect -1095 -3895 -1093 -3891
rect -1087 -3895 -1085 -3891
rect -1077 -3895 -1075 -3891
rect -1069 -3895 -1067 -3891
rect -1053 -3895 -1051 -3891
rect -1045 -3895 -1043 -3891
rect -929 -3895 -927 -3891
rect -919 -3895 -917 -3891
rect -903 -3895 -901 -3891
rect -895 -3895 -893 -3891
rect -879 -3895 -877 -3891
rect -871 -3895 -869 -3891
rect -861 -3895 -859 -3891
rect -853 -3895 -851 -3891
rect -837 -3895 -835 -3891
rect -829 -3895 -827 -3891
rect -819 -3895 -817 -3891
rect -811 -3895 -809 -3891
rect -795 -3895 -793 -3891
rect -787 -3895 -785 -3891
rect -777 -3895 -775 -3891
rect -769 -3895 -767 -3891
rect -753 -3895 -751 -3891
rect -745 -3895 -743 -3891
rect -572 -3895 -570 -3891
rect -562 -3895 -560 -3891
rect -546 -3895 -544 -3891
rect -538 -3895 -536 -3891
rect -522 -3895 -520 -3891
rect -514 -3895 -512 -3891
rect -504 -3895 -502 -3891
rect -496 -3895 -494 -3891
rect -480 -3895 -478 -3891
rect -472 -3895 -470 -3891
rect -462 -3895 -460 -3891
rect -454 -3895 -452 -3891
rect -438 -3895 -436 -3891
rect -430 -3895 -428 -3891
rect -420 -3895 -418 -3891
rect -412 -3895 -410 -3891
rect -396 -3895 -394 -3891
rect -388 -3895 -386 -3891
rect -214 -3895 -212 -3891
rect -204 -3895 -202 -3891
rect -188 -3895 -186 -3891
rect -180 -3895 -178 -3891
rect -164 -3895 -162 -3891
rect -156 -3895 -154 -3891
rect -146 -3895 -144 -3891
rect -138 -3895 -136 -3891
rect -122 -3895 -120 -3891
rect -114 -3895 -112 -3891
rect -104 -3895 -102 -3891
rect -96 -3895 -94 -3891
rect -80 -3895 -78 -3891
rect -72 -3895 -70 -3891
rect -62 -3895 -60 -3891
rect -54 -3895 -52 -3891
rect -38 -3895 -36 -3891
rect -30 -3895 -28 -3891
rect 144 -3895 146 -3891
rect 154 -3895 156 -3891
rect 170 -3895 172 -3891
rect 178 -3895 180 -3891
rect 194 -3895 196 -3891
rect 202 -3895 204 -3891
rect 212 -3895 214 -3891
rect 220 -3895 222 -3891
rect 236 -3895 238 -3891
rect 244 -3895 246 -3891
rect 254 -3895 256 -3891
rect 262 -3895 264 -3891
rect 278 -3895 280 -3891
rect 286 -3895 288 -3891
rect 296 -3895 298 -3891
rect 304 -3895 306 -3891
rect 320 -3895 322 -3891
rect 328 -3895 330 -3891
rect 500 -3895 502 -3891
rect 510 -3895 512 -3891
rect 526 -3895 528 -3891
rect 534 -3895 536 -3891
rect 550 -3895 552 -3891
rect 558 -3895 560 -3891
rect 568 -3895 570 -3891
rect 576 -3895 578 -3891
rect 592 -3895 594 -3891
rect 600 -3895 602 -3891
rect 610 -3895 612 -3891
rect 618 -3895 620 -3891
rect 634 -3895 636 -3891
rect 642 -3895 644 -3891
rect 652 -3895 654 -3891
rect 660 -3895 662 -3891
rect 676 -3895 678 -3891
rect 684 -3895 686 -3891
rect 858 -3895 860 -3891
rect 868 -3895 870 -3891
rect 884 -3895 886 -3891
rect 892 -3895 894 -3891
rect 908 -3895 910 -3891
rect 916 -3895 918 -3891
rect 926 -3895 928 -3891
rect 934 -3895 936 -3891
rect 950 -3895 952 -3891
rect 958 -3895 960 -3891
rect 968 -3895 970 -3891
rect 976 -3895 978 -3891
rect 992 -3895 994 -3891
rect 1000 -3895 1002 -3891
rect 1010 -3895 1012 -3891
rect 1018 -3895 1020 -3891
rect 1034 -3895 1036 -3891
rect 1042 -3895 1044 -3891
rect 1216 -3895 1218 -3891
rect 1226 -3895 1228 -3891
rect 1242 -3895 1244 -3891
rect 1250 -3895 1252 -3891
rect 1266 -3895 1268 -3891
rect 1274 -3895 1276 -3891
rect 1284 -3895 1286 -3891
rect 1292 -3895 1294 -3891
rect 1308 -3895 1310 -3891
rect 1316 -3895 1318 -3891
rect 1326 -3895 1328 -3891
rect 1334 -3895 1336 -3891
rect 1350 -3895 1352 -3891
rect 1358 -3895 1360 -3891
rect 1368 -3895 1370 -3891
rect 1376 -3895 1378 -3891
rect 1392 -3895 1394 -3891
rect 1400 -3895 1402 -3891
rect -1554 -4070 -1552 -4066
rect -1544 -4070 -1542 -4066
rect -1528 -4070 -1526 -4066
rect -1520 -4070 -1518 -4066
rect -1504 -4070 -1502 -4066
rect -1496 -4070 -1494 -4066
rect -1486 -4070 -1484 -4066
rect -1478 -4070 -1476 -4066
rect -1462 -4070 -1460 -4066
rect -1454 -4070 -1452 -4066
rect -1444 -4070 -1442 -4066
rect -1436 -4070 -1434 -4066
rect -1420 -4070 -1418 -4066
rect -1412 -4070 -1410 -4066
rect -1402 -4070 -1400 -4066
rect -1394 -4070 -1392 -4066
rect -1378 -4070 -1376 -4066
rect -1370 -4070 -1368 -4066
rect -1229 -4070 -1227 -4066
rect -1219 -4070 -1217 -4066
rect -1203 -4070 -1201 -4066
rect -1195 -4070 -1193 -4066
rect -1179 -4070 -1177 -4066
rect -1171 -4070 -1169 -4066
rect -1161 -4070 -1159 -4066
rect -1153 -4070 -1151 -4066
rect -1137 -4070 -1135 -4066
rect -1129 -4070 -1127 -4066
rect -1119 -4070 -1117 -4066
rect -1111 -4070 -1109 -4066
rect -1095 -4070 -1093 -4066
rect -1087 -4070 -1085 -4066
rect -1077 -4070 -1075 -4066
rect -1069 -4070 -1067 -4066
rect -1053 -4070 -1051 -4066
rect -1045 -4070 -1043 -4066
rect -930 -4070 -928 -4066
rect -920 -4070 -918 -4066
rect -904 -4070 -902 -4066
rect -896 -4070 -894 -4066
rect -880 -4070 -878 -4066
rect -872 -4070 -870 -4066
rect -862 -4070 -860 -4066
rect -854 -4070 -852 -4066
rect -838 -4070 -836 -4066
rect -830 -4070 -828 -4066
rect -820 -4070 -818 -4066
rect -812 -4070 -810 -4066
rect -796 -4070 -794 -4066
rect -788 -4070 -786 -4066
rect -778 -4070 -776 -4066
rect -770 -4070 -768 -4066
rect -754 -4070 -752 -4066
rect -746 -4070 -744 -4066
rect -572 -4070 -570 -4066
rect -562 -4070 -560 -4066
rect -546 -4070 -544 -4066
rect -538 -4070 -536 -4066
rect -522 -4070 -520 -4066
rect -514 -4070 -512 -4066
rect -504 -4070 -502 -4066
rect -496 -4070 -494 -4066
rect -480 -4070 -478 -4066
rect -472 -4070 -470 -4066
rect -462 -4070 -460 -4066
rect -454 -4070 -452 -4066
rect -438 -4070 -436 -4066
rect -430 -4070 -428 -4066
rect -420 -4070 -418 -4066
rect -412 -4070 -410 -4066
rect -396 -4070 -394 -4066
rect -388 -4070 -386 -4066
rect -214 -4070 -212 -4066
rect -204 -4070 -202 -4066
rect -188 -4070 -186 -4066
rect -180 -4070 -178 -4066
rect -164 -4070 -162 -4066
rect -156 -4070 -154 -4066
rect -146 -4070 -144 -4066
rect -138 -4070 -136 -4066
rect -122 -4070 -120 -4066
rect -114 -4070 -112 -4066
rect -104 -4070 -102 -4066
rect -96 -4070 -94 -4066
rect -80 -4070 -78 -4066
rect -72 -4070 -70 -4066
rect -62 -4070 -60 -4066
rect -54 -4070 -52 -4066
rect -38 -4070 -36 -4066
rect -30 -4070 -28 -4066
rect 144 -4070 146 -4066
rect 154 -4070 156 -4066
rect 170 -4070 172 -4066
rect 178 -4070 180 -4066
rect 194 -4070 196 -4066
rect 202 -4070 204 -4066
rect 212 -4070 214 -4066
rect 220 -4070 222 -4066
rect 236 -4070 238 -4066
rect 244 -4070 246 -4066
rect 254 -4070 256 -4066
rect 262 -4070 264 -4066
rect 278 -4070 280 -4066
rect 286 -4070 288 -4066
rect 296 -4070 298 -4066
rect 304 -4070 306 -4066
rect 320 -4070 322 -4066
rect 328 -4070 330 -4066
rect 500 -4070 502 -4066
rect 510 -4070 512 -4066
rect 526 -4070 528 -4066
rect 534 -4070 536 -4066
rect 550 -4070 552 -4066
rect 558 -4070 560 -4066
rect 568 -4070 570 -4066
rect 576 -4070 578 -4066
rect 592 -4070 594 -4066
rect 600 -4070 602 -4066
rect 610 -4070 612 -4066
rect 618 -4070 620 -4066
rect 634 -4070 636 -4066
rect 642 -4070 644 -4066
rect 652 -4070 654 -4066
rect 660 -4070 662 -4066
rect 676 -4070 678 -4066
rect 684 -4070 686 -4066
rect 858 -4070 860 -4066
rect 868 -4070 870 -4066
rect 884 -4070 886 -4066
rect 892 -4070 894 -4066
rect 908 -4070 910 -4066
rect 916 -4070 918 -4066
rect 926 -4070 928 -4066
rect 934 -4070 936 -4066
rect 950 -4070 952 -4066
rect 958 -4070 960 -4066
rect 968 -4070 970 -4066
rect 976 -4070 978 -4066
rect 992 -4070 994 -4066
rect 1000 -4070 1002 -4066
rect 1010 -4070 1012 -4066
rect 1018 -4070 1020 -4066
rect 1034 -4070 1036 -4066
rect 1042 -4070 1044 -4066
rect 1216 -4070 1218 -4066
rect 1226 -4070 1228 -4066
rect 1242 -4070 1244 -4066
rect 1250 -4070 1252 -4066
rect 1266 -4070 1268 -4066
rect 1274 -4070 1276 -4066
rect 1284 -4070 1286 -4066
rect 1292 -4070 1294 -4066
rect 1308 -4070 1310 -4066
rect 1316 -4070 1318 -4066
rect 1326 -4070 1328 -4066
rect 1334 -4070 1336 -4066
rect 1350 -4070 1352 -4066
rect 1358 -4070 1360 -4066
rect 1368 -4070 1370 -4066
rect 1376 -4070 1378 -4066
rect 1392 -4070 1394 -4066
rect 1400 -4070 1402 -4066
rect -1304 -4185 -1302 -4181
rect -1296 -4185 -1294 -4181
rect -1286 -4185 -1284 -4181
rect -930 -4185 -928 -4181
rect -922 -4185 -920 -4181
rect -912 -4185 -910 -4181
rect -572 -4185 -570 -4181
rect -564 -4185 -562 -4181
rect -554 -4185 -552 -4181
rect -214 -4185 -212 -4181
rect -206 -4185 -204 -4181
rect -196 -4185 -194 -4181
rect 144 -4185 146 -4181
rect 152 -4185 154 -4181
rect 162 -4185 164 -4181
rect 500 -4185 502 -4181
rect 508 -4185 510 -4181
rect 518 -4185 520 -4181
rect 858 -4185 860 -4181
rect 866 -4185 868 -4181
rect 876 -4185 878 -4181
rect 1216 -4185 1218 -4181
rect 1224 -4185 1226 -4181
rect 1234 -4185 1236 -4181
rect -1229 -4344 -1227 -4340
rect -1219 -4344 -1217 -4340
rect -1203 -4344 -1201 -4340
rect -1193 -4344 -1191 -4340
rect -1185 -4344 -1183 -4340
rect -1175 -4344 -1173 -4340
rect -1159 -4344 -1157 -4340
rect -1151 -4344 -1149 -4340
rect -1141 -4344 -1139 -4340
rect -930 -4344 -928 -4340
rect -920 -4344 -918 -4340
rect -904 -4344 -902 -4340
rect -894 -4344 -892 -4340
rect -878 -4344 -876 -4340
rect -868 -4344 -866 -4340
rect -860 -4344 -858 -4340
rect -850 -4344 -848 -4340
rect -834 -4344 -832 -4340
rect -826 -4344 -824 -4340
rect -816 -4344 -814 -4340
rect -800 -4344 -798 -4340
rect -790 -4344 -788 -4340
rect -782 -4344 -780 -4340
rect -772 -4344 -770 -4340
rect -756 -4344 -754 -4340
rect -748 -4344 -746 -4340
rect -732 -4344 -730 -4340
rect -716 -4344 -714 -4340
rect -708 -4344 -706 -4340
rect -698 -4344 -696 -4340
rect -572 -4344 -570 -4340
rect -562 -4344 -560 -4340
rect -546 -4344 -544 -4340
rect -536 -4344 -534 -4340
rect -520 -4344 -518 -4340
rect -510 -4344 -508 -4340
rect -502 -4344 -500 -4340
rect -492 -4344 -490 -4340
rect -476 -4344 -474 -4340
rect -468 -4344 -466 -4340
rect -458 -4344 -456 -4340
rect -442 -4344 -440 -4340
rect -432 -4344 -430 -4340
rect -424 -4344 -422 -4340
rect -414 -4344 -412 -4340
rect -398 -4344 -396 -4340
rect -390 -4344 -388 -4340
rect -374 -4344 -372 -4340
rect -358 -4344 -356 -4340
rect -350 -4344 -348 -4340
rect -340 -4344 -338 -4340
rect -214 -4344 -212 -4340
rect -204 -4344 -202 -4340
rect -188 -4344 -186 -4340
rect -178 -4344 -176 -4340
rect -162 -4344 -160 -4340
rect -152 -4344 -150 -4340
rect -144 -4344 -142 -4340
rect -134 -4344 -132 -4340
rect -118 -4344 -116 -4340
rect -110 -4344 -108 -4340
rect -100 -4344 -98 -4340
rect -84 -4344 -82 -4340
rect -74 -4344 -72 -4340
rect -66 -4344 -64 -4340
rect -56 -4344 -54 -4340
rect -40 -4344 -38 -4340
rect -32 -4344 -30 -4340
rect -16 -4344 -14 -4340
rect 0 -4344 2 -4340
rect 8 -4344 10 -4340
rect 18 -4344 20 -4340
rect 144 -4344 146 -4340
rect 154 -4344 156 -4340
rect 170 -4344 172 -4340
rect 180 -4344 182 -4340
rect 196 -4344 198 -4340
rect 206 -4344 208 -4340
rect 214 -4344 216 -4340
rect 224 -4344 226 -4340
rect 240 -4344 242 -4340
rect 248 -4344 250 -4340
rect 258 -4344 260 -4340
rect 274 -4344 276 -4340
rect 284 -4344 286 -4340
rect 292 -4344 294 -4340
rect 302 -4344 304 -4340
rect 318 -4344 320 -4340
rect 326 -4344 328 -4340
rect 342 -4344 344 -4340
rect 358 -4344 360 -4340
rect 366 -4344 368 -4340
rect 376 -4344 378 -4340
rect 500 -4344 502 -4340
rect 510 -4344 512 -4340
rect 526 -4344 528 -4340
rect 536 -4344 538 -4340
rect 552 -4344 554 -4340
rect 562 -4344 564 -4340
rect 570 -4344 572 -4340
rect 580 -4344 582 -4340
rect 596 -4344 598 -4340
rect 604 -4344 606 -4340
rect 614 -4344 616 -4340
rect 630 -4344 632 -4340
rect 640 -4344 642 -4340
rect 648 -4344 650 -4340
rect 658 -4344 660 -4340
rect 674 -4344 676 -4340
rect 682 -4344 684 -4340
rect 698 -4344 700 -4340
rect 714 -4344 716 -4340
rect 722 -4344 724 -4340
rect 732 -4344 734 -4340
rect 858 -4344 860 -4340
rect 868 -4344 870 -4340
rect 884 -4344 886 -4340
rect 894 -4344 896 -4340
rect 910 -4344 912 -4340
rect 920 -4344 922 -4340
rect 928 -4344 930 -4340
rect 938 -4344 940 -4340
rect 954 -4344 956 -4340
rect 962 -4344 964 -4340
rect 972 -4344 974 -4340
rect 988 -4344 990 -4340
rect 998 -4344 1000 -4340
rect 1006 -4344 1008 -4340
rect 1016 -4344 1018 -4340
rect 1032 -4344 1034 -4340
rect 1040 -4344 1042 -4340
rect 1056 -4344 1058 -4340
rect 1072 -4344 1074 -4340
rect 1080 -4344 1082 -4340
rect 1090 -4344 1092 -4340
rect 1216 -4344 1218 -4340
rect 1226 -4344 1228 -4340
rect 1242 -4344 1244 -4340
rect 1252 -4344 1254 -4340
rect 1268 -4344 1270 -4340
rect 1278 -4344 1280 -4340
rect 1286 -4344 1288 -4340
rect 1296 -4344 1298 -4340
rect 1312 -4344 1314 -4340
rect 1320 -4344 1322 -4340
rect 1330 -4344 1332 -4340
rect 1346 -4344 1348 -4340
rect 1356 -4344 1358 -4340
rect 1364 -4344 1366 -4340
rect 1374 -4344 1376 -4340
rect 1390 -4344 1392 -4340
rect 1398 -4344 1400 -4340
rect 1414 -4344 1416 -4340
rect 1430 -4344 1432 -4340
rect 1438 -4344 1440 -4340
rect 1448 -4344 1450 -4340
rect -1809 -4467 -1807 -4463
rect -1799 -4467 -1797 -4463
rect -1783 -4467 -1781 -4463
rect -1775 -4467 -1773 -4463
rect -1759 -4467 -1757 -4463
rect -1751 -4467 -1749 -4463
rect -1741 -4467 -1739 -4463
rect -1733 -4467 -1731 -4463
rect -1717 -4467 -1715 -4463
rect -1709 -4467 -1707 -4463
rect -1699 -4467 -1697 -4463
rect -1691 -4467 -1689 -4463
rect -1675 -4467 -1673 -4463
rect -1667 -4467 -1665 -4463
rect -1657 -4467 -1655 -4463
rect -1649 -4467 -1647 -4463
rect -1633 -4467 -1631 -4463
rect -1625 -4467 -1623 -4463
rect -1546 -4467 -1544 -4463
rect -1536 -4467 -1534 -4463
rect -1520 -4467 -1518 -4463
rect -1512 -4467 -1510 -4463
rect -1496 -4467 -1494 -4463
rect -1488 -4467 -1486 -4463
rect -1478 -4467 -1476 -4463
rect -1470 -4467 -1468 -4463
rect -1454 -4467 -1452 -4463
rect -1446 -4467 -1444 -4463
rect -1436 -4467 -1434 -4463
rect -1428 -4467 -1426 -4463
rect -1412 -4467 -1410 -4463
rect -1404 -4467 -1402 -4463
rect -1394 -4467 -1392 -4463
rect -1386 -4467 -1384 -4463
rect -1370 -4467 -1368 -4463
rect -1362 -4467 -1360 -4463
rect -1229 -4467 -1227 -4463
rect -1219 -4467 -1217 -4463
rect -1203 -4467 -1201 -4463
rect -1195 -4467 -1193 -4463
rect -1179 -4467 -1177 -4463
rect -1171 -4467 -1169 -4463
rect -1161 -4467 -1159 -4463
rect -1153 -4467 -1151 -4463
rect -1137 -4467 -1135 -4463
rect -1129 -4467 -1127 -4463
rect -1119 -4467 -1117 -4463
rect -1111 -4467 -1109 -4463
rect -1095 -4467 -1093 -4463
rect -1087 -4467 -1085 -4463
rect -1077 -4467 -1075 -4463
rect -1069 -4467 -1067 -4463
rect -1053 -4467 -1051 -4463
rect -1045 -4467 -1043 -4463
rect -930 -4467 -928 -4463
rect -920 -4467 -918 -4463
rect -904 -4467 -902 -4463
rect -896 -4467 -894 -4463
rect -880 -4467 -878 -4463
rect -872 -4467 -870 -4463
rect -862 -4467 -860 -4463
rect -854 -4467 -852 -4463
rect -838 -4467 -836 -4463
rect -830 -4467 -828 -4463
rect -820 -4467 -818 -4463
rect -812 -4467 -810 -4463
rect -796 -4467 -794 -4463
rect -788 -4467 -786 -4463
rect -778 -4467 -776 -4463
rect -770 -4467 -768 -4463
rect -754 -4467 -752 -4463
rect -746 -4467 -744 -4463
rect -572 -4467 -570 -4463
rect -562 -4467 -560 -4463
rect -546 -4467 -544 -4463
rect -538 -4467 -536 -4463
rect -522 -4467 -520 -4463
rect -514 -4467 -512 -4463
rect -504 -4467 -502 -4463
rect -496 -4467 -494 -4463
rect -480 -4467 -478 -4463
rect -472 -4467 -470 -4463
rect -462 -4467 -460 -4463
rect -454 -4467 -452 -4463
rect -438 -4467 -436 -4463
rect -430 -4467 -428 -4463
rect -420 -4467 -418 -4463
rect -412 -4467 -410 -4463
rect -396 -4467 -394 -4463
rect -388 -4467 -386 -4463
rect -1809 -4638 -1807 -4634
rect -1799 -4638 -1797 -4634
rect -1783 -4638 -1781 -4634
rect -1775 -4638 -1773 -4634
rect -1759 -4638 -1757 -4634
rect -1751 -4638 -1749 -4634
rect -1741 -4638 -1739 -4634
rect -1733 -4638 -1731 -4634
rect -1717 -4638 -1715 -4634
rect -1709 -4638 -1707 -4634
rect -1699 -4638 -1697 -4634
rect -1691 -4638 -1689 -4634
rect -1675 -4638 -1673 -4634
rect -1667 -4638 -1665 -4634
rect -1657 -4638 -1655 -4634
rect -1649 -4638 -1647 -4634
rect -1633 -4638 -1631 -4634
rect -1625 -4638 -1623 -4634
rect -1546 -4638 -1544 -4634
rect -1536 -4638 -1534 -4634
rect -1520 -4638 -1518 -4634
rect -1512 -4638 -1510 -4634
rect -1496 -4638 -1494 -4634
rect -1488 -4638 -1486 -4634
rect -1478 -4638 -1476 -4634
rect -1470 -4638 -1468 -4634
rect -1454 -4638 -1452 -4634
rect -1446 -4638 -1444 -4634
rect -1436 -4638 -1434 -4634
rect -1428 -4638 -1426 -4634
rect -1412 -4638 -1410 -4634
rect -1404 -4638 -1402 -4634
rect -1394 -4638 -1392 -4634
rect -1386 -4638 -1384 -4634
rect -1370 -4638 -1368 -4634
rect -1362 -4638 -1360 -4634
rect -1229 -4638 -1227 -4634
rect -1219 -4638 -1217 -4634
rect -1203 -4638 -1201 -4634
rect -1195 -4638 -1193 -4634
rect -1179 -4638 -1177 -4634
rect -1171 -4638 -1169 -4634
rect -1161 -4638 -1159 -4634
rect -1153 -4638 -1151 -4634
rect -1137 -4638 -1135 -4634
rect -1129 -4638 -1127 -4634
rect -1119 -4638 -1117 -4634
rect -1111 -4638 -1109 -4634
rect -1095 -4638 -1093 -4634
rect -1087 -4638 -1085 -4634
rect -1077 -4638 -1075 -4634
rect -1069 -4638 -1067 -4634
rect -1053 -4638 -1051 -4634
rect -1045 -4638 -1043 -4634
rect -930 -4638 -928 -4634
rect -920 -4638 -918 -4634
rect -904 -4638 -902 -4634
rect -896 -4638 -894 -4634
rect -880 -4638 -878 -4634
rect -872 -4638 -870 -4634
rect -862 -4638 -860 -4634
rect -854 -4638 -852 -4634
rect -838 -4638 -836 -4634
rect -830 -4638 -828 -4634
rect -820 -4638 -818 -4634
rect -812 -4638 -810 -4634
rect -796 -4638 -794 -4634
rect -788 -4638 -786 -4634
rect -778 -4638 -776 -4634
rect -770 -4638 -768 -4634
rect -754 -4638 -752 -4634
rect -746 -4638 -744 -4634
rect -572 -4638 -570 -4634
rect -562 -4638 -560 -4634
rect -546 -4638 -544 -4634
rect -538 -4638 -536 -4634
rect -522 -4638 -520 -4634
rect -514 -4638 -512 -4634
rect -504 -4638 -502 -4634
rect -496 -4638 -494 -4634
rect -480 -4638 -478 -4634
rect -472 -4638 -470 -4634
rect -462 -4638 -460 -4634
rect -454 -4638 -452 -4634
rect -438 -4638 -436 -4634
rect -430 -4638 -428 -4634
rect -420 -4638 -418 -4634
rect -412 -4638 -410 -4634
rect -396 -4638 -394 -4634
rect -388 -4638 -386 -4634
rect -214 -4638 -212 -4634
rect -204 -4638 -202 -4634
rect -188 -4638 -186 -4634
rect -180 -4638 -178 -4634
rect -164 -4638 -162 -4634
rect -156 -4638 -154 -4634
rect -146 -4638 -144 -4634
rect -138 -4638 -136 -4634
rect -122 -4638 -120 -4634
rect -114 -4638 -112 -4634
rect -104 -4638 -102 -4634
rect -96 -4638 -94 -4634
rect -80 -4638 -78 -4634
rect -72 -4638 -70 -4634
rect -62 -4638 -60 -4634
rect -54 -4638 -52 -4634
rect -38 -4638 -36 -4634
rect -30 -4638 -28 -4634
rect 144 -4638 146 -4634
rect 154 -4638 156 -4634
rect 170 -4638 172 -4634
rect 178 -4638 180 -4634
rect 194 -4638 196 -4634
rect 202 -4638 204 -4634
rect 212 -4638 214 -4634
rect 220 -4638 222 -4634
rect 236 -4638 238 -4634
rect 244 -4638 246 -4634
rect 254 -4638 256 -4634
rect 262 -4638 264 -4634
rect 278 -4638 280 -4634
rect 286 -4638 288 -4634
rect 296 -4638 298 -4634
rect 304 -4638 306 -4634
rect 320 -4638 322 -4634
rect 328 -4638 330 -4634
rect 500 -4638 502 -4634
rect 510 -4638 512 -4634
rect 526 -4638 528 -4634
rect 534 -4638 536 -4634
rect 550 -4638 552 -4634
rect 558 -4638 560 -4634
rect 568 -4638 570 -4634
rect 576 -4638 578 -4634
rect 592 -4638 594 -4634
rect 600 -4638 602 -4634
rect 610 -4638 612 -4634
rect 618 -4638 620 -4634
rect 634 -4638 636 -4634
rect 642 -4638 644 -4634
rect 652 -4638 654 -4634
rect 660 -4638 662 -4634
rect 676 -4638 678 -4634
rect 684 -4638 686 -4634
rect 858 -4638 860 -4634
rect 868 -4638 870 -4634
rect 884 -4638 886 -4634
rect 892 -4638 894 -4634
rect 908 -4638 910 -4634
rect 916 -4638 918 -4634
rect 926 -4638 928 -4634
rect 934 -4638 936 -4634
rect 950 -4638 952 -4634
rect 958 -4638 960 -4634
rect 968 -4638 970 -4634
rect 976 -4638 978 -4634
rect 992 -4638 994 -4634
rect 1000 -4638 1002 -4634
rect 1010 -4638 1012 -4634
rect 1018 -4638 1020 -4634
rect 1034 -4638 1036 -4634
rect 1042 -4638 1044 -4634
rect 1216 -4638 1218 -4634
rect 1226 -4638 1228 -4634
rect 1242 -4638 1244 -4634
rect 1250 -4638 1252 -4634
rect 1266 -4638 1268 -4634
rect 1274 -4638 1276 -4634
rect 1284 -4638 1286 -4634
rect 1292 -4638 1294 -4634
rect 1308 -4638 1310 -4634
rect 1316 -4638 1318 -4634
rect 1326 -4638 1328 -4634
rect 1334 -4638 1336 -4634
rect 1350 -4638 1352 -4634
rect 1358 -4638 1360 -4634
rect 1368 -4638 1370 -4634
rect 1376 -4638 1378 -4634
rect 1392 -4638 1394 -4634
rect 1400 -4638 1402 -4634
rect -1546 -4809 -1544 -4805
rect -1536 -4809 -1534 -4805
rect -1520 -4809 -1518 -4805
rect -1512 -4809 -1510 -4805
rect -1496 -4809 -1494 -4805
rect -1488 -4809 -1486 -4805
rect -1478 -4809 -1476 -4805
rect -1470 -4809 -1468 -4805
rect -1454 -4809 -1452 -4805
rect -1446 -4809 -1444 -4805
rect -1436 -4809 -1434 -4805
rect -1428 -4809 -1426 -4805
rect -1412 -4809 -1410 -4805
rect -1404 -4809 -1402 -4805
rect -1394 -4809 -1392 -4805
rect -1386 -4809 -1384 -4805
rect -1370 -4809 -1368 -4805
rect -1362 -4809 -1360 -4805
rect -1229 -4809 -1227 -4805
rect -1219 -4809 -1217 -4805
rect -1203 -4809 -1201 -4805
rect -1195 -4809 -1193 -4805
rect -1179 -4809 -1177 -4805
rect -1171 -4809 -1169 -4805
rect -1161 -4809 -1159 -4805
rect -1153 -4809 -1151 -4805
rect -1137 -4809 -1135 -4805
rect -1129 -4809 -1127 -4805
rect -1119 -4809 -1117 -4805
rect -1111 -4809 -1109 -4805
rect -1095 -4809 -1093 -4805
rect -1087 -4809 -1085 -4805
rect -1077 -4809 -1075 -4805
rect -1069 -4809 -1067 -4805
rect -1053 -4809 -1051 -4805
rect -1045 -4809 -1043 -4805
rect -930 -4809 -928 -4805
rect -920 -4809 -918 -4805
rect -904 -4809 -902 -4805
rect -896 -4809 -894 -4805
rect -880 -4809 -878 -4805
rect -872 -4809 -870 -4805
rect -862 -4809 -860 -4805
rect -854 -4809 -852 -4805
rect -838 -4809 -836 -4805
rect -830 -4809 -828 -4805
rect -820 -4809 -818 -4805
rect -812 -4809 -810 -4805
rect -796 -4809 -794 -4805
rect -788 -4809 -786 -4805
rect -778 -4809 -776 -4805
rect -770 -4809 -768 -4805
rect -754 -4809 -752 -4805
rect -746 -4809 -744 -4805
rect -572 -4809 -570 -4805
rect -562 -4809 -560 -4805
rect -546 -4809 -544 -4805
rect -538 -4809 -536 -4805
rect -522 -4809 -520 -4805
rect -514 -4809 -512 -4805
rect -504 -4809 -502 -4805
rect -496 -4809 -494 -4805
rect -480 -4809 -478 -4805
rect -472 -4809 -470 -4805
rect -462 -4809 -460 -4805
rect -454 -4809 -452 -4805
rect -438 -4809 -436 -4805
rect -430 -4809 -428 -4805
rect -420 -4809 -418 -4805
rect -412 -4809 -410 -4805
rect -396 -4809 -394 -4805
rect -388 -4809 -386 -4805
rect -214 -4809 -212 -4805
rect -204 -4809 -202 -4805
rect -188 -4809 -186 -4805
rect -180 -4809 -178 -4805
rect -164 -4809 -162 -4805
rect -156 -4809 -154 -4805
rect -146 -4809 -144 -4805
rect -138 -4809 -136 -4805
rect -122 -4809 -120 -4805
rect -114 -4809 -112 -4805
rect -104 -4809 -102 -4805
rect -96 -4809 -94 -4805
rect -80 -4809 -78 -4805
rect -72 -4809 -70 -4805
rect -62 -4809 -60 -4805
rect -54 -4809 -52 -4805
rect -38 -4809 -36 -4805
rect -30 -4809 -28 -4805
rect 144 -4809 146 -4805
rect 154 -4809 156 -4805
rect 170 -4809 172 -4805
rect 178 -4809 180 -4805
rect 194 -4809 196 -4805
rect 202 -4809 204 -4805
rect 212 -4809 214 -4805
rect 220 -4809 222 -4805
rect 236 -4809 238 -4805
rect 244 -4809 246 -4805
rect 254 -4809 256 -4805
rect 262 -4809 264 -4805
rect 278 -4809 280 -4805
rect 286 -4809 288 -4805
rect 296 -4809 298 -4805
rect 304 -4809 306 -4805
rect 320 -4809 322 -4805
rect 328 -4809 330 -4805
rect 500 -4809 502 -4805
rect 510 -4809 512 -4805
rect 526 -4809 528 -4805
rect 534 -4809 536 -4805
rect 550 -4809 552 -4805
rect 558 -4809 560 -4805
rect 568 -4809 570 -4805
rect 576 -4809 578 -4805
rect 592 -4809 594 -4805
rect 600 -4809 602 -4805
rect 610 -4809 612 -4805
rect 618 -4809 620 -4805
rect 634 -4809 636 -4805
rect 642 -4809 644 -4805
rect 652 -4809 654 -4805
rect 660 -4809 662 -4805
rect 676 -4809 678 -4805
rect 684 -4809 686 -4805
rect 858 -4809 860 -4805
rect 868 -4809 870 -4805
rect 884 -4809 886 -4805
rect 892 -4809 894 -4805
rect 908 -4809 910 -4805
rect 916 -4809 918 -4805
rect 926 -4809 928 -4805
rect 934 -4809 936 -4805
rect 950 -4809 952 -4805
rect 958 -4809 960 -4805
rect 968 -4809 970 -4805
rect 976 -4809 978 -4805
rect 992 -4809 994 -4805
rect 1000 -4809 1002 -4805
rect 1010 -4809 1012 -4805
rect 1018 -4809 1020 -4805
rect 1034 -4809 1036 -4805
rect 1042 -4809 1044 -4805
rect 1216 -4809 1218 -4805
rect 1226 -4809 1228 -4805
rect 1242 -4809 1244 -4805
rect 1250 -4809 1252 -4805
rect 1266 -4809 1268 -4805
rect 1274 -4809 1276 -4805
rect 1284 -4809 1286 -4805
rect 1292 -4809 1294 -4805
rect 1308 -4809 1310 -4805
rect 1316 -4809 1318 -4805
rect 1326 -4809 1328 -4805
rect 1334 -4809 1336 -4805
rect 1350 -4809 1352 -4805
rect 1358 -4809 1360 -4805
rect 1368 -4809 1370 -4805
rect 1376 -4809 1378 -4805
rect 1392 -4809 1394 -4805
rect 1400 -4809 1402 -4805
rect -1304 -4924 -1302 -4920
rect -1296 -4924 -1294 -4920
rect -1286 -4924 -1284 -4920
rect -930 -4924 -928 -4920
rect -922 -4924 -920 -4920
rect -912 -4924 -910 -4920
rect -572 -4924 -570 -4920
rect -564 -4924 -562 -4920
rect -554 -4924 -552 -4920
rect -214 -4924 -212 -4920
rect -206 -4924 -204 -4920
rect -196 -4924 -194 -4920
rect 144 -4924 146 -4920
rect 152 -4924 154 -4920
rect 162 -4924 164 -4920
rect 500 -4924 502 -4920
rect 508 -4924 510 -4920
rect 518 -4924 520 -4920
rect 858 -4924 860 -4920
rect 866 -4924 868 -4920
rect 876 -4924 878 -4920
rect 1216 -4924 1218 -4920
rect 1224 -4924 1226 -4920
rect 1234 -4924 1236 -4920
rect -1229 -5083 -1227 -5079
rect -1219 -5083 -1217 -5079
rect -1203 -5083 -1201 -5079
rect -1193 -5083 -1191 -5079
rect -1185 -5083 -1183 -5079
rect -1175 -5083 -1173 -5079
rect -1159 -5083 -1157 -5079
rect -1151 -5083 -1149 -5079
rect -1141 -5083 -1139 -5079
rect -930 -5083 -928 -5079
rect -920 -5083 -918 -5079
rect -904 -5083 -902 -5079
rect -894 -5083 -892 -5079
rect -878 -5083 -876 -5079
rect -868 -5083 -866 -5079
rect -860 -5083 -858 -5079
rect -850 -5083 -848 -5079
rect -834 -5083 -832 -5079
rect -826 -5083 -824 -5079
rect -816 -5083 -814 -5079
rect -800 -5083 -798 -5079
rect -790 -5083 -788 -5079
rect -782 -5083 -780 -5079
rect -772 -5083 -770 -5079
rect -756 -5083 -754 -5079
rect -748 -5083 -746 -5079
rect -732 -5083 -730 -5079
rect -716 -5083 -714 -5079
rect -708 -5083 -706 -5079
rect -698 -5083 -696 -5079
rect -572 -5083 -570 -5079
rect -562 -5083 -560 -5079
rect -546 -5083 -544 -5079
rect -536 -5083 -534 -5079
rect -520 -5083 -518 -5079
rect -510 -5083 -508 -5079
rect -502 -5083 -500 -5079
rect -492 -5083 -490 -5079
rect -476 -5083 -474 -5079
rect -468 -5083 -466 -5079
rect -458 -5083 -456 -5079
rect -442 -5083 -440 -5079
rect -432 -5083 -430 -5079
rect -424 -5083 -422 -5079
rect -414 -5083 -412 -5079
rect -398 -5083 -396 -5079
rect -390 -5083 -388 -5079
rect -374 -5083 -372 -5079
rect -358 -5083 -356 -5079
rect -350 -5083 -348 -5079
rect -340 -5083 -338 -5079
rect -214 -5083 -212 -5079
rect -204 -5083 -202 -5079
rect -188 -5083 -186 -5079
rect -178 -5083 -176 -5079
rect -162 -5083 -160 -5079
rect -152 -5083 -150 -5079
rect -144 -5083 -142 -5079
rect -134 -5083 -132 -5079
rect -118 -5083 -116 -5079
rect -110 -5083 -108 -5079
rect -100 -5083 -98 -5079
rect -84 -5083 -82 -5079
rect -74 -5083 -72 -5079
rect -66 -5083 -64 -5079
rect -56 -5083 -54 -5079
rect -40 -5083 -38 -5079
rect -32 -5083 -30 -5079
rect -16 -5083 -14 -5079
rect 0 -5083 2 -5079
rect 8 -5083 10 -5079
rect 18 -5083 20 -5079
rect 144 -5083 146 -5079
rect 154 -5083 156 -5079
rect 170 -5083 172 -5079
rect 180 -5083 182 -5079
rect 196 -5083 198 -5079
rect 206 -5083 208 -5079
rect 214 -5083 216 -5079
rect 224 -5083 226 -5079
rect 240 -5083 242 -5079
rect 248 -5083 250 -5079
rect 258 -5083 260 -5079
rect 274 -5083 276 -5079
rect 284 -5083 286 -5079
rect 292 -5083 294 -5079
rect 302 -5083 304 -5079
rect 318 -5083 320 -5079
rect 326 -5083 328 -5079
rect 342 -5083 344 -5079
rect 358 -5083 360 -5079
rect 366 -5083 368 -5079
rect 376 -5083 378 -5079
rect 500 -5083 502 -5079
rect 510 -5083 512 -5079
rect 526 -5083 528 -5079
rect 536 -5083 538 -5079
rect 552 -5083 554 -5079
rect 562 -5083 564 -5079
rect 570 -5083 572 -5079
rect 580 -5083 582 -5079
rect 596 -5083 598 -5079
rect 604 -5083 606 -5079
rect 614 -5083 616 -5079
rect 630 -5083 632 -5079
rect 640 -5083 642 -5079
rect 648 -5083 650 -5079
rect 658 -5083 660 -5079
rect 674 -5083 676 -5079
rect 682 -5083 684 -5079
rect 698 -5083 700 -5079
rect 714 -5083 716 -5079
rect 722 -5083 724 -5079
rect 732 -5083 734 -5079
rect 858 -5083 860 -5079
rect 868 -5083 870 -5079
rect 884 -5083 886 -5079
rect 894 -5083 896 -5079
rect 910 -5083 912 -5079
rect 920 -5083 922 -5079
rect 928 -5083 930 -5079
rect 938 -5083 940 -5079
rect 954 -5083 956 -5079
rect 962 -5083 964 -5079
rect 972 -5083 974 -5079
rect 988 -5083 990 -5079
rect 998 -5083 1000 -5079
rect 1006 -5083 1008 -5079
rect 1016 -5083 1018 -5079
rect 1032 -5083 1034 -5079
rect 1040 -5083 1042 -5079
rect 1056 -5083 1058 -5079
rect 1072 -5083 1074 -5079
rect 1080 -5083 1082 -5079
rect 1090 -5083 1092 -5079
rect 1216 -5083 1218 -5079
rect 1226 -5083 1228 -5079
rect 1242 -5083 1244 -5079
rect 1252 -5083 1254 -5079
rect 1268 -5083 1270 -5079
rect 1278 -5083 1280 -5079
rect 1286 -5083 1288 -5079
rect 1296 -5083 1298 -5079
rect 1312 -5083 1314 -5079
rect 1320 -5083 1322 -5079
rect 1330 -5083 1332 -5079
rect 1346 -5083 1348 -5079
rect 1356 -5083 1358 -5079
rect 1364 -5083 1366 -5079
rect 1374 -5083 1376 -5079
rect 1390 -5083 1392 -5079
rect 1398 -5083 1400 -5079
rect 1414 -5083 1416 -5079
rect 1430 -5083 1432 -5079
rect 1438 -5083 1440 -5079
rect 1448 -5083 1450 -5079
rect -1805 -5202 -1803 -5198
rect -1795 -5202 -1793 -5198
rect -1779 -5202 -1777 -5198
rect -1771 -5202 -1769 -5198
rect -1755 -5202 -1753 -5198
rect -1747 -5202 -1745 -5198
rect -1737 -5202 -1735 -5198
rect -1729 -5202 -1727 -5198
rect -1713 -5202 -1711 -5198
rect -1705 -5202 -1703 -5198
rect -1695 -5202 -1693 -5198
rect -1687 -5202 -1685 -5198
rect -1671 -5202 -1669 -5198
rect -1663 -5202 -1661 -5198
rect -1653 -5202 -1651 -5198
rect -1645 -5202 -1643 -5198
rect -1629 -5202 -1627 -5198
rect -1621 -5202 -1619 -5198
rect -1542 -5202 -1540 -5198
rect -1532 -5202 -1530 -5198
rect -1516 -5202 -1514 -5198
rect -1508 -5202 -1506 -5198
rect -1492 -5202 -1490 -5198
rect -1484 -5202 -1482 -5198
rect -1474 -5202 -1472 -5198
rect -1466 -5202 -1464 -5198
rect -1450 -5202 -1448 -5198
rect -1442 -5202 -1440 -5198
rect -1432 -5202 -1430 -5198
rect -1424 -5202 -1422 -5198
rect -1408 -5202 -1406 -5198
rect -1400 -5202 -1398 -5198
rect -1390 -5202 -1388 -5198
rect -1382 -5202 -1380 -5198
rect -1366 -5202 -1364 -5198
rect -1358 -5202 -1356 -5198
rect -1229 -5202 -1227 -5198
rect -1219 -5202 -1217 -5198
rect -1203 -5202 -1201 -5198
rect -1195 -5202 -1193 -5198
rect -1179 -5202 -1177 -5198
rect -1171 -5202 -1169 -5198
rect -1161 -5202 -1159 -5198
rect -1153 -5202 -1151 -5198
rect -1137 -5202 -1135 -5198
rect -1129 -5202 -1127 -5198
rect -1119 -5202 -1117 -5198
rect -1111 -5202 -1109 -5198
rect -1095 -5202 -1093 -5198
rect -1087 -5202 -1085 -5198
rect -1077 -5202 -1075 -5198
rect -1069 -5202 -1067 -5198
rect -1053 -5202 -1051 -5198
rect -1045 -5202 -1043 -5198
rect -930 -5202 -928 -5198
rect -920 -5202 -918 -5198
rect -904 -5202 -902 -5198
rect -896 -5202 -894 -5198
rect -880 -5202 -878 -5198
rect -872 -5202 -870 -5198
rect -862 -5202 -860 -5198
rect -854 -5202 -852 -5198
rect -838 -5202 -836 -5198
rect -830 -5202 -828 -5198
rect -820 -5202 -818 -5198
rect -812 -5202 -810 -5198
rect -796 -5202 -794 -5198
rect -788 -5202 -786 -5198
rect -778 -5202 -776 -5198
rect -770 -5202 -768 -5198
rect -754 -5202 -752 -5198
rect -746 -5202 -744 -5198
rect -1805 -5373 -1803 -5369
rect -1795 -5373 -1793 -5369
rect -1779 -5373 -1777 -5369
rect -1771 -5373 -1769 -5369
rect -1755 -5373 -1753 -5369
rect -1747 -5373 -1745 -5369
rect -1737 -5373 -1735 -5369
rect -1729 -5373 -1727 -5369
rect -1713 -5373 -1711 -5369
rect -1705 -5373 -1703 -5369
rect -1695 -5373 -1693 -5369
rect -1687 -5373 -1685 -5369
rect -1671 -5373 -1669 -5369
rect -1663 -5373 -1661 -5369
rect -1653 -5373 -1651 -5369
rect -1645 -5373 -1643 -5369
rect -1629 -5373 -1627 -5369
rect -1621 -5373 -1619 -5369
rect -1542 -5373 -1540 -5369
rect -1532 -5373 -1530 -5369
rect -1516 -5373 -1514 -5369
rect -1508 -5373 -1506 -5369
rect -1492 -5373 -1490 -5369
rect -1484 -5373 -1482 -5369
rect -1474 -5373 -1472 -5369
rect -1466 -5373 -1464 -5369
rect -1450 -5373 -1448 -5369
rect -1442 -5373 -1440 -5369
rect -1432 -5373 -1430 -5369
rect -1424 -5373 -1422 -5369
rect -1408 -5373 -1406 -5369
rect -1400 -5373 -1398 -5369
rect -1390 -5373 -1388 -5369
rect -1382 -5373 -1380 -5369
rect -1366 -5373 -1364 -5369
rect -1358 -5373 -1356 -5369
rect -1229 -5373 -1227 -5369
rect -1219 -5373 -1217 -5369
rect -1203 -5373 -1201 -5369
rect -1195 -5373 -1193 -5369
rect -1179 -5373 -1177 -5369
rect -1171 -5373 -1169 -5369
rect -1161 -5373 -1159 -5369
rect -1153 -5373 -1151 -5369
rect -1137 -5373 -1135 -5369
rect -1129 -5373 -1127 -5369
rect -1119 -5373 -1117 -5369
rect -1111 -5373 -1109 -5369
rect -1095 -5373 -1093 -5369
rect -1087 -5373 -1085 -5369
rect -1077 -5373 -1075 -5369
rect -1069 -5373 -1067 -5369
rect -1053 -5373 -1051 -5369
rect -1045 -5373 -1043 -5369
rect -930 -5373 -928 -5369
rect -920 -5373 -918 -5369
rect -904 -5373 -902 -5369
rect -896 -5373 -894 -5369
rect -880 -5373 -878 -5369
rect -872 -5373 -870 -5369
rect -862 -5373 -860 -5369
rect -854 -5373 -852 -5369
rect -838 -5373 -836 -5369
rect -830 -5373 -828 -5369
rect -820 -5373 -818 -5369
rect -812 -5373 -810 -5369
rect -796 -5373 -794 -5369
rect -788 -5373 -786 -5369
rect -778 -5373 -776 -5369
rect -770 -5373 -768 -5369
rect -754 -5373 -752 -5369
rect -746 -5373 -744 -5369
rect -572 -5373 -570 -5369
rect -562 -5373 -560 -5369
rect -546 -5373 -544 -5369
rect -538 -5373 -536 -5369
rect -522 -5373 -520 -5369
rect -514 -5373 -512 -5369
rect -504 -5373 -502 -5369
rect -496 -5373 -494 -5369
rect -480 -5373 -478 -5369
rect -472 -5373 -470 -5369
rect -462 -5373 -460 -5369
rect -454 -5373 -452 -5369
rect -438 -5373 -436 -5369
rect -430 -5373 -428 -5369
rect -420 -5373 -418 -5369
rect -412 -5373 -410 -5369
rect -396 -5373 -394 -5369
rect -388 -5373 -386 -5369
rect -214 -5373 -212 -5369
rect -204 -5373 -202 -5369
rect -188 -5373 -186 -5369
rect -180 -5373 -178 -5369
rect -164 -5373 -162 -5369
rect -156 -5373 -154 -5369
rect -146 -5373 -144 -5369
rect -138 -5373 -136 -5369
rect -122 -5373 -120 -5369
rect -114 -5373 -112 -5369
rect -104 -5373 -102 -5369
rect -96 -5373 -94 -5369
rect -80 -5373 -78 -5369
rect -72 -5373 -70 -5369
rect -62 -5373 -60 -5369
rect -54 -5373 -52 -5369
rect -38 -5373 -36 -5369
rect -30 -5373 -28 -5369
rect 144 -5373 146 -5369
rect 154 -5373 156 -5369
rect 170 -5373 172 -5369
rect 178 -5373 180 -5369
rect 194 -5373 196 -5369
rect 202 -5373 204 -5369
rect 212 -5373 214 -5369
rect 220 -5373 222 -5369
rect 236 -5373 238 -5369
rect 244 -5373 246 -5369
rect 254 -5373 256 -5369
rect 262 -5373 264 -5369
rect 278 -5373 280 -5369
rect 286 -5373 288 -5369
rect 296 -5373 298 -5369
rect 304 -5373 306 -5369
rect 320 -5373 322 -5369
rect 328 -5373 330 -5369
rect 500 -5373 502 -5369
rect 510 -5373 512 -5369
rect 526 -5373 528 -5369
rect 534 -5373 536 -5369
rect 550 -5373 552 -5369
rect 558 -5373 560 -5369
rect 568 -5373 570 -5369
rect 576 -5373 578 -5369
rect 592 -5373 594 -5369
rect 600 -5373 602 -5369
rect 610 -5373 612 -5369
rect 618 -5373 620 -5369
rect 634 -5373 636 -5369
rect 642 -5373 644 -5369
rect 652 -5373 654 -5369
rect 660 -5373 662 -5369
rect 676 -5373 678 -5369
rect 684 -5373 686 -5369
rect 858 -5373 860 -5369
rect 868 -5373 870 -5369
rect 884 -5373 886 -5369
rect 892 -5373 894 -5369
rect 908 -5373 910 -5369
rect 916 -5373 918 -5369
rect 926 -5373 928 -5369
rect 934 -5373 936 -5369
rect 950 -5373 952 -5369
rect 958 -5373 960 -5369
rect 968 -5373 970 -5369
rect 976 -5373 978 -5369
rect 992 -5373 994 -5369
rect 1000 -5373 1002 -5369
rect 1010 -5373 1012 -5369
rect 1018 -5373 1020 -5369
rect 1034 -5373 1036 -5369
rect 1042 -5373 1044 -5369
rect 1216 -5373 1218 -5369
rect 1226 -5373 1228 -5369
rect 1242 -5373 1244 -5369
rect 1250 -5373 1252 -5369
rect 1266 -5373 1268 -5369
rect 1274 -5373 1276 -5369
rect 1284 -5373 1286 -5369
rect 1292 -5373 1294 -5369
rect 1308 -5373 1310 -5369
rect 1316 -5373 1318 -5369
rect 1326 -5373 1328 -5369
rect 1334 -5373 1336 -5369
rect 1350 -5373 1352 -5369
rect 1358 -5373 1360 -5369
rect 1368 -5373 1370 -5369
rect 1376 -5373 1378 -5369
rect 1392 -5373 1394 -5369
rect 1400 -5373 1402 -5369
rect -1805 -5533 -1803 -5529
rect -1795 -5533 -1793 -5529
rect -1779 -5533 -1777 -5529
rect -1771 -5533 -1769 -5529
rect -1755 -5533 -1753 -5529
rect -1747 -5533 -1745 -5529
rect -1737 -5533 -1735 -5529
rect -1729 -5533 -1727 -5529
rect -1713 -5533 -1711 -5529
rect -1705 -5533 -1703 -5529
rect -1695 -5533 -1693 -5529
rect -1687 -5533 -1685 -5529
rect -1671 -5533 -1669 -5529
rect -1663 -5533 -1661 -5529
rect -1653 -5533 -1651 -5529
rect -1645 -5533 -1643 -5529
rect -1629 -5533 -1627 -5529
rect -1621 -5533 -1619 -5529
rect -1542 -5533 -1540 -5529
rect -1532 -5533 -1530 -5529
rect -1516 -5533 -1514 -5529
rect -1508 -5533 -1506 -5529
rect -1492 -5533 -1490 -5529
rect -1484 -5533 -1482 -5529
rect -1474 -5533 -1472 -5529
rect -1466 -5533 -1464 -5529
rect -1450 -5533 -1448 -5529
rect -1442 -5533 -1440 -5529
rect -1432 -5533 -1430 -5529
rect -1424 -5533 -1422 -5529
rect -1408 -5533 -1406 -5529
rect -1400 -5533 -1398 -5529
rect -1390 -5533 -1388 -5529
rect -1382 -5533 -1380 -5529
rect -1366 -5533 -1364 -5529
rect -1358 -5533 -1356 -5529
rect -1229 -5533 -1227 -5529
rect -1219 -5533 -1217 -5529
rect -1203 -5533 -1201 -5529
rect -1195 -5533 -1193 -5529
rect -1179 -5533 -1177 -5529
rect -1171 -5533 -1169 -5529
rect -1161 -5533 -1159 -5529
rect -1153 -5533 -1151 -5529
rect -1137 -5533 -1135 -5529
rect -1129 -5533 -1127 -5529
rect -1119 -5533 -1117 -5529
rect -1111 -5533 -1109 -5529
rect -1095 -5533 -1093 -5529
rect -1087 -5533 -1085 -5529
rect -1077 -5533 -1075 -5529
rect -1069 -5533 -1067 -5529
rect -1053 -5533 -1051 -5529
rect -1045 -5533 -1043 -5529
rect -930 -5533 -928 -5529
rect -920 -5533 -918 -5529
rect -904 -5533 -902 -5529
rect -896 -5533 -894 -5529
rect -880 -5533 -878 -5529
rect -872 -5533 -870 -5529
rect -862 -5533 -860 -5529
rect -854 -5533 -852 -5529
rect -838 -5533 -836 -5529
rect -830 -5533 -828 -5529
rect -820 -5533 -818 -5529
rect -812 -5533 -810 -5529
rect -796 -5533 -794 -5529
rect -788 -5533 -786 -5529
rect -778 -5533 -776 -5529
rect -770 -5533 -768 -5529
rect -754 -5533 -752 -5529
rect -746 -5533 -744 -5529
rect -572 -5533 -570 -5529
rect -562 -5533 -560 -5529
rect -546 -5533 -544 -5529
rect -538 -5533 -536 -5529
rect -522 -5533 -520 -5529
rect -514 -5533 -512 -5529
rect -504 -5533 -502 -5529
rect -496 -5533 -494 -5529
rect -480 -5533 -478 -5529
rect -472 -5533 -470 -5529
rect -462 -5533 -460 -5529
rect -454 -5533 -452 -5529
rect -438 -5533 -436 -5529
rect -430 -5533 -428 -5529
rect -420 -5533 -418 -5529
rect -412 -5533 -410 -5529
rect -396 -5533 -394 -5529
rect -388 -5533 -386 -5529
rect -214 -5533 -212 -5529
rect -204 -5533 -202 -5529
rect -188 -5533 -186 -5529
rect -180 -5533 -178 -5529
rect -164 -5533 -162 -5529
rect -156 -5533 -154 -5529
rect -146 -5533 -144 -5529
rect -138 -5533 -136 -5529
rect -122 -5533 -120 -5529
rect -114 -5533 -112 -5529
rect -104 -5533 -102 -5529
rect -96 -5533 -94 -5529
rect -80 -5533 -78 -5529
rect -72 -5533 -70 -5529
rect -62 -5533 -60 -5529
rect -54 -5533 -52 -5529
rect -38 -5533 -36 -5529
rect -30 -5533 -28 -5529
rect 144 -5533 146 -5529
rect 154 -5533 156 -5529
rect 170 -5533 172 -5529
rect 178 -5533 180 -5529
rect 194 -5533 196 -5529
rect 202 -5533 204 -5529
rect 212 -5533 214 -5529
rect 220 -5533 222 -5529
rect 236 -5533 238 -5529
rect 244 -5533 246 -5529
rect 254 -5533 256 -5529
rect 262 -5533 264 -5529
rect 278 -5533 280 -5529
rect 286 -5533 288 -5529
rect 296 -5533 298 -5529
rect 304 -5533 306 -5529
rect 320 -5533 322 -5529
rect 328 -5533 330 -5529
rect 500 -5533 502 -5529
rect 510 -5533 512 -5529
rect 526 -5533 528 -5529
rect 534 -5533 536 -5529
rect 550 -5533 552 -5529
rect 558 -5533 560 -5529
rect 568 -5533 570 -5529
rect 576 -5533 578 -5529
rect 592 -5533 594 -5529
rect 600 -5533 602 -5529
rect 610 -5533 612 -5529
rect 618 -5533 620 -5529
rect 634 -5533 636 -5529
rect 642 -5533 644 -5529
rect 652 -5533 654 -5529
rect 660 -5533 662 -5529
rect 676 -5533 678 -5529
rect 684 -5533 686 -5529
rect 858 -5533 860 -5529
rect 868 -5533 870 -5529
rect 884 -5533 886 -5529
rect 892 -5533 894 -5529
rect 908 -5533 910 -5529
rect 916 -5533 918 -5529
rect 926 -5533 928 -5529
rect 934 -5533 936 -5529
rect 950 -5533 952 -5529
rect 958 -5533 960 -5529
rect 968 -5533 970 -5529
rect 976 -5533 978 -5529
rect 992 -5533 994 -5529
rect 1000 -5533 1002 -5529
rect 1010 -5533 1012 -5529
rect 1018 -5533 1020 -5529
rect 1034 -5533 1036 -5529
rect 1042 -5533 1044 -5529
rect 1216 -5533 1218 -5529
rect 1226 -5533 1228 -5529
rect 1242 -5533 1244 -5529
rect 1250 -5533 1252 -5529
rect 1266 -5533 1268 -5529
rect 1274 -5533 1276 -5529
rect 1284 -5533 1286 -5529
rect 1292 -5533 1294 -5529
rect 1308 -5533 1310 -5529
rect 1316 -5533 1318 -5529
rect 1326 -5533 1328 -5529
rect 1334 -5533 1336 -5529
rect 1350 -5533 1352 -5529
rect 1358 -5533 1360 -5529
rect 1368 -5533 1370 -5529
rect 1376 -5533 1378 -5529
rect 1392 -5533 1394 -5529
rect 1400 -5533 1402 -5529
rect -1304 -5647 -1302 -5643
rect -1296 -5647 -1294 -5643
rect -1286 -5647 -1284 -5643
rect -930 -5647 -928 -5643
rect -922 -5647 -920 -5643
rect -912 -5647 -910 -5643
rect -572 -5647 -570 -5643
rect -564 -5647 -562 -5643
rect -554 -5647 -552 -5643
rect -214 -5647 -212 -5643
rect -206 -5647 -204 -5643
rect -196 -5647 -194 -5643
rect 144 -5647 146 -5643
rect 152 -5647 154 -5643
rect 162 -5647 164 -5643
rect 500 -5647 502 -5643
rect 508 -5647 510 -5643
rect 518 -5647 520 -5643
rect 858 -5647 860 -5643
rect 866 -5647 868 -5643
rect 876 -5647 878 -5643
rect 1216 -5647 1218 -5643
rect 1224 -5647 1226 -5643
rect 1234 -5647 1236 -5643
rect -1229 -5806 -1227 -5802
rect -1219 -5806 -1217 -5802
rect -1203 -5806 -1201 -5802
rect -1193 -5806 -1191 -5802
rect -1185 -5806 -1183 -5802
rect -1175 -5806 -1173 -5802
rect -1159 -5806 -1157 -5802
rect -1151 -5806 -1149 -5802
rect -1141 -5806 -1139 -5802
rect -930 -5806 -928 -5802
rect -920 -5806 -918 -5802
rect -904 -5806 -902 -5802
rect -894 -5806 -892 -5802
rect -878 -5806 -876 -5802
rect -868 -5806 -866 -5802
rect -860 -5806 -858 -5802
rect -850 -5806 -848 -5802
rect -834 -5806 -832 -5802
rect -826 -5806 -824 -5802
rect -816 -5806 -814 -5802
rect -800 -5806 -798 -5802
rect -790 -5806 -788 -5802
rect -782 -5806 -780 -5802
rect -772 -5806 -770 -5802
rect -756 -5806 -754 -5802
rect -748 -5806 -746 -5802
rect -732 -5806 -730 -5802
rect -716 -5806 -714 -5802
rect -708 -5806 -706 -5802
rect -698 -5806 -696 -5802
rect -572 -5806 -570 -5802
rect -562 -5806 -560 -5802
rect -546 -5806 -544 -5802
rect -536 -5806 -534 -5802
rect -520 -5806 -518 -5802
rect -510 -5806 -508 -5802
rect -502 -5806 -500 -5802
rect -492 -5806 -490 -5802
rect -476 -5806 -474 -5802
rect -468 -5806 -466 -5802
rect -458 -5806 -456 -5802
rect -442 -5806 -440 -5802
rect -432 -5806 -430 -5802
rect -424 -5806 -422 -5802
rect -414 -5806 -412 -5802
rect -398 -5806 -396 -5802
rect -390 -5806 -388 -5802
rect -374 -5806 -372 -5802
rect -358 -5806 -356 -5802
rect -350 -5806 -348 -5802
rect -340 -5806 -338 -5802
rect -214 -5806 -212 -5802
rect -204 -5806 -202 -5802
rect -188 -5806 -186 -5802
rect -178 -5806 -176 -5802
rect -162 -5806 -160 -5802
rect -152 -5806 -150 -5802
rect -144 -5806 -142 -5802
rect -134 -5806 -132 -5802
rect -118 -5806 -116 -5802
rect -110 -5806 -108 -5802
rect -100 -5806 -98 -5802
rect -84 -5806 -82 -5802
rect -74 -5806 -72 -5802
rect -66 -5806 -64 -5802
rect -56 -5806 -54 -5802
rect -40 -5806 -38 -5802
rect -32 -5806 -30 -5802
rect -16 -5806 -14 -5802
rect 0 -5806 2 -5802
rect 8 -5806 10 -5802
rect 18 -5806 20 -5802
rect 144 -5806 146 -5802
rect 154 -5806 156 -5802
rect 170 -5806 172 -5802
rect 180 -5806 182 -5802
rect 196 -5806 198 -5802
rect 206 -5806 208 -5802
rect 214 -5806 216 -5802
rect 224 -5806 226 -5802
rect 240 -5806 242 -5802
rect 248 -5806 250 -5802
rect 258 -5806 260 -5802
rect 274 -5806 276 -5802
rect 284 -5806 286 -5802
rect 292 -5806 294 -5802
rect 302 -5806 304 -5802
rect 318 -5806 320 -5802
rect 326 -5806 328 -5802
rect 342 -5806 344 -5802
rect 358 -5806 360 -5802
rect 366 -5806 368 -5802
rect 376 -5806 378 -5802
rect 500 -5806 502 -5802
rect 510 -5806 512 -5802
rect 526 -5806 528 -5802
rect 536 -5806 538 -5802
rect 552 -5806 554 -5802
rect 562 -5806 564 -5802
rect 570 -5806 572 -5802
rect 580 -5806 582 -5802
rect 596 -5806 598 -5802
rect 604 -5806 606 -5802
rect 614 -5806 616 -5802
rect 630 -5806 632 -5802
rect 640 -5806 642 -5802
rect 648 -5806 650 -5802
rect 658 -5806 660 -5802
rect 674 -5806 676 -5802
rect 682 -5806 684 -5802
rect 698 -5806 700 -5802
rect 714 -5806 716 -5802
rect 722 -5806 724 -5802
rect 732 -5806 734 -5802
rect 858 -5806 860 -5802
rect 868 -5806 870 -5802
rect 884 -5806 886 -5802
rect 894 -5806 896 -5802
rect 910 -5806 912 -5802
rect 920 -5806 922 -5802
rect 928 -5806 930 -5802
rect 938 -5806 940 -5802
rect 954 -5806 956 -5802
rect 962 -5806 964 -5802
rect 972 -5806 974 -5802
rect 988 -5806 990 -5802
rect 998 -5806 1000 -5802
rect 1006 -5806 1008 -5802
rect 1016 -5806 1018 -5802
rect 1032 -5806 1034 -5802
rect 1040 -5806 1042 -5802
rect 1056 -5806 1058 -5802
rect 1072 -5806 1074 -5802
rect 1080 -5806 1082 -5802
rect 1090 -5806 1092 -5802
rect 1216 -5806 1218 -5802
rect 1226 -5806 1228 -5802
rect 1242 -5806 1244 -5802
rect 1252 -5806 1254 -5802
rect 1268 -5806 1270 -5802
rect 1278 -5806 1280 -5802
rect 1286 -5806 1288 -5802
rect 1296 -5806 1298 -5802
rect 1312 -5806 1314 -5802
rect 1320 -5806 1322 -5802
rect 1330 -5806 1332 -5802
rect 1346 -5806 1348 -5802
rect 1356 -5806 1358 -5802
rect 1364 -5806 1366 -5802
rect 1374 -5806 1376 -5802
rect 1390 -5806 1392 -5802
rect 1398 -5806 1400 -5802
rect 1414 -5806 1416 -5802
rect 1430 -5806 1432 -5802
rect 1438 -5806 1440 -5802
rect 1448 -5806 1450 -5802
rect -1229 -5929 -1227 -5925
rect -1219 -5929 -1217 -5925
rect -1203 -5929 -1201 -5925
rect -1195 -5929 -1193 -5925
rect -1179 -5929 -1177 -5925
rect -1171 -5929 -1169 -5925
rect -1161 -5929 -1159 -5925
rect -1153 -5929 -1151 -5925
rect -1137 -5929 -1135 -5925
rect -1129 -5929 -1127 -5925
rect -1119 -5929 -1117 -5925
rect -1111 -5929 -1109 -5925
rect -1095 -5929 -1093 -5925
rect -1087 -5929 -1085 -5925
rect -1077 -5929 -1075 -5925
rect -1069 -5929 -1067 -5925
rect -1053 -5929 -1051 -5925
rect -1045 -5929 -1043 -5925
rect -930 -5929 -928 -5925
rect -920 -5929 -918 -5925
rect -904 -5929 -902 -5925
rect -896 -5929 -894 -5925
rect -880 -5929 -878 -5925
rect -872 -5929 -870 -5925
rect -862 -5929 -860 -5925
rect -854 -5929 -852 -5925
rect -838 -5929 -836 -5925
rect -830 -5929 -828 -5925
rect -820 -5929 -818 -5925
rect -812 -5929 -810 -5925
rect -796 -5929 -794 -5925
rect -788 -5929 -786 -5925
rect -778 -5929 -776 -5925
rect -770 -5929 -768 -5925
rect -754 -5929 -752 -5925
rect -746 -5929 -744 -5925
rect -572 -5929 -570 -5925
rect -562 -5929 -560 -5925
rect -546 -5929 -544 -5925
rect -538 -5929 -536 -5925
rect -522 -5929 -520 -5925
rect -514 -5929 -512 -5925
rect -504 -5929 -502 -5925
rect -496 -5929 -494 -5925
rect -480 -5929 -478 -5925
rect -472 -5929 -470 -5925
rect -462 -5929 -460 -5925
rect -454 -5929 -452 -5925
rect -438 -5929 -436 -5925
rect -430 -5929 -428 -5925
rect -420 -5929 -418 -5925
rect -412 -5929 -410 -5925
rect -396 -5929 -394 -5925
rect -388 -5929 -386 -5925
rect -214 -5929 -212 -5925
rect -204 -5929 -202 -5925
rect -188 -5929 -186 -5925
rect -180 -5929 -178 -5925
rect -164 -5929 -162 -5925
rect -156 -5929 -154 -5925
rect -146 -5929 -144 -5925
rect -138 -5929 -136 -5925
rect -122 -5929 -120 -5925
rect -114 -5929 -112 -5925
rect -104 -5929 -102 -5925
rect -96 -5929 -94 -5925
rect -80 -5929 -78 -5925
rect -72 -5929 -70 -5925
rect -62 -5929 -60 -5925
rect -54 -5929 -52 -5925
rect -38 -5929 -36 -5925
rect -30 -5929 -28 -5925
rect 144 -5929 146 -5925
rect 154 -5929 156 -5925
rect 170 -5929 172 -5925
rect 178 -5929 180 -5925
rect 194 -5929 196 -5925
rect 202 -5929 204 -5925
rect 212 -5929 214 -5925
rect 220 -5929 222 -5925
rect 236 -5929 238 -5925
rect 244 -5929 246 -5925
rect 254 -5929 256 -5925
rect 262 -5929 264 -5925
rect 278 -5929 280 -5925
rect 286 -5929 288 -5925
rect 296 -5929 298 -5925
rect 304 -5929 306 -5925
rect 320 -5929 322 -5925
rect 328 -5929 330 -5925
rect 500 -5929 502 -5925
rect 510 -5929 512 -5925
rect 526 -5929 528 -5925
rect 534 -5929 536 -5925
rect 550 -5929 552 -5925
rect 558 -5929 560 -5925
rect 568 -5929 570 -5925
rect 576 -5929 578 -5925
rect 592 -5929 594 -5925
rect 600 -5929 602 -5925
rect 610 -5929 612 -5925
rect 618 -5929 620 -5925
rect 634 -5929 636 -5925
rect 642 -5929 644 -5925
rect 652 -5929 654 -5925
rect 660 -5929 662 -5925
rect 676 -5929 678 -5925
rect 684 -5929 686 -5925
rect 858 -5929 860 -5925
rect 868 -5929 870 -5925
rect 884 -5929 886 -5925
rect 892 -5929 894 -5925
rect 908 -5929 910 -5925
rect 916 -5929 918 -5925
rect 926 -5929 928 -5925
rect 934 -5929 936 -5925
rect 950 -5929 952 -5925
rect 958 -5929 960 -5925
rect 968 -5929 970 -5925
rect 976 -5929 978 -5925
rect 992 -5929 994 -5925
rect 1000 -5929 1002 -5925
rect 1010 -5929 1012 -5925
rect 1018 -5929 1020 -5925
rect 1034 -5929 1036 -5925
rect 1042 -5929 1044 -5925
rect 1216 -5929 1218 -5925
rect 1226 -5929 1228 -5925
rect 1242 -5929 1244 -5925
rect 1250 -5929 1252 -5925
rect 1266 -5929 1268 -5925
rect 1274 -5929 1276 -5925
rect 1284 -5929 1286 -5925
rect 1292 -5929 1294 -5925
rect 1308 -5929 1310 -5925
rect 1316 -5929 1318 -5925
rect 1326 -5929 1328 -5925
rect 1334 -5929 1336 -5925
rect 1350 -5929 1352 -5925
rect 1358 -5929 1360 -5925
rect 1368 -5929 1370 -5925
rect 1376 -5929 1378 -5925
rect 1392 -5929 1394 -5925
rect 1400 -5929 1402 -5925
rect 1560 -5929 1562 -5925
rect 1570 -5929 1572 -5925
rect 1586 -5929 1588 -5925
rect 1594 -5929 1596 -5925
rect 1610 -5929 1612 -5925
rect 1618 -5929 1620 -5925
rect 1628 -5929 1630 -5925
rect 1636 -5929 1638 -5925
rect 1652 -5929 1654 -5925
rect 1660 -5929 1662 -5925
rect 1670 -5929 1672 -5925
rect 1678 -5929 1680 -5925
rect 1694 -5929 1696 -5925
rect 1702 -5929 1704 -5925
rect 1712 -5929 1714 -5925
rect 1720 -5929 1722 -5925
rect 1736 -5929 1738 -5925
rect 1744 -5929 1746 -5925
<< ptransistor >>
rect -1302 -796 -1300 -788
rect -1294 -796 -1292 -788
rect -1284 -796 -1282 -788
rect -931 -796 -929 -788
rect -923 -796 -921 -788
rect -913 -796 -911 -788
rect -572 -796 -570 -788
rect -564 -796 -562 -788
rect -554 -796 -552 -788
rect -214 -796 -212 -788
rect -206 -796 -204 -788
rect -196 -796 -194 -788
rect 143 -796 145 -788
rect 151 -796 153 -788
rect 161 -796 163 -788
rect 500 -796 502 -788
rect 508 -796 510 -788
rect 518 -796 520 -788
rect 858 -796 860 -788
rect 866 -796 868 -788
rect 876 -796 878 -788
rect 1216 -796 1218 -788
rect 1224 -796 1226 -788
rect 1234 -796 1236 -788
rect -1225 -1030 -1223 -1022
rect -1215 -1030 -1213 -1022
rect -1199 -1030 -1197 -1022
rect -1191 -1030 -1189 -1022
rect -1175 -1030 -1173 -1022
rect -1167 -1030 -1165 -1022
rect -1157 -1030 -1155 -1022
rect -1149 -1030 -1147 -1022
rect -1133 -1030 -1131 -1022
rect -1125 -1030 -1123 -1022
rect -1115 -1030 -1113 -1022
rect -1107 -1030 -1105 -1022
rect -1091 -1030 -1089 -1022
rect -1083 -1030 -1081 -1022
rect -1073 -1030 -1071 -1022
rect -1065 -1030 -1063 -1022
rect -1049 -1030 -1047 -1022
rect -1041 -1030 -1039 -1022
rect -930 -1030 -928 -1022
rect -920 -1030 -918 -1022
rect -904 -1030 -902 -1022
rect -896 -1030 -894 -1022
rect -880 -1030 -878 -1022
rect -872 -1030 -870 -1022
rect -862 -1030 -860 -1022
rect -854 -1030 -852 -1022
rect -838 -1030 -836 -1022
rect -830 -1030 -828 -1022
rect -820 -1030 -818 -1022
rect -812 -1030 -810 -1022
rect -796 -1030 -794 -1022
rect -788 -1030 -786 -1022
rect -778 -1030 -776 -1022
rect -770 -1030 -768 -1022
rect -754 -1030 -752 -1022
rect -746 -1030 -744 -1022
rect -572 -1030 -570 -1022
rect -562 -1030 -560 -1022
rect -546 -1030 -544 -1022
rect -538 -1030 -536 -1022
rect -522 -1030 -520 -1022
rect -514 -1030 -512 -1022
rect -504 -1030 -502 -1022
rect -496 -1030 -494 -1022
rect -480 -1030 -478 -1022
rect -472 -1030 -470 -1022
rect -462 -1030 -460 -1022
rect -454 -1030 -452 -1022
rect -438 -1030 -436 -1022
rect -430 -1030 -428 -1022
rect -420 -1030 -418 -1022
rect -412 -1030 -410 -1022
rect -396 -1030 -394 -1022
rect -388 -1030 -386 -1022
rect -214 -1030 -212 -1022
rect -204 -1030 -202 -1022
rect -188 -1030 -186 -1022
rect -180 -1030 -178 -1022
rect -164 -1030 -162 -1022
rect -156 -1030 -154 -1022
rect -146 -1030 -144 -1022
rect -138 -1030 -136 -1022
rect -122 -1030 -120 -1022
rect -114 -1030 -112 -1022
rect -104 -1030 -102 -1022
rect -96 -1030 -94 -1022
rect -80 -1030 -78 -1022
rect -72 -1030 -70 -1022
rect -62 -1030 -60 -1022
rect -54 -1030 -52 -1022
rect -38 -1030 -36 -1022
rect -30 -1030 -28 -1022
rect 144 -1030 146 -1022
rect 154 -1030 156 -1022
rect 170 -1030 172 -1022
rect 178 -1030 180 -1022
rect 194 -1030 196 -1022
rect 202 -1030 204 -1022
rect 212 -1030 214 -1022
rect 220 -1030 222 -1022
rect 236 -1030 238 -1022
rect 244 -1030 246 -1022
rect 254 -1030 256 -1022
rect 262 -1030 264 -1022
rect 278 -1030 280 -1022
rect 286 -1030 288 -1022
rect 296 -1030 298 -1022
rect 304 -1030 306 -1022
rect 320 -1030 322 -1022
rect 328 -1030 330 -1022
rect 500 -1030 502 -1022
rect 510 -1030 512 -1022
rect 526 -1030 528 -1022
rect 534 -1030 536 -1022
rect 550 -1030 552 -1022
rect 558 -1030 560 -1022
rect 568 -1030 570 -1022
rect 576 -1030 578 -1022
rect 592 -1030 594 -1022
rect 600 -1030 602 -1022
rect 610 -1030 612 -1022
rect 618 -1030 620 -1022
rect 634 -1030 636 -1022
rect 642 -1030 644 -1022
rect 652 -1030 654 -1022
rect 660 -1030 662 -1022
rect 676 -1030 678 -1022
rect 684 -1030 686 -1022
rect 858 -1030 860 -1022
rect 868 -1030 870 -1022
rect 884 -1030 886 -1022
rect 892 -1030 894 -1022
rect 908 -1030 910 -1022
rect 916 -1030 918 -1022
rect 926 -1030 928 -1022
rect 934 -1030 936 -1022
rect 950 -1030 952 -1022
rect 958 -1030 960 -1022
rect 968 -1030 970 -1022
rect 976 -1030 978 -1022
rect 992 -1030 994 -1022
rect 1000 -1030 1002 -1022
rect 1010 -1030 1012 -1022
rect 1018 -1030 1020 -1022
rect 1034 -1030 1036 -1022
rect 1042 -1030 1044 -1022
rect -1304 -1146 -1302 -1138
rect -1296 -1146 -1294 -1138
rect -1286 -1146 -1284 -1138
rect -930 -1146 -928 -1138
rect -922 -1146 -920 -1138
rect -912 -1146 -910 -1138
rect -572 -1146 -570 -1138
rect -564 -1146 -562 -1138
rect -554 -1146 -552 -1138
rect -214 -1146 -212 -1138
rect -206 -1146 -204 -1138
rect -196 -1146 -194 -1138
rect 144 -1146 146 -1138
rect 152 -1146 154 -1138
rect 162 -1146 164 -1138
rect 500 -1146 502 -1138
rect 508 -1146 510 -1138
rect 518 -1146 520 -1138
rect 858 -1146 860 -1138
rect 866 -1146 868 -1138
rect 876 -1146 878 -1138
rect 1216 -1146 1218 -1138
rect 1224 -1146 1226 -1138
rect 1234 -1146 1236 -1138
rect -1225 -1310 -1223 -1302
rect -1215 -1310 -1213 -1302
rect -1199 -1310 -1197 -1302
rect -1189 -1310 -1187 -1302
rect -1181 -1310 -1179 -1302
rect -1171 -1310 -1169 -1302
rect -1155 -1310 -1153 -1302
rect -1147 -1310 -1145 -1302
rect -1137 -1310 -1135 -1302
rect -930 -1310 -928 -1302
rect -920 -1310 -918 -1302
rect -904 -1310 -902 -1302
rect -894 -1310 -892 -1302
rect -878 -1310 -876 -1302
rect -868 -1310 -866 -1302
rect -860 -1310 -858 -1302
rect -850 -1310 -848 -1302
rect -834 -1310 -832 -1302
rect -826 -1310 -824 -1302
rect -816 -1310 -814 -1302
rect -800 -1310 -798 -1302
rect -790 -1310 -788 -1302
rect -782 -1310 -780 -1302
rect -772 -1310 -770 -1302
rect -756 -1310 -754 -1302
rect -748 -1310 -746 -1302
rect -732 -1310 -730 -1302
rect -716 -1310 -714 -1302
rect -708 -1310 -706 -1302
rect -698 -1310 -696 -1302
rect -572 -1310 -570 -1302
rect -562 -1310 -560 -1302
rect -546 -1310 -544 -1302
rect -536 -1310 -534 -1302
rect -520 -1310 -518 -1302
rect -510 -1310 -508 -1302
rect -502 -1310 -500 -1302
rect -492 -1310 -490 -1302
rect -476 -1310 -474 -1302
rect -468 -1310 -466 -1302
rect -458 -1310 -456 -1302
rect -442 -1310 -440 -1302
rect -432 -1310 -430 -1302
rect -424 -1310 -422 -1302
rect -414 -1310 -412 -1302
rect -398 -1310 -396 -1302
rect -390 -1310 -388 -1302
rect -374 -1310 -372 -1302
rect -358 -1310 -356 -1302
rect -350 -1310 -348 -1302
rect -340 -1310 -338 -1302
rect -214 -1310 -212 -1302
rect -204 -1310 -202 -1302
rect -188 -1310 -186 -1302
rect -178 -1310 -176 -1302
rect -162 -1310 -160 -1302
rect -152 -1310 -150 -1302
rect -144 -1310 -142 -1302
rect -134 -1310 -132 -1302
rect -118 -1310 -116 -1302
rect -110 -1310 -108 -1302
rect -100 -1310 -98 -1302
rect -84 -1310 -82 -1302
rect -74 -1310 -72 -1302
rect -66 -1310 -64 -1302
rect -56 -1310 -54 -1302
rect -40 -1310 -38 -1302
rect -32 -1310 -30 -1302
rect -16 -1310 -14 -1302
rect 0 -1310 2 -1302
rect 8 -1310 10 -1302
rect 18 -1310 20 -1302
rect 144 -1310 146 -1302
rect 154 -1310 156 -1302
rect 170 -1310 172 -1302
rect 180 -1310 182 -1302
rect 196 -1310 198 -1302
rect 206 -1310 208 -1302
rect 214 -1310 216 -1302
rect 224 -1310 226 -1302
rect 240 -1310 242 -1302
rect 248 -1310 250 -1302
rect 258 -1310 260 -1302
rect 274 -1310 276 -1302
rect 284 -1310 286 -1302
rect 292 -1310 294 -1302
rect 302 -1310 304 -1302
rect 318 -1310 320 -1302
rect 326 -1310 328 -1302
rect 342 -1310 344 -1302
rect 358 -1310 360 -1302
rect 366 -1310 368 -1302
rect 376 -1310 378 -1302
rect 500 -1310 502 -1302
rect 510 -1310 512 -1302
rect 526 -1310 528 -1302
rect 536 -1310 538 -1302
rect 552 -1310 554 -1302
rect 562 -1310 564 -1302
rect 570 -1310 572 -1302
rect 580 -1310 582 -1302
rect 596 -1310 598 -1302
rect 604 -1310 606 -1302
rect 614 -1310 616 -1302
rect 630 -1310 632 -1302
rect 640 -1310 642 -1302
rect 648 -1310 650 -1302
rect 658 -1310 660 -1302
rect 674 -1310 676 -1302
rect 682 -1310 684 -1302
rect 698 -1310 700 -1302
rect 714 -1310 716 -1302
rect 722 -1310 724 -1302
rect 732 -1310 734 -1302
rect 858 -1310 860 -1302
rect 868 -1310 870 -1302
rect 884 -1310 886 -1302
rect 894 -1310 896 -1302
rect 910 -1310 912 -1302
rect 920 -1310 922 -1302
rect 928 -1310 930 -1302
rect 938 -1310 940 -1302
rect 954 -1310 956 -1302
rect 962 -1310 964 -1302
rect 972 -1310 974 -1302
rect 988 -1310 990 -1302
rect 998 -1310 1000 -1302
rect 1006 -1310 1008 -1302
rect 1016 -1310 1018 -1302
rect 1032 -1310 1034 -1302
rect 1040 -1310 1042 -1302
rect 1056 -1310 1058 -1302
rect 1072 -1310 1074 -1302
rect 1080 -1310 1082 -1302
rect 1090 -1310 1092 -1302
rect 1216 -1310 1218 -1302
rect 1226 -1310 1228 -1302
rect 1242 -1310 1244 -1302
rect 1252 -1310 1254 -1302
rect 1260 -1310 1262 -1302
rect 1270 -1310 1272 -1302
rect 1286 -1310 1288 -1302
rect 1294 -1310 1296 -1302
rect 1304 -1310 1306 -1302
rect -1225 -1433 -1223 -1425
rect -1215 -1433 -1213 -1425
rect -1199 -1433 -1197 -1425
rect -1191 -1433 -1189 -1425
rect -1175 -1433 -1173 -1425
rect -1167 -1433 -1165 -1425
rect -1157 -1433 -1155 -1425
rect -1149 -1433 -1147 -1425
rect -1133 -1433 -1131 -1425
rect -1125 -1433 -1123 -1425
rect -1115 -1433 -1113 -1425
rect -1107 -1433 -1105 -1425
rect -1091 -1433 -1089 -1425
rect -1083 -1433 -1081 -1425
rect -1073 -1433 -1071 -1425
rect -1065 -1433 -1063 -1425
rect -1049 -1433 -1047 -1425
rect -1041 -1433 -1039 -1425
rect -930 -1433 -928 -1425
rect -920 -1433 -918 -1425
rect -904 -1433 -902 -1425
rect -896 -1433 -894 -1425
rect -880 -1433 -878 -1425
rect -872 -1433 -870 -1425
rect -862 -1433 -860 -1425
rect -854 -1433 -852 -1425
rect -838 -1433 -836 -1425
rect -830 -1433 -828 -1425
rect -820 -1433 -818 -1425
rect -812 -1433 -810 -1425
rect -796 -1433 -794 -1425
rect -788 -1433 -786 -1425
rect -778 -1433 -776 -1425
rect -770 -1433 -768 -1425
rect -754 -1433 -752 -1425
rect -746 -1433 -744 -1425
rect -572 -1433 -570 -1425
rect -562 -1433 -560 -1425
rect -546 -1433 -544 -1425
rect -538 -1433 -536 -1425
rect -522 -1433 -520 -1425
rect -514 -1433 -512 -1425
rect -504 -1433 -502 -1425
rect -496 -1433 -494 -1425
rect -480 -1433 -478 -1425
rect -472 -1433 -470 -1425
rect -462 -1433 -460 -1425
rect -454 -1433 -452 -1425
rect -438 -1433 -436 -1425
rect -430 -1433 -428 -1425
rect -420 -1433 -418 -1425
rect -412 -1433 -410 -1425
rect -396 -1433 -394 -1425
rect -388 -1433 -386 -1425
rect -214 -1433 -212 -1425
rect -204 -1433 -202 -1425
rect -188 -1433 -186 -1425
rect -180 -1433 -178 -1425
rect -164 -1433 -162 -1425
rect -156 -1433 -154 -1425
rect -146 -1433 -144 -1425
rect -138 -1433 -136 -1425
rect -122 -1433 -120 -1425
rect -114 -1433 -112 -1425
rect -104 -1433 -102 -1425
rect -96 -1433 -94 -1425
rect -80 -1433 -78 -1425
rect -72 -1433 -70 -1425
rect -62 -1433 -60 -1425
rect -54 -1433 -52 -1425
rect -38 -1433 -36 -1425
rect -30 -1433 -28 -1425
rect 144 -1433 146 -1425
rect 154 -1433 156 -1425
rect 170 -1433 172 -1425
rect 178 -1433 180 -1425
rect 194 -1433 196 -1425
rect 202 -1433 204 -1425
rect 212 -1433 214 -1425
rect 220 -1433 222 -1425
rect 236 -1433 238 -1425
rect 244 -1433 246 -1425
rect 254 -1433 256 -1425
rect 262 -1433 264 -1425
rect 278 -1433 280 -1425
rect 286 -1433 288 -1425
rect 296 -1433 298 -1425
rect 304 -1433 306 -1425
rect 320 -1433 322 -1425
rect 328 -1433 330 -1425
rect 500 -1433 502 -1425
rect 510 -1433 512 -1425
rect 526 -1433 528 -1425
rect 534 -1433 536 -1425
rect 550 -1433 552 -1425
rect 558 -1433 560 -1425
rect 568 -1433 570 -1425
rect 576 -1433 578 -1425
rect 592 -1433 594 -1425
rect 600 -1433 602 -1425
rect 610 -1433 612 -1425
rect 618 -1433 620 -1425
rect 634 -1433 636 -1425
rect 642 -1433 644 -1425
rect 652 -1433 654 -1425
rect 660 -1433 662 -1425
rect 676 -1433 678 -1425
rect 684 -1433 686 -1425
rect 858 -1433 860 -1425
rect 868 -1433 870 -1425
rect 884 -1433 886 -1425
rect 892 -1433 894 -1425
rect 908 -1433 910 -1425
rect 916 -1433 918 -1425
rect 926 -1433 928 -1425
rect 934 -1433 936 -1425
rect 950 -1433 952 -1425
rect 958 -1433 960 -1425
rect 968 -1433 970 -1425
rect 976 -1433 978 -1425
rect 992 -1433 994 -1425
rect 1000 -1433 1002 -1425
rect 1010 -1433 1012 -1425
rect 1018 -1433 1020 -1425
rect 1034 -1433 1036 -1425
rect 1042 -1433 1044 -1425
rect -1225 -1604 -1223 -1596
rect -1215 -1604 -1213 -1596
rect -1199 -1604 -1197 -1596
rect -1191 -1604 -1189 -1596
rect -1175 -1604 -1173 -1596
rect -1167 -1604 -1165 -1596
rect -1157 -1604 -1155 -1596
rect -1149 -1604 -1147 -1596
rect -1133 -1604 -1131 -1596
rect -1125 -1604 -1123 -1596
rect -1115 -1604 -1113 -1596
rect -1107 -1604 -1105 -1596
rect -1091 -1604 -1089 -1596
rect -1083 -1604 -1081 -1596
rect -1073 -1604 -1071 -1596
rect -1065 -1604 -1063 -1596
rect -1049 -1604 -1047 -1596
rect -1041 -1604 -1039 -1596
rect -930 -1604 -928 -1596
rect -920 -1604 -918 -1596
rect -904 -1604 -902 -1596
rect -896 -1604 -894 -1596
rect -880 -1604 -878 -1596
rect -872 -1604 -870 -1596
rect -862 -1604 -860 -1596
rect -854 -1604 -852 -1596
rect -838 -1604 -836 -1596
rect -830 -1604 -828 -1596
rect -820 -1604 -818 -1596
rect -812 -1604 -810 -1596
rect -796 -1604 -794 -1596
rect -788 -1604 -786 -1596
rect -778 -1604 -776 -1596
rect -770 -1604 -768 -1596
rect -754 -1604 -752 -1596
rect -746 -1604 -744 -1596
rect -572 -1604 -570 -1596
rect -562 -1604 -560 -1596
rect -546 -1604 -544 -1596
rect -538 -1604 -536 -1596
rect -522 -1604 -520 -1596
rect -514 -1604 -512 -1596
rect -504 -1604 -502 -1596
rect -496 -1604 -494 -1596
rect -480 -1604 -478 -1596
rect -472 -1604 -470 -1596
rect -462 -1604 -460 -1596
rect -454 -1604 -452 -1596
rect -438 -1604 -436 -1596
rect -430 -1604 -428 -1596
rect -420 -1604 -418 -1596
rect -412 -1604 -410 -1596
rect -396 -1604 -394 -1596
rect -388 -1604 -386 -1596
rect -214 -1604 -212 -1596
rect -204 -1604 -202 -1596
rect -188 -1604 -186 -1596
rect -180 -1604 -178 -1596
rect -164 -1604 -162 -1596
rect -156 -1604 -154 -1596
rect -146 -1604 -144 -1596
rect -138 -1604 -136 -1596
rect -122 -1604 -120 -1596
rect -114 -1604 -112 -1596
rect -104 -1604 -102 -1596
rect -96 -1604 -94 -1596
rect -80 -1604 -78 -1596
rect -72 -1604 -70 -1596
rect -62 -1604 -60 -1596
rect -54 -1604 -52 -1596
rect -38 -1604 -36 -1596
rect -30 -1604 -28 -1596
rect 144 -1604 146 -1596
rect 154 -1604 156 -1596
rect 170 -1604 172 -1596
rect 178 -1604 180 -1596
rect 194 -1604 196 -1596
rect 202 -1604 204 -1596
rect 212 -1604 214 -1596
rect 220 -1604 222 -1596
rect 236 -1604 238 -1596
rect 244 -1604 246 -1596
rect 254 -1604 256 -1596
rect 262 -1604 264 -1596
rect 278 -1604 280 -1596
rect 286 -1604 288 -1596
rect 296 -1604 298 -1596
rect 304 -1604 306 -1596
rect 320 -1604 322 -1596
rect 328 -1604 330 -1596
rect 500 -1604 502 -1596
rect 510 -1604 512 -1596
rect 526 -1604 528 -1596
rect 534 -1604 536 -1596
rect 550 -1604 552 -1596
rect 558 -1604 560 -1596
rect 568 -1604 570 -1596
rect 576 -1604 578 -1596
rect 592 -1604 594 -1596
rect 600 -1604 602 -1596
rect 610 -1604 612 -1596
rect 618 -1604 620 -1596
rect 634 -1604 636 -1596
rect 642 -1604 644 -1596
rect 652 -1604 654 -1596
rect 660 -1604 662 -1596
rect 676 -1604 678 -1596
rect 684 -1604 686 -1596
rect 858 -1604 860 -1596
rect 868 -1604 870 -1596
rect 884 -1604 886 -1596
rect 892 -1604 894 -1596
rect 908 -1604 910 -1596
rect 916 -1604 918 -1596
rect 926 -1604 928 -1596
rect 934 -1604 936 -1596
rect 950 -1604 952 -1596
rect 958 -1604 960 -1596
rect 968 -1604 970 -1596
rect 976 -1604 978 -1596
rect 992 -1604 994 -1596
rect 1000 -1604 1002 -1596
rect 1010 -1604 1012 -1596
rect 1018 -1604 1020 -1596
rect 1034 -1604 1036 -1596
rect 1042 -1604 1044 -1596
rect 1216 -1604 1218 -1596
rect 1226 -1604 1228 -1596
rect 1242 -1604 1244 -1596
rect 1250 -1604 1252 -1596
rect 1266 -1604 1268 -1596
rect 1274 -1604 1276 -1596
rect 1284 -1604 1286 -1596
rect 1292 -1604 1294 -1596
rect 1308 -1604 1310 -1596
rect 1316 -1604 1318 -1596
rect 1326 -1604 1328 -1596
rect 1334 -1604 1336 -1596
rect 1350 -1604 1352 -1596
rect 1358 -1604 1360 -1596
rect 1368 -1604 1370 -1596
rect 1376 -1604 1378 -1596
rect 1392 -1604 1394 -1596
rect 1400 -1604 1402 -1596
rect -1554 -1775 -1552 -1767
rect -1544 -1775 -1542 -1767
rect -1528 -1775 -1526 -1767
rect -1520 -1775 -1518 -1767
rect -1504 -1775 -1502 -1767
rect -1496 -1775 -1494 -1767
rect -1486 -1775 -1484 -1767
rect -1478 -1775 -1476 -1767
rect -1462 -1775 -1460 -1767
rect -1454 -1775 -1452 -1767
rect -1444 -1775 -1442 -1767
rect -1436 -1775 -1434 -1767
rect -1420 -1775 -1418 -1767
rect -1412 -1775 -1410 -1767
rect -1402 -1775 -1400 -1767
rect -1394 -1775 -1392 -1767
rect -1378 -1775 -1376 -1767
rect -1370 -1775 -1368 -1767
rect -1225 -1775 -1223 -1767
rect -1215 -1775 -1213 -1767
rect -1199 -1775 -1197 -1767
rect -1191 -1775 -1189 -1767
rect -1175 -1775 -1173 -1767
rect -1167 -1775 -1165 -1767
rect -1157 -1775 -1155 -1767
rect -1149 -1775 -1147 -1767
rect -1133 -1775 -1131 -1767
rect -1125 -1775 -1123 -1767
rect -1115 -1775 -1113 -1767
rect -1107 -1775 -1105 -1767
rect -1091 -1775 -1089 -1767
rect -1083 -1775 -1081 -1767
rect -1073 -1775 -1071 -1767
rect -1065 -1775 -1063 -1767
rect -1049 -1775 -1047 -1767
rect -1041 -1775 -1039 -1767
rect -930 -1775 -928 -1767
rect -920 -1775 -918 -1767
rect -904 -1775 -902 -1767
rect -896 -1775 -894 -1767
rect -880 -1775 -878 -1767
rect -872 -1775 -870 -1767
rect -862 -1775 -860 -1767
rect -854 -1775 -852 -1767
rect -838 -1775 -836 -1767
rect -830 -1775 -828 -1767
rect -820 -1775 -818 -1767
rect -812 -1775 -810 -1767
rect -796 -1775 -794 -1767
rect -788 -1775 -786 -1767
rect -778 -1775 -776 -1767
rect -770 -1775 -768 -1767
rect -754 -1775 -752 -1767
rect -746 -1775 -744 -1767
rect -572 -1775 -570 -1767
rect -562 -1775 -560 -1767
rect -546 -1775 -544 -1767
rect -538 -1775 -536 -1767
rect -522 -1775 -520 -1767
rect -514 -1775 -512 -1767
rect -504 -1775 -502 -1767
rect -496 -1775 -494 -1767
rect -480 -1775 -478 -1767
rect -472 -1775 -470 -1767
rect -462 -1775 -460 -1767
rect -454 -1775 -452 -1767
rect -438 -1775 -436 -1767
rect -430 -1775 -428 -1767
rect -420 -1775 -418 -1767
rect -412 -1775 -410 -1767
rect -396 -1775 -394 -1767
rect -388 -1775 -386 -1767
rect -214 -1775 -212 -1767
rect -204 -1775 -202 -1767
rect -188 -1775 -186 -1767
rect -180 -1775 -178 -1767
rect -164 -1775 -162 -1767
rect -156 -1775 -154 -1767
rect -146 -1775 -144 -1767
rect -138 -1775 -136 -1767
rect -122 -1775 -120 -1767
rect -114 -1775 -112 -1767
rect -104 -1775 -102 -1767
rect -96 -1775 -94 -1767
rect -80 -1775 -78 -1767
rect -72 -1775 -70 -1767
rect -62 -1775 -60 -1767
rect -54 -1775 -52 -1767
rect -38 -1775 -36 -1767
rect -30 -1775 -28 -1767
rect 144 -1775 146 -1767
rect 154 -1775 156 -1767
rect 170 -1775 172 -1767
rect 178 -1775 180 -1767
rect 194 -1775 196 -1767
rect 202 -1775 204 -1767
rect 212 -1775 214 -1767
rect 220 -1775 222 -1767
rect 236 -1775 238 -1767
rect 244 -1775 246 -1767
rect 254 -1775 256 -1767
rect 262 -1775 264 -1767
rect 278 -1775 280 -1767
rect 286 -1775 288 -1767
rect 296 -1775 298 -1767
rect 304 -1775 306 -1767
rect 320 -1775 322 -1767
rect 328 -1775 330 -1767
rect 500 -1775 502 -1767
rect 510 -1775 512 -1767
rect 526 -1775 528 -1767
rect 534 -1775 536 -1767
rect 550 -1775 552 -1767
rect 558 -1775 560 -1767
rect 568 -1775 570 -1767
rect 576 -1775 578 -1767
rect 592 -1775 594 -1767
rect 600 -1775 602 -1767
rect 610 -1775 612 -1767
rect 618 -1775 620 -1767
rect 634 -1775 636 -1767
rect 642 -1775 644 -1767
rect 652 -1775 654 -1767
rect 660 -1775 662 -1767
rect 676 -1775 678 -1767
rect 684 -1775 686 -1767
rect 858 -1775 860 -1767
rect 868 -1775 870 -1767
rect 884 -1775 886 -1767
rect 892 -1775 894 -1767
rect 908 -1775 910 -1767
rect 916 -1775 918 -1767
rect 926 -1775 928 -1767
rect 934 -1775 936 -1767
rect 950 -1775 952 -1767
rect 958 -1775 960 -1767
rect 968 -1775 970 -1767
rect 976 -1775 978 -1767
rect 992 -1775 994 -1767
rect 1000 -1775 1002 -1767
rect 1010 -1775 1012 -1767
rect 1018 -1775 1020 -1767
rect 1034 -1775 1036 -1767
rect 1042 -1775 1044 -1767
rect 1216 -1775 1218 -1767
rect 1226 -1775 1228 -1767
rect 1242 -1775 1244 -1767
rect 1250 -1775 1252 -1767
rect 1266 -1775 1268 -1767
rect 1274 -1775 1276 -1767
rect 1284 -1775 1286 -1767
rect 1292 -1775 1294 -1767
rect 1308 -1775 1310 -1767
rect 1316 -1775 1318 -1767
rect 1326 -1775 1328 -1767
rect 1334 -1775 1336 -1767
rect 1350 -1775 1352 -1767
rect 1358 -1775 1360 -1767
rect 1368 -1775 1370 -1767
rect 1376 -1775 1378 -1767
rect 1392 -1775 1394 -1767
rect 1400 -1775 1402 -1767
rect -1304 -1882 -1302 -1874
rect -1296 -1882 -1294 -1874
rect -1286 -1882 -1284 -1874
rect -930 -1882 -928 -1874
rect -922 -1882 -920 -1874
rect -912 -1882 -910 -1874
rect -572 -1882 -570 -1874
rect -564 -1882 -562 -1874
rect -554 -1882 -552 -1874
rect -214 -1882 -212 -1874
rect -206 -1882 -204 -1874
rect -196 -1882 -194 -1874
rect 144 -1882 146 -1874
rect 152 -1882 154 -1874
rect 162 -1882 164 -1874
rect 500 -1882 502 -1874
rect 508 -1882 510 -1874
rect 518 -1882 520 -1874
rect 858 -1882 860 -1874
rect 866 -1882 868 -1874
rect 876 -1882 878 -1874
rect 1216 -1882 1218 -1874
rect 1224 -1882 1226 -1874
rect 1234 -1882 1236 -1874
rect -1229 -2041 -1227 -2033
rect -1219 -2041 -1217 -2033
rect -1203 -2041 -1201 -2033
rect -1193 -2041 -1191 -2033
rect -1185 -2041 -1183 -2033
rect -1175 -2041 -1173 -2033
rect -1159 -2041 -1157 -2033
rect -1151 -2041 -1149 -2033
rect -1141 -2041 -1139 -2033
rect -930 -2041 -928 -2033
rect -920 -2041 -918 -2033
rect -904 -2041 -902 -2033
rect -894 -2041 -892 -2033
rect -878 -2041 -876 -2033
rect -868 -2041 -866 -2033
rect -860 -2041 -858 -2033
rect -850 -2041 -848 -2033
rect -834 -2041 -832 -2033
rect -826 -2041 -824 -2033
rect -816 -2041 -814 -2033
rect -800 -2041 -798 -2033
rect -790 -2041 -788 -2033
rect -782 -2041 -780 -2033
rect -772 -2041 -770 -2033
rect -756 -2041 -754 -2033
rect -748 -2041 -746 -2033
rect -732 -2041 -730 -2033
rect -716 -2041 -714 -2033
rect -708 -2041 -706 -2033
rect -698 -2041 -696 -2033
rect -572 -2041 -570 -2033
rect -562 -2041 -560 -2033
rect -546 -2041 -544 -2033
rect -536 -2041 -534 -2033
rect -520 -2041 -518 -2033
rect -510 -2041 -508 -2033
rect -502 -2041 -500 -2033
rect -492 -2041 -490 -2033
rect -476 -2041 -474 -2033
rect -468 -2041 -466 -2033
rect -458 -2041 -456 -2033
rect -442 -2041 -440 -2033
rect -432 -2041 -430 -2033
rect -424 -2041 -422 -2033
rect -414 -2041 -412 -2033
rect -398 -2041 -396 -2033
rect -390 -2041 -388 -2033
rect -374 -2041 -372 -2033
rect -358 -2041 -356 -2033
rect -350 -2041 -348 -2033
rect -340 -2041 -338 -2033
rect -214 -2041 -212 -2033
rect -204 -2041 -202 -2033
rect -188 -2041 -186 -2033
rect -178 -2041 -176 -2033
rect -162 -2041 -160 -2033
rect -152 -2041 -150 -2033
rect -144 -2041 -142 -2033
rect -134 -2041 -132 -2033
rect -118 -2041 -116 -2033
rect -110 -2041 -108 -2033
rect -100 -2041 -98 -2033
rect -84 -2041 -82 -2033
rect -74 -2041 -72 -2033
rect -66 -2041 -64 -2033
rect -56 -2041 -54 -2033
rect -40 -2041 -38 -2033
rect -32 -2041 -30 -2033
rect -16 -2041 -14 -2033
rect 0 -2041 2 -2033
rect 8 -2041 10 -2033
rect 18 -2041 20 -2033
rect 144 -2041 146 -2033
rect 154 -2041 156 -2033
rect 170 -2041 172 -2033
rect 180 -2041 182 -2033
rect 196 -2041 198 -2033
rect 206 -2041 208 -2033
rect 214 -2041 216 -2033
rect 224 -2041 226 -2033
rect 240 -2041 242 -2033
rect 248 -2041 250 -2033
rect 258 -2041 260 -2033
rect 274 -2041 276 -2033
rect 284 -2041 286 -2033
rect 292 -2041 294 -2033
rect 302 -2041 304 -2033
rect 318 -2041 320 -2033
rect 326 -2041 328 -2033
rect 342 -2041 344 -2033
rect 358 -2041 360 -2033
rect 366 -2041 368 -2033
rect 376 -2041 378 -2033
rect 500 -2041 502 -2033
rect 510 -2041 512 -2033
rect 526 -2041 528 -2033
rect 536 -2041 538 -2033
rect 552 -2041 554 -2033
rect 562 -2041 564 -2033
rect 570 -2041 572 -2033
rect 580 -2041 582 -2033
rect 596 -2041 598 -2033
rect 604 -2041 606 -2033
rect 614 -2041 616 -2033
rect 630 -2041 632 -2033
rect 640 -2041 642 -2033
rect 648 -2041 650 -2033
rect 658 -2041 660 -2033
rect 674 -2041 676 -2033
rect 682 -2041 684 -2033
rect 698 -2041 700 -2033
rect 714 -2041 716 -2033
rect 722 -2041 724 -2033
rect 732 -2041 734 -2033
rect 858 -2041 860 -2033
rect 868 -2041 870 -2033
rect 884 -2041 886 -2033
rect 894 -2041 896 -2033
rect 910 -2041 912 -2033
rect 920 -2041 922 -2033
rect 928 -2041 930 -2033
rect 938 -2041 940 -2033
rect 954 -2041 956 -2033
rect 962 -2041 964 -2033
rect 972 -2041 974 -2033
rect 988 -2041 990 -2033
rect 998 -2041 1000 -2033
rect 1006 -2041 1008 -2033
rect 1016 -2041 1018 -2033
rect 1032 -2041 1034 -2033
rect 1040 -2041 1042 -2033
rect 1056 -2041 1058 -2033
rect 1072 -2041 1074 -2033
rect 1080 -2041 1082 -2033
rect 1090 -2041 1092 -2033
rect 1216 -2041 1218 -2033
rect 1226 -2041 1228 -2033
rect 1242 -2041 1244 -2033
rect 1252 -2041 1254 -2033
rect 1268 -2041 1270 -2033
rect 1278 -2041 1280 -2033
rect 1286 -2041 1288 -2033
rect 1296 -2041 1298 -2033
rect 1312 -2041 1314 -2033
rect 1320 -2041 1322 -2033
rect 1330 -2041 1332 -2033
rect 1346 -2041 1348 -2033
rect 1356 -2041 1358 -2033
rect 1364 -2041 1366 -2033
rect 1374 -2041 1376 -2033
rect 1390 -2041 1392 -2033
rect 1398 -2041 1400 -2033
rect 1414 -2041 1416 -2033
rect 1430 -2041 1432 -2033
rect 1438 -2041 1440 -2033
rect 1448 -2041 1450 -2033
rect -1229 -2185 -1227 -2177
rect -1219 -2185 -1217 -2177
rect -1203 -2185 -1201 -2177
rect -1195 -2185 -1193 -2177
rect -1179 -2185 -1177 -2177
rect -1171 -2185 -1169 -2177
rect -1161 -2185 -1159 -2177
rect -1153 -2185 -1151 -2177
rect -1137 -2185 -1135 -2177
rect -1129 -2185 -1127 -2177
rect -1119 -2185 -1117 -2177
rect -1111 -2185 -1109 -2177
rect -1095 -2185 -1093 -2177
rect -1087 -2185 -1085 -2177
rect -1077 -2185 -1075 -2177
rect -1069 -2185 -1067 -2177
rect -1053 -2185 -1051 -2177
rect -1045 -2185 -1043 -2177
rect -930 -2185 -928 -2177
rect -920 -2185 -918 -2177
rect -904 -2185 -902 -2177
rect -896 -2185 -894 -2177
rect -880 -2185 -878 -2177
rect -872 -2185 -870 -2177
rect -862 -2185 -860 -2177
rect -854 -2185 -852 -2177
rect -838 -2185 -836 -2177
rect -830 -2185 -828 -2177
rect -820 -2185 -818 -2177
rect -812 -2185 -810 -2177
rect -796 -2185 -794 -2177
rect -788 -2185 -786 -2177
rect -778 -2185 -776 -2177
rect -770 -2185 -768 -2177
rect -754 -2185 -752 -2177
rect -746 -2185 -744 -2177
rect -572 -2185 -570 -2177
rect -562 -2185 -560 -2177
rect -546 -2185 -544 -2177
rect -538 -2185 -536 -2177
rect -522 -2185 -520 -2177
rect -514 -2185 -512 -2177
rect -504 -2185 -502 -2177
rect -496 -2185 -494 -2177
rect -480 -2185 -478 -2177
rect -472 -2185 -470 -2177
rect -462 -2185 -460 -2177
rect -454 -2185 -452 -2177
rect -438 -2185 -436 -2177
rect -430 -2185 -428 -2177
rect -420 -2185 -418 -2177
rect -412 -2185 -410 -2177
rect -396 -2185 -394 -2177
rect -388 -2185 -386 -2177
rect -214 -2185 -212 -2177
rect -204 -2185 -202 -2177
rect -188 -2185 -186 -2177
rect -180 -2185 -178 -2177
rect -164 -2185 -162 -2177
rect -156 -2185 -154 -2177
rect -146 -2185 -144 -2177
rect -138 -2185 -136 -2177
rect -122 -2185 -120 -2177
rect -114 -2185 -112 -2177
rect -104 -2185 -102 -2177
rect -96 -2185 -94 -2177
rect -80 -2185 -78 -2177
rect -72 -2185 -70 -2177
rect -62 -2185 -60 -2177
rect -54 -2185 -52 -2177
rect -38 -2185 -36 -2177
rect -30 -2185 -28 -2177
rect 144 -2185 146 -2177
rect 154 -2185 156 -2177
rect 170 -2185 172 -2177
rect 178 -2185 180 -2177
rect 194 -2185 196 -2177
rect 202 -2185 204 -2177
rect 212 -2185 214 -2177
rect 220 -2185 222 -2177
rect 236 -2185 238 -2177
rect 244 -2185 246 -2177
rect 254 -2185 256 -2177
rect 262 -2185 264 -2177
rect 278 -2185 280 -2177
rect 286 -2185 288 -2177
rect 296 -2185 298 -2177
rect 304 -2185 306 -2177
rect 320 -2185 322 -2177
rect 328 -2185 330 -2177
rect 500 -2185 502 -2177
rect 510 -2185 512 -2177
rect 526 -2185 528 -2177
rect 534 -2185 536 -2177
rect 550 -2185 552 -2177
rect 558 -2185 560 -2177
rect 568 -2185 570 -2177
rect 576 -2185 578 -2177
rect 592 -2185 594 -2177
rect 600 -2185 602 -2177
rect 610 -2185 612 -2177
rect 618 -2185 620 -2177
rect 634 -2185 636 -2177
rect 642 -2185 644 -2177
rect 652 -2185 654 -2177
rect 660 -2185 662 -2177
rect 676 -2185 678 -2177
rect 684 -2185 686 -2177
rect -1554 -2356 -1552 -2348
rect -1544 -2356 -1542 -2348
rect -1528 -2356 -1526 -2348
rect -1520 -2356 -1518 -2348
rect -1504 -2356 -1502 -2348
rect -1496 -2356 -1494 -2348
rect -1486 -2356 -1484 -2348
rect -1478 -2356 -1476 -2348
rect -1462 -2356 -1460 -2348
rect -1454 -2356 -1452 -2348
rect -1444 -2356 -1442 -2348
rect -1436 -2356 -1434 -2348
rect -1420 -2356 -1418 -2348
rect -1412 -2356 -1410 -2348
rect -1402 -2356 -1400 -2348
rect -1394 -2356 -1392 -2348
rect -1378 -2356 -1376 -2348
rect -1370 -2356 -1368 -2348
rect -1229 -2356 -1227 -2348
rect -1219 -2356 -1217 -2348
rect -1203 -2356 -1201 -2348
rect -1195 -2356 -1193 -2348
rect -1179 -2356 -1177 -2348
rect -1171 -2356 -1169 -2348
rect -1161 -2356 -1159 -2348
rect -1153 -2356 -1151 -2348
rect -1137 -2356 -1135 -2348
rect -1129 -2356 -1127 -2348
rect -1119 -2356 -1117 -2348
rect -1111 -2356 -1109 -2348
rect -1095 -2356 -1093 -2348
rect -1087 -2356 -1085 -2348
rect -1077 -2356 -1075 -2348
rect -1069 -2356 -1067 -2348
rect -1053 -2356 -1051 -2348
rect -1045 -2356 -1043 -2348
rect -930 -2356 -928 -2348
rect -920 -2356 -918 -2348
rect -904 -2356 -902 -2348
rect -896 -2356 -894 -2348
rect -880 -2356 -878 -2348
rect -872 -2356 -870 -2348
rect -862 -2356 -860 -2348
rect -854 -2356 -852 -2348
rect -838 -2356 -836 -2348
rect -830 -2356 -828 -2348
rect -820 -2356 -818 -2348
rect -812 -2356 -810 -2348
rect -796 -2356 -794 -2348
rect -788 -2356 -786 -2348
rect -778 -2356 -776 -2348
rect -770 -2356 -768 -2348
rect -754 -2356 -752 -2348
rect -746 -2356 -744 -2348
rect -572 -2356 -570 -2348
rect -562 -2356 -560 -2348
rect -546 -2356 -544 -2348
rect -538 -2356 -536 -2348
rect -522 -2356 -520 -2348
rect -514 -2356 -512 -2348
rect -504 -2356 -502 -2348
rect -496 -2356 -494 -2348
rect -480 -2356 -478 -2348
rect -472 -2356 -470 -2348
rect -462 -2356 -460 -2348
rect -454 -2356 -452 -2348
rect -438 -2356 -436 -2348
rect -430 -2356 -428 -2348
rect -420 -2356 -418 -2348
rect -412 -2356 -410 -2348
rect -396 -2356 -394 -2348
rect -388 -2356 -386 -2348
rect -214 -2356 -212 -2348
rect -204 -2356 -202 -2348
rect -188 -2356 -186 -2348
rect -180 -2356 -178 -2348
rect -164 -2356 -162 -2348
rect -156 -2356 -154 -2348
rect -146 -2356 -144 -2348
rect -138 -2356 -136 -2348
rect -122 -2356 -120 -2348
rect -114 -2356 -112 -2348
rect -104 -2356 -102 -2348
rect -96 -2356 -94 -2348
rect -80 -2356 -78 -2348
rect -72 -2356 -70 -2348
rect -62 -2356 -60 -2348
rect -54 -2356 -52 -2348
rect -38 -2356 -36 -2348
rect -30 -2356 -28 -2348
rect 144 -2356 146 -2348
rect 154 -2356 156 -2348
rect 170 -2356 172 -2348
rect 178 -2356 180 -2348
rect 194 -2356 196 -2348
rect 202 -2356 204 -2348
rect 212 -2356 214 -2348
rect 220 -2356 222 -2348
rect 236 -2356 238 -2348
rect 244 -2356 246 -2348
rect 254 -2356 256 -2348
rect 262 -2356 264 -2348
rect 278 -2356 280 -2348
rect 286 -2356 288 -2348
rect 296 -2356 298 -2348
rect 304 -2356 306 -2348
rect 320 -2356 322 -2348
rect 328 -2356 330 -2348
rect 500 -2356 502 -2348
rect 510 -2356 512 -2348
rect 526 -2356 528 -2348
rect 534 -2356 536 -2348
rect 550 -2356 552 -2348
rect 558 -2356 560 -2348
rect 568 -2356 570 -2348
rect 576 -2356 578 -2348
rect 592 -2356 594 -2348
rect 600 -2356 602 -2348
rect 610 -2356 612 -2348
rect 618 -2356 620 -2348
rect 634 -2356 636 -2348
rect 642 -2356 644 -2348
rect 652 -2356 654 -2348
rect 660 -2356 662 -2348
rect 676 -2356 678 -2348
rect 684 -2356 686 -2348
rect 858 -2356 860 -2348
rect 868 -2356 870 -2348
rect 884 -2356 886 -2348
rect 892 -2356 894 -2348
rect 908 -2356 910 -2348
rect 916 -2356 918 -2348
rect 926 -2356 928 -2348
rect 934 -2356 936 -2348
rect 950 -2356 952 -2348
rect 958 -2356 960 -2348
rect 968 -2356 970 -2348
rect 976 -2356 978 -2348
rect 992 -2356 994 -2348
rect 1000 -2356 1002 -2348
rect 1010 -2356 1012 -2348
rect 1018 -2356 1020 -2348
rect 1034 -2356 1036 -2348
rect 1042 -2356 1044 -2348
rect 1216 -2356 1218 -2348
rect 1226 -2356 1228 -2348
rect 1242 -2356 1244 -2348
rect 1250 -2356 1252 -2348
rect 1266 -2356 1268 -2348
rect 1274 -2356 1276 -2348
rect 1284 -2356 1286 -2348
rect 1292 -2356 1294 -2348
rect 1308 -2356 1310 -2348
rect 1316 -2356 1318 -2348
rect 1326 -2356 1328 -2348
rect 1334 -2356 1336 -2348
rect 1350 -2356 1352 -2348
rect 1358 -2356 1360 -2348
rect 1368 -2356 1370 -2348
rect 1376 -2356 1378 -2348
rect 1392 -2356 1394 -2348
rect 1400 -2356 1402 -2348
rect -1554 -2527 -1552 -2519
rect -1544 -2527 -1542 -2519
rect -1528 -2527 -1526 -2519
rect -1520 -2527 -1518 -2519
rect -1504 -2527 -1502 -2519
rect -1496 -2527 -1494 -2519
rect -1486 -2527 -1484 -2519
rect -1478 -2527 -1476 -2519
rect -1462 -2527 -1460 -2519
rect -1454 -2527 -1452 -2519
rect -1444 -2527 -1442 -2519
rect -1436 -2527 -1434 -2519
rect -1420 -2527 -1418 -2519
rect -1412 -2527 -1410 -2519
rect -1402 -2527 -1400 -2519
rect -1394 -2527 -1392 -2519
rect -1378 -2527 -1376 -2519
rect -1370 -2527 -1368 -2519
rect -1229 -2527 -1227 -2519
rect -1219 -2527 -1217 -2519
rect -1203 -2527 -1201 -2519
rect -1195 -2527 -1193 -2519
rect -1179 -2527 -1177 -2519
rect -1171 -2527 -1169 -2519
rect -1161 -2527 -1159 -2519
rect -1153 -2527 -1151 -2519
rect -1137 -2527 -1135 -2519
rect -1129 -2527 -1127 -2519
rect -1119 -2527 -1117 -2519
rect -1111 -2527 -1109 -2519
rect -1095 -2527 -1093 -2519
rect -1087 -2527 -1085 -2519
rect -1077 -2527 -1075 -2519
rect -1069 -2527 -1067 -2519
rect -1053 -2527 -1051 -2519
rect -1045 -2527 -1043 -2519
rect -930 -2527 -928 -2519
rect -920 -2527 -918 -2519
rect -904 -2527 -902 -2519
rect -896 -2527 -894 -2519
rect -880 -2527 -878 -2519
rect -872 -2527 -870 -2519
rect -862 -2527 -860 -2519
rect -854 -2527 -852 -2519
rect -838 -2527 -836 -2519
rect -830 -2527 -828 -2519
rect -820 -2527 -818 -2519
rect -812 -2527 -810 -2519
rect -796 -2527 -794 -2519
rect -788 -2527 -786 -2519
rect -778 -2527 -776 -2519
rect -770 -2527 -768 -2519
rect -754 -2527 -752 -2519
rect -746 -2527 -744 -2519
rect -572 -2527 -570 -2519
rect -562 -2527 -560 -2519
rect -546 -2527 -544 -2519
rect -538 -2527 -536 -2519
rect -522 -2527 -520 -2519
rect -514 -2527 -512 -2519
rect -504 -2527 -502 -2519
rect -496 -2527 -494 -2519
rect -480 -2527 -478 -2519
rect -472 -2527 -470 -2519
rect -462 -2527 -460 -2519
rect -454 -2527 -452 -2519
rect -438 -2527 -436 -2519
rect -430 -2527 -428 -2519
rect -420 -2527 -418 -2519
rect -412 -2527 -410 -2519
rect -396 -2527 -394 -2519
rect -388 -2527 -386 -2519
rect -215 -2527 -213 -2519
rect -205 -2527 -203 -2519
rect -189 -2527 -187 -2519
rect -181 -2527 -179 -2519
rect -165 -2527 -163 -2519
rect -157 -2527 -155 -2519
rect -147 -2527 -145 -2519
rect -139 -2527 -137 -2519
rect -123 -2527 -121 -2519
rect -115 -2527 -113 -2519
rect -105 -2527 -103 -2519
rect -97 -2527 -95 -2519
rect -81 -2527 -79 -2519
rect -73 -2527 -71 -2519
rect -63 -2527 -61 -2519
rect -55 -2527 -53 -2519
rect -39 -2527 -37 -2519
rect -31 -2527 -29 -2519
rect 144 -2527 146 -2519
rect 154 -2527 156 -2519
rect 170 -2527 172 -2519
rect 178 -2527 180 -2519
rect 194 -2527 196 -2519
rect 202 -2527 204 -2519
rect 212 -2527 214 -2519
rect 220 -2527 222 -2519
rect 236 -2527 238 -2519
rect 244 -2527 246 -2519
rect 254 -2527 256 -2519
rect 262 -2527 264 -2519
rect 278 -2527 280 -2519
rect 286 -2527 288 -2519
rect 296 -2527 298 -2519
rect 304 -2527 306 -2519
rect 320 -2527 322 -2519
rect 328 -2527 330 -2519
rect 500 -2527 502 -2519
rect 510 -2527 512 -2519
rect 526 -2527 528 -2519
rect 534 -2527 536 -2519
rect 550 -2527 552 -2519
rect 558 -2527 560 -2519
rect 568 -2527 570 -2519
rect 576 -2527 578 -2519
rect 592 -2527 594 -2519
rect 600 -2527 602 -2519
rect 610 -2527 612 -2519
rect 618 -2527 620 -2519
rect 634 -2527 636 -2519
rect 642 -2527 644 -2519
rect 652 -2527 654 -2519
rect 660 -2527 662 -2519
rect 676 -2527 678 -2519
rect 684 -2527 686 -2519
rect 858 -2527 860 -2519
rect 868 -2527 870 -2519
rect 884 -2527 886 -2519
rect 892 -2527 894 -2519
rect 908 -2527 910 -2519
rect 916 -2527 918 -2519
rect 926 -2527 928 -2519
rect 934 -2527 936 -2519
rect 950 -2527 952 -2519
rect 958 -2527 960 -2519
rect 968 -2527 970 -2519
rect 976 -2527 978 -2519
rect 992 -2527 994 -2519
rect 1000 -2527 1002 -2519
rect 1010 -2527 1012 -2519
rect 1018 -2527 1020 -2519
rect 1034 -2527 1036 -2519
rect 1042 -2527 1044 -2519
rect 1216 -2527 1218 -2519
rect 1226 -2527 1228 -2519
rect 1242 -2527 1244 -2519
rect 1250 -2527 1252 -2519
rect 1266 -2527 1268 -2519
rect 1274 -2527 1276 -2519
rect 1284 -2527 1286 -2519
rect 1292 -2527 1294 -2519
rect 1308 -2527 1310 -2519
rect 1316 -2527 1318 -2519
rect 1326 -2527 1328 -2519
rect 1334 -2527 1336 -2519
rect 1350 -2527 1352 -2519
rect 1358 -2527 1360 -2519
rect 1368 -2527 1370 -2519
rect 1376 -2527 1378 -2519
rect 1392 -2527 1394 -2519
rect 1400 -2527 1402 -2519
rect -1304 -2632 -1302 -2624
rect -1296 -2632 -1294 -2624
rect -1286 -2632 -1284 -2624
rect -930 -2632 -928 -2624
rect -922 -2632 -920 -2624
rect -912 -2632 -910 -2624
rect -572 -2632 -570 -2624
rect -564 -2632 -562 -2624
rect -554 -2632 -552 -2624
rect -214 -2632 -212 -2624
rect -206 -2632 -204 -2624
rect -196 -2632 -194 -2624
rect 144 -2632 146 -2624
rect 152 -2632 154 -2624
rect 162 -2632 164 -2624
rect 500 -2632 502 -2624
rect 508 -2632 510 -2624
rect 518 -2632 520 -2624
rect 858 -2632 860 -2624
rect 866 -2632 868 -2624
rect 876 -2632 878 -2624
rect 1216 -2632 1218 -2624
rect 1224 -2632 1226 -2624
rect 1234 -2632 1236 -2624
rect -1229 -2791 -1227 -2783
rect -1219 -2791 -1217 -2783
rect -1203 -2791 -1201 -2783
rect -1193 -2791 -1191 -2783
rect -1185 -2791 -1183 -2783
rect -1175 -2791 -1173 -2783
rect -1159 -2791 -1157 -2783
rect -1151 -2791 -1149 -2783
rect -1141 -2791 -1139 -2783
rect -930 -2791 -928 -2783
rect -920 -2791 -918 -2783
rect -904 -2791 -902 -2783
rect -894 -2791 -892 -2783
rect -878 -2791 -876 -2783
rect -868 -2791 -866 -2783
rect -860 -2791 -858 -2783
rect -850 -2791 -848 -2783
rect -834 -2791 -832 -2783
rect -826 -2791 -824 -2783
rect -816 -2791 -814 -2783
rect -800 -2791 -798 -2783
rect -790 -2791 -788 -2783
rect -782 -2791 -780 -2783
rect -772 -2791 -770 -2783
rect -756 -2791 -754 -2783
rect -748 -2791 -746 -2783
rect -732 -2791 -730 -2783
rect -716 -2791 -714 -2783
rect -708 -2791 -706 -2783
rect -698 -2791 -696 -2783
rect -572 -2791 -570 -2783
rect -562 -2791 -560 -2783
rect -546 -2791 -544 -2783
rect -536 -2791 -534 -2783
rect -520 -2791 -518 -2783
rect -510 -2791 -508 -2783
rect -502 -2791 -500 -2783
rect -492 -2791 -490 -2783
rect -476 -2791 -474 -2783
rect -468 -2791 -466 -2783
rect -458 -2791 -456 -2783
rect -442 -2791 -440 -2783
rect -432 -2791 -430 -2783
rect -424 -2791 -422 -2783
rect -414 -2791 -412 -2783
rect -398 -2791 -396 -2783
rect -390 -2791 -388 -2783
rect -374 -2791 -372 -2783
rect -358 -2791 -356 -2783
rect -350 -2791 -348 -2783
rect -340 -2791 -338 -2783
rect -214 -2791 -212 -2783
rect -204 -2791 -202 -2783
rect -188 -2791 -186 -2783
rect -178 -2791 -176 -2783
rect -162 -2791 -160 -2783
rect -152 -2791 -150 -2783
rect -144 -2791 -142 -2783
rect -134 -2791 -132 -2783
rect -118 -2791 -116 -2783
rect -110 -2791 -108 -2783
rect -100 -2791 -98 -2783
rect -84 -2791 -82 -2783
rect -74 -2791 -72 -2783
rect -66 -2791 -64 -2783
rect -56 -2791 -54 -2783
rect -40 -2791 -38 -2783
rect -32 -2791 -30 -2783
rect -16 -2791 -14 -2783
rect 0 -2791 2 -2783
rect 8 -2791 10 -2783
rect 18 -2791 20 -2783
rect 144 -2791 146 -2783
rect 154 -2791 156 -2783
rect 170 -2791 172 -2783
rect 180 -2791 182 -2783
rect 196 -2791 198 -2783
rect 206 -2791 208 -2783
rect 214 -2791 216 -2783
rect 224 -2791 226 -2783
rect 240 -2791 242 -2783
rect 248 -2791 250 -2783
rect 258 -2791 260 -2783
rect 274 -2791 276 -2783
rect 284 -2791 286 -2783
rect 292 -2791 294 -2783
rect 302 -2791 304 -2783
rect 318 -2791 320 -2783
rect 326 -2791 328 -2783
rect 342 -2791 344 -2783
rect 358 -2791 360 -2783
rect 366 -2791 368 -2783
rect 376 -2791 378 -2783
rect 500 -2791 502 -2783
rect 510 -2791 512 -2783
rect 526 -2791 528 -2783
rect 536 -2791 538 -2783
rect 552 -2791 554 -2783
rect 562 -2791 564 -2783
rect 570 -2791 572 -2783
rect 580 -2791 582 -2783
rect 596 -2791 598 -2783
rect 604 -2791 606 -2783
rect 614 -2791 616 -2783
rect 630 -2791 632 -2783
rect 640 -2791 642 -2783
rect 648 -2791 650 -2783
rect 658 -2791 660 -2783
rect 674 -2791 676 -2783
rect 682 -2791 684 -2783
rect 698 -2791 700 -2783
rect 714 -2791 716 -2783
rect 722 -2791 724 -2783
rect 732 -2791 734 -2783
rect 858 -2791 860 -2783
rect 868 -2791 870 -2783
rect 884 -2791 886 -2783
rect 894 -2791 896 -2783
rect 910 -2791 912 -2783
rect 920 -2791 922 -2783
rect 928 -2791 930 -2783
rect 938 -2791 940 -2783
rect 954 -2791 956 -2783
rect 962 -2791 964 -2783
rect 972 -2791 974 -2783
rect 988 -2791 990 -2783
rect 998 -2791 1000 -2783
rect 1006 -2791 1008 -2783
rect 1016 -2791 1018 -2783
rect 1032 -2791 1034 -2783
rect 1040 -2791 1042 -2783
rect 1056 -2791 1058 -2783
rect 1072 -2791 1074 -2783
rect 1080 -2791 1082 -2783
rect 1090 -2791 1092 -2783
rect 1216 -2791 1218 -2783
rect 1226 -2791 1228 -2783
rect 1242 -2791 1244 -2783
rect 1252 -2791 1254 -2783
rect 1268 -2791 1270 -2783
rect 1278 -2791 1280 -2783
rect 1286 -2791 1288 -2783
rect 1296 -2791 1298 -2783
rect 1312 -2791 1314 -2783
rect 1320 -2791 1322 -2783
rect 1330 -2791 1332 -2783
rect 1346 -2791 1348 -2783
rect 1356 -2791 1358 -2783
rect 1364 -2791 1366 -2783
rect 1374 -2791 1376 -2783
rect 1390 -2791 1392 -2783
rect 1398 -2791 1400 -2783
rect 1414 -2791 1416 -2783
rect 1430 -2791 1432 -2783
rect 1438 -2791 1440 -2783
rect 1448 -2791 1450 -2783
rect -1554 -2910 -1552 -2902
rect -1544 -2910 -1542 -2902
rect -1528 -2910 -1526 -2902
rect -1520 -2910 -1518 -2902
rect -1504 -2910 -1502 -2902
rect -1496 -2910 -1494 -2902
rect -1486 -2910 -1484 -2902
rect -1478 -2910 -1476 -2902
rect -1462 -2910 -1460 -2902
rect -1454 -2910 -1452 -2902
rect -1444 -2910 -1442 -2902
rect -1436 -2910 -1434 -2902
rect -1420 -2910 -1418 -2902
rect -1412 -2910 -1410 -2902
rect -1402 -2910 -1400 -2902
rect -1394 -2910 -1392 -2902
rect -1378 -2910 -1376 -2902
rect -1370 -2910 -1368 -2902
rect -1229 -2910 -1227 -2902
rect -1219 -2910 -1217 -2902
rect -1203 -2910 -1201 -2902
rect -1195 -2910 -1193 -2902
rect -1179 -2910 -1177 -2902
rect -1171 -2910 -1169 -2902
rect -1161 -2910 -1159 -2902
rect -1153 -2910 -1151 -2902
rect -1137 -2910 -1135 -2902
rect -1129 -2910 -1127 -2902
rect -1119 -2910 -1117 -2902
rect -1111 -2910 -1109 -2902
rect -1095 -2910 -1093 -2902
rect -1087 -2910 -1085 -2902
rect -1077 -2910 -1075 -2902
rect -1069 -2910 -1067 -2902
rect -1053 -2910 -1051 -2902
rect -1045 -2910 -1043 -2902
rect -930 -2910 -928 -2902
rect -920 -2910 -918 -2902
rect -904 -2910 -902 -2902
rect -896 -2910 -894 -2902
rect -880 -2910 -878 -2902
rect -872 -2910 -870 -2902
rect -862 -2910 -860 -2902
rect -854 -2910 -852 -2902
rect -838 -2910 -836 -2902
rect -830 -2910 -828 -2902
rect -820 -2910 -818 -2902
rect -812 -2910 -810 -2902
rect -796 -2910 -794 -2902
rect -788 -2910 -786 -2902
rect -778 -2910 -776 -2902
rect -770 -2910 -768 -2902
rect -754 -2910 -752 -2902
rect -746 -2910 -744 -2902
rect -572 -2910 -570 -2902
rect -562 -2910 -560 -2902
rect -546 -2910 -544 -2902
rect -538 -2910 -536 -2902
rect -522 -2910 -520 -2902
rect -514 -2910 -512 -2902
rect -504 -2910 -502 -2902
rect -496 -2910 -494 -2902
rect -480 -2910 -478 -2902
rect -472 -2910 -470 -2902
rect -462 -2910 -460 -2902
rect -454 -2910 -452 -2902
rect -438 -2910 -436 -2902
rect -430 -2910 -428 -2902
rect -420 -2910 -418 -2902
rect -412 -2910 -410 -2902
rect -396 -2910 -394 -2902
rect -388 -2910 -386 -2902
rect -214 -2910 -212 -2902
rect -204 -2910 -202 -2902
rect -188 -2910 -186 -2902
rect -180 -2910 -178 -2902
rect -164 -2910 -162 -2902
rect -156 -2910 -154 -2902
rect -146 -2910 -144 -2902
rect -138 -2910 -136 -2902
rect -122 -2910 -120 -2902
rect -114 -2910 -112 -2902
rect -104 -2910 -102 -2902
rect -96 -2910 -94 -2902
rect -80 -2910 -78 -2902
rect -72 -2910 -70 -2902
rect -62 -2910 -60 -2902
rect -54 -2910 -52 -2902
rect -38 -2910 -36 -2902
rect -30 -2910 -28 -2902
rect 144 -2910 146 -2902
rect 154 -2910 156 -2902
rect 170 -2910 172 -2902
rect 178 -2910 180 -2902
rect 194 -2910 196 -2902
rect 202 -2910 204 -2902
rect 212 -2910 214 -2902
rect 220 -2910 222 -2902
rect 236 -2910 238 -2902
rect 244 -2910 246 -2902
rect 254 -2910 256 -2902
rect 262 -2910 264 -2902
rect 278 -2910 280 -2902
rect 286 -2910 288 -2902
rect 296 -2910 298 -2902
rect 304 -2910 306 -2902
rect 320 -2910 322 -2902
rect 328 -2910 330 -2902
rect -1554 -3081 -1552 -3073
rect -1544 -3081 -1542 -3073
rect -1528 -3081 -1526 -3073
rect -1520 -3081 -1518 -3073
rect -1504 -3081 -1502 -3073
rect -1496 -3081 -1494 -3073
rect -1486 -3081 -1484 -3073
rect -1478 -3081 -1476 -3073
rect -1462 -3081 -1460 -3073
rect -1454 -3081 -1452 -3073
rect -1444 -3081 -1442 -3073
rect -1436 -3081 -1434 -3073
rect -1420 -3081 -1418 -3073
rect -1412 -3081 -1410 -3073
rect -1402 -3081 -1400 -3073
rect -1394 -3081 -1392 -3073
rect -1378 -3081 -1376 -3073
rect -1370 -3081 -1368 -3073
rect -1229 -3081 -1227 -3073
rect -1219 -3081 -1217 -3073
rect -1203 -3081 -1201 -3073
rect -1195 -3081 -1193 -3073
rect -1179 -3081 -1177 -3073
rect -1171 -3081 -1169 -3073
rect -1161 -3081 -1159 -3073
rect -1153 -3081 -1151 -3073
rect -1137 -3081 -1135 -3073
rect -1129 -3081 -1127 -3073
rect -1119 -3081 -1117 -3073
rect -1111 -3081 -1109 -3073
rect -1095 -3081 -1093 -3073
rect -1087 -3081 -1085 -3073
rect -1077 -3081 -1075 -3073
rect -1069 -3081 -1067 -3073
rect -1053 -3081 -1051 -3073
rect -1045 -3081 -1043 -3073
rect -930 -3081 -928 -3073
rect -920 -3081 -918 -3073
rect -904 -3081 -902 -3073
rect -896 -3081 -894 -3073
rect -880 -3081 -878 -3073
rect -872 -3081 -870 -3073
rect -862 -3081 -860 -3073
rect -854 -3081 -852 -3073
rect -838 -3081 -836 -3073
rect -830 -3081 -828 -3073
rect -820 -3081 -818 -3073
rect -812 -3081 -810 -3073
rect -796 -3081 -794 -3073
rect -788 -3081 -786 -3073
rect -778 -3081 -776 -3073
rect -770 -3081 -768 -3073
rect -754 -3081 -752 -3073
rect -746 -3081 -744 -3073
rect -572 -3081 -570 -3073
rect -562 -3081 -560 -3073
rect -546 -3081 -544 -3073
rect -538 -3081 -536 -3073
rect -522 -3081 -520 -3073
rect -514 -3081 -512 -3073
rect -504 -3081 -502 -3073
rect -496 -3081 -494 -3073
rect -480 -3081 -478 -3073
rect -472 -3081 -470 -3073
rect -462 -3081 -460 -3073
rect -454 -3081 -452 -3073
rect -438 -3081 -436 -3073
rect -430 -3081 -428 -3073
rect -420 -3081 -418 -3073
rect -412 -3081 -410 -3073
rect -396 -3081 -394 -3073
rect -388 -3081 -386 -3073
rect -214 -3081 -212 -3073
rect -204 -3081 -202 -3073
rect -188 -3081 -186 -3073
rect -180 -3081 -178 -3073
rect -164 -3081 -162 -3073
rect -156 -3081 -154 -3073
rect -146 -3081 -144 -3073
rect -138 -3081 -136 -3073
rect -122 -3081 -120 -3073
rect -114 -3081 -112 -3073
rect -104 -3081 -102 -3073
rect -96 -3081 -94 -3073
rect -80 -3081 -78 -3073
rect -72 -3081 -70 -3073
rect -62 -3081 -60 -3073
rect -54 -3081 -52 -3073
rect -38 -3081 -36 -3073
rect -30 -3081 -28 -3073
rect 144 -3081 146 -3073
rect 154 -3081 156 -3073
rect 170 -3081 172 -3073
rect 178 -3081 180 -3073
rect 194 -3081 196 -3073
rect 202 -3081 204 -3073
rect 212 -3081 214 -3073
rect 220 -3081 222 -3073
rect 236 -3081 238 -3073
rect 244 -3081 246 -3073
rect 254 -3081 256 -3073
rect 262 -3081 264 -3073
rect 278 -3081 280 -3073
rect 286 -3081 288 -3073
rect 296 -3081 298 -3073
rect 304 -3081 306 -3073
rect 320 -3081 322 -3073
rect 328 -3081 330 -3073
rect 500 -3081 502 -3073
rect 510 -3081 512 -3073
rect 526 -3081 528 -3073
rect 534 -3081 536 -3073
rect 550 -3081 552 -3073
rect 558 -3081 560 -3073
rect 568 -3081 570 -3073
rect 576 -3081 578 -3073
rect 592 -3081 594 -3073
rect 600 -3081 602 -3073
rect 610 -3081 612 -3073
rect 618 -3081 620 -3073
rect 634 -3081 636 -3073
rect 642 -3081 644 -3073
rect 652 -3081 654 -3073
rect 660 -3081 662 -3073
rect 676 -3081 678 -3073
rect 684 -3081 686 -3073
rect 858 -3081 860 -3073
rect 868 -3081 870 -3073
rect 884 -3081 886 -3073
rect 892 -3081 894 -3073
rect 908 -3081 910 -3073
rect 916 -3081 918 -3073
rect 926 -3081 928 -3073
rect 934 -3081 936 -3073
rect 950 -3081 952 -3073
rect 958 -3081 960 -3073
rect 968 -3081 970 -3073
rect 976 -3081 978 -3073
rect 992 -3081 994 -3073
rect 1000 -3081 1002 -3073
rect 1010 -3081 1012 -3073
rect 1018 -3081 1020 -3073
rect 1034 -3081 1036 -3073
rect 1042 -3081 1044 -3073
rect 1216 -3081 1218 -3073
rect 1226 -3081 1228 -3073
rect 1242 -3081 1244 -3073
rect 1250 -3081 1252 -3073
rect 1266 -3081 1268 -3073
rect 1274 -3081 1276 -3073
rect 1284 -3081 1286 -3073
rect 1292 -3081 1294 -3073
rect 1308 -3081 1310 -3073
rect 1316 -3081 1318 -3073
rect 1326 -3081 1328 -3073
rect 1334 -3081 1336 -3073
rect 1350 -3081 1352 -3073
rect 1358 -3081 1360 -3073
rect 1368 -3081 1370 -3073
rect 1376 -3081 1378 -3073
rect 1392 -3081 1394 -3073
rect 1400 -3081 1402 -3073
rect -1554 -3252 -1552 -3244
rect -1544 -3252 -1542 -3244
rect -1528 -3252 -1526 -3244
rect -1520 -3252 -1518 -3244
rect -1504 -3252 -1502 -3244
rect -1496 -3252 -1494 -3244
rect -1486 -3252 -1484 -3244
rect -1478 -3252 -1476 -3244
rect -1462 -3252 -1460 -3244
rect -1454 -3252 -1452 -3244
rect -1444 -3252 -1442 -3244
rect -1436 -3252 -1434 -3244
rect -1420 -3252 -1418 -3244
rect -1412 -3252 -1410 -3244
rect -1402 -3252 -1400 -3244
rect -1394 -3252 -1392 -3244
rect -1378 -3252 -1376 -3244
rect -1370 -3252 -1368 -3244
rect -1229 -3252 -1227 -3244
rect -1219 -3252 -1217 -3244
rect -1203 -3252 -1201 -3244
rect -1195 -3252 -1193 -3244
rect -1179 -3252 -1177 -3244
rect -1171 -3252 -1169 -3244
rect -1161 -3252 -1159 -3244
rect -1153 -3252 -1151 -3244
rect -1137 -3252 -1135 -3244
rect -1129 -3252 -1127 -3244
rect -1119 -3252 -1117 -3244
rect -1111 -3252 -1109 -3244
rect -1095 -3252 -1093 -3244
rect -1087 -3252 -1085 -3244
rect -1077 -3252 -1075 -3244
rect -1069 -3252 -1067 -3244
rect -1053 -3252 -1051 -3244
rect -1045 -3252 -1043 -3244
rect -930 -3252 -928 -3244
rect -920 -3252 -918 -3244
rect -904 -3252 -902 -3244
rect -896 -3252 -894 -3244
rect -880 -3252 -878 -3244
rect -872 -3252 -870 -3244
rect -862 -3252 -860 -3244
rect -854 -3252 -852 -3244
rect -838 -3252 -836 -3244
rect -830 -3252 -828 -3244
rect -820 -3252 -818 -3244
rect -812 -3252 -810 -3244
rect -796 -3252 -794 -3244
rect -788 -3252 -786 -3244
rect -778 -3252 -776 -3244
rect -770 -3252 -768 -3244
rect -754 -3252 -752 -3244
rect -746 -3252 -744 -3244
rect -572 -3252 -570 -3244
rect -562 -3252 -560 -3244
rect -546 -3252 -544 -3244
rect -538 -3252 -536 -3244
rect -522 -3252 -520 -3244
rect -514 -3252 -512 -3244
rect -504 -3252 -502 -3244
rect -496 -3252 -494 -3244
rect -480 -3252 -478 -3244
rect -472 -3252 -470 -3244
rect -462 -3252 -460 -3244
rect -454 -3252 -452 -3244
rect -438 -3252 -436 -3244
rect -430 -3252 -428 -3244
rect -420 -3252 -418 -3244
rect -412 -3252 -410 -3244
rect -396 -3252 -394 -3244
rect -388 -3252 -386 -3244
rect -214 -3252 -212 -3244
rect -204 -3252 -202 -3244
rect -188 -3252 -186 -3244
rect -180 -3252 -178 -3244
rect -164 -3252 -162 -3244
rect -156 -3252 -154 -3244
rect -146 -3252 -144 -3244
rect -138 -3252 -136 -3244
rect -122 -3252 -120 -3244
rect -114 -3252 -112 -3244
rect -104 -3252 -102 -3244
rect -96 -3252 -94 -3244
rect -80 -3252 -78 -3244
rect -72 -3252 -70 -3244
rect -62 -3252 -60 -3244
rect -54 -3252 -52 -3244
rect -38 -3252 -36 -3244
rect -30 -3252 -28 -3244
rect 144 -3252 146 -3244
rect 154 -3252 156 -3244
rect 170 -3252 172 -3244
rect 178 -3252 180 -3244
rect 194 -3252 196 -3244
rect 202 -3252 204 -3244
rect 212 -3252 214 -3244
rect 220 -3252 222 -3244
rect 236 -3252 238 -3244
rect 244 -3252 246 -3244
rect 254 -3252 256 -3244
rect 262 -3252 264 -3244
rect 278 -3252 280 -3244
rect 286 -3252 288 -3244
rect 296 -3252 298 -3244
rect 304 -3252 306 -3244
rect 320 -3252 322 -3244
rect 328 -3252 330 -3244
rect 500 -3252 502 -3244
rect 510 -3252 512 -3244
rect 526 -3252 528 -3244
rect 534 -3252 536 -3244
rect 550 -3252 552 -3244
rect 558 -3252 560 -3244
rect 568 -3252 570 -3244
rect 576 -3252 578 -3244
rect 592 -3252 594 -3244
rect 600 -3252 602 -3244
rect 610 -3252 612 -3244
rect 618 -3252 620 -3244
rect 634 -3252 636 -3244
rect 642 -3252 644 -3244
rect 652 -3252 654 -3244
rect 660 -3252 662 -3244
rect 676 -3252 678 -3244
rect 684 -3252 686 -3244
rect 858 -3252 860 -3244
rect 868 -3252 870 -3244
rect 884 -3252 886 -3244
rect 892 -3252 894 -3244
rect 908 -3252 910 -3244
rect 916 -3252 918 -3244
rect 926 -3252 928 -3244
rect 934 -3252 936 -3244
rect 950 -3252 952 -3244
rect 958 -3252 960 -3244
rect 968 -3252 970 -3244
rect 976 -3252 978 -3244
rect 992 -3252 994 -3244
rect 1000 -3252 1002 -3244
rect 1010 -3252 1012 -3244
rect 1018 -3252 1020 -3244
rect 1034 -3252 1036 -3244
rect 1042 -3252 1044 -3244
rect 1216 -3252 1218 -3244
rect 1226 -3252 1228 -3244
rect 1242 -3252 1244 -3244
rect 1250 -3252 1252 -3244
rect 1266 -3252 1268 -3244
rect 1274 -3252 1276 -3244
rect 1284 -3252 1286 -3244
rect 1292 -3252 1294 -3244
rect 1308 -3252 1310 -3244
rect 1316 -3252 1318 -3244
rect 1326 -3252 1328 -3244
rect 1334 -3252 1336 -3244
rect 1350 -3252 1352 -3244
rect 1358 -3252 1360 -3244
rect 1368 -3252 1370 -3244
rect 1376 -3252 1378 -3244
rect 1392 -3252 1394 -3244
rect 1400 -3252 1402 -3244
rect -1304 -3363 -1302 -3355
rect -1296 -3363 -1294 -3355
rect -1286 -3363 -1284 -3355
rect -930 -3363 -928 -3355
rect -922 -3363 -920 -3355
rect -912 -3363 -910 -3355
rect -572 -3363 -570 -3355
rect -564 -3363 -562 -3355
rect -554 -3363 -552 -3355
rect -214 -3363 -212 -3355
rect -206 -3363 -204 -3355
rect -196 -3363 -194 -3355
rect 144 -3363 146 -3355
rect 152 -3363 154 -3355
rect 162 -3363 164 -3355
rect 500 -3363 502 -3355
rect 508 -3363 510 -3355
rect 518 -3363 520 -3355
rect 858 -3363 860 -3355
rect 866 -3363 868 -3355
rect 876 -3363 878 -3355
rect 1216 -3363 1218 -3355
rect 1224 -3363 1226 -3355
rect 1234 -3363 1236 -3355
rect -1229 -3522 -1227 -3514
rect -1219 -3522 -1217 -3514
rect -1203 -3522 -1201 -3514
rect -1193 -3522 -1191 -3514
rect -1185 -3522 -1183 -3514
rect -1175 -3522 -1173 -3514
rect -1159 -3522 -1157 -3514
rect -1151 -3522 -1149 -3514
rect -1141 -3522 -1139 -3514
rect -930 -3522 -928 -3514
rect -920 -3522 -918 -3514
rect -904 -3522 -902 -3514
rect -894 -3522 -892 -3514
rect -878 -3522 -876 -3514
rect -868 -3522 -866 -3514
rect -860 -3522 -858 -3514
rect -850 -3522 -848 -3514
rect -834 -3522 -832 -3514
rect -826 -3522 -824 -3514
rect -816 -3522 -814 -3514
rect -800 -3522 -798 -3514
rect -790 -3522 -788 -3514
rect -782 -3522 -780 -3514
rect -772 -3522 -770 -3514
rect -756 -3522 -754 -3514
rect -748 -3522 -746 -3514
rect -732 -3522 -730 -3514
rect -716 -3522 -714 -3514
rect -708 -3522 -706 -3514
rect -698 -3522 -696 -3514
rect -572 -3522 -570 -3514
rect -562 -3522 -560 -3514
rect -546 -3522 -544 -3514
rect -536 -3522 -534 -3514
rect -520 -3522 -518 -3514
rect -510 -3522 -508 -3514
rect -502 -3522 -500 -3514
rect -492 -3522 -490 -3514
rect -476 -3522 -474 -3514
rect -468 -3522 -466 -3514
rect -458 -3522 -456 -3514
rect -442 -3522 -440 -3514
rect -432 -3522 -430 -3514
rect -424 -3522 -422 -3514
rect -414 -3522 -412 -3514
rect -398 -3522 -396 -3514
rect -390 -3522 -388 -3514
rect -374 -3522 -372 -3514
rect -358 -3522 -356 -3514
rect -350 -3522 -348 -3514
rect -340 -3522 -338 -3514
rect -214 -3522 -212 -3514
rect -204 -3522 -202 -3514
rect -188 -3522 -186 -3514
rect -178 -3522 -176 -3514
rect -162 -3522 -160 -3514
rect -152 -3522 -150 -3514
rect -144 -3522 -142 -3514
rect -134 -3522 -132 -3514
rect -118 -3522 -116 -3514
rect -110 -3522 -108 -3514
rect -100 -3522 -98 -3514
rect -84 -3522 -82 -3514
rect -74 -3522 -72 -3514
rect -66 -3522 -64 -3514
rect -56 -3522 -54 -3514
rect -40 -3522 -38 -3514
rect -32 -3522 -30 -3514
rect -16 -3522 -14 -3514
rect 0 -3522 2 -3514
rect 8 -3522 10 -3514
rect 18 -3522 20 -3514
rect 144 -3522 146 -3514
rect 154 -3522 156 -3514
rect 170 -3522 172 -3514
rect 180 -3522 182 -3514
rect 196 -3522 198 -3514
rect 206 -3522 208 -3514
rect 214 -3522 216 -3514
rect 224 -3522 226 -3514
rect 240 -3522 242 -3514
rect 248 -3522 250 -3514
rect 258 -3522 260 -3514
rect 274 -3522 276 -3514
rect 284 -3522 286 -3514
rect 292 -3522 294 -3514
rect 302 -3522 304 -3514
rect 318 -3522 320 -3514
rect 326 -3522 328 -3514
rect 342 -3522 344 -3514
rect 358 -3522 360 -3514
rect 366 -3522 368 -3514
rect 376 -3522 378 -3514
rect 500 -3522 502 -3514
rect 510 -3522 512 -3514
rect 526 -3522 528 -3514
rect 536 -3522 538 -3514
rect 552 -3522 554 -3514
rect 562 -3522 564 -3514
rect 570 -3522 572 -3514
rect 580 -3522 582 -3514
rect 596 -3522 598 -3514
rect 604 -3522 606 -3514
rect 614 -3522 616 -3514
rect 630 -3522 632 -3514
rect 640 -3522 642 -3514
rect 648 -3522 650 -3514
rect 658 -3522 660 -3514
rect 674 -3522 676 -3514
rect 682 -3522 684 -3514
rect 698 -3522 700 -3514
rect 714 -3522 716 -3514
rect 722 -3522 724 -3514
rect 732 -3522 734 -3514
rect 858 -3522 860 -3514
rect 868 -3522 870 -3514
rect 884 -3522 886 -3514
rect 894 -3522 896 -3514
rect 910 -3522 912 -3514
rect 920 -3522 922 -3514
rect 928 -3522 930 -3514
rect 938 -3522 940 -3514
rect 954 -3522 956 -3514
rect 962 -3522 964 -3514
rect 972 -3522 974 -3514
rect 988 -3522 990 -3514
rect 998 -3522 1000 -3514
rect 1006 -3522 1008 -3514
rect 1016 -3522 1018 -3514
rect 1032 -3522 1034 -3514
rect 1040 -3522 1042 -3514
rect 1056 -3522 1058 -3514
rect 1072 -3522 1074 -3514
rect 1080 -3522 1082 -3514
rect 1090 -3522 1092 -3514
rect 1216 -3522 1218 -3514
rect 1226 -3522 1228 -3514
rect 1242 -3522 1244 -3514
rect 1252 -3522 1254 -3514
rect 1268 -3522 1270 -3514
rect 1278 -3522 1280 -3514
rect 1286 -3522 1288 -3514
rect 1296 -3522 1298 -3514
rect 1312 -3522 1314 -3514
rect 1320 -3522 1322 -3514
rect 1330 -3522 1332 -3514
rect 1346 -3522 1348 -3514
rect 1356 -3522 1358 -3514
rect 1364 -3522 1366 -3514
rect 1374 -3522 1376 -3514
rect 1390 -3522 1392 -3514
rect 1398 -3522 1400 -3514
rect 1414 -3522 1416 -3514
rect 1430 -3522 1432 -3514
rect 1438 -3522 1440 -3514
rect 1448 -3522 1450 -3514
rect -1817 -3652 -1815 -3644
rect -1807 -3652 -1805 -3644
rect -1791 -3652 -1789 -3644
rect -1783 -3652 -1781 -3644
rect -1767 -3652 -1765 -3644
rect -1759 -3652 -1757 -3644
rect -1749 -3652 -1747 -3644
rect -1741 -3652 -1739 -3644
rect -1725 -3652 -1723 -3644
rect -1717 -3652 -1715 -3644
rect -1707 -3652 -1705 -3644
rect -1699 -3652 -1697 -3644
rect -1683 -3652 -1681 -3644
rect -1675 -3652 -1673 -3644
rect -1665 -3652 -1663 -3644
rect -1657 -3652 -1655 -3644
rect -1641 -3652 -1639 -3644
rect -1633 -3652 -1631 -3644
rect -1554 -3652 -1552 -3644
rect -1544 -3652 -1542 -3644
rect -1528 -3652 -1526 -3644
rect -1520 -3652 -1518 -3644
rect -1504 -3652 -1502 -3644
rect -1496 -3652 -1494 -3644
rect -1486 -3652 -1484 -3644
rect -1478 -3652 -1476 -3644
rect -1462 -3652 -1460 -3644
rect -1454 -3652 -1452 -3644
rect -1444 -3652 -1442 -3644
rect -1436 -3652 -1434 -3644
rect -1420 -3652 -1418 -3644
rect -1412 -3652 -1410 -3644
rect -1402 -3652 -1400 -3644
rect -1394 -3652 -1392 -3644
rect -1378 -3652 -1376 -3644
rect -1370 -3652 -1368 -3644
rect -1229 -3652 -1227 -3644
rect -1219 -3652 -1217 -3644
rect -1203 -3652 -1201 -3644
rect -1195 -3652 -1193 -3644
rect -1179 -3652 -1177 -3644
rect -1171 -3652 -1169 -3644
rect -1161 -3652 -1159 -3644
rect -1153 -3652 -1151 -3644
rect -1137 -3652 -1135 -3644
rect -1129 -3652 -1127 -3644
rect -1119 -3652 -1117 -3644
rect -1111 -3652 -1109 -3644
rect -1095 -3652 -1093 -3644
rect -1087 -3652 -1085 -3644
rect -1077 -3652 -1075 -3644
rect -1069 -3652 -1067 -3644
rect -1053 -3652 -1051 -3644
rect -1045 -3652 -1043 -3644
rect -929 -3652 -927 -3644
rect -919 -3652 -917 -3644
rect -903 -3652 -901 -3644
rect -895 -3652 -893 -3644
rect -879 -3652 -877 -3644
rect -871 -3652 -869 -3644
rect -861 -3652 -859 -3644
rect -853 -3652 -851 -3644
rect -837 -3652 -835 -3644
rect -829 -3652 -827 -3644
rect -819 -3652 -817 -3644
rect -811 -3652 -809 -3644
rect -795 -3652 -793 -3644
rect -787 -3652 -785 -3644
rect -777 -3652 -775 -3644
rect -769 -3652 -767 -3644
rect -753 -3652 -751 -3644
rect -745 -3652 -743 -3644
rect -572 -3652 -570 -3644
rect -562 -3652 -560 -3644
rect -546 -3652 -544 -3644
rect -538 -3652 -536 -3644
rect -522 -3652 -520 -3644
rect -514 -3652 -512 -3644
rect -504 -3652 -502 -3644
rect -496 -3652 -494 -3644
rect -480 -3652 -478 -3644
rect -472 -3652 -470 -3644
rect -462 -3652 -460 -3644
rect -454 -3652 -452 -3644
rect -438 -3652 -436 -3644
rect -430 -3652 -428 -3644
rect -420 -3652 -418 -3644
rect -412 -3652 -410 -3644
rect -396 -3652 -394 -3644
rect -388 -3652 -386 -3644
rect -214 -3652 -212 -3644
rect -204 -3652 -202 -3644
rect -188 -3652 -186 -3644
rect -180 -3652 -178 -3644
rect -164 -3652 -162 -3644
rect -156 -3652 -154 -3644
rect -146 -3652 -144 -3644
rect -138 -3652 -136 -3644
rect -122 -3652 -120 -3644
rect -114 -3652 -112 -3644
rect -104 -3652 -102 -3644
rect -96 -3652 -94 -3644
rect -80 -3652 -78 -3644
rect -72 -3652 -70 -3644
rect -62 -3652 -60 -3644
rect -54 -3652 -52 -3644
rect -38 -3652 -36 -3644
rect -30 -3652 -28 -3644
rect -1554 -3823 -1552 -3815
rect -1544 -3823 -1542 -3815
rect -1528 -3823 -1526 -3815
rect -1520 -3823 -1518 -3815
rect -1504 -3823 -1502 -3815
rect -1496 -3823 -1494 -3815
rect -1486 -3823 -1484 -3815
rect -1478 -3823 -1476 -3815
rect -1462 -3823 -1460 -3815
rect -1454 -3823 -1452 -3815
rect -1444 -3823 -1442 -3815
rect -1436 -3823 -1434 -3815
rect -1420 -3823 -1418 -3815
rect -1412 -3823 -1410 -3815
rect -1402 -3823 -1400 -3815
rect -1394 -3823 -1392 -3815
rect -1378 -3823 -1376 -3815
rect -1370 -3823 -1368 -3815
rect -1229 -3823 -1227 -3815
rect -1219 -3823 -1217 -3815
rect -1203 -3823 -1201 -3815
rect -1195 -3823 -1193 -3815
rect -1179 -3823 -1177 -3815
rect -1171 -3823 -1169 -3815
rect -1161 -3823 -1159 -3815
rect -1153 -3823 -1151 -3815
rect -1137 -3823 -1135 -3815
rect -1129 -3823 -1127 -3815
rect -1119 -3823 -1117 -3815
rect -1111 -3823 -1109 -3815
rect -1095 -3823 -1093 -3815
rect -1087 -3823 -1085 -3815
rect -1077 -3823 -1075 -3815
rect -1069 -3823 -1067 -3815
rect -1053 -3823 -1051 -3815
rect -1045 -3823 -1043 -3815
rect -929 -3823 -927 -3815
rect -919 -3823 -917 -3815
rect -903 -3823 -901 -3815
rect -895 -3823 -893 -3815
rect -879 -3823 -877 -3815
rect -871 -3823 -869 -3815
rect -861 -3823 -859 -3815
rect -853 -3823 -851 -3815
rect -837 -3823 -835 -3815
rect -829 -3823 -827 -3815
rect -819 -3823 -817 -3815
rect -811 -3823 -809 -3815
rect -795 -3823 -793 -3815
rect -787 -3823 -785 -3815
rect -777 -3823 -775 -3815
rect -769 -3823 -767 -3815
rect -753 -3823 -751 -3815
rect -745 -3823 -743 -3815
rect -572 -3823 -570 -3815
rect -562 -3823 -560 -3815
rect -546 -3823 -544 -3815
rect -538 -3823 -536 -3815
rect -522 -3823 -520 -3815
rect -514 -3823 -512 -3815
rect -504 -3823 -502 -3815
rect -496 -3823 -494 -3815
rect -480 -3823 -478 -3815
rect -472 -3823 -470 -3815
rect -462 -3823 -460 -3815
rect -454 -3823 -452 -3815
rect -438 -3823 -436 -3815
rect -430 -3823 -428 -3815
rect -420 -3823 -418 -3815
rect -412 -3823 -410 -3815
rect -396 -3823 -394 -3815
rect -388 -3823 -386 -3815
rect -214 -3823 -212 -3815
rect -204 -3823 -202 -3815
rect -188 -3823 -186 -3815
rect -180 -3823 -178 -3815
rect -164 -3823 -162 -3815
rect -156 -3823 -154 -3815
rect -146 -3823 -144 -3815
rect -138 -3823 -136 -3815
rect -122 -3823 -120 -3815
rect -114 -3823 -112 -3815
rect -104 -3823 -102 -3815
rect -96 -3823 -94 -3815
rect -80 -3823 -78 -3815
rect -72 -3823 -70 -3815
rect -62 -3823 -60 -3815
rect -54 -3823 -52 -3815
rect -38 -3823 -36 -3815
rect -30 -3823 -28 -3815
rect 144 -3823 146 -3815
rect 154 -3823 156 -3815
rect 170 -3823 172 -3815
rect 178 -3823 180 -3815
rect 194 -3823 196 -3815
rect 202 -3823 204 -3815
rect 212 -3823 214 -3815
rect 220 -3823 222 -3815
rect 236 -3823 238 -3815
rect 244 -3823 246 -3815
rect 254 -3823 256 -3815
rect 262 -3823 264 -3815
rect 278 -3823 280 -3815
rect 286 -3823 288 -3815
rect 296 -3823 298 -3815
rect 304 -3823 306 -3815
rect 320 -3823 322 -3815
rect 328 -3823 330 -3815
rect 500 -3823 502 -3815
rect 510 -3823 512 -3815
rect 526 -3823 528 -3815
rect 534 -3823 536 -3815
rect 550 -3823 552 -3815
rect 558 -3823 560 -3815
rect 568 -3823 570 -3815
rect 576 -3823 578 -3815
rect 592 -3823 594 -3815
rect 600 -3823 602 -3815
rect 610 -3823 612 -3815
rect 618 -3823 620 -3815
rect 634 -3823 636 -3815
rect 642 -3823 644 -3815
rect 652 -3823 654 -3815
rect 660 -3823 662 -3815
rect 676 -3823 678 -3815
rect 684 -3823 686 -3815
rect 858 -3823 860 -3815
rect 868 -3823 870 -3815
rect 884 -3823 886 -3815
rect 892 -3823 894 -3815
rect 908 -3823 910 -3815
rect 916 -3823 918 -3815
rect 926 -3823 928 -3815
rect 934 -3823 936 -3815
rect 950 -3823 952 -3815
rect 958 -3823 960 -3815
rect 968 -3823 970 -3815
rect 976 -3823 978 -3815
rect 992 -3823 994 -3815
rect 1000 -3823 1002 -3815
rect 1010 -3823 1012 -3815
rect 1018 -3823 1020 -3815
rect 1034 -3823 1036 -3815
rect 1042 -3823 1044 -3815
rect 1216 -3823 1218 -3815
rect 1226 -3823 1228 -3815
rect 1242 -3823 1244 -3815
rect 1250 -3823 1252 -3815
rect 1266 -3823 1268 -3815
rect 1274 -3823 1276 -3815
rect 1284 -3823 1286 -3815
rect 1292 -3823 1294 -3815
rect 1308 -3823 1310 -3815
rect 1316 -3823 1318 -3815
rect 1326 -3823 1328 -3815
rect 1334 -3823 1336 -3815
rect 1350 -3823 1352 -3815
rect 1358 -3823 1360 -3815
rect 1368 -3823 1370 -3815
rect 1376 -3823 1378 -3815
rect 1392 -3823 1394 -3815
rect 1400 -3823 1402 -3815
rect -1554 -3998 -1552 -3990
rect -1544 -3998 -1542 -3990
rect -1528 -3998 -1526 -3990
rect -1520 -3998 -1518 -3990
rect -1504 -3998 -1502 -3990
rect -1496 -3998 -1494 -3990
rect -1486 -3998 -1484 -3990
rect -1478 -3998 -1476 -3990
rect -1462 -3998 -1460 -3990
rect -1454 -3998 -1452 -3990
rect -1444 -3998 -1442 -3990
rect -1436 -3998 -1434 -3990
rect -1420 -3998 -1418 -3990
rect -1412 -3998 -1410 -3990
rect -1402 -3998 -1400 -3990
rect -1394 -3998 -1392 -3990
rect -1378 -3998 -1376 -3990
rect -1370 -3998 -1368 -3990
rect -1229 -3998 -1227 -3990
rect -1219 -3998 -1217 -3990
rect -1203 -3998 -1201 -3990
rect -1195 -3998 -1193 -3990
rect -1179 -3998 -1177 -3990
rect -1171 -3998 -1169 -3990
rect -1161 -3998 -1159 -3990
rect -1153 -3998 -1151 -3990
rect -1137 -3998 -1135 -3990
rect -1129 -3998 -1127 -3990
rect -1119 -3998 -1117 -3990
rect -1111 -3998 -1109 -3990
rect -1095 -3998 -1093 -3990
rect -1087 -3998 -1085 -3990
rect -1077 -3998 -1075 -3990
rect -1069 -3998 -1067 -3990
rect -1053 -3998 -1051 -3990
rect -1045 -3998 -1043 -3990
rect -930 -3998 -928 -3990
rect -920 -3998 -918 -3990
rect -904 -3998 -902 -3990
rect -896 -3998 -894 -3990
rect -880 -3998 -878 -3990
rect -872 -3998 -870 -3990
rect -862 -3998 -860 -3990
rect -854 -3998 -852 -3990
rect -838 -3998 -836 -3990
rect -830 -3998 -828 -3990
rect -820 -3998 -818 -3990
rect -812 -3998 -810 -3990
rect -796 -3998 -794 -3990
rect -788 -3998 -786 -3990
rect -778 -3998 -776 -3990
rect -770 -3998 -768 -3990
rect -754 -3998 -752 -3990
rect -746 -3998 -744 -3990
rect -572 -3998 -570 -3990
rect -562 -3998 -560 -3990
rect -546 -3998 -544 -3990
rect -538 -3998 -536 -3990
rect -522 -3998 -520 -3990
rect -514 -3998 -512 -3990
rect -504 -3998 -502 -3990
rect -496 -3998 -494 -3990
rect -480 -3998 -478 -3990
rect -472 -3998 -470 -3990
rect -462 -3998 -460 -3990
rect -454 -3998 -452 -3990
rect -438 -3998 -436 -3990
rect -430 -3998 -428 -3990
rect -420 -3998 -418 -3990
rect -412 -3998 -410 -3990
rect -396 -3998 -394 -3990
rect -388 -3998 -386 -3990
rect -214 -3998 -212 -3990
rect -204 -3998 -202 -3990
rect -188 -3998 -186 -3990
rect -180 -3998 -178 -3990
rect -164 -3998 -162 -3990
rect -156 -3998 -154 -3990
rect -146 -3998 -144 -3990
rect -138 -3998 -136 -3990
rect -122 -3998 -120 -3990
rect -114 -3998 -112 -3990
rect -104 -3998 -102 -3990
rect -96 -3998 -94 -3990
rect -80 -3998 -78 -3990
rect -72 -3998 -70 -3990
rect -62 -3998 -60 -3990
rect -54 -3998 -52 -3990
rect -38 -3998 -36 -3990
rect -30 -3998 -28 -3990
rect 144 -3998 146 -3990
rect 154 -3998 156 -3990
rect 170 -3998 172 -3990
rect 178 -3998 180 -3990
rect 194 -3998 196 -3990
rect 202 -3998 204 -3990
rect 212 -3998 214 -3990
rect 220 -3998 222 -3990
rect 236 -3998 238 -3990
rect 244 -3998 246 -3990
rect 254 -3998 256 -3990
rect 262 -3998 264 -3990
rect 278 -3998 280 -3990
rect 286 -3998 288 -3990
rect 296 -3998 298 -3990
rect 304 -3998 306 -3990
rect 320 -3998 322 -3990
rect 328 -3998 330 -3990
rect 500 -3998 502 -3990
rect 510 -3998 512 -3990
rect 526 -3998 528 -3990
rect 534 -3998 536 -3990
rect 550 -3998 552 -3990
rect 558 -3998 560 -3990
rect 568 -3998 570 -3990
rect 576 -3998 578 -3990
rect 592 -3998 594 -3990
rect 600 -3998 602 -3990
rect 610 -3998 612 -3990
rect 618 -3998 620 -3990
rect 634 -3998 636 -3990
rect 642 -3998 644 -3990
rect 652 -3998 654 -3990
rect 660 -3998 662 -3990
rect 676 -3998 678 -3990
rect 684 -3998 686 -3990
rect 858 -3998 860 -3990
rect 868 -3998 870 -3990
rect 884 -3998 886 -3990
rect 892 -3998 894 -3990
rect 908 -3998 910 -3990
rect 916 -3998 918 -3990
rect 926 -3998 928 -3990
rect 934 -3998 936 -3990
rect 950 -3998 952 -3990
rect 958 -3998 960 -3990
rect 968 -3998 970 -3990
rect 976 -3998 978 -3990
rect 992 -3998 994 -3990
rect 1000 -3998 1002 -3990
rect 1010 -3998 1012 -3990
rect 1018 -3998 1020 -3990
rect 1034 -3998 1036 -3990
rect 1042 -3998 1044 -3990
rect 1216 -3998 1218 -3990
rect 1226 -3998 1228 -3990
rect 1242 -3998 1244 -3990
rect 1250 -3998 1252 -3990
rect 1266 -3998 1268 -3990
rect 1274 -3998 1276 -3990
rect 1284 -3998 1286 -3990
rect 1292 -3998 1294 -3990
rect 1308 -3998 1310 -3990
rect 1316 -3998 1318 -3990
rect 1326 -3998 1328 -3990
rect 1334 -3998 1336 -3990
rect 1350 -3998 1352 -3990
rect 1358 -3998 1360 -3990
rect 1368 -3998 1370 -3990
rect 1376 -3998 1378 -3990
rect 1392 -3998 1394 -3990
rect 1400 -3998 1402 -3990
rect -1304 -4113 -1302 -4105
rect -1296 -4113 -1294 -4105
rect -1286 -4113 -1284 -4105
rect -930 -4113 -928 -4105
rect -922 -4113 -920 -4105
rect -912 -4113 -910 -4105
rect -572 -4113 -570 -4105
rect -564 -4113 -562 -4105
rect -554 -4113 -552 -4105
rect -214 -4113 -212 -4105
rect -206 -4113 -204 -4105
rect -196 -4113 -194 -4105
rect 144 -4113 146 -4105
rect 152 -4113 154 -4105
rect 162 -4113 164 -4105
rect 500 -4113 502 -4105
rect 508 -4113 510 -4105
rect 518 -4113 520 -4105
rect 858 -4113 860 -4105
rect 866 -4113 868 -4105
rect 876 -4113 878 -4105
rect 1216 -4113 1218 -4105
rect 1224 -4113 1226 -4105
rect 1234 -4113 1236 -4105
rect -1229 -4272 -1227 -4264
rect -1219 -4272 -1217 -4264
rect -1203 -4272 -1201 -4264
rect -1193 -4272 -1191 -4264
rect -1185 -4272 -1183 -4264
rect -1175 -4272 -1173 -4264
rect -1159 -4272 -1157 -4264
rect -1151 -4272 -1149 -4264
rect -1141 -4272 -1139 -4264
rect -930 -4272 -928 -4264
rect -920 -4272 -918 -4264
rect -904 -4272 -902 -4264
rect -894 -4272 -892 -4264
rect -878 -4272 -876 -4264
rect -868 -4272 -866 -4264
rect -860 -4272 -858 -4264
rect -850 -4272 -848 -4264
rect -834 -4272 -832 -4264
rect -826 -4272 -824 -4264
rect -816 -4272 -814 -4264
rect -800 -4272 -798 -4264
rect -790 -4272 -788 -4264
rect -782 -4272 -780 -4264
rect -772 -4272 -770 -4264
rect -756 -4272 -754 -4264
rect -748 -4272 -746 -4264
rect -732 -4272 -730 -4264
rect -716 -4272 -714 -4264
rect -708 -4272 -706 -4264
rect -698 -4272 -696 -4264
rect -572 -4272 -570 -4264
rect -562 -4272 -560 -4264
rect -546 -4272 -544 -4264
rect -536 -4272 -534 -4264
rect -520 -4272 -518 -4264
rect -510 -4272 -508 -4264
rect -502 -4272 -500 -4264
rect -492 -4272 -490 -4264
rect -476 -4272 -474 -4264
rect -468 -4272 -466 -4264
rect -458 -4272 -456 -4264
rect -442 -4272 -440 -4264
rect -432 -4272 -430 -4264
rect -424 -4272 -422 -4264
rect -414 -4272 -412 -4264
rect -398 -4272 -396 -4264
rect -390 -4272 -388 -4264
rect -374 -4272 -372 -4264
rect -358 -4272 -356 -4264
rect -350 -4272 -348 -4264
rect -340 -4272 -338 -4264
rect -214 -4272 -212 -4264
rect -204 -4272 -202 -4264
rect -188 -4272 -186 -4264
rect -178 -4272 -176 -4264
rect -162 -4272 -160 -4264
rect -152 -4272 -150 -4264
rect -144 -4272 -142 -4264
rect -134 -4272 -132 -4264
rect -118 -4272 -116 -4264
rect -110 -4272 -108 -4264
rect -100 -4272 -98 -4264
rect -84 -4272 -82 -4264
rect -74 -4272 -72 -4264
rect -66 -4272 -64 -4264
rect -56 -4272 -54 -4264
rect -40 -4272 -38 -4264
rect -32 -4272 -30 -4264
rect -16 -4272 -14 -4264
rect 0 -4272 2 -4264
rect 8 -4272 10 -4264
rect 18 -4272 20 -4264
rect 144 -4272 146 -4264
rect 154 -4272 156 -4264
rect 170 -4272 172 -4264
rect 180 -4272 182 -4264
rect 196 -4272 198 -4264
rect 206 -4272 208 -4264
rect 214 -4272 216 -4264
rect 224 -4272 226 -4264
rect 240 -4272 242 -4264
rect 248 -4272 250 -4264
rect 258 -4272 260 -4264
rect 274 -4272 276 -4264
rect 284 -4272 286 -4264
rect 292 -4272 294 -4264
rect 302 -4272 304 -4264
rect 318 -4272 320 -4264
rect 326 -4272 328 -4264
rect 342 -4272 344 -4264
rect 358 -4272 360 -4264
rect 366 -4272 368 -4264
rect 376 -4272 378 -4264
rect 500 -4272 502 -4264
rect 510 -4272 512 -4264
rect 526 -4272 528 -4264
rect 536 -4272 538 -4264
rect 552 -4272 554 -4264
rect 562 -4272 564 -4264
rect 570 -4272 572 -4264
rect 580 -4272 582 -4264
rect 596 -4272 598 -4264
rect 604 -4272 606 -4264
rect 614 -4272 616 -4264
rect 630 -4272 632 -4264
rect 640 -4272 642 -4264
rect 648 -4272 650 -4264
rect 658 -4272 660 -4264
rect 674 -4272 676 -4264
rect 682 -4272 684 -4264
rect 698 -4272 700 -4264
rect 714 -4272 716 -4264
rect 722 -4272 724 -4264
rect 732 -4272 734 -4264
rect 858 -4272 860 -4264
rect 868 -4272 870 -4264
rect 884 -4272 886 -4264
rect 894 -4272 896 -4264
rect 910 -4272 912 -4264
rect 920 -4272 922 -4264
rect 928 -4272 930 -4264
rect 938 -4272 940 -4264
rect 954 -4272 956 -4264
rect 962 -4272 964 -4264
rect 972 -4272 974 -4264
rect 988 -4272 990 -4264
rect 998 -4272 1000 -4264
rect 1006 -4272 1008 -4264
rect 1016 -4272 1018 -4264
rect 1032 -4272 1034 -4264
rect 1040 -4272 1042 -4264
rect 1056 -4272 1058 -4264
rect 1072 -4272 1074 -4264
rect 1080 -4272 1082 -4264
rect 1090 -4272 1092 -4264
rect 1216 -4272 1218 -4264
rect 1226 -4272 1228 -4264
rect 1242 -4272 1244 -4264
rect 1252 -4272 1254 -4264
rect 1268 -4272 1270 -4264
rect 1278 -4272 1280 -4264
rect 1286 -4272 1288 -4264
rect 1296 -4272 1298 -4264
rect 1312 -4272 1314 -4264
rect 1320 -4272 1322 -4264
rect 1330 -4272 1332 -4264
rect 1346 -4272 1348 -4264
rect 1356 -4272 1358 -4264
rect 1364 -4272 1366 -4264
rect 1374 -4272 1376 -4264
rect 1390 -4272 1392 -4264
rect 1398 -4272 1400 -4264
rect 1414 -4272 1416 -4264
rect 1430 -4272 1432 -4264
rect 1438 -4272 1440 -4264
rect 1448 -4272 1450 -4264
rect -1809 -4395 -1807 -4387
rect -1799 -4395 -1797 -4387
rect -1783 -4395 -1781 -4387
rect -1775 -4395 -1773 -4387
rect -1759 -4395 -1757 -4387
rect -1751 -4395 -1749 -4387
rect -1741 -4395 -1739 -4387
rect -1733 -4395 -1731 -4387
rect -1717 -4395 -1715 -4387
rect -1709 -4395 -1707 -4387
rect -1699 -4395 -1697 -4387
rect -1691 -4395 -1689 -4387
rect -1675 -4395 -1673 -4387
rect -1667 -4395 -1665 -4387
rect -1657 -4395 -1655 -4387
rect -1649 -4395 -1647 -4387
rect -1633 -4395 -1631 -4387
rect -1625 -4395 -1623 -4387
rect -1546 -4395 -1544 -4387
rect -1536 -4395 -1534 -4387
rect -1520 -4395 -1518 -4387
rect -1512 -4395 -1510 -4387
rect -1496 -4395 -1494 -4387
rect -1488 -4395 -1486 -4387
rect -1478 -4395 -1476 -4387
rect -1470 -4395 -1468 -4387
rect -1454 -4395 -1452 -4387
rect -1446 -4395 -1444 -4387
rect -1436 -4395 -1434 -4387
rect -1428 -4395 -1426 -4387
rect -1412 -4395 -1410 -4387
rect -1404 -4395 -1402 -4387
rect -1394 -4395 -1392 -4387
rect -1386 -4395 -1384 -4387
rect -1370 -4395 -1368 -4387
rect -1362 -4395 -1360 -4387
rect -1229 -4395 -1227 -4387
rect -1219 -4395 -1217 -4387
rect -1203 -4395 -1201 -4387
rect -1195 -4395 -1193 -4387
rect -1179 -4395 -1177 -4387
rect -1171 -4395 -1169 -4387
rect -1161 -4395 -1159 -4387
rect -1153 -4395 -1151 -4387
rect -1137 -4395 -1135 -4387
rect -1129 -4395 -1127 -4387
rect -1119 -4395 -1117 -4387
rect -1111 -4395 -1109 -4387
rect -1095 -4395 -1093 -4387
rect -1087 -4395 -1085 -4387
rect -1077 -4395 -1075 -4387
rect -1069 -4395 -1067 -4387
rect -1053 -4395 -1051 -4387
rect -1045 -4395 -1043 -4387
rect -930 -4395 -928 -4387
rect -920 -4395 -918 -4387
rect -904 -4395 -902 -4387
rect -896 -4395 -894 -4387
rect -880 -4395 -878 -4387
rect -872 -4395 -870 -4387
rect -862 -4395 -860 -4387
rect -854 -4395 -852 -4387
rect -838 -4395 -836 -4387
rect -830 -4395 -828 -4387
rect -820 -4395 -818 -4387
rect -812 -4395 -810 -4387
rect -796 -4395 -794 -4387
rect -788 -4395 -786 -4387
rect -778 -4395 -776 -4387
rect -770 -4395 -768 -4387
rect -754 -4395 -752 -4387
rect -746 -4395 -744 -4387
rect -572 -4395 -570 -4387
rect -562 -4395 -560 -4387
rect -546 -4395 -544 -4387
rect -538 -4395 -536 -4387
rect -522 -4395 -520 -4387
rect -514 -4395 -512 -4387
rect -504 -4395 -502 -4387
rect -496 -4395 -494 -4387
rect -480 -4395 -478 -4387
rect -472 -4395 -470 -4387
rect -462 -4395 -460 -4387
rect -454 -4395 -452 -4387
rect -438 -4395 -436 -4387
rect -430 -4395 -428 -4387
rect -420 -4395 -418 -4387
rect -412 -4395 -410 -4387
rect -396 -4395 -394 -4387
rect -388 -4395 -386 -4387
rect -1809 -4566 -1807 -4558
rect -1799 -4566 -1797 -4558
rect -1783 -4566 -1781 -4558
rect -1775 -4566 -1773 -4558
rect -1759 -4566 -1757 -4558
rect -1751 -4566 -1749 -4558
rect -1741 -4566 -1739 -4558
rect -1733 -4566 -1731 -4558
rect -1717 -4566 -1715 -4558
rect -1709 -4566 -1707 -4558
rect -1699 -4566 -1697 -4558
rect -1691 -4566 -1689 -4558
rect -1675 -4566 -1673 -4558
rect -1667 -4566 -1665 -4558
rect -1657 -4566 -1655 -4558
rect -1649 -4566 -1647 -4558
rect -1633 -4566 -1631 -4558
rect -1625 -4566 -1623 -4558
rect -1546 -4566 -1544 -4558
rect -1536 -4566 -1534 -4558
rect -1520 -4566 -1518 -4558
rect -1512 -4566 -1510 -4558
rect -1496 -4566 -1494 -4558
rect -1488 -4566 -1486 -4558
rect -1478 -4566 -1476 -4558
rect -1470 -4566 -1468 -4558
rect -1454 -4566 -1452 -4558
rect -1446 -4566 -1444 -4558
rect -1436 -4566 -1434 -4558
rect -1428 -4566 -1426 -4558
rect -1412 -4566 -1410 -4558
rect -1404 -4566 -1402 -4558
rect -1394 -4566 -1392 -4558
rect -1386 -4566 -1384 -4558
rect -1370 -4566 -1368 -4558
rect -1362 -4566 -1360 -4558
rect -1229 -4566 -1227 -4558
rect -1219 -4566 -1217 -4558
rect -1203 -4566 -1201 -4558
rect -1195 -4566 -1193 -4558
rect -1179 -4566 -1177 -4558
rect -1171 -4566 -1169 -4558
rect -1161 -4566 -1159 -4558
rect -1153 -4566 -1151 -4558
rect -1137 -4566 -1135 -4558
rect -1129 -4566 -1127 -4558
rect -1119 -4566 -1117 -4558
rect -1111 -4566 -1109 -4558
rect -1095 -4566 -1093 -4558
rect -1087 -4566 -1085 -4558
rect -1077 -4566 -1075 -4558
rect -1069 -4566 -1067 -4558
rect -1053 -4566 -1051 -4558
rect -1045 -4566 -1043 -4558
rect -930 -4566 -928 -4558
rect -920 -4566 -918 -4558
rect -904 -4566 -902 -4558
rect -896 -4566 -894 -4558
rect -880 -4566 -878 -4558
rect -872 -4566 -870 -4558
rect -862 -4566 -860 -4558
rect -854 -4566 -852 -4558
rect -838 -4566 -836 -4558
rect -830 -4566 -828 -4558
rect -820 -4566 -818 -4558
rect -812 -4566 -810 -4558
rect -796 -4566 -794 -4558
rect -788 -4566 -786 -4558
rect -778 -4566 -776 -4558
rect -770 -4566 -768 -4558
rect -754 -4566 -752 -4558
rect -746 -4566 -744 -4558
rect -572 -4566 -570 -4558
rect -562 -4566 -560 -4558
rect -546 -4566 -544 -4558
rect -538 -4566 -536 -4558
rect -522 -4566 -520 -4558
rect -514 -4566 -512 -4558
rect -504 -4566 -502 -4558
rect -496 -4566 -494 -4558
rect -480 -4566 -478 -4558
rect -472 -4566 -470 -4558
rect -462 -4566 -460 -4558
rect -454 -4566 -452 -4558
rect -438 -4566 -436 -4558
rect -430 -4566 -428 -4558
rect -420 -4566 -418 -4558
rect -412 -4566 -410 -4558
rect -396 -4566 -394 -4558
rect -388 -4566 -386 -4558
rect -214 -4566 -212 -4558
rect -204 -4566 -202 -4558
rect -188 -4566 -186 -4558
rect -180 -4566 -178 -4558
rect -164 -4566 -162 -4558
rect -156 -4566 -154 -4558
rect -146 -4566 -144 -4558
rect -138 -4566 -136 -4558
rect -122 -4566 -120 -4558
rect -114 -4566 -112 -4558
rect -104 -4566 -102 -4558
rect -96 -4566 -94 -4558
rect -80 -4566 -78 -4558
rect -72 -4566 -70 -4558
rect -62 -4566 -60 -4558
rect -54 -4566 -52 -4558
rect -38 -4566 -36 -4558
rect -30 -4566 -28 -4558
rect 144 -4566 146 -4558
rect 154 -4566 156 -4558
rect 170 -4566 172 -4558
rect 178 -4566 180 -4558
rect 194 -4566 196 -4558
rect 202 -4566 204 -4558
rect 212 -4566 214 -4558
rect 220 -4566 222 -4558
rect 236 -4566 238 -4558
rect 244 -4566 246 -4558
rect 254 -4566 256 -4558
rect 262 -4566 264 -4558
rect 278 -4566 280 -4558
rect 286 -4566 288 -4558
rect 296 -4566 298 -4558
rect 304 -4566 306 -4558
rect 320 -4566 322 -4558
rect 328 -4566 330 -4558
rect 500 -4566 502 -4558
rect 510 -4566 512 -4558
rect 526 -4566 528 -4558
rect 534 -4566 536 -4558
rect 550 -4566 552 -4558
rect 558 -4566 560 -4558
rect 568 -4566 570 -4558
rect 576 -4566 578 -4558
rect 592 -4566 594 -4558
rect 600 -4566 602 -4558
rect 610 -4566 612 -4558
rect 618 -4566 620 -4558
rect 634 -4566 636 -4558
rect 642 -4566 644 -4558
rect 652 -4566 654 -4558
rect 660 -4566 662 -4558
rect 676 -4566 678 -4558
rect 684 -4566 686 -4558
rect 858 -4566 860 -4558
rect 868 -4566 870 -4558
rect 884 -4566 886 -4558
rect 892 -4566 894 -4558
rect 908 -4566 910 -4558
rect 916 -4566 918 -4558
rect 926 -4566 928 -4558
rect 934 -4566 936 -4558
rect 950 -4566 952 -4558
rect 958 -4566 960 -4558
rect 968 -4566 970 -4558
rect 976 -4566 978 -4558
rect 992 -4566 994 -4558
rect 1000 -4566 1002 -4558
rect 1010 -4566 1012 -4558
rect 1018 -4566 1020 -4558
rect 1034 -4566 1036 -4558
rect 1042 -4566 1044 -4558
rect 1216 -4566 1218 -4558
rect 1226 -4566 1228 -4558
rect 1242 -4566 1244 -4558
rect 1250 -4566 1252 -4558
rect 1266 -4566 1268 -4558
rect 1274 -4566 1276 -4558
rect 1284 -4566 1286 -4558
rect 1292 -4566 1294 -4558
rect 1308 -4566 1310 -4558
rect 1316 -4566 1318 -4558
rect 1326 -4566 1328 -4558
rect 1334 -4566 1336 -4558
rect 1350 -4566 1352 -4558
rect 1358 -4566 1360 -4558
rect 1368 -4566 1370 -4558
rect 1376 -4566 1378 -4558
rect 1392 -4566 1394 -4558
rect 1400 -4566 1402 -4558
rect -1546 -4737 -1544 -4729
rect -1536 -4737 -1534 -4729
rect -1520 -4737 -1518 -4729
rect -1512 -4737 -1510 -4729
rect -1496 -4737 -1494 -4729
rect -1488 -4737 -1486 -4729
rect -1478 -4737 -1476 -4729
rect -1470 -4737 -1468 -4729
rect -1454 -4737 -1452 -4729
rect -1446 -4737 -1444 -4729
rect -1436 -4737 -1434 -4729
rect -1428 -4737 -1426 -4729
rect -1412 -4737 -1410 -4729
rect -1404 -4737 -1402 -4729
rect -1394 -4737 -1392 -4729
rect -1386 -4737 -1384 -4729
rect -1370 -4737 -1368 -4729
rect -1362 -4737 -1360 -4729
rect -1229 -4737 -1227 -4729
rect -1219 -4737 -1217 -4729
rect -1203 -4737 -1201 -4729
rect -1195 -4737 -1193 -4729
rect -1179 -4737 -1177 -4729
rect -1171 -4737 -1169 -4729
rect -1161 -4737 -1159 -4729
rect -1153 -4737 -1151 -4729
rect -1137 -4737 -1135 -4729
rect -1129 -4737 -1127 -4729
rect -1119 -4737 -1117 -4729
rect -1111 -4737 -1109 -4729
rect -1095 -4737 -1093 -4729
rect -1087 -4737 -1085 -4729
rect -1077 -4737 -1075 -4729
rect -1069 -4737 -1067 -4729
rect -1053 -4737 -1051 -4729
rect -1045 -4737 -1043 -4729
rect -930 -4737 -928 -4729
rect -920 -4737 -918 -4729
rect -904 -4737 -902 -4729
rect -896 -4737 -894 -4729
rect -880 -4737 -878 -4729
rect -872 -4737 -870 -4729
rect -862 -4737 -860 -4729
rect -854 -4737 -852 -4729
rect -838 -4737 -836 -4729
rect -830 -4737 -828 -4729
rect -820 -4737 -818 -4729
rect -812 -4737 -810 -4729
rect -796 -4737 -794 -4729
rect -788 -4737 -786 -4729
rect -778 -4737 -776 -4729
rect -770 -4737 -768 -4729
rect -754 -4737 -752 -4729
rect -746 -4737 -744 -4729
rect -572 -4737 -570 -4729
rect -562 -4737 -560 -4729
rect -546 -4737 -544 -4729
rect -538 -4737 -536 -4729
rect -522 -4737 -520 -4729
rect -514 -4737 -512 -4729
rect -504 -4737 -502 -4729
rect -496 -4737 -494 -4729
rect -480 -4737 -478 -4729
rect -472 -4737 -470 -4729
rect -462 -4737 -460 -4729
rect -454 -4737 -452 -4729
rect -438 -4737 -436 -4729
rect -430 -4737 -428 -4729
rect -420 -4737 -418 -4729
rect -412 -4737 -410 -4729
rect -396 -4737 -394 -4729
rect -388 -4737 -386 -4729
rect -214 -4737 -212 -4729
rect -204 -4737 -202 -4729
rect -188 -4737 -186 -4729
rect -180 -4737 -178 -4729
rect -164 -4737 -162 -4729
rect -156 -4737 -154 -4729
rect -146 -4737 -144 -4729
rect -138 -4737 -136 -4729
rect -122 -4737 -120 -4729
rect -114 -4737 -112 -4729
rect -104 -4737 -102 -4729
rect -96 -4737 -94 -4729
rect -80 -4737 -78 -4729
rect -72 -4737 -70 -4729
rect -62 -4737 -60 -4729
rect -54 -4737 -52 -4729
rect -38 -4737 -36 -4729
rect -30 -4737 -28 -4729
rect 144 -4737 146 -4729
rect 154 -4737 156 -4729
rect 170 -4737 172 -4729
rect 178 -4737 180 -4729
rect 194 -4737 196 -4729
rect 202 -4737 204 -4729
rect 212 -4737 214 -4729
rect 220 -4737 222 -4729
rect 236 -4737 238 -4729
rect 244 -4737 246 -4729
rect 254 -4737 256 -4729
rect 262 -4737 264 -4729
rect 278 -4737 280 -4729
rect 286 -4737 288 -4729
rect 296 -4737 298 -4729
rect 304 -4737 306 -4729
rect 320 -4737 322 -4729
rect 328 -4737 330 -4729
rect 500 -4737 502 -4729
rect 510 -4737 512 -4729
rect 526 -4737 528 -4729
rect 534 -4737 536 -4729
rect 550 -4737 552 -4729
rect 558 -4737 560 -4729
rect 568 -4737 570 -4729
rect 576 -4737 578 -4729
rect 592 -4737 594 -4729
rect 600 -4737 602 -4729
rect 610 -4737 612 -4729
rect 618 -4737 620 -4729
rect 634 -4737 636 -4729
rect 642 -4737 644 -4729
rect 652 -4737 654 -4729
rect 660 -4737 662 -4729
rect 676 -4737 678 -4729
rect 684 -4737 686 -4729
rect 858 -4737 860 -4729
rect 868 -4737 870 -4729
rect 884 -4737 886 -4729
rect 892 -4737 894 -4729
rect 908 -4737 910 -4729
rect 916 -4737 918 -4729
rect 926 -4737 928 -4729
rect 934 -4737 936 -4729
rect 950 -4737 952 -4729
rect 958 -4737 960 -4729
rect 968 -4737 970 -4729
rect 976 -4737 978 -4729
rect 992 -4737 994 -4729
rect 1000 -4737 1002 -4729
rect 1010 -4737 1012 -4729
rect 1018 -4737 1020 -4729
rect 1034 -4737 1036 -4729
rect 1042 -4737 1044 -4729
rect 1216 -4737 1218 -4729
rect 1226 -4737 1228 -4729
rect 1242 -4737 1244 -4729
rect 1250 -4737 1252 -4729
rect 1266 -4737 1268 -4729
rect 1274 -4737 1276 -4729
rect 1284 -4737 1286 -4729
rect 1292 -4737 1294 -4729
rect 1308 -4737 1310 -4729
rect 1316 -4737 1318 -4729
rect 1326 -4737 1328 -4729
rect 1334 -4737 1336 -4729
rect 1350 -4737 1352 -4729
rect 1358 -4737 1360 -4729
rect 1368 -4737 1370 -4729
rect 1376 -4737 1378 -4729
rect 1392 -4737 1394 -4729
rect 1400 -4737 1402 -4729
rect -1304 -4852 -1302 -4844
rect -1296 -4852 -1294 -4844
rect -1286 -4852 -1284 -4844
rect -930 -4852 -928 -4844
rect -922 -4852 -920 -4844
rect -912 -4852 -910 -4844
rect -572 -4852 -570 -4844
rect -564 -4852 -562 -4844
rect -554 -4852 -552 -4844
rect -214 -4852 -212 -4844
rect -206 -4852 -204 -4844
rect -196 -4852 -194 -4844
rect 144 -4852 146 -4844
rect 152 -4852 154 -4844
rect 162 -4852 164 -4844
rect 500 -4852 502 -4844
rect 508 -4852 510 -4844
rect 518 -4852 520 -4844
rect 858 -4852 860 -4844
rect 866 -4852 868 -4844
rect 876 -4852 878 -4844
rect 1216 -4852 1218 -4844
rect 1224 -4852 1226 -4844
rect 1234 -4852 1236 -4844
rect -1229 -5011 -1227 -5003
rect -1219 -5011 -1217 -5003
rect -1203 -5011 -1201 -5003
rect -1193 -5011 -1191 -5003
rect -1185 -5011 -1183 -5003
rect -1175 -5011 -1173 -5003
rect -1159 -5011 -1157 -5003
rect -1151 -5011 -1149 -5003
rect -1141 -5011 -1139 -5003
rect -930 -5011 -928 -5003
rect -920 -5011 -918 -5003
rect -904 -5011 -902 -5003
rect -894 -5011 -892 -5003
rect -878 -5011 -876 -5003
rect -868 -5011 -866 -5003
rect -860 -5011 -858 -5003
rect -850 -5011 -848 -5003
rect -834 -5011 -832 -5003
rect -826 -5011 -824 -5003
rect -816 -5011 -814 -5003
rect -800 -5011 -798 -5003
rect -790 -5011 -788 -5003
rect -782 -5011 -780 -5003
rect -772 -5011 -770 -5003
rect -756 -5011 -754 -5003
rect -748 -5011 -746 -5003
rect -732 -5011 -730 -5003
rect -716 -5011 -714 -5003
rect -708 -5011 -706 -5003
rect -698 -5011 -696 -5003
rect -572 -5011 -570 -5003
rect -562 -5011 -560 -5003
rect -546 -5011 -544 -5003
rect -536 -5011 -534 -5003
rect -520 -5011 -518 -5003
rect -510 -5011 -508 -5003
rect -502 -5011 -500 -5003
rect -492 -5011 -490 -5003
rect -476 -5011 -474 -5003
rect -468 -5011 -466 -5003
rect -458 -5011 -456 -5003
rect -442 -5011 -440 -5003
rect -432 -5011 -430 -5003
rect -424 -5011 -422 -5003
rect -414 -5011 -412 -5003
rect -398 -5011 -396 -5003
rect -390 -5011 -388 -5003
rect -374 -5011 -372 -5003
rect -358 -5011 -356 -5003
rect -350 -5011 -348 -5003
rect -340 -5011 -338 -5003
rect -214 -5011 -212 -5003
rect -204 -5011 -202 -5003
rect -188 -5011 -186 -5003
rect -178 -5011 -176 -5003
rect -162 -5011 -160 -5003
rect -152 -5011 -150 -5003
rect -144 -5011 -142 -5003
rect -134 -5011 -132 -5003
rect -118 -5011 -116 -5003
rect -110 -5011 -108 -5003
rect -100 -5011 -98 -5003
rect -84 -5011 -82 -5003
rect -74 -5011 -72 -5003
rect -66 -5011 -64 -5003
rect -56 -5011 -54 -5003
rect -40 -5011 -38 -5003
rect -32 -5011 -30 -5003
rect -16 -5011 -14 -5003
rect 0 -5011 2 -5003
rect 8 -5011 10 -5003
rect 18 -5011 20 -5003
rect 144 -5011 146 -5003
rect 154 -5011 156 -5003
rect 170 -5011 172 -5003
rect 180 -5011 182 -5003
rect 196 -5011 198 -5003
rect 206 -5011 208 -5003
rect 214 -5011 216 -5003
rect 224 -5011 226 -5003
rect 240 -5011 242 -5003
rect 248 -5011 250 -5003
rect 258 -5011 260 -5003
rect 274 -5011 276 -5003
rect 284 -5011 286 -5003
rect 292 -5011 294 -5003
rect 302 -5011 304 -5003
rect 318 -5011 320 -5003
rect 326 -5011 328 -5003
rect 342 -5011 344 -5003
rect 358 -5011 360 -5003
rect 366 -5011 368 -5003
rect 376 -5011 378 -5003
rect 500 -5011 502 -5003
rect 510 -5011 512 -5003
rect 526 -5011 528 -5003
rect 536 -5011 538 -5003
rect 552 -5011 554 -5003
rect 562 -5011 564 -5003
rect 570 -5011 572 -5003
rect 580 -5011 582 -5003
rect 596 -5011 598 -5003
rect 604 -5011 606 -5003
rect 614 -5011 616 -5003
rect 630 -5011 632 -5003
rect 640 -5011 642 -5003
rect 648 -5011 650 -5003
rect 658 -5011 660 -5003
rect 674 -5011 676 -5003
rect 682 -5011 684 -5003
rect 698 -5011 700 -5003
rect 714 -5011 716 -5003
rect 722 -5011 724 -5003
rect 732 -5011 734 -5003
rect 858 -5011 860 -5003
rect 868 -5011 870 -5003
rect 884 -5011 886 -5003
rect 894 -5011 896 -5003
rect 910 -5011 912 -5003
rect 920 -5011 922 -5003
rect 928 -5011 930 -5003
rect 938 -5011 940 -5003
rect 954 -5011 956 -5003
rect 962 -5011 964 -5003
rect 972 -5011 974 -5003
rect 988 -5011 990 -5003
rect 998 -5011 1000 -5003
rect 1006 -5011 1008 -5003
rect 1016 -5011 1018 -5003
rect 1032 -5011 1034 -5003
rect 1040 -5011 1042 -5003
rect 1056 -5011 1058 -5003
rect 1072 -5011 1074 -5003
rect 1080 -5011 1082 -5003
rect 1090 -5011 1092 -5003
rect 1216 -5011 1218 -5003
rect 1226 -5011 1228 -5003
rect 1242 -5011 1244 -5003
rect 1252 -5011 1254 -5003
rect 1268 -5011 1270 -5003
rect 1278 -5011 1280 -5003
rect 1286 -5011 1288 -5003
rect 1296 -5011 1298 -5003
rect 1312 -5011 1314 -5003
rect 1320 -5011 1322 -5003
rect 1330 -5011 1332 -5003
rect 1346 -5011 1348 -5003
rect 1356 -5011 1358 -5003
rect 1364 -5011 1366 -5003
rect 1374 -5011 1376 -5003
rect 1390 -5011 1392 -5003
rect 1398 -5011 1400 -5003
rect 1414 -5011 1416 -5003
rect 1430 -5011 1432 -5003
rect 1438 -5011 1440 -5003
rect 1448 -5011 1450 -5003
rect -1805 -5130 -1803 -5122
rect -1795 -5130 -1793 -5122
rect -1779 -5130 -1777 -5122
rect -1771 -5130 -1769 -5122
rect -1755 -5130 -1753 -5122
rect -1747 -5130 -1745 -5122
rect -1737 -5130 -1735 -5122
rect -1729 -5130 -1727 -5122
rect -1713 -5130 -1711 -5122
rect -1705 -5130 -1703 -5122
rect -1695 -5130 -1693 -5122
rect -1687 -5130 -1685 -5122
rect -1671 -5130 -1669 -5122
rect -1663 -5130 -1661 -5122
rect -1653 -5130 -1651 -5122
rect -1645 -5130 -1643 -5122
rect -1629 -5130 -1627 -5122
rect -1621 -5130 -1619 -5122
rect -1542 -5130 -1540 -5122
rect -1532 -5130 -1530 -5122
rect -1516 -5130 -1514 -5122
rect -1508 -5130 -1506 -5122
rect -1492 -5130 -1490 -5122
rect -1484 -5130 -1482 -5122
rect -1474 -5130 -1472 -5122
rect -1466 -5130 -1464 -5122
rect -1450 -5130 -1448 -5122
rect -1442 -5130 -1440 -5122
rect -1432 -5130 -1430 -5122
rect -1424 -5130 -1422 -5122
rect -1408 -5130 -1406 -5122
rect -1400 -5130 -1398 -5122
rect -1390 -5130 -1388 -5122
rect -1382 -5130 -1380 -5122
rect -1366 -5130 -1364 -5122
rect -1358 -5130 -1356 -5122
rect -1229 -5130 -1227 -5122
rect -1219 -5130 -1217 -5122
rect -1203 -5130 -1201 -5122
rect -1195 -5130 -1193 -5122
rect -1179 -5130 -1177 -5122
rect -1171 -5130 -1169 -5122
rect -1161 -5130 -1159 -5122
rect -1153 -5130 -1151 -5122
rect -1137 -5130 -1135 -5122
rect -1129 -5130 -1127 -5122
rect -1119 -5130 -1117 -5122
rect -1111 -5130 -1109 -5122
rect -1095 -5130 -1093 -5122
rect -1087 -5130 -1085 -5122
rect -1077 -5130 -1075 -5122
rect -1069 -5130 -1067 -5122
rect -1053 -5130 -1051 -5122
rect -1045 -5130 -1043 -5122
rect -930 -5130 -928 -5122
rect -920 -5130 -918 -5122
rect -904 -5130 -902 -5122
rect -896 -5130 -894 -5122
rect -880 -5130 -878 -5122
rect -872 -5130 -870 -5122
rect -862 -5130 -860 -5122
rect -854 -5130 -852 -5122
rect -838 -5130 -836 -5122
rect -830 -5130 -828 -5122
rect -820 -5130 -818 -5122
rect -812 -5130 -810 -5122
rect -796 -5130 -794 -5122
rect -788 -5130 -786 -5122
rect -778 -5130 -776 -5122
rect -770 -5130 -768 -5122
rect -754 -5130 -752 -5122
rect -746 -5130 -744 -5122
rect -1805 -5301 -1803 -5293
rect -1795 -5301 -1793 -5293
rect -1779 -5301 -1777 -5293
rect -1771 -5301 -1769 -5293
rect -1755 -5301 -1753 -5293
rect -1747 -5301 -1745 -5293
rect -1737 -5301 -1735 -5293
rect -1729 -5301 -1727 -5293
rect -1713 -5301 -1711 -5293
rect -1705 -5301 -1703 -5293
rect -1695 -5301 -1693 -5293
rect -1687 -5301 -1685 -5293
rect -1671 -5301 -1669 -5293
rect -1663 -5301 -1661 -5293
rect -1653 -5301 -1651 -5293
rect -1645 -5301 -1643 -5293
rect -1629 -5301 -1627 -5293
rect -1621 -5301 -1619 -5293
rect -1542 -5301 -1540 -5293
rect -1532 -5301 -1530 -5293
rect -1516 -5301 -1514 -5293
rect -1508 -5301 -1506 -5293
rect -1492 -5301 -1490 -5293
rect -1484 -5301 -1482 -5293
rect -1474 -5301 -1472 -5293
rect -1466 -5301 -1464 -5293
rect -1450 -5301 -1448 -5293
rect -1442 -5301 -1440 -5293
rect -1432 -5301 -1430 -5293
rect -1424 -5301 -1422 -5293
rect -1408 -5301 -1406 -5293
rect -1400 -5301 -1398 -5293
rect -1390 -5301 -1388 -5293
rect -1382 -5301 -1380 -5293
rect -1366 -5301 -1364 -5293
rect -1358 -5301 -1356 -5293
rect -1229 -5301 -1227 -5293
rect -1219 -5301 -1217 -5293
rect -1203 -5301 -1201 -5293
rect -1195 -5301 -1193 -5293
rect -1179 -5301 -1177 -5293
rect -1171 -5301 -1169 -5293
rect -1161 -5301 -1159 -5293
rect -1153 -5301 -1151 -5293
rect -1137 -5301 -1135 -5293
rect -1129 -5301 -1127 -5293
rect -1119 -5301 -1117 -5293
rect -1111 -5301 -1109 -5293
rect -1095 -5301 -1093 -5293
rect -1087 -5301 -1085 -5293
rect -1077 -5301 -1075 -5293
rect -1069 -5301 -1067 -5293
rect -1053 -5301 -1051 -5293
rect -1045 -5301 -1043 -5293
rect -930 -5301 -928 -5293
rect -920 -5301 -918 -5293
rect -904 -5301 -902 -5293
rect -896 -5301 -894 -5293
rect -880 -5301 -878 -5293
rect -872 -5301 -870 -5293
rect -862 -5301 -860 -5293
rect -854 -5301 -852 -5293
rect -838 -5301 -836 -5293
rect -830 -5301 -828 -5293
rect -820 -5301 -818 -5293
rect -812 -5301 -810 -5293
rect -796 -5301 -794 -5293
rect -788 -5301 -786 -5293
rect -778 -5301 -776 -5293
rect -770 -5301 -768 -5293
rect -754 -5301 -752 -5293
rect -746 -5301 -744 -5293
rect -572 -5301 -570 -5293
rect -562 -5301 -560 -5293
rect -546 -5301 -544 -5293
rect -538 -5301 -536 -5293
rect -522 -5301 -520 -5293
rect -514 -5301 -512 -5293
rect -504 -5301 -502 -5293
rect -496 -5301 -494 -5293
rect -480 -5301 -478 -5293
rect -472 -5301 -470 -5293
rect -462 -5301 -460 -5293
rect -454 -5301 -452 -5293
rect -438 -5301 -436 -5293
rect -430 -5301 -428 -5293
rect -420 -5301 -418 -5293
rect -412 -5301 -410 -5293
rect -396 -5301 -394 -5293
rect -388 -5301 -386 -5293
rect -214 -5301 -212 -5293
rect -204 -5301 -202 -5293
rect -188 -5301 -186 -5293
rect -180 -5301 -178 -5293
rect -164 -5301 -162 -5293
rect -156 -5301 -154 -5293
rect -146 -5301 -144 -5293
rect -138 -5301 -136 -5293
rect -122 -5301 -120 -5293
rect -114 -5301 -112 -5293
rect -104 -5301 -102 -5293
rect -96 -5301 -94 -5293
rect -80 -5301 -78 -5293
rect -72 -5301 -70 -5293
rect -62 -5301 -60 -5293
rect -54 -5301 -52 -5293
rect -38 -5301 -36 -5293
rect -30 -5301 -28 -5293
rect 144 -5301 146 -5293
rect 154 -5301 156 -5293
rect 170 -5301 172 -5293
rect 178 -5301 180 -5293
rect 194 -5301 196 -5293
rect 202 -5301 204 -5293
rect 212 -5301 214 -5293
rect 220 -5301 222 -5293
rect 236 -5301 238 -5293
rect 244 -5301 246 -5293
rect 254 -5301 256 -5293
rect 262 -5301 264 -5293
rect 278 -5301 280 -5293
rect 286 -5301 288 -5293
rect 296 -5301 298 -5293
rect 304 -5301 306 -5293
rect 320 -5301 322 -5293
rect 328 -5301 330 -5293
rect 500 -5301 502 -5293
rect 510 -5301 512 -5293
rect 526 -5301 528 -5293
rect 534 -5301 536 -5293
rect 550 -5301 552 -5293
rect 558 -5301 560 -5293
rect 568 -5301 570 -5293
rect 576 -5301 578 -5293
rect 592 -5301 594 -5293
rect 600 -5301 602 -5293
rect 610 -5301 612 -5293
rect 618 -5301 620 -5293
rect 634 -5301 636 -5293
rect 642 -5301 644 -5293
rect 652 -5301 654 -5293
rect 660 -5301 662 -5293
rect 676 -5301 678 -5293
rect 684 -5301 686 -5293
rect 858 -5301 860 -5293
rect 868 -5301 870 -5293
rect 884 -5301 886 -5293
rect 892 -5301 894 -5293
rect 908 -5301 910 -5293
rect 916 -5301 918 -5293
rect 926 -5301 928 -5293
rect 934 -5301 936 -5293
rect 950 -5301 952 -5293
rect 958 -5301 960 -5293
rect 968 -5301 970 -5293
rect 976 -5301 978 -5293
rect 992 -5301 994 -5293
rect 1000 -5301 1002 -5293
rect 1010 -5301 1012 -5293
rect 1018 -5301 1020 -5293
rect 1034 -5301 1036 -5293
rect 1042 -5301 1044 -5293
rect 1216 -5301 1218 -5293
rect 1226 -5301 1228 -5293
rect 1242 -5301 1244 -5293
rect 1250 -5301 1252 -5293
rect 1266 -5301 1268 -5293
rect 1274 -5301 1276 -5293
rect 1284 -5301 1286 -5293
rect 1292 -5301 1294 -5293
rect 1308 -5301 1310 -5293
rect 1316 -5301 1318 -5293
rect 1326 -5301 1328 -5293
rect 1334 -5301 1336 -5293
rect 1350 -5301 1352 -5293
rect 1358 -5301 1360 -5293
rect 1368 -5301 1370 -5293
rect 1376 -5301 1378 -5293
rect 1392 -5301 1394 -5293
rect 1400 -5301 1402 -5293
rect -1805 -5461 -1803 -5453
rect -1795 -5461 -1793 -5453
rect -1779 -5461 -1777 -5453
rect -1771 -5461 -1769 -5453
rect -1755 -5461 -1753 -5453
rect -1747 -5461 -1745 -5453
rect -1737 -5461 -1735 -5453
rect -1729 -5461 -1727 -5453
rect -1713 -5461 -1711 -5453
rect -1705 -5461 -1703 -5453
rect -1695 -5461 -1693 -5453
rect -1687 -5461 -1685 -5453
rect -1671 -5461 -1669 -5453
rect -1663 -5461 -1661 -5453
rect -1653 -5461 -1651 -5453
rect -1645 -5461 -1643 -5453
rect -1629 -5461 -1627 -5453
rect -1621 -5461 -1619 -5453
rect -1542 -5461 -1540 -5453
rect -1532 -5461 -1530 -5453
rect -1516 -5461 -1514 -5453
rect -1508 -5461 -1506 -5453
rect -1492 -5461 -1490 -5453
rect -1484 -5461 -1482 -5453
rect -1474 -5461 -1472 -5453
rect -1466 -5461 -1464 -5453
rect -1450 -5461 -1448 -5453
rect -1442 -5461 -1440 -5453
rect -1432 -5461 -1430 -5453
rect -1424 -5461 -1422 -5453
rect -1408 -5461 -1406 -5453
rect -1400 -5461 -1398 -5453
rect -1390 -5461 -1388 -5453
rect -1382 -5461 -1380 -5453
rect -1366 -5461 -1364 -5453
rect -1358 -5461 -1356 -5453
rect -1229 -5461 -1227 -5453
rect -1219 -5461 -1217 -5453
rect -1203 -5461 -1201 -5453
rect -1195 -5461 -1193 -5453
rect -1179 -5461 -1177 -5453
rect -1171 -5461 -1169 -5453
rect -1161 -5461 -1159 -5453
rect -1153 -5461 -1151 -5453
rect -1137 -5461 -1135 -5453
rect -1129 -5461 -1127 -5453
rect -1119 -5461 -1117 -5453
rect -1111 -5461 -1109 -5453
rect -1095 -5461 -1093 -5453
rect -1087 -5461 -1085 -5453
rect -1077 -5461 -1075 -5453
rect -1069 -5461 -1067 -5453
rect -1053 -5461 -1051 -5453
rect -1045 -5461 -1043 -5453
rect -930 -5461 -928 -5453
rect -920 -5461 -918 -5453
rect -904 -5461 -902 -5453
rect -896 -5461 -894 -5453
rect -880 -5461 -878 -5453
rect -872 -5461 -870 -5453
rect -862 -5461 -860 -5453
rect -854 -5461 -852 -5453
rect -838 -5461 -836 -5453
rect -830 -5461 -828 -5453
rect -820 -5461 -818 -5453
rect -812 -5461 -810 -5453
rect -796 -5461 -794 -5453
rect -788 -5461 -786 -5453
rect -778 -5461 -776 -5453
rect -770 -5461 -768 -5453
rect -754 -5461 -752 -5453
rect -746 -5461 -744 -5453
rect -572 -5461 -570 -5453
rect -562 -5461 -560 -5453
rect -546 -5461 -544 -5453
rect -538 -5461 -536 -5453
rect -522 -5461 -520 -5453
rect -514 -5461 -512 -5453
rect -504 -5461 -502 -5453
rect -496 -5461 -494 -5453
rect -480 -5461 -478 -5453
rect -472 -5461 -470 -5453
rect -462 -5461 -460 -5453
rect -454 -5461 -452 -5453
rect -438 -5461 -436 -5453
rect -430 -5461 -428 -5453
rect -420 -5461 -418 -5453
rect -412 -5461 -410 -5453
rect -396 -5461 -394 -5453
rect -388 -5461 -386 -5453
rect -214 -5461 -212 -5453
rect -204 -5461 -202 -5453
rect -188 -5461 -186 -5453
rect -180 -5461 -178 -5453
rect -164 -5461 -162 -5453
rect -156 -5461 -154 -5453
rect -146 -5461 -144 -5453
rect -138 -5461 -136 -5453
rect -122 -5461 -120 -5453
rect -114 -5461 -112 -5453
rect -104 -5461 -102 -5453
rect -96 -5461 -94 -5453
rect -80 -5461 -78 -5453
rect -72 -5461 -70 -5453
rect -62 -5461 -60 -5453
rect -54 -5461 -52 -5453
rect -38 -5461 -36 -5453
rect -30 -5461 -28 -5453
rect 144 -5461 146 -5453
rect 154 -5461 156 -5453
rect 170 -5461 172 -5453
rect 178 -5461 180 -5453
rect 194 -5461 196 -5453
rect 202 -5461 204 -5453
rect 212 -5461 214 -5453
rect 220 -5461 222 -5453
rect 236 -5461 238 -5453
rect 244 -5461 246 -5453
rect 254 -5461 256 -5453
rect 262 -5461 264 -5453
rect 278 -5461 280 -5453
rect 286 -5461 288 -5453
rect 296 -5461 298 -5453
rect 304 -5461 306 -5453
rect 320 -5461 322 -5453
rect 328 -5461 330 -5453
rect 500 -5461 502 -5453
rect 510 -5461 512 -5453
rect 526 -5461 528 -5453
rect 534 -5461 536 -5453
rect 550 -5461 552 -5453
rect 558 -5461 560 -5453
rect 568 -5461 570 -5453
rect 576 -5461 578 -5453
rect 592 -5461 594 -5453
rect 600 -5461 602 -5453
rect 610 -5461 612 -5453
rect 618 -5461 620 -5453
rect 634 -5461 636 -5453
rect 642 -5461 644 -5453
rect 652 -5461 654 -5453
rect 660 -5461 662 -5453
rect 676 -5461 678 -5453
rect 684 -5461 686 -5453
rect 858 -5461 860 -5453
rect 868 -5461 870 -5453
rect 884 -5461 886 -5453
rect 892 -5461 894 -5453
rect 908 -5461 910 -5453
rect 916 -5461 918 -5453
rect 926 -5461 928 -5453
rect 934 -5461 936 -5453
rect 950 -5461 952 -5453
rect 958 -5461 960 -5453
rect 968 -5461 970 -5453
rect 976 -5461 978 -5453
rect 992 -5461 994 -5453
rect 1000 -5461 1002 -5453
rect 1010 -5461 1012 -5453
rect 1018 -5461 1020 -5453
rect 1034 -5461 1036 -5453
rect 1042 -5461 1044 -5453
rect 1216 -5461 1218 -5453
rect 1226 -5461 1228 -5453
rect 1242 -5461 1244 -5453
rect 1250 -5461 1252 -5453
rect 1266 -5461 1268 -5453
rect 1274 -5461 1276 -5453
rect 1284 -5461 1286 -5453
rect 1292 -5461 1294 -5453
rect 1308 -5461 1310 -5453
rect 1316 -5461 1318 -5453
rect 1326 -5461 1328 -5453
rect 1334 -5461 1336 -5453
rect 1350 -5461 1352 -5453
rect 1358 -5461 1360 -5453
rect 1368 -5461 1370 -5453
rect 1376 -5461 1378 -5453
rect 1392 -5461 1394 -5453
rect 1400 -5461 1402 -5453
rect -1304 -5575 -1302 -5567
rect -1296 -5575 -1294 -5567
rect -1286 -5575 -1284 -5567
rect -930 -5575 -928 -5567
rect -922 -5575 -920 -5567
rect -912 -5575 -910 -5567
rect -572 -5575 -570 -5567
rect -564 -5575 -562 -5567
rect -554 -5575 -552 -5567
rect -214 -5575 -212 -5567
rect -206 -5575 -204 -5567
rect -196 -5575 -194 -5567
rect 144 -5575 146 -5567
rect 152 -5575 154 -5567
rect 162 -5575 164 -5567
rect 500 -5575 502 -5567
rect 508 -5575 510 -5567
rect 518 -5575 520 -5567
rect 858 -5575 860 -5567
rect 866 -5575 868 -5567
rect 876 -5575 878 -5567
rect 1216 -5575 1218 -5567
rect 1224 -5575 1226 -5567
rect 1234 -5575 1236 -5567
rect -1229 -5734 -1227 -5726
rect -1219 -5734 -1217 -5726
rect -1203 -5734 -1201 -5726
rect -1193 -5734 -1191 -5726
rect -1185 -5734 -1183 -5726
rect -1175 -5734 -1173 -5726
rect -1159 -5734 -1157 -5726
rect -1151 -5734 -1149 -5726
rect -1141 -5734 -1139 -5726
rect -930 -5734 -928 -5726
rect -920 -5734 -918 -5726
rect -904 -5734 -902 -5726
rect -894 -5734 -892 -5726
rect -878 -5734 -876 -5726
rect -868 -5734 -866 -5726
rect -860 -5734 -858 -5726
rect -850 -5734 -848 -5726
rect -834 -5734 -832 -5726
rect -826 -5734 -824 -5726
rect -816 -5734 -814 -5726
rect -800 -5734 -798 -5726
rect -790 -5734 -788 -5726
rect -782 -5734 -780 -5726
rect -772 -5734 -770 -5726
rect -756 -5734 -754 -5726
rect -748 -5734 -746 -5726
rect -732 -5734 -730 -5726
rect -716 -5734 -714 -5726
rect -708 -5734 -706 -5726
rect -698 -5734 -696 -5726
rect -572 -5734 -570 -5726
rect -562 -5734 -560 -5726
rect -546 -5734 -544 -5726
rect -536 -5734 -534 -5726
rect -520 -5734 -518 -5726
rect -510 -5734 -508 -5726
rect -502 -5734 -500 -5726
rect -492 -5734 -490 -5726
rect -476 -5734 -474 -5726
rect -468 -5734 -466 -5726
rect -458 -5734 -456 -5726
rect -442 -5734 -440 -5726
rect -432 -5734 -430 -5726
rect -424 -5734 -422 -5726
rect -414 -5734 -412 -5726
rect -398 -5734 -396 -5726
rect -390 -5734 -388 -5726
rect -374 -5734 -372 -5726
rect -358 -5734 -356 -5726
rect -350 -5734 -348 -5726
rect -340 -5734 -338 -5726
rect -214 -5734 -212 -5726
rect -204 -5734 -202 -5726
rect -188 -5734 -186 -5726
rect -178 -5734 -176 -5726
rect -162 -5734 -160 -5726
rect -152 -5734 -150 -5726
rect -144 -5734 -142 -5726
rect -134 -5734 -132 -5726
rect -118 -5734 -116 -5726
rect -110 -5734 -108 -5726
rect -100 -5734 -98 -5726
rect -84 -5734 -82 -5726
rect -74 -5734 -72 -5726
rect -66 -5734 -64 -5726
rect -56 -5734 -54 -5726
rect -40 -5734 -38 -5726
rect -32 -5734 -30 -5726
rect -16 -5734 -14 -5726
rect 0 -5734 2 -5726
rect 8 -5734 10 -5726
rect 18 -5734 20 -5726
rect 144 -5734 146 -5726
rect 154 -5734 156 -5726
rect 170 -5734 172 -5726
rect 180 -5734 182 -5726
rect 196 -5734 198 -5726
rect 206 -5734 208 -5726
rect 214 -5734 216 -5726
rect 224 -5734 226 -5726
rect 240 -5734 242 -5726
rect 248 -5734 250 -5726
rect 258 -5734 260 -5726
rect 274 -5734 276 -5726
rect 284 -5734 286 -5726
rect 292 -5734 294 -5726
rect 302 -5734 304 -5726
rect 318 -5734 320 -5726
rect 326 -5734 328 -5726
rect 342 -5734 344 -5726
rect 358 -5734 360 -5726
rect 366 -5734 368 -5726
rect 376 -5734 378 -5726
rect 500 -5734 502 -5726
rect 510 -5734 512 -5726
rect 526 -5734 528 -5726
rect 536 -5734 538 -5726
rect 552 -5734 554 -5726
rect 562 -5734 564 -5726
rect 570 -5734 572 -5726
rect 580 -5734 582 -5726
rect 596 -5734 598 -5726
rect 604 -5734 606 -5726
rect 614 -5734 616 -5726
rect 630 -5734 632 -5726
rect 640 -5734 642 -5726
rect 648 -5734 650 -5726
rect 658 -5734 660 -5726
rect 674 -5734 676 -5726
rect 682 -5734 684 -5726
rect 698 -5734 700 -5726
rect 714 -5734 716 -5726
rect 722 -5734 724 -5726
rect 732 -5734 734 -5726
rect 858 -5734 860 -5726
rect 868 -5734 870 -5726
rect 884 -5734 886 -5726
rect 894 -5734 896 -5726
rect 910 -5734 912 -5726
rect 920 -5734 922 -5726
rect 928 -5734 930 -5726
rect 938 -5734 940 -5726
rect 954 -5734 956 -5726
rect 962 -5734 964 -5726
rect 972 -5734 974 -5726
rect 988 -5734 990 -5726
rect 998 -5734 1000 -5726
rect 1006 -5734 1008 -5726
rect 1016 -5734 1018 -5726
rect 1032 -5734 1034 -5726
rect 1040 -5734 1042 -5726
rect 1056 -5734 1058 -5726
rect 1072 -5734 1074 -5726
rect 1080 -5734 1082 -5726
rect 1090 -5734 1092 -5726
rect 1216 -5734 1218 -5726
rect 1226 -5734 1228 -5726
rect 1242 -5734 1244 -5726
rect 1252 -5734 1254 -5726
rect 1268 -5734 1270 -5726
rect 1278 -5734 1280 -5726
rect 1286 -5734 1288 -5726
rect 1296 -5734 1298 -5726
rect 1312 -5734 1314 -5726
rect 1320 -5734 1322 -5726
rect 1330 -5734 1332 -5726
rect 1346 -5734 1348 -5726
rect 1356 -5734 1358 -5726
rect 1364 -5734 1366 -5726
rect 1374 -5734 1376 -5726
rect 1390 -5734 1392 -5726
rect 1398 -5734 1400 -5726
rect 1414 -5734 1416 -5726
rect 1430 -5734 1432 -5726
rect 1438 -5734 1440 -5726
rect 1448 -5734 1450 -5726
rect -1229 -5857 -1227 -5849
rect -1219 -5857 -1217 -5849
rect -1203 -5857 -1201 -5849
rect -1195 -5857 -1193 -5849
rect -1179 -5857 -1177 -5849
rect -1171 -5857 -1169 -5849
rect -1161 -5857 -1159 -5849
rect -1153 -5857 -1151 -5849
rect -1137 -5857 -1135 -5849
rect -1129 -5857 -1127 -5849
rect -1119 -5857 -1117 -5849
rect -1111 -5857 -1109 -5849
rect -1095 -5857 -1093 -5849
rect -1087 -5857 -1085 -5849
rect -1077 -5857 -1075 -5849
rect -1069 -5857 -1067 -5849
rect -1053 -5857 -1051 -5849
rect -1045 -5857 -1043 -5849
rect -930 -5857 -928 -5849
rect -920 -5857 -918 -5849
rect -904 -5857 -902 -5849
rect -896 -5857 -894 -5849
rect -880 -5857 -878 -5849
rect -872 -5857 -870 -5849
rect -862 -5857 -860 -5849
rect -854 -5857 -852 -5849
rect -838 -5857 -836 -5849
rect -830 -5857 -828 -5849
rect -820 -5857 -818 -5849
rect -812 -5857 -810 -5849
rect -796 -5857 -794 -5849
rect -788 -5857 -786 -5849
rect -778 -5857 -776 -5849
rect -770 -5857 -768 -5849
rect -754 -5857 -752 -5849
rect -746 -5857 -744 -5849
rect -572 -5857 -570 -5849
rect -562 -5857 -560 -5849
rect -546 -5857 -544 -5849
rect -538 -5857 -536 -5849
rect -522 -5857 -520 -5849
rect -514 -5857 -512 -5849
rect -504 -5857 -502 -5849
rect -496 -5857 -494 -5849
rect -480 -5857 -478 -5849
rect -472 -5857 -470 -5849
rect -462 -5857 -460 -5849
rect -454 -5857 -452 -5849
rect -438 -5857 -436 -5849
rect -430 -5857 -428 -5849
rect -420 -5857 -418 -5849
rect -412 -5857 -410 -5849
rect -396 -5857 -394 -5849
rect -388 -5857 -386 -5849
rect -214 -5857 -212 -5849
rect -204 -5857 -202 -5849
rect -188 -5857 -186 -5849
rect -180 -5857 -178 -5849
rect -164 -5857 -162 -5849
rect -156 -5857 -154 -5849
rect -146 -5857 -144 -5849
rect -138 -5857 -136 -5849
rect -122 -5857 -120 -5849
rect -114 -5857 -112 -5849
rect -104 -5857 -102 -5849
rect -96 -5857 -94 -5849
rect -80 -5857 -78 -5849
rect -72 -5857 -70 -5849
rect -62 -5857 -60 -5849
rect -54 -5857 -52 -5849
rect -38 -5857 -36 -5849
rect -30 -5857 -28 -5849
rect 144 -5857 146 -5849
rect 154 -5857 156 -5849
rect 170 -5857 172 -5849
rect 178 -5857 180 -5849
rect 194 -5857 196 -5849
rect 202 -5857 204 -5849
rect 212 -5857 214 -5849
rect 220 -5857 222 -5849
rect 236 -5857 238 -5849
rect 244 -5857 246 -5849
rect 254 -5857 256 -5849
rect 262 -5857 264 -5849
rect 278 -5857 280 -5849
rect 286 -5857 288 -5849
rect 296 -5857 298 -5849
rect 304 -5857 306 -5849
rect 320 -5857 322 -5849
rect 328 -5857 330 -5849
rect 500 -5857 502 -5849
rect 510 -5857 512 -5849
rect 526 -5857 528 -5849
rect 534 -5857 536 -5849
rect 550 -5857 552 -5849
rect 558 -5857 560 -5849
rect 568 -5857 570 -5849
rect 576 -5857 578 -5849
rect 592 -5857 594 -5849
rect 600 -5857 602 -5849
rect 610 -5857 612 -5849
rect 618 -5857 620 -5849
rect 634 -5857 636 -5849
rect 642 -5857 644 -5849
rect 652 -5857 654 -5849
rect 660 -5857 662 -5849
rect 676 -5857 678 -5849
rect 684 -5857 686 -5849
rect 858 -5857 860 -5849
rect 868 -5857 870 -5849
rect 884 -5857 886 -5849
rect 892 -5857 894 -5849
rect 908 -5857 910 -5849
rect 916 -5857 918 -5849
rect 926 -5857 928 -5849
rect 934 -5857 936 -5849
rect 950 -5857 952 -5849
rect 958 -5857 960 -5849
rect 968 -5857 970 -5849
rect 976 -5857 978 -5849
rect 992 -5857 994 -5849
rect 1000 -5857 1002 -5849
rect 1010 -5857 1012 -5849
rect 1018 -5857 1020 -5849
rect 1034 -5857 1036 -5849
rect 1042 -5857 1044 -5849
rect 1216 -5857 1218 -5849
rect 1226 -5857 1228 -5849
rect 1242 -5857 1244 -5849
rect 1250 -5857 1252 -5849
rect 1266 -5857 1268 -5849
rect 1274 -5857 1276 -5849
rect 1284 -5857 1286 -5849
rect 1292 -5857 1294 -5849
rect 1308 -5857 1310 -5849
rect 1316 -5857 1318 -5849
rect 1326 -5857 1328 -5849
rect 1334 -5857 1336 -5849
rect 1350 -5857 1352 -5849
rect 1358 -5857 1360 -5849
rect 1368 -5857 1370 -5849
rect 1376 -5857 1378 -5849
rect 1392 -5857 1394 -5849
rect 1400 -5857 1402 -5849
rect 1560 -5857 1562 -5849
rect 1570 -5857 1572 -5849
rect 1586 -5857 1588 -5849
rect 1594 -5857 1596 -5849
rect 1610 -5857 1612 -5849
rect 1618 -5857 1620 -5849
rect 1628 -5857 1630 -5849
rect 1636 -5857 1638 -5849
rect 1652 -5857 1654 -5849
rect 1660 -5857 1662 -5849
rect 1670 -5857 1672 -5849
rect 1678 -5857 1680 -5849
rect 1694 -5857 1696 -5849
rect 1702 -5857 1704 -5849
rect 1712 -5857 1714 -5849
rect 1720 -5857 1722 -5849
rect 1736 -5857 1738 -5849
rect 1744 -5857 1746 -5849
<< polycontact >>
rect -1306 -816 -1302 -812
rect -1295 -824 -1291 -820
rect -1288 -846 -1284 -842
rect -935 -816 -931 -812
rect -924 -824 -920 -820
rect -917 -848 -913 -844
rect -576 -816 -572 -812
rect -565 -824 -561 -820
rect -558 -848 -554 -844
rect -218 -816 -214 -812
rect -207 -824 -203 -820
rect -200 -848 -196 -844
rect 139 -816 143 -812
rect 150 -824 154 -820
rect 157 -861 161 -857
rect 496 -816 500 -812
rect 507 -824 511 -820
rect 514 -861 518 -857
rect 854 -816 858 -812
rect 865 -824 869 -820
rect 872 -861 876 -857
rect 1212 -816 1216 -812
rect 1223 -824 1227 -820
rect 1230 -861 1234 -857
rect -1223 -1074 -1219 -1070
rect -1219 -1088 -1215 -1084
rect -1203 -1066 -1199 -1062
rect -1203 -1095 -1199 -1091
rect -1189 -1074 -1185 -1070
rect -1179 -1081 -1175 -1077
rect -1165 -1066 -1161 -1062
rect -1161 -1095 -1157 -1091
rect -1137 -1074 -1133 -1070
rect -1147 -1081 -1143 -1077
rect -1123 -1095 -1119 -1091
rect -1105 -1066 -1101 -1062
rect -1095 -1081 -1091 -1077
rect -1105 -1088 -1101 -1084
rect -1081 -1066 -1077 -1062
rect -1077 -1074 -1073 -1070
rect -1063 -1081 -1059 -1077
rect -1053 -1088 -1049 -1084
rect -1039 -1074 -1035 -1070
rect -928 -1074 -924 -1070
rect -924 -1088 -920 -1084
rect -908 -1066 -904 -1062
rect -908 -1095 -904 -1091
rect -894 -1074 -890 -1070
rect -884 -1081 -880 -1077
rect -870 -1066 -866 -1062
rect -866 -1095 -862 -1091
rect -842 -1074 -838 -1070
rect -852 -1081 -848 -1077
rect -828 -1095 -824 -1091
rect -810 -1066 -806 -1062
rect -800 -1081 -796 -1077
rect -810 -1088 -806 -1084
rect -786 -1066 -782 -1062
rect -782 -1074 -778 -1070
rect -768 -1081 -764 -1077
rect -758 -1088 -754 -1084
rect -744 -1074 -740 -1070
rect -570 -1074 -566 -1070
rect -566 -1088 -562 -1084
rect -550 -1066 -546 -1062
rect -550 -1095 -546 -1091
rect -536 -1074 -532 -1070
rect -526 -1081 -522 -1077
rect -512 -1066 -508 -1062
rect -508 -1095 -504 -1091
rect -484 -1074 -480 -1070
rect -494 -1081 -490 -1077
rect -470 -1095 -466 -1091
rect -452 -1066 -448 -1062
rect -442 -1081 -438 -1077
rect -452 -1088 -448 -1084
rect -428 -1066 -424 -1062
rect -424 -1074 -420 -1070
rect -410 -1081 -406 -1077
rect -400 -1088 -396 -1084
rect -386 -1074 -382 -1070
rect -212 -1074 -208 -1070
rect -208 -1088 -204 -1084
rect -192 -1066 -188 -1062
rect -192 -1095 -188 -1091
rect -178 -1074 -174 -1070
rect -168 -1081 -164 -1077
rect -154 -1066 -150 -1062
rect -150 -1095 -146 -1091
rect -126 -1074 -122 -1070
rect -136 -1081 -132 -1077
rect -112 -1095 -108 -1091
rect -94 -1066 -90 -1062
rect -84 -1081 -80 -1077
rect -94 -1088 -90 -1084
rect -70 -1066 -66 -1062
rect -66 -1074 -62 -1070
rect -52 -1081 -48 -1077
rect -42 -1088 -38 -1084
rect -28 -1074 -24 -1070
rect 146 -1074 150 -1070
rect 150 -1088 154 -1084
rect 166 -1066 170 -1062
rect 166 -1095 170 -1091
rect 180 -1074 184 -1070
rect 190 -1081 194 -1077
rect 204 -1066 208 -1062
rect 208 -1095 212 -1091
rect 232 -1074 236 -1070
rect 222 -1081 226 -1077
rect 246 -1095 250 -1091
rect 264 -1066 268 -1062
rect 274 -1081 278 -1077
rect 264 -1088 268 -1084
rect 288 -1066 292 -1062
rect 292 -1074 296 -1070
rect 306 -1081 310 -1077
rect 316 -1088 320 -1084
rect 330 -1074 334 -1070
rect 502 -1074 506 -1070
rect 506 -1088 510 -1084
rect 522 -1066 526 -1062
rect 522 -1095 526 -1091
rect 536 -1074 540 -1070
rect 546 -1081 550 -1077
rect 560 -1066 564 -1062
rect 564 -1095 568 -1091
rect 588 -1074 592 -1070
rect 578 -1081 582 -1077
rect 602 -1095 606 -1091
rect 620 -1066 624 -1062
rect 630 -1081 634 -1077
rect 620 -1088 624 -1084
rect 644 -1066 648 -1062
rect 648 -1074 652 -1070
rect 662 -1081 666 -1077
rect 672 -1088 676 -1084
rect 686 -1074 690 -1070
rect 860 -1074 864 -1070
rect 864 -1088 868 -1084
rect 880 -1066 884 -1062
rect 880 -1095 884 -1091
rect 894 -1074 898 -1070
rect 904 -1081 908 -1077
rect 918 -1066 922 -1062
rect 922 -1095 926 -1091
rect 946 -1074 950 -1070
rect 936 -1081 940 -1077
rect 960 -1095 964 -1091
rect 978 -1066 982 -1062
rect 988 -1081 992 -1077
rect 978 -1088 982 -1084
rect 1002 -1066 1006 -1062
rect 1006 -1074 1010 -1070
rect 1020 -1081 1024 -1077
rect 1030 -1088 1034 -1084
rect 1044 -1074 1048 -1070
rect -1308 -1166 -1304 -1162
rect -1297 -1174 -1293 -1170
rect -1290 -1196 -1286 -1192
rect -934 -1166 -930 -1162
rect -923 -1174 -919 -1170
rect -916 -1196 -912 -1192
rect -576 -1166 -572 -1162
rect -565 -1174 -561 -1170
rect -558 -1196 -554 -1192
rect -218 -1166 -214 -1162
rect -207 -1174 -203 -1170
rect -200 -1196 -196 -1192
rect 140 -1166 144 -1162
rect 151 -1174 155 -1170
rect 158 -1196 162 -1192
rect 496 -1166 500 -1162
rect 507 -1174 511 -1170
rect 514 -1196 518 -1192
rect 854 -1166 858 -1162
rect 865 -1174 869 -1170
rect 872 -1196 876 -1192
rect 1212 -1166 1216 -1162
rect 1223 -1174 1227 -1170
rect 1230 -1196 1234 -1192
rect -1219 -1354 -1215 -1350
rect -1223 -1361 -1219 -1357
rect -1203 -1341 -1199 -1337
rect -1193 -1361 -1189 -1357
rect -1179 -1354 -1175 -1350
rect -1169 -1347 -1165 -1343
rect -1159 -1354 -1155 -1350
rect -1145 -1361 -1141 -1357
rect -1141 -1375 -1137 -1371
rect -924 -1317 -920 -1313
rect -928 -1338 -924 -1334
rect -924 -1353 -920 -1349
rect -928 -1367 -924 -1363
rect -898 -1338 -894 -1334
rect -902 -1346 -898 -1342
rect -902 -1360 -898 -1356
rect -882 -1324 -878 -1320
rect -872 -1367 -868 -1363
rect -858 -1317 -854 -1313
rect -848 -1331 -844 -1327
rect -838 -1367 -834 -1363
rect -824 -1317 -820 -1313
rect -820 -1375 -816 -1371
rect -804 -1346 -800 -1342
rect -794 -1360 -790 -1356
rect -780 -1317 -776 -1313
rect -780 -1338 -776 -1334
rect -776 -1353 -772 -1349
rect -760 -1360 -756 -1356
rect -746 -1317 -742 -1313
rect -736 -1368 -732 -1364
rect -720 -1375 -716 -1371
rect -706 -1331 -702 -1327
rect -702 -1368 -698 -1364
rect -566 -1317 -562 -1313
rect -570 -1338 -566 -1334
rect -566 -1353 -562 -1349
rect -570 -1367 -566 -1363
rect -540 -1338 -536 -1334
rect -544 -1346 -540 -1342
rect -544 -1360 -540 -1356
rect -524 -1324 -520 -1320
rect -514 -1367 -510 -1363
rect -500 -1317 -496 -1313
rect -490 -1331 -486 -1327
rect -480 -1367 -476 -1363
rect -466 -1317 -462 -1313
rect -462 -1375 -458 -1371
rect -446 -1346 -442 -1342
rect -436 -1360 -432 -1356
rect -422 -1317 -418 -1313
rect -422 -1338 -418 -1334
rect -418 -1353 -414 -1349
rect -402 -1360 -398 -1356
rect -388 -1317 -384 -1313
rect -378 -1368 -374 -1364
rect -362 -1375 -358 -1371
rect -348 -1331 -344 -1327
rect -344 -1368 -340 -1364
rect -208 -1317 -204 -1313
rect -212 -1338 -208 -1334
rect -208 -1353 -204 -1349
rect -212 -1367 -208 -1363
rect -182 -1338 -178 -1334
rect -186 -1346 -182 -1342
rect -186 -1360 -182 -1356
rect -166 -1324 -162 -1320
rect -156 -1367 -152 -1363
rect -142 -1317 -138 -1313
rect -132 -1331 -128 -1327
rect -122 -1367 -118 -1363
rect -108 -1317 -104 -1313
rect -104 -1375 -100 -1371
rect -88 -1346 -84 -1342
rect -78 -1360 -74 -1356
rect -64 -1317 -60 -1313
rect -64 -1338 -60 -1334
rect -60 -1353 -56 -1349
rect -44 -1360 -40 -1356
rect -30 -1317 -26 -1313
rect -20 -1368 -16 -1364
rect -4 -1375 0 -1371
rect 10 -1331 14 -1327
rect 14 -1368 18 -1364
rect 150 -1317 154 -1313
rect 146 -1338 150 -1334
rect 150 -1353 154 -1349
rect 146 -1367 150 -1363
rect 176 -1338 180 -1334
rect 172 -1346 176 -1342
rect 172 -1360 176 -1356
rect 192 -1324 196 -1320
rect 202 -1367 206 -1363
rect 216 -1317 220 -1313
rect 226 -1331 230 -1327
rect 236 -1367 240 -1363
rect 250 -1317 254 -1313
rect 254 -1375 258 -1371
rect 270 -1346 274 -1342
rect 280 -1360 284 -1356
rect 294 -1317 298 -1313
rect 294 -1338 298 -1334
rect 298 -1353 302 -1349
rect 314 -1360 318 -1356
rect 328 -1317 332 -1313
rect 338 -1368 342 -1364
rect 354 -1375 358 -1371
rect 368 -1331 372 -1327
rect 372 -1368 376 -1364
rect 506 -1317 510 -1313
rect 502 -1338 506 -1334
rect 506 -1353 510 -1349
rect 502 -1367 506 -1363
rect 532 -1338 536 -1334
rect 528 -1346 532 -1342
rect 528 -1360 532 -1356
rect 548 -1324 552 -1320
rect 558 -1367 562 -1363
rect 572 -1317 576 -1313
rect 582 -1331 586 -1327
rect 592 -1367 596 -1363
rect 606 -1317 610 -1313
rect 610 -1375 614 -1371
rect 626 -1346 630 -1342
rect 636 -1360 640 -1356
rect 650 -1317 654 -1313
rect 650 -1338 654 -1334
rect 654 -1353 658 -1349
rect 670 -1360 674 -1356
rect 684 -1317 688 -1313
rect 694 -1368 698 -1364
rect 710 -1375 714 -1371
rect 724 -1331 728 -1327
rect 728 -1368 732 -1364
rect 864 -1317 868 -1313
rect 860 -1338 864 -1334
rect 864 -1353 868 -1349
rect 860 -1367 864 -1363
rect 890 -1338 894 -1334
rect 886 -1346 890 -1342
rect 886 -1360 890 -1356
rect 906 -1324 910 -1320
rect 916 -1367 920 -1363
rect 930 -1317 934 -1313
rect 940 -1331 944 -1327
rect 950 -1367 954 -1363
rect 964 -1317 968 -1313
rect 968 -1375 972 -1371
rect 984 -1346 988 -1342
rect 994 -1360 998 -1356
rect 1008 -1317 1012 -1313
rect 1008 -1338 1012 -1334
rect 1012 -1353 1016 -1349
rect 1028 -1360 1032 -1356
rect 1042 -1317 1046 -1313
rect 1052 -1368 1056 -1364
rect 1068 -1375 1072 -1371
rect 1082 -1331 1086 -1327
rect 1086 -1368 1090 -1364
rect 1222 -1354 1226 -1350
rect 1218 -1361 1222 -1357
rect 1238 -1341 1242 -1337
rect 1248 -1361 1252 -1357
rect 1262 -1354 1266 -1350
rect 1272 -1347 1276 -1343
rect 1282 -1354 1286 -1350
rect 1296 -1361 1300 -1357
rect 1300 -1375 1304 -1371
rect -1223 -1477 -1219 -1473
rect -1219 -1491 -1215 -1487
rect -1203 -1469 -1199 -1465
rect -1203 -1498 -1199 -1494
rect -1189 -1477 -1185 -1473
rect -1179 -1484 -1175 -1480
rect -1165 -1469 -1161 -1465
rect -1161 -1498 -1157 -1494
rect -1137 -1477 -1133 -1473
rect -1147 -1484 -1143 -1480
rect -1123 -1498 -1119 -1494
rect -1105 -1469 -1101 -1465
rect -1095 -1484 -1091 -1480
rect -1105 -1491 -1101 -1487
rect -1081 -1469 -1077 -1465
rect -1077 -1477 -1073 -1473
rect -1063 -1484 -1059 -1480
rect -1053 -1491 -1049 -1487
rect -1039 -1477 -1035 -1473
rect -928 -1477 -924 -1473
rect -924 -1491 -920 -1487
rect -908 -1469 -904 -1465
rect -908 -1498 -904 -1494
rect -894 -1477 -890 -1473
rect -884 -1484 -880 -1480
rect -870 -1469 -866 -1465
rect -866 -1498 -862 -1494
rect -842 -1477 -838 -1473
rect -852 -1484 -848 -1480
rect -828 -1498 -824 -1494
rect -810 -1469 -806 -1465
rect -800 -1484 -796 -1480
rect -810 -1491 -806 -1487
rect -786 -1469 -782 -1465
rect -782 -1477 -778 -1473
rect -768 -1484 -764 -1480
rect -758 -1491 -754 -1487
rect -744 -1477 -740 -1473
rect -570 -1477 -566 -1473
rect -566 -1491 -562 -1487
rect -550 -1469 -546 -1465
rect -550 -1498 -546 -1494
rect -536 -1477 -532 -1473
rect -526 -1484 -522 -1480
rect -512 -1469 -508 -1465
rect -508 -1498 -504 -1494
rect -484 -1477 -480 -1473
rect -494 -1484 -490 -1480
rect -470 -1498 -466 -1494
rect -452 -1469 -448 -1465
rect -442 -1484 -438 -1480
rect -452 -1491 -448 -1487
rect -428 -1469 -424 -1465
rect -424 -1477 -420 -1473
rect -410 -1484 -406 -1480
rect -400 -1491 -396 -1487
rect -386 -1477 -382 -1473
rect -212 -1477 -208 -1473
rect -208 -1491 -204 -1487
rect -192 -1469 -188 -1465
rect -192 -1498 -188 -1494
rect -178 -1477 -174 -1473
rect -168 -1484 -164 -1480
rect -154 -1469 -150 -1465
rect -150 -1498 -146 -1494
rect -126 -1477 -122 -1473
rect -136 -1484 -132 -1480
rect -112 -1498 -108 -1494
rect -94 -1469 -90 -1465
rect -84 -1484 -80 -1480
rect -94 -1491 -90 -1487
rect -70 -1469 -66 -1465
rect -66 -1477 -62 -1473
rect -52 -1484 -48 -1480
rect -42 -1491 -38 -1487
rect -28 -1477 -24 -1473
rect 146 -1477 150 -1473
rect 150 -1491 154 -1487
rect 166 -1469 170 -1465
rect 166 -1498 170 -1494
rect 180 -1477 184 -1473
rect 190 -1484 194 -1480
rect 204 -1469 208 -1465
rect 208 -1498 212 -1494
rect 232 -1477 236 -1473
rect 222 -1484 226 -1480
rect 246 -1498 250 -1494
rect 264 -1469 268 -1465
rect 274 -1484 278 -1480
rect 264 -1491 268 -1487
rect 288 -1469 292 -1465
rect 292 -1477 296 -1473
rect 306 -1484 310 -1480
rect 316 -1491 320 -1487
rect 330 -1477 334 -1473
rect 502 -1477 506 -1473
rect 506 -1491 510 -1487
rect 522 -1469 526 -1465
rect 522 -1498 526 -1494
rect 536 -1477 540 -1473
rect 546 -1484 550 -1480
rect 560 -1469 564 -1465
rect 564 -1498 568 -1494
rect 588 -1477 592 -1473
rect 578 -1484 582 -1480
rect 602 -1498 606 -1494
rect 620 -1469 624 -1465
rect 630 -1484 634 -1480
rect 620 -1491 624 -1487
rect 644 -1469 648 -1465
rect 648 -1477 652 -1473
rect 662 -1484 666 -1480
rect 672 -1491 676 -1487
rect 686 -1477 690 -1473
rect 860 -1477 864 -1473
rect 864 -1491 868 -1487
rect 880 -1469 884 -1465
rect 880 -1498 884 -1494
rect 894 -1477 898 -1473
rect 904 -1484 908 -1480
rect 918 -1469 922 -1465
rect 922 -1498 926 -1494
rect 946 -1477 950 -1473
rect 936 -1484 940 -1480
rect 960 -1498 964 -1494
rect 978 -1469 982 -1465
rect 988 -1484 992 -1480
rect 978 -1491 982 -1487
rect 1002 -1469 1006 -1465
rect 1006 -1477 1010 -1473
rect 1020 -1484 1024 -1480
rect 1030 -1491 1034 -1487
rect 1044 -1477 1048 -1473
rect -1223 -1648 -1219 -1644
rect -1219 -1662 -1215 -1658
rect -1203 -1640 -1199 -1636
rect -1203 -1669 -1199 -1665
rect -1189 -1648 -1185 -1644
rect -1179 -1655 -1175 -1651
rect -1165 -1640 -1161 -1636
rect -1161 -1669 -1157 -1665
rect -1137 -1648 -1133 -1644
rect -1147 -1655 -1143 -1651
rect -1123 -1669 -1119 -1665
rect -1105 -1640 -1101 -1636
rect -1095 -1655 -1091 -1651
rect -1105 -1662 -1101 -1658
rect -1081 -1640 -1077 -1636
rect -1077 -1648 -1073 -1644
rect -1063 -1655 -1059 -1651
rect -1053 -1662 -1049 -1658
rect -1039 -1648 -1035 -1644
rect -928 -1648 -924 -1644
rect -924 -1662 -920 -1658
rect -908 -1640 -904 -1636
rect -908 -1669 -904 -1665
rect -894 -1648 -890 -1644
rect -884 -1655 -880 -1651
rect -870 -1640 -866 -1636
rect -866 -1669 -862 -1665
rect -842 -1648 -838 -1644
rect -852 -1655 -848 -1651
rect -828 -1669 -824 -1665
rect -810 -1640 -806 -1636
rect -800 -1655 -796 -1651
rect -810 -1662 -806 -1658
rect -786 -1640 -782 -1636
rect -782 -1648 -778 -1644
rect -768 -1655 -764 -1651
rect -758 -1662 -754 -1658
rect -744 -1648 -740 -1644
rect -570 -1648 -566 -1644
rect -566 -1662 -562 -1658
rect -550 -1640 -546 -1636
rect -550 -1669 -546 -1665
rect -536 -1648 -532 -1644
rect -526 -1655 -522 -1651
rect -512 -1640 -508 -1636
rect -508 -1669 -504 -1665
rect -484 -1648 -480 -1644
rect -494 -1655 -490 -1651
rect -470 -1669 -466 -1665
rect -452 -1640 -448 -1636
rect -442 -1655 -438 -1651
rect -452 -1662 -448 -1658
rect -428 -1640 -424 -1636
rect -424 -1648 -420 -1644
rect -410 -1655 -406 -1651
rect -400 -1662 -396 -1658
rect -386 -1648 -382 -1644
rect -212 -1648 -208 -1644
rect -208 -1662 -204 -1658
rect -192 -1640 -188 -1636
rect -192 -1669 -188 -1665
rect -178 -1648 -174 -1644
rect -168 -1655 -164 -1651
rect -154 -1640 -150 -1636
rect -150 -1669 -146 -1665
rect -126 -1648 -122 -1644
rect -136 -1655 -132 -1651
rect -112 -1669 -108 -1665
rect -94 -1640 -90 -1636
rect -84 -1655 -80 -1651
rect -94 -1662 -90 -1658
rect -70 -1640 -66 -1636
rect -66 -1648 -62 -1644
rect -52 -1655 -48 -1651
rect -42 -1662 -38 -1658
rect -28 -1648 -24 -1644
rect 146 -1648 150 -1644
rect 150 -1662 154 -1658
rect 166 -1640 170 -1636
rect 166 -1669 170 -1665
rect 180 -1648 184 -1644
rect 190 -1655 194 -1651
rect 204 -1640 208 -1636
rect 208 -1669 212 -1665
rect 232 -1648 236 -1644
rect 222 -1655 226 -1651
rect 246 -1669 250 -1665
rect 264 -1640 268 -1636
rect 274 -1655 278 -1651
rect 264 -1662 268 -1658
rect 288 -1640 292 -1636
rect 292 -1648 296 -1644
rect 306 -1655 310 -1651
rect 316 -1662 320 -1658
rect 330 -1648 334 -1644
rect 502 -1648 506 -1644
rect 506 -1662 510 -1658
rect 522 -1640 526 -1636
rect 522 -1669 526 -1665
rect 536 -1648 540 -1644
rect 546 -1655 550 -1651
rect 560 -1640 564 -1636
rect 564 -1669 568 -1665
rect 588 -1648 592 -1644
rect 578 -1655 582 -1651
rect 602 -1669 606 -1665
rect 620 -1640 624 -1636
rect 630 -1655 634 -1651
rect 620 -1662 624 -1658
rect 644 -1640 648 -1636
rect 648 -1648 652 -1644
rect 662 -1655 666 -1651
rect 672 -1662 676 -1658
rect 686 -1648 690 -1644
rect 860 -1648 864 -1644
rect 864 -1662 868 -1658
rect 880 -1640 884 -1636
rect 880 -1669 884 -1665
rect 894 -1648 898 -1644
rect 904 -1655 908 -1651
rect 918 -1640 922 -1636
rect 922 -1669 926 -1665
rect 946 -1648 950 -1644
rect 936 -1655 940 -1651
rect 960 -1669 964 -1665
rect 978 -1640 982 -1636
rect 988 -1655 992 -1651
rect 978 -1662 982 -1658
rect 1002 -1640 1006 -1636
rect 1006 -1648 1010 -1644
rect 1020 -1655 1024 -1651
rect 1030 -1662 1034 -1658
rect 1044 -1648 1048 -1644
rect 1218 -1648 1222 -1644
rect 1222 -1662 1226 -1658
rect 1238 -1640 1242 -1636
rect 1238 -1669 1242 -1665
rect 1252 -1648 1256 -1644
rect 1262 -1655 1266 -1651
rect 1276 -1640 1280 -1636
rect 1280 -1669 1284 -1665
rect 1304 -1648 1308 -1644
rect 1294 -1655 1298 -1651
rect 1318 -1669 1322 -1665
rect 1336 -1640 1340 -1636
rect 1346 -1655 1350 -1651
rect 1336 -1662 1340 -1658
rect 1360 -1640 1364 -1636
rect 1364 -1648 1368 -1644
rect 1378 -1655 1382 -1651
rect 1388 -1662 1392 -1658
rect 1402 -1648 1406 -1644
rect -1552 -1819 -1548 -1815
rect -1548 -1833 -1544 -1829
rect -1532 -1811 -1528 -1807
rect -1532 -1840 -1528 -1836
rect -1518 -1819 -1514 -1815
rect -1508 -1826 -1504 -1822
rect -1494 -1811 -1490 -1807
rect -1490 -1840 -1486 -1836
rect -1466 -1819 -1462 -1815
rect -1476 -1826 -1472 -1822
rect -1452 -1840 -1448 -1836
rect -1434 -1811 -1430 -1807
rect -1424 -1826 -1420 -1822
rect -1434 -1833 -1430 -1829
rect -1410 -1811 -1406 -1807
rect -1406 -1819 -1402 -1815
rect -1392 -1826 -1388 -1822
rect -1382 -1833 -1378 -1829
rect -1368 -1819 -1364 -1815
rect -1223 -1819 -1219 -1815
rect -1219 -1833 -1215 -1829
rect -1203 -1811 -1199 -1807
rect -1203 -1840 -1199 -1836
rect -1189 -1819 -1185 -1815
rect -1179 -1826 -1175 -1822
rect -1165 -1811 -1161 -1807
rect -1161 -1840 -1157 -1836
rect -1137 -1819 -1133 -1815
rect -1147 -1826 -1143 -1822
rect -1123 -1840 -1119 -1836
rect -1105 -1811 -1101 -1807
rect -1095 -1826 -1091 -1822
rect -1105 -1833 -1101 -1829
rect -1081 -1811 -1077 -1807
rect -1077 -1819 -1073 -1815
rect -1063 -1826 -1059 -1822
rect -1053 -1833 -1049 -1829
rect -1039 -1819 -1035 -1815
rect -928 -1819 -924 -1815
rect -924 -1833 -920 -1829
rect -908 -1811 -904 -1807
rect -908 -1840 -904 -1836
rect -894 -1819 -890 -1815
rect -884 -1826 -880 -1822
rect -870 -1811 -866 -1807
rect -866 -1840 -862 -1836
rect -842 -1819 -838 -1815
rect -852 -1826 -848 -1822
rect -828 -1840 -824 -1836
rect -810 -1811 -806 -1807
rect -800 -1826 -796 -1822
rect -810 -1833 -806 -1829
rect -786 -1811 -782 -1807
rect -782 -1819 -778 -1815
rect -768 -1826 -764 -1822
rect -758 -1833 -754 -1829
rect -744 -1819 -740 -1815
rect -570 -1819 -566 -1815
rect -566 -1833 -562 -1829
rect -550 -1811 -546 -1807
rect -550 -1840 -546 -1836
rect -536 -1819 -532 -1815
rect -526 -1826 -522 -1822
rect -512 -1811 -508 -1807
rect -508 -1840 -504 -1836
rect -484 -1819 -480 -1815
rect -494 -1826 -490 -1822
rect -470 -1840 -466 -1836
rect -452 -1811 -448 -1807
rect -442 -1826 -438 -1822
rect -452 -1833 -448 -1829
rect -428 -1811 -424 -1807
rect -424 -1819 -420 -1815
rect -410 -1826 -406 -1822
rect -400 -1833 -396 -1829
rect -386 -1819 -382 -1815
rect -212 -1819 -208 -1815
rect -208 -1833 -204 -1829
rect -192 -1811 -188 -1807
rect -192 -1840 -188 -1836
rect -178 -1819 -174 -1815
rect -168 -1826 -164 -1822
rect -154 -1811 -150 -1807
rect -150 -1840 -146 -1836
rect -126 -1819 -122 -1815
rect -136 -1826 -132 -1822
rect -112 -1840 -108 -1836
rect -94 -1811 -90 -1807
rect -84 -1826 -80 -1822
rect -94 -1833 -90 -1829
rect -70 -1811 -66 -1807
rect -66 -1819 -62 -1815
rect -52 -1826 -48 -1822
rect -42 -1833 -38 -1829
rect -28 -1819 -24 -1815
rect 146 -1819 150 -1815
rect 150 -1833 154 -1829
rect 166 -1811 170 -1807
rect 166 -1840 170 -1836
rect 180 -1819 184 -1815
rect 190 -1826 194 -1822
rect 204 -1811 208 -1807
rect 208 -1840 212 -1836
rect 232 -1819 236 -1815
rect 222 -1826 226 -1822
rect 246 -1840 250 -1836
rect 264 -1811 268 -1807
rect 274 -1826 278 -1822
rect 264 -1833 268 -1829
rect 288 -1811 292 -1807
rect 292 -1819 296 -1815
rect 306 -1826 310 -1822
rect 316 -1833 320 -1829
rect 330 -1819 334 -1815
rect 502 -1819 506 -1815
rect 506 -1833 510 -1829
rect 522 -1811 526 -1807
rect 522 -1840 526 -1836
rect 536 -1819 540 -1815
rect 546 -1826 550 -1822
rect 560 -1811 564 -1807
rect 564 -1840 568 -1836
rect 588 -1819 592 -1815
rect 578 -1826 582 -1822
rect 602 -1840 606 -1836
rect 620 -1811 624 -1807
rect 630 -1826 634 -1822
rect 620 -1833 624 -1829
rect 644 -1811 648 -1807
rect 648 -1819 652 -1815
rect 662 -1826 666 -1822
rect 672 -1833 676 -1829
rect 686 -1819 690 -1815
rect 860 -1819 864 -1815
rect 864 -1833 868 -1829
rect 880 -1811 884 -1807
rect 880 -1840 884 -1836
rect 894 -1819 898 -1815
rect 904 -1826 908 -1822
rect 918 -1811 922 -1807
rect 922 -1840 926 -1836
rect 946 -1819 950 -1815
rect 936 -1826 940 -1822
rect 960 -1840 964 -1836
rect 978 -1811 982 -1807
rect 988 -1826 992 -1822
rect 978 -1833 982 -1829
rect 1002 -1811 1006 -1807
rect 1006 -1819 1010 -1815
rect 1020 -1826 1024 -1822
rect 1030 -1833 1034 -1829
rect 1044 -1819 1048 -1815
rect 1218 -1819 1222 -1815
rect 1222 -1833 1226 -1829
rect 1238 -1811 1242 -1807
rect 1238 -1840 1242 -1836
rect 1252 -1819 1256 -1815
rect 1262 -1826 1266 -1822
rect 1276 -1811 1280 -1807
rect 1280 -1840 1284 -1836
rect 1304 -1819 1308 -1815
rect 1294 -1826 1298 -1822
rect 1318 -1840 1322 -1836
rect 1336 -1811 1340 -1807
rect 1346 -1826 1350 -1822
rect 1336 -1833 1340 -1829
rect 1360 -1811 1364 -1807
rect 1364 -1819 1368 -1815
rect 1378 -1826 1382 -1822
rect 1388 -1833 1392 -1829
rect 1402 -1819 1406 -1815
rect -1308 -1902 -1304 -1898
rect -1297 -1910 -1293 -1906
rect -1290 -1932 -1286 -1928
rect -934 -1902 -930 -1898
rect -923 -1910 -919 -1906
rect -916 -1932 -912 -1928
rect -576 -1902 -572 -1898
rect -565 -1910 -561 -1906
rect -558 -1932 -554 -1928
rect -218 -1902 -214 -1898
rect -207 -1910 -203 -1906
rect -200 -1932 -196 -1928
rect 140 -1902 144 -1898
rect 151 -1910 155 -1906
rect 158 -1932 162 -1928
rect 496 -1902 500 -1898
rect 507 -1910 511 -1906
rect 514 -1932 518 -1928
rect 854 -1902 858 -1898
rect 865 -1910 869 -1906
rect 872 -1932 876 -1928
rect 1212 -1902 1216 -1898
rect 1223 -1910 1227 -1906
rect 1230 -1932 1234 -1928
rect -1223 -2085 -1219 -2081
rect -1227 -2092 -1223 -2088
rect -1207 -2072 -1203 -2068
rect -1197 -2092 -1193 -2088
rect -1183 -2085 -1179 -2081
rect -1173 -2078 -1169 -2074
rect -1163 -2085 -1159 -2081
rect -1149 -2092 -1145 -2088
rect -1145 -2106 -1141 -2102
rect -924 -2048 -920 -2044
rect -928 -2069 -924 -2065
rect -924 -2084 -920 -2080
rect -928 -2098 -924 -2094
rect -898 -2069 -894 -2065
rect -902 -2077 -898 -2073
rect -902 -2091 -898 -2087
rect -882 -2055 -878 -2051
rect -872 -2098 -868 -2094
rect -858 -2048 -854 -2044
rect -848 -2062 -844 -2058
rect -838 -2098 -834 -2094
rect -824 -2048 -820 -2044
rect -820 -2106 -816 -2102
rect -804 -2077 -800 -2073
rect -794 -2091 -790 -2087
rect -780 -2048 -776 -2044
rect -780 -2069 -776 -2065
rect -776 -2084 -772 -2080
rect -760 -2091 -756 -2087
rect -746 -2048 -742 -2044
rect -736 -2099 -732 -2095
rect -720 -2106 -716 -2102
rect -706 -2062 -702 -2058
rect -702 -2099 -698 -2095
rect -566 -2048 -562 -2044
rect -570 -2069 -566 -2065
rect -566 -2084 -562 -2080
rect -570 -2098 -566 -2094
rect -540 -2069 -536 -2065
rect -544 -2077 -540 -2073
rect -544 -2091 -540 -2087
rect -524 -2055 -520 -2051
rect -514 -2098 -510 -2094
rect -500 -2048 -496 -2044
rect -490 -2062 -486 -2058
rect -480 -2098 -476 -2094
rect -466 -2048 -462 -2044
rect -462 -2106 -458 -2102
rect -446 -2077 -442 -2073
rect -436 -2091 -432 -2087
rect -422 -2048 -418 -2044
rect -422 -2069 -418 -2065
rect -418 -2084 -414 -2080
rect -402 -2091 -398 -2087
rect -388 -2048 -384 -2044
rect -378 -2099 -374 -2095
rect -362 -2106 -358 -2102
rect -348 -2062 -344 -2058
rect -344 -2099 -340 -2095
rect -208 -2048 -204 -2044
rect -212 -2069 -208 -2065
rect -208 -2084 -204 -2080
rect -212 -2098 -208 -2094
rect -182 -2069 -178 -2065
rect -186 -2077 -182 -2073
rect -186 -2091 -182 -2087
rect -166 -2055 -162 -2051
rect -156 -2098 -152 -2094
rect -142 -2048 -138 -2044
rect -132 -2062 -128 -2058
rect -122 -2098 -118 -2094
rect -108 -2048 -104 -2044
rect -104 -2106 -100 -2102
rect -88 -2077 -84 -2073
rect -78 -2091 -74 -2087
rect -64 -2048 -60 -2044
rect -64 -2069 -60 -2065
rect -60 -2084 -56 -2080
rect -44 -2091 -40 -2087
rect -30 -2048 -26 -2044
rect -20 -2099 -16 -2095
rect -4 -2106 0 -2102
rect 10 -2062 14 -2058
rect 14 -2099 18 -2095
rect 150 -2048 154 -2044
rect 146 -2069 150 -2065
rect 150 -2084 154 -2080
rect 146 -2098 150 -2094
rect 176 -2069 180 -2065
rect 172 -2077 176 -2073
rect 172 -2091 176 -2087
rect 192 -2055 196 -2051
rect 202 -2098 206 -2094
rect 216 -2048 220 -2044
rect 226 -2062 230 -2058
rect 236 -2098 240 -2094
rect 250 -2048 254 -2044
rect 254 -2106 258 -2102
rect 270 -2077 274 -2073
rect 280 -2091 284 -2087
rect 294 -2048 298 -2044
rect 294 -2069 298 -2065
rect 298 -2084 302 -2080
rect 314 -2091 318 -2087
rect 328 -2048 332 -2044
rect 338 -2099 342 -2095
rect 354 -2106 358 -2102
rect 368 -2062 372 -2058
rect 372 -2099 376 -2095
rect 506 -2048 510 -2044
rect 502 -2069 506 -2065
rect 506 -2084 510 -2080
rect 502 -2098 506 -2094
rect 532 -2069 536 -2065
rect 528 -2077 532 -2073
rect 528 -2091 532 -2087
rect 548 -2055 552 -2051
rect 558 -2098 562 -2094
rect 572 -2048 576 -2044
rect 582 -2062 586 -2058
rect 592 -2098 596 -2094
rect 606 -2048 610 -2044
rect 610 -2106 614 -2102
rect 626 -2077 630 -2073
rect 636 -2091 640 -2087
rect 650 -2048 654 -2044
rect 650 -2069 654 -2065
rect 654 -2084 658 -2080
rect 670 -2091 674 -2087
rect 684 -2048 688 -2044
rect 694 -2099 698 -2095
rect 710 -2106 714 -2102
rect 724 -2062 728 -2058
rect 728 -2099 732 -2095
rect 864 -2048 868 -2044
rect 860 -2069 864 -2065
rect 864 -2084 868 -2080
rect 860 -2098 864 -2094
rect 890 -2069 894 -2065
rect 886 -2077 890 -2073
rect 886 -2091 890 -2087
rect 906 -2055 910 -2051
rect 916 -2098 920 -2094
rect 930 -2048 934 -2044
rect 940 -2062 944 -2058
rect 950 -2098 954 -2094
rect 964 -2048 968 -2044
rect 968 -2106 972 -2102
rect 984 -2077 988 -2073
rect 994 -2091 998 -2087
rect 1008 -2048 1012 -2044
rect 1008 -2069 1012 -2065
rect 1012 -2084 1016 -2080
rect 1028 -2091 1032 -2087
rect 1042 -2048 1046 -2044
rect 1052 -2099 1056 -2095
rect 1068 -2106 1072 -2102
rect 1082 -2062 1086 -2058
rect 1086 -2099 1090 -2095
rect 1222 -2048 1226 -2044
rect 1218 -2069 1222 -2065
rect 1222 -2084 1226 -2080
rect 1218 -2098 1222 -2094
rect 1248 -2069 1252 -2065
rect 1244 -2077 1248 -2073
rect 1244 -2091 1248 -2087
rect 1264 -2055 1268 -2051
rect 1274 -2098 1278 -2094
rect 1288 -2048 1292 -2044
rect 1298 -2062 1302 -2058
rect 1308 -2098 1312 -2094
rect 1322 -2048 1326 -2044
rect 1326 -2106 1330 -2102
rect 1342 -2077 1346 -2073
rect 1352 -2091 1356 -2087
rect 1366 -2048 1370 -2044
rect 1366 -2069 1370 -2065
rect 1370 -2084 1374 -2080
rect 1386 -2091 1390 -2087
rect 1400 -2048 1404 -2044
rect 1410 -2099 1414 -2095
rect 1426 -2106 1430 -2102
rect 1440 -2062 1444 -2058
rect 1444 -2099 1448 -2095
rect -1227 -2229 -1223 -2225
rect -1223 -2243 -1219 -2239
rect -1207 -2221 -1203 -2217
rect -1207 -2250 -1203 -2246
rect -1193 -2229 -1189 -2225
rect -1183 -2236 -1179 -2232
rect -1169 -2221 -1165 -2217
rect -1165 -2250 -1161 -2246
rect -1141 -2229 -1137 -2225
rect -1151 -2236 -1147 -2232
rect -1127 -2250 -1123 -2246
rect -1109 -2221 -1105 -2217
rect -1099 -2236 -1095 -2232
rect -1109 -2243 -1105 -2239
rect -1085 -2221 -1081 -2217
rect -1081 -2229 -1077 -2225
rect -1067 -2236 -1063 -2232
rect -1057 -2243 -1053 -2239
rect -1043 -2229 -1039 -2225
rect -928 -2229 -924 -2225
rect -924 -2243 -920 -2239
rect -908 -2221 -904 -2217
rect -908 -2250 -904 -2246
rect -894 -2229 -890 -2225
rect -884 -2236 -880 -2232
rect -870 -2221 -866 -2217
rect -866 -2250 -862 -2246
rect -842 -2229 -838 -2225
rect -852 -2236 -848 -2232
rect -828 -2250 -824 -2246
rect -810 -2221 -806 -2217
rect -800 -2236 -796 -2232
rect -810 -2243 -806 -2239
rect -786 -2221 -782 -2217
rect -782 -2229 -778 -2225
rect -768 -2236 -764 -2232
rect -758 -2243 -754 -2239
rect -744 -2229 -740 -2225
rect -570 -2229 -566 -2225
rect -566 -2243 -562 -2239
rect -550 -2221 -546 -2217
rect -550 -2250 -546 -2246
rect -536 -2229 -532 -2225
rect -526 -2236 -522 -2232
rect -512 -2221 -508 -2217
rect -508 -2250 -504 -2246
rect -484 -2229 -480 -2225
rect -494 -2236 -490 -2232
rect -470 -2250 -466 -2246
rect -452 -2221 -448 -2217
rect -442 -2236 -438 -2232
rect -452 -2243 -448 -2239
rect -428 -2221 -424 -2217
rect -424 -2229 -420 -2225
rect -410 -2236 -406 -2232
rect -400 -2243 -396 -2239
rect -386 -2229 -382 -2225
rect -212 -2229 -208 -2225
rect -208 -2243 -204 -2239
rect -192 -2221 -188 -2217
rect -192 -2250 -188 -2246
rect -178 -2229 -174 -2225
rect -168 -2236 -164 -2232
rect -154 -2221 -150 -2217
rect -150 -2250 -146 -2246
rect -126 -2229 -122 -2225
rect -136 -2236 -132 -2232
rect -112 -2250 -108 -2246
rect -94 -2221 -90 -2217
rect -84 -2236 -80 -2232
rect -94 -2243 -90 -2239
rect -70 -2221 -66 -2217
rect -66 -2229 -62 -2225
rect -52 -2236 -48 -2232
rect -42 -2243 -38 -2239
rect -28 -2229 -24 -2225
rect 146 -2229 150 -2225
rect 150 -2243 154 -2239
rect 166 -2221 170 -2217
rect 166 -2250 170 -2246
rect 180 -2229 184 -2225
rect 190 -2236 194 -2232
rect 204 -2221 208 -2217
rect 208 -2250 212 -2246
rect 232 -2229 236 -2225
rect 222 -2236 226 -2232
rect 246 -2250 250 -2246
rect 264 -2221 268 -2217
rect 274 -2236 278 -2232
rect 264 -2243 268 -2239
rect 288 -2221 292 -2217
rect 292 -2229 296 -2225
rect 306 -2236 310 -2232
rect 316 -2243 320 -2239
rect 330 -2229 334 -2225
rect 502 -2229 506 -2225
rect 506 -2243 510 -2239
rect 522 -2221 526 -2217
rect 522 -2250 526 -2246
rect 536 -2229 540 -2225
rect 546 -2236 550 -2232
rect 560 -2221 564 -2217
rect 564 -2250 568 -2246
rect 588 -2229 592 -2225
rect 578 -2236 582 -2232
rect 602 -2250 606 -2246
rect 620 -2221 624 -2217
rect 630 -2236 634 -2232
rect 620 -2243 624 -2239
rect 644 -2221 648 -2217
rect 648 -2229 652 -2225
rect 662 -2236 666 -2232
rect 672 -2243 676 -2239
rect 686 -2229 690 -2225
rect -1552 -2400 -1548 -2396
rect -1548 -2414 -1544 -2410
rect -1532 -2392 -1528 -2388
rect -1532 -2421 -1528 -2417
rect -1518 -2400 -1514 -2396
rect -1508 -2407 -1504 -2403
rect -1494 -2392 -1490 -2388
rect -1490 -2421 -1486 -2417
rect -1466 -2400 -1462 -2396
rect -1476 -2407 -1472 -2403
rect -1452 -2421 -1448 -2417
rect -1434 -2392 -1430 -2388
rect -1424 -2407 -1420 -2403
rect -1434 -2414 -1430 -2410
rect -1410 -2392 -1406 -2388
rect -1406 -2400 -1402 -2396
rect -1392 -2407 -1388 -2403
rect -1382 -2414 -1378 -2410
rect -1368 -2400 -1364 -2396
rect -1227 -2400 -1223 -2396
rect -1223 -2414 -1219 -2410
rect -1207 -2392 -1203 -2388
rect -1207 -2421 -1203 -2417
rect -1193 -2400 -1189 -2396
rect -1183 -2407 -1179 -2403
rect -1169 -2392 -1165 -2388
rect -1165 -2421 -1161 -2417
rect -1141 -2400 -1137 -2396
rect -1151 -2407 -1147 -2403
rect -1127 -2421 -1123 -2417
rect -1109 -2392 -1105 -2388
rect -1099 -2407 -1095 -2403
rect -1109 -2414 -1105 -2410
rect -1085 -2392 -1081 -2388
rect -1081 -2400 -1077 -2396
rect -1067 -2407 -1063 -2403
rect -1057 -2414 -1053 -2410
rect -1043 -2400 -1039 -2396
rect -928 -2400 -924 -2396
rect -924 -2414 -920 -2410
rect -908 -2392 -904 -2388
rect -908 -2421 -904 -2417
rect -894 -2400 -890 -2396
rect -884 -2407 -880 -2403
rect -870 -2392 -866 -2388
rect -866 -2421 -862 -2417
rect -842 -2400 -838 -2396
rect -852 -2407 -848 -2403
rect -828 -2421 -824 -2417
rect -810 -2392 -806 -2388
rect -800 -2407 -796 -2403
rect -810 -2414 -806 -2410
rect -786 -2392 -782 -2388
rect -782 -2400 -778 -2396
rect -768 -2407 -764 -2403
rect -758 -2414 -754 -2410
rect -744 -2400 -740 -2396
rect -570 -2400 -566 -2396
rect -566 -2414 -562 -2410
rect -550 -2392 -546 -2388
rect -550 -2421 -546 -2417
rect -536 -2400 -532 -2396
rect -526 -2407 -522 -2403
rect -512 -2392 -508 -2388
rect -508 -2421 -504 -2417
rect -484 -2400 -480 -2396
rect -494 -2407 -490 -2403
rect -470 -2421 -466 -2417
rect -452 -2392 -448 -2388
rect -442 -2407 -438 -2403
rect -452 -2414 -448 -2410
rect -428 -2392 -424 -2388
rect -424 -2400 -420 -2396
rect -410 -2407 -406 -2403
rect -400 -2414 -396 -2410
rect -386 -2400 -382 -2396
rect -212 -2400 -208 -2396
rect -208 -2414 -204 -2410
rect -192 -2392 -188 -2388
rect -192 -2421 -188 -2417
rect -178 -2400 -174 -2396
rect -168 -2407 -164 -2403
rect -154 -2392 -150 -2388
rect -150 -2421 -146 -2417
rect -126 -2400 -122 -2396
rect -136 -2407 -132 -2403
rect -112 -2421 -108 -2417
rect -94 -2392 -90 -2388
rect -84 -2407 -80 -2403
rect -94 -2414 -90 -2410
rect -70 -2392 -66 -2388
rect -66 -2400 -62 -2396
rect -52 -2407 -48 -2403
rect -42 -2414 -38 -2410
rect -28 -2400 -24 -2396
rect 146 -2400 150 -2396
rect 150 -2414 154 -2410
rect 166 -2392 170 -2388
rect 166 -2421 170 -2417
rect 180 -2400 184 -2396
rect 190 -2407 194 -2403
rect 204 -2392 208 -2388
rect 208 -2421 212 -2417
rect 232 -2400 236 -2396
rect 222 -2407 226 -2403
rect 246 -2421 250 -2417
rect 264 -2392 268 -2388
rect 274 -2407 278 -2403
rect 264 -2414 268 -2410
rect 288 -2392 292 -2388
rect 292 -2400 296 -2396
rect 306 -2407 310 -2403
rect 316 -2414 320 -2410
rect 330 -2400 334 -2396
rect 502 -2400 506 -2396
rect 506 -2414 510 -2410
rect 522 -2392 526 -2388
rect 522 -2421 526 -2417
rect 536 -2400 540 -2396
rect 546 -2407 550 -2403
rect 560 -2392 564 -2388
rect 564 -2421 568 -2417
rect 588 -2400 592 -2396
rect 578 -2407 582 -2403
rect 602 -2421 606 -2417
rect 620 -2392 624 -2388
rect 630 -2407 634 -2403
rect 620 -2414 624 -2410
rect 644 -2392 648 -2388
rect 648 -2400 652 -2396
rect 662 -2407 666 -2403
rect 672 -2414 676 -2410
rect 686 -2400 690 -2396
rect 860 -2400 864 -2396
rect 864 -2414 868 -2410
rect 880 -2392 884 -2388
rect 880 -2421 884 -2417
rect 894 -2400 898 -2396
rect 904 -2407 908 -2403
rect 918 -2392 922 -2388
rect 922 -2421 926 -2417
rect 946 -2400 950 -2396
rect 936 -2407 940 -2403
rect 960 -2421 964 -2417
rect 978 -2392 982 -2388
rect 988 -2407 992 -2403
rect 978 -2414 982 -2410
rect 1002 -2392 1006 -2388
rect 1006 -2400 1010 -2396
rect 1020 -2407 1024 -2403
rect 1030 -2414 1034 -2410
rect 1044 -2400 1048 -2396
rect 1218 -2400 1222 -2396
rect 1222 -2414 1226 -2410
rect 1238 -2392 1242 -2388
rect 1238 -2421 1242 -2417
rect 1252 -2400 1256 -2396
rect 1262 -2407 1266 -2403
rect 1276 -2392 1280 -2388
rect 1280 -2421 1284 -2417
rect 1304 -2400 1308 -2396
rect 1294 -2407 1298 -2403
rect 1318 -2421 1322 -2417
rect 1336 -2392 1340 -2388
rect 1346 -2407 1350 -2403
rect 1336 -2414 1340 -2410
rect 1360 -2392 1364 -2388
rect 1364 -2400 1368 -2396
rect 1378 -2407 1382 -2403
rect 1388 -2414 1392 -2410
rect 1402 -2400 1406 -2396
rect -1552 -2571 -1548 -2567
rect -1548 -2585 -1544 -2581
rect -1532 -2563 -1528 -2559
rect -1532 -2592 -1528 -2588
rect -1518 -2571 -1514 -2567
rect -1508 -2578 -1504 -2574
rect -1494 -2563 -1490 -2559
rect -1490 -2592 -1486 -2588
rect -1466 -2571 -1462 -2567
rect -1476 -2578 -1472 -2574
rect -1452 -2592 -1448 -2588
rect -1434 -2563 -1430 -2559
rect -1424 -2578 -1420 -2574
rect -1434 -2585 -1430 -2581
rect -1410 -2563 -1406 -2559
rect -1406 -2571 -1402 -2567
rect -1392 -2578 -1388 -2574
rect -1382 -2585 -1378 -2581
rect -1368 -2571 -1364 -2567
rect -1227 -2571 -1223 -2567
rect -1223 -2585 -1219 -2581
rect -1207 -2563 -1203 -2559
rect -1207 -2592 -1203 -2588
rect -1193 -2571 -1189 -2567
rect -1183 -2578 -1179 -2574
rect -1169 -2563 -1165 -2559
rect -1165 -2592 -1161 -2588
rect -1141 -2571 -1137 -2567
rect -1151 -2578 -1147 -2574
rect -1127 -2592 -1123 -2588
rect -1109 -2563 -1105 -2559
rect -1099 -2578 -1095 -2574
rect -1109 -2585 -1105 -2581
rect -1085 -2563 -1081 -2559
rect -1081 -2571 -1077 -2567
rect -1067 -2578 -1063 -2574
rect -1057 -2585 -1053 -2581
rect -1043 -2571 -1039 -2567
rect -928 -2571 -924 -2567
rect -924 -2585 -920 -2581
rect -908 -2563 -904 -2559
rect -908 -2592 -904 -2588
rect -894 -2571 -890 -2567
rect -884 -2578 -880 -2574
rect -870 -2563 -866 -2559
rect -866 -2592 -862 -2588
rect -842 -2571 -838 -2567
rect -852 -2578 -848 -2574
rect -828 -2592 -824 -2588
rect -810 -2563 -806 -2559
rect -800 -2578 -796 -2574
rect -810 -2585 -806 -2581
rect -786 -2563 -782 -2559
rect -782 -2571 -778 -2567
rect -768 -2578 -764 -2574
rect -758 -2585 -754 -2581
rect -744 -2571 -740 -2567
rect -570 -2571 -566 -2567
rect -566 -2585 -562 -2581
rect -550 -2563 -546 -2559
rect -550 -2592 -546 -2588
rect -536 -2571 -532 -2567
rect -526 -2578 -522 -2574
rect -512 -2563 -508 -2559
rect -508 -2592 -504 -2588
rect -484 -2571 -480 -2567
rect -494 -2578 -490 -2574
rect -470 -2592 -466 -2588
rect -452 -2563 -448 -2559
rect -442 -2578 -438 -2574
rect -452 -2585 -448 -2581
rect -428 -2563 -424 -2559
rect -424 -2571 -420 -2567
rect -410 -2578 -406 -2574
rect -400 -2585 -396 -2581
rect -386 -2571 -382 -2567
rect -213 -2571 -209 -2567
rect -209 -2585 -205 -2581
rect -193 -2563 -189 -2559
rect -193 -2592 -189 -2588
rect -179 -2571 -175 -2567
rect -169 -2578 -165 -2574
rect -155 -2563 -151 -2559
rect -151 -2592 -147 -2588
rect -127 -2571 -123 -2567
rect -137 -2578 -133 -2574
rect -113 -2592 -109 -2588
rect -95 -2563 -91 -2559
rect -85 -2578 -81 -2574
rect -95 -2585 -91 -2581
rect -71 -2563 -67 -2559
rect -67 -2571 -63 -2567
rect -53 -2578 -49 -2574
rect -43 -2585 -39 -2581
rect -29 -2571 -25 -2567
rect 146 -2571 150 -2567
rect 150 -2585 154 -2581
rect 166 -2563 170 -2559
rect 166 -2592 170 -2588
rect 180 -2571 184 -2567
rect 190 -2578 194 -2574
rect 204 -2563 208 -2559
rect 208 -2592 212 -2588
rect 232 -2571 236 -2567
rect 222 -2578 226 -2574
rect 246 -2592 250 -2588
rect 264 -2563 268 -2559
rect 274 -2578 278 -2574
rect 264 -2585 268 -2581
rect 288 -2563 292 -2559
rect 292 -2571 296 -2567
rect 306 -2578 310 -2574
rect 316 -2585 320 -2581
rect 330 -2571 334 -2567
rect 502 -2571 506 -2567
rect 506 -2585 510 -2581
rect 522 -2563 526 -2559
rect 522 -2592 526 -2588
rect 536 -2571 540 -2567
rect 546 -2578 550 -2574
rect 560 -2563 564 -2559
rect 564 -2592 568 -2588
rect 588 -2571 592 -2567
rect 578 -2578 582 -2574
rect 602 -2592 606 -2588
rect 620 -2563 624 -2559
rect 630 -2578 634 -2574
rect 620 -2585 624 -2581
rect 644 -2563 648 -2559
rect 648 -2571 652 -2567
rect 662 -2578 666 -2574
rect 672 -2585 676 -2581
rect 686 -2571 690 -2567
rect 860 -2571 864 -2567
rect 864 -2585 868 -2581
rect 880 -2563 884 -2559
rect 880 -2592 884 -2588
rect 894 -2571 898 -2567
rect 904 -2578 908 -2574
rect 918 -2563 922 -2559
rect 922 -2592 926 -2588
rect 946 -2571 950 -2567
rect 936 -2578 940 -2574
rect 960 -2592 964 -2588
rect 978 -2563 982 -2559
rect 988 -2578 992 -2574
rect 978 -2585 982 -2581
rect 1002 -2563 1006 -2559
rect 1006 -2571 1010 -2567
rect 1020 -2578 1024 -2574
rect 1030 -2585 1034 -2581
rect 1044 -2571 1048 -2567
rect 1218 -2571 1222 -2567
rect 1222 -2585 1226 -2581
rect 1238 -2563 1242 -2559
rect 1238 -2592 1242 -2588
rect 1252 -2571 1256 -2567
rect 1262 -2578 1266 -2574
rect 1276 -2563 1280 -2559
rect 1280 -2592 1284 -2588
rect 1304 -2571 1308 -2567
rect 1294 -2578 1298 -2574
rect 1318 -2592 1322 -2588
rect 1336 -2563 1340 -2559
rect 1346 -2578 1350 -2574
rect 1336 -2585 1340 -2581
rect 1360 -2563 1364 -2559
rect 1364 -2571 1368 -2567
rect 1378 -2578 1382 -2574
rect 1388 -2585 1392 -2581
rect 1402 -2571 1406 -2567
rect -1308 -2652 -1304 -2648
rect -1297 -2660 -1293 -2656
rect -1290 -2682 -1286 -2678
rect -934 -2652 -930 -2648
rect -923 -2660 -919 -2656
rect -916 -2682 -912 -2678
rect -576 -2652 -572 -2648
rect -565 -2660 -561 -2656
rect -558 -2682 -554 -2678
rect -218 -2652 -214 -2648
rect -207 -2660 -203 -2656
rect -200 -2682 -196 -2678
rect 140 -2652 144 -2648
rect 151 -2660 155 -2656
rect 158 -2682 162 -2678
rect 496 -2652 500 -2648
rect 507 -2660 511 -2656
rect 514 -2682 518 -2678
rect 854 -2652 858 -2648
rect 865 -2660 869 -2656
rect 872 -2682 876 -2678
rect 1212 -2652 1216 -2648
rect 1223 -2660 1227 -2656
rect 1230 -2682 1234 -2678
rect -1223 -2835 -1219 -2831
rect -1227 -2842 -1223 -2838
rect -1207 -2822 -1203 -2818
rect -1197 -2842 -1193 -2838
rect -1183 -2835 -1179 -2831
rect -1173 -2828 -1169 -2824
rect -1163 -2835 -1159 -2831
rect -1149 -2842 -1145 -2838
rect -1145 -2856 -1141 -2852
rect -924 -2798 -920 -2794
rect -928 -2819 -924 -2815
rect -924 -2834 -920 -2830
rect -928 -2848 -924 -2844
rect -898 -2819 -894 -2815
rect -902 -2827 -898 -2823
rect -902 -2841 -898 -2837
rect -882 -2805 -878 -2801
rect -872 -2848 -868 -2844
rect -858 -2798 -854 -2794
rect -848 -2812 -844 -2808
rect -838 -2848 -834 -2844
rect -824 -2798 -820 -2794
rect -820 -2856 -816 -2852
rect -804 -2827 -800 -2823
rect -794 -2841 -790 -2837
rect -780 -2798 -776 -2794
rect -780 -2819 -776 -2815
rect -776 -2834 -772 -2830
rect -760 -2841 -756 -2837
rect -746 -2798 -742 -2794
rect -736 -2849 -732 -2845
rect -720 -2856 -716 -2852
rect -706 -2812 -702 -2808
rect -702 -2849 -698 -2845
rect -566 -2798 -562 -2794
rect -570 -2819 -566 -2815
rect -566 -2834 -562 -2830
rect -570 -2848 -566 -2844
rect -540 -2819 -536 -2815
rect -544 -2827 -540 -2823
rect -544 -2841 -540 -2837
rect -524 -2805 -520 -2801
rect -514 -2848 -510 -2844
rect -500 -2798 -496 -2794
rect -490 -2812 -486 -2808
rect -480 -2848 -476 -2844
rect -466 -2798 -462 -2794
rect -462 -2856 -458 -2852
rect -446 -2827 -442 -2823
rect -436 -2841 -432 -2837
rect -422 -2798 -418 -2794
rect -422 -2819 -418 -2815
rect -418 -2834 -414 -2830
rect -402 -2841 -398 -2837
rect -388 -2798 -384 -2794
rect -378 -2849 -374 -2845
rect -362 -2856 -358 -2852
rect -348 -2812 -344 -2808
rect -344 -2849 -340 -2845
rect -208 -2798 -204 -2794
rect -212 -2819 -208 -2815
rect -208 -2834 -204 -2830
rect -212 -2848 -208 -2844
rect -182 -2819 -178 -2815
rect -186 -2827 -182 -2823
rect -186 -2841 -182 -2837
rect -166 -2805 -162 -2801
rect -156 -2848 -152 -2844
rect -142 -2798 -138 -2794
rect -132 -2812 -128 -2808
rect -122 -2848 -118 -2844
rect -108 -2798 -104 -2794
rect -104 -2856 -100 -2852
rect -88 -2827 -84 -2823
rect -78 -2841 -74 -2837
rect -64 -2798 -60 -2794
rect -64 -2819 -60 -2815
rect -60 -2834 -56 -2830
rect -44 -2841 -40 -2837
rect -30 -2798 -26 -2794
rect -20 -2849 -16 -2845
rect -4 -2856 0 -2852
rect 10 -2812 14 -2808
rect 14 -2849 18 -2845
rect 150 -2798 154 -2794
rect 146 -2819 150 -2815
rect 150 -2834 154 -2830
rect 146 -2848 150 -2844
rect 176 -2819 180 -2815
rect 172 -2827 176 -2823
rect 172 -2841 176 -2837
rect 192 -2805 196 -2801
rect 202 -2848 206 -2844
rect 216 -2798 220 -2794
rect 226 -2812 230 -2808
rect 236 -2848 240 -2844
rect 250 -2798 254 -2794
rect 254 -2856 258 -2852
rect 270 -2827 274 -2823
rect 280 -2841 284 -2837
rect 294 -2798 298 -2794
rect 294 -2819 298 -2815
rect 298 -2834 302 -2830
rect 314 -2841 318 -2837
rect 328 -2798 332 -2794
rect 338 -2849 342 -2845
rect 354 -2856 358 -2852
rect 368 -2812 372 -2808
rect 372 -2849 376 -2845
rect 506 -2798 510 -2794
rect 502 -2819 506 -2815
rect 506 -2834 510 -2830
rect 502 -2848 506 -2844
rect 532 -2819 536 -2815
rect 528 -2827 532 -2823
rect 528 -2841 532 -2837
rect 548 -2805 552 -2801
rect 558 -2848 562 -2844
rect 572 -2798 576 -2794
rect 582 -2812 586 -2808
rect 592 -2848 596 -2844
rect 606 -2798 610 -2794
rect 610 -2856 614 -2852
rect 626 -2827 630 -2823
rect 636 -2841 640 -2837
rect 650 -2798 654 -2794
rect 650 -2819 654 -2815
rect 654 -2834 658 -2830
rect 670 -2841 674 -2837
rect 684 -2798 688 -2794
rect 694 -2849 698 -2845
rect 710 -2856 714 -2852
rect 724 -2812 728 -2808
rect 728 -2849 732 -2845
rect 864 -2798 868 -2794
rect 860 -2819 864 -2815
rect 864 -2834 868 -2830
rect 860 -2848 864 -2844
rect 890 -2819 894 -2815
rect 886 -2827 890 -2823
rect 886 -2841 890 -2837
rect 906 -2805 910 -2801
rect 916 -2848 920 -2844
rect 930 -2798 934 -2794
rect 940 -2812 944 -2808
rect 950 -2848 954 -2844
rect 964 -2798 968 -2794
rect 968 -2856 972 -2852
rect 984 -2827 988 -2823
rect 994 -2841 998 -2837
rect 1008 -2798 1012 -2794
rect 1008 -2819 1012 -2815
rect 1012 -2834 1016 -2830
rect 1028 -2841 1032 -2837
rect 1042 -2798 1046 -2794
rect 1052 -2849 1056 -2845
rect 1068 -2856 1072 -2852
rect 1082 -2812 1086 -2808
rect 1086 -2849 1090 -2845
rect 1222 -2798 1226 -2794
rect 1218 -2819 1222 -2815
rect 1222 -2834 1226 -2830
rect 1218 -2848 1222 -2844
rect 1248 -2819 1252 -2815
rect 1244 -2827 1248 -2823
rect 1244 -2841 1248 -2837
rect 1264 -2805 1268 -2801
rect 1274 -2848 1278 -2844
rect 1288 -2798 1292 -2794
rect 1298 -2812 1302 -2808
rect 1308 -2848 1312 -2844
rect 1322 -2798 1326 -2794
rect 1326 -2856 1330 -2852
rect 1342 -2827 1346 -2823
rect 1352 -2841 1356 -2837
rect 1366 -2798 1370 -2794
rect 1366 -2819 1370 -2815
rect 1370 -2834 1374 -2830
rect 1386 -2841 1390 -2837
rect 1400 -2798 1404 -2794
rect 1410 -2849 1414 -2845
rect 1426 -2856 1430 -2852
rect 1440 -2812 1444 -2808
rect 1444 -2849 1448 -2845
rect -1552 -2954 -1548 -2950
rect -1548 -2968 -1544 -2964
rect -1532 -2946 -1528 -2942
rect -1532 -2975 -1528 -2971
rect -1518 -2954 -1514 -2950
rect -1508 -2961 -1504 -2957
rect -1494 -2946 -1490 -2942
rect -1490 -2975 -1486 -2971
rect -1466 -2954 -1462 -2950
rect -1476 -2961 -1472 -2957
rect -1452 -2975 -1448 -2971
rect -1434 -2946 -1430 -2942
rect -1424 -2961 -1420 -2957
rect -1434 -2968 -1430 -2964
rect -1410 -2946 -1406 -2942
rect -1406 -2954 -1402 -2950
rect -1392 -2961 -1388 -2957
rect -1382 -2968 -1378 -2964
rect -1368 -2954 -1364 -2950
rect -1227 -2954 -1223 -2950
rect -1223 -2968 -1219 -2964
rect -1207 -2946 -1203 -2942
rect -1207 -2975 -1203 -2971
rect -1193 -2954 -1189 -2950
rect -1183 -2961 -1179 -2957
rect -1169 -2946 -1165 -2942
rect -1165 -2975 -1161 -2971
rect -1141 -2954 -1137 -2950
rect -1151 -2961 -1147 -2957
rect -1127 -2975 -1123 -2971
rect -1109 -2946 -1105 -2942
rect -1099 -2961 -1095 -2957
rect -1109 -2968 -1105 -2964
rect -1085 -2946 -1081 -2942
rect -1081 -2954 -1077 -2950
rect -1067 -2961 -1063 -2957
rect -1057 -2968 -1053 -2964
rect -1043 -2954 -1039 -2950
rect -928 -2954 -924 -2950
rect -924 -2968 -920 -2964
rect -908 -2946 -904 -2942
rect -908 -2975 -904 -2971
rect -894 -2954 -890 -2950
rect -884 -2961 -880 -2957
rect -870 -2946 -866 -2942
rect -866 -2975 -862 -2971
rect -842 -2954 -838 -2950
rect -852 -2961 -848 -2957
rect -828 -2975 -824 -2971
rect -810 -2946 -806 -2942
rect -800 -2961 -796 -2957
rect -810 -2968 -806 -2964
rect -786 -2946 -782 -2942
rect -782 -2954 -778 -2950
rect -768 -2961 -764 -2957
rect -758 -2968 -754 -2964
rect -744 -2954 -740 -2950
rect -570 -2954 -566 -2950
rect -566 -2968 -562 -2964
rect -550 -2946 -546 -2942
rect -550 -2975 -546 -2971
rect -536 -2954 -532 -2950
rect -526 -2961 -522 -2957
rect -512 -2946 -508 -2942
rect -508 -2975 -504 -2971
rect -484 -2954 -480 -2950
rect -494 -2961 -490 -2957
rect -470 -2975 -466 -2971
rect -452 -2946 -448 -2942
rect -442 -2961 -438 -2957
rect -452 -2968 -448 -2964
rect -428 -2946 -424 -2942
rect -424 -2954 -420 -2950
rect -410 -2961 -406 -2957
rect -400 -2968 -396 -2964
rect -386 -2954 -382 -2950
rect -212 -2954 -208 -2950
rect -208 -2968 -204 -2964
rect -192 -2946 -188 -2942
rect -192 -2975 -188 -2971
rect -178 -2954 -174 -2950
rect -168 -2961 -164 -2957
rect -154 -2946 -150 -2942
rect -150 -2975 -146 -2971
rect -126 -2954 -122 -2950
rect -136 -2961 -132 -2957
rect -112 -2975 -108 -2971
rect -94 -2946 -90 -2942
rect -84 -2961 -80 -2957
rect -94 -2968 -90 -2964
rect -70 -2946 -66 -2942
rect -66 -2954 -62 -2950
rect -52 -2961 -48 -2957
rect -42 -2968 -38 -2964
rect -28 -2954 -24 -2950
rect 146 -2954 150 -2950
rect 150 -2968 154 -2964
rect 166 -2946 170 -2942
rect 166 -2975 170 -2971
rect 180 -2954 184 -2950
rect 190 -2961 194 -2957
rect 204 -2946 208 -2942
rect 208 -2975 212 -2971
rect 232 -2954 236 -2950
rect 222 -2961 226 -2957
rect 246 -2975 250 -2971
rect 264 -2946 268 -2942
rect 274 -2961 278 -2957
rect 264 -2968 268 -2964
rect 288 -2946 292 -2942
rect 292 -2954 296 -2950
rect 306 -2961 310 -2957
rect 316 -2968 320 -2964
rect 330 -2954 334 -2950
rect -1552 -3125 -1548 -3121
rect -1548 -3139 -1544 -3135
rect -1532 -3117 -1528 -3113
rect -1532 -3146 -1528 -3142
rect -1518 -3125 -1514 -3121
rect -1508 -3132 -1504 -3128
rect -1494 -3117 -1490 -3113
rect -1490 -3146 -1486 -3142
rect -1466 -3125 -1462 -3121
rect -1476 -3132 -1472 -3128
rect -1452 -3146 -1448 -3142
rect -1434 -3117 -1430 -3113
rect -1424 -3132 -1420 -3128
rect -1434 -3139 -1430 -3135
rect -1410 -3117 -1406 -3113
rect -1406 -3125 -1402 -3121
rect -1392 -3132 -1388 -3128
rect -1382 -3139 -1378 -3135
rect -1368 -3125 -1364 -3121
rect -1227 -3125 -1223 -3121
rect -1223 -3139 -1219 -3135
rect -1207 -3117 -1203 -3113
rect -1207 -3146 -1203 -3142
rect -1193 -3125 -1189 -3121
rect -1183 -3132 -1179 -3128
rect -1169 -3117 -1165 -3113
rect -1165 -3146 -1161 -3142
rect -1141 -3125 -1137 -3121
rect -1151 -3132 -1147 -3128
rect -1127 -3146 -1123 -3142
rect -1109 -3117 -1105 -3113
rect -1099 -3132 -1095 -3128
rect -1109 -3139 -1105 -3135
rect -1085 -3117 -1081 -3113
rect -1081 -3125 -1077 -3121
rect -1067 -3132 -1063 -3128
rect -1057 -3139 -1053 -3135
rect -1043 -3125 -1039 -3121
rect -928 -3125 -924 -3121
rect -924 -3139 -920 -3135
rect -908 -3117 -904 -3113
rect -908 -3146 -904 -3142
rect -894 -3125 -890 -3121
rect -884 -3132 -880 -3128
rect -870 -3117 -866 -3113
rect -866 -3146 -862 -3142
rect -842 -3125 -838 -3121
rect -852 -3132 -848 -3128
rect -828 -3146 -824 -3142
rect -810 -3117 -806 -3113
rect -800 -3132 -796 -3128
rect -810 -3139 -806 -3135
rect -786 -3117 -782 -3113
rect -782 -3125 -778 -3121
rect -768 -3132 -764 -3128
rect -758 -3139 -754 -3135
rect -744 -3125 -740 -3121
rect -570 -3125 -566 -3121
rect -566 -3139 -562 -3135
rect -550 -3117 -546 -3113
rect -550 -3146 -546 -3142
rect -536 -3125 -532 -3121
rect -526 -3132 -522 -3128
rect -512 -3117 -508 -3113
rect -508 -3146 -504 -3142
rect -484 -3125 -480 -3121
rect -494 -3132 -490 -3128
rect -470 -3146 -466 -3142
rect -452 -3117 -448 -3113
rect -442 -3132 -438 -3128
rect -452 -3139 -448 -3135
rect -428 -3117 -424 -3113
rect -424 -3125 -420 -3121
rect -410 -3132 -406 -3128
rect -400 -3139 -396 -3135
rect -386 -3125 -382 -3121
rect -212 -3125 -208 -3121
rect -208 -3139 -204 -3135
rect -192 -3117 -188 -3113
rect -192 -3146 -188 -3142
rect -178 -3125 -174 -3121
rect -168 -3132 -164 -3128
rect -154 -3117 -150 -3113
rect -150 -3146 -146 -3142
rect -126 -3125 -122 -3121
rect -136 -3132 -132 -3128
rect -112 -3146 -108 -3142
rect -94 -3117 -90 -3113
rect -84 -3132 -80 -3128
rect -94 -3139 -90 -3135
rect -70 -3117 -66 -3113
rect -66 -3125 -62 -3121
rect -52 -3132 -48 -3128
rect -42 -3139 -38 -3135
rect -28 -3125 -24 -3121
rect 146 -3125 150 -3121
rect 150 -3139 154 -3135
rect 166 -3117 170 -3113
rect 166 -3146 170 -3142
rect 180 -3125 184 -3121
rect 190 -3132 194 -3128
rect 204 -3117 208 -3113
rect 208 -3146 212 -3142
rect 232 -3125 236 -3121
rect 222 -3132 226 -3128
rect 246 -3146 250 -3142
rect 264 -3117 268 -3113
rect 274 -3132 278 -3128
rect 264 -3139 268 -3135
rect 288 -3117 292 -3113
rect 292 -3125 296 -3121
rect 306 -3132 310 -3128
rect 316 -3139 320 -3135
rect 330 -3125 334 -3121
rect 502 -3125 506 -3121
rect 506 -3139 510 -3135
rect 522 -3117 526 -3113
rect 522 -3146 526 -3142
rect 536 -3125 540 -3121
rect 546 -3132 550 -3128
rect 560 -3117 564 -3113
rect 564 -3146 568 -3142
rect 588 -3125 592 -3121
rect 578 -3132 582 -3128
rect 602 -3146 606 -3142
rect 620 -3117 624 -3113
rect 630 -3132 634 -3128
rect 620 -3139 624 -3135
rect 644 -3117 648 -3113
rect 648 -3125 652 -3121
rect 662 -3132 666 -3128
rect 672 -3139 676 -3135
rect 686 -3125 690 -3121
rect 860 -3125 864 -3121
rect 864 -3139 868 -3135
rect 880 -3117 884 -3113
rect 880 -3146 884 -3142
rect 894 -3125 898 -3121
rect 904 -3132 908 -3128
rect 918 -3117 922 -3113
rect 922 -3146 926 -3142
rect 946 -3125 950 -3121
rect 936 -3132 940 -3128
rect 960 -3146 964 -3142
rect 978 -3117 982 -3113
rect 988 -3132 992 -3128
rect 978 -3139 982 -3135
rect 1002 -3117 1006 -3113
rect 1006 -3125 1010 -3121
rect 1020 -3132 1024 -3128
rect 1030 -3139 1034 -3135
rect 1044 -3125 1048 -3121
rect 1218 -3125 1222 -3121
rect 1222 -3139 1226 -3135
rect 1238 -3117 1242 -3113
rect 1238 -3146 1242 -3142
rect 1252 -3125 1256 -3121
rect 1262 -3132 1266 -3128
rect 1276 -3117 1280 -3113
rect 1280 -3146 1284 -3142
rect 1304 -3125 1308 -3121
rect 1294 -3132 1298 -3128
rect 1318 -3146 1322 -3142
rect 1336 -3117 1340 -3113
rect 1346 -3132 1350 -3128
rect 1336 -3139 1340 -3135
rect 1360 -3117 1364 -3113
rect 1364 -3125 1368 -3121
rect 1378 -3132 1382 -3128
rect 1388 -3139 1392 -3135
rect 1402 -3125 1406 -3121
rect -1552 -3296 -1548 -3292
rect -1548 -3310 -1544 -3306
rect -1532 -3288 -1528 -3284
rect -1532 -3317 -1528 -3313
rect -1518 -3296 -1514 -3292
rect -1508 -3303 -1504 -3299
rect -1494 -3288 -1490 -3284
rect -1490 -3317 -1486 -3313
rect -1466 -3296 -1462 -3292
rect -1476 -3303 -1472 -3299
rect -1452 -3317 -1448 -3313
rect -1434 -3288 -1430 -3284
rect -1424 -3303 -1420 -3299
rect -1434 -3310 -1430 -3306
rect -1410 -3288 -1406 -3284
rect -1406 -3296 -1402 -3292
rect -1392 -3303 -1388 -3299
rect -1382 -3310 -1378 -3306
rect -1368 -3296 -1364 -3292
rect -1227 -3296 -1223 -3292
rect -1223 -3310 -1219 -3306
rect -1207 -3288 -1203 -3284
rect -1207 -3317 -1203 -3313
rect -1193 -3296 -1189 -3292
rect -1183 -3303 -1179 -3299
rect -1169 -3288 -1165 -3284
rect -1165 -3317 -1161 -3313
rect -1141 -3296 -1137 -3292
rect -1151 -3303 -1147 -3299
rect -1127 -3317 -1123 -3313
rect -1109 -3288 -1105 -3284
rect -1099 -3303 -1095 -3299
rect -1109 -3310 -1105 -3306
rect -1085 -3288 -1081 -3284
rect -1081 -3296 -1077 -3292
rect -1067 -3303 -1063 -3299
rect -1057 -3310 -1053 -3306
rect -1043 -3296 -1039 -3292
rect -928 -3296 -924 -3292
rect -924 -3310 -920 -3306
rect -908 -3288 -904 -3284
rect -908 -3317 -904 -3313
rect -894 -3296 -890 -3292
rect -884 -3303 -880 -3299
rect -870 -3288 -866 -3284
rect -866 -3317 -862 -3313
rect -842 -3296 -838 -3292
rect -852 -3303 -848 -3299
rect -828 -3317 -824 -3313
rect -810 -3288 -806 -3284
rect -800 -3303 -796 -3299
rect -810 -3310 -806 -3306
rect -786 -3288 -782 -3284
rect -782 -3296 -778 -3292
rect -768 -3303 -764 -3299
rect -758 -3310 -754 -3306
rect -744 -3296 -740 -3292
rect -570 -3296 -566 -3292
rect -566 -3310 -562 -3306
rect -550 -3288 -546 -3284
rect -550 -3317 -546 -3313
rect -536 -3296 -532 -3292
rect -526 -3303 -522 -3299
rect -512 -3288 -508 -3284
rect -508 -3317 -504 -3313
rect -484 -3296 -480 -3292
rect -494 -3303 -490 -3299
rect -470 -3317 -466 -3313
rect -452 -3288 -448 -3284
rect -442 -3303 -438 -3299
rect -452 -3310 -448 -3306
rect -428 -3288 -424 -3284
rect -424 -3296 -420 -3292
rect -410 -3303 -406 -3299
rect -400 -3310 -396 -3306
rect -386 -3296 -382 -3292
rect -212 -3296 -208 -3292
rect -208 -3310 -204 -3306
rect -192 -3288 -188 -3284
rect -192 -3317 -188 -3313
rect -178 -3296 -174 -3292
rect -168 -3303 -164 -3299
rect -154 -3288 -150 -3284
rect -150 -3317 -146 -3313
rect -126 -3296 -122 -3292
rect -136 -3303 -132 -3299
rect -112 -3317 -108 -3313
rect -94 -3288 -90 -3284
rect -84 -3303 -80 -3299
rect -94 -3310 -90 -3306
rect -70 -3288 -66 -3284
rect -66 -3296 -62 -3292
rect -52 -3303 -48 -3299
rect -42 -3310 -38 -3306
rect -28 -3296 -24 -3292
rect 146 -3296 150 -3292
rect 150 -3310 154 -3306
rect 166 -3288 170 -3284
rect 166 -3317 170 -3313
rect 180 -3296 184 -3292
rect 190 -3303 194 -3299
rect 204 -3288 208 -3284
rect 208 -3317 212 -3313
rect 232 -3296 236 -3292
rect 222 -3303 226 -3299
rect 246 -3317 250 -3313
rect 264 -3288 268 -3284
rect 274 -3303 278 -3299
rect 264 -3310 268 -3306
rect 288 -3288 292 -3284
rect 292 -3296 296 -3292
rect 306 -3303 310 -3299
rect 316 -3310 320 -3306
rect 330 -3296 334 -3292
rect 502 -3296 506 -3292
rect 506 -3310 510 -3306
rect 522 -3288 526 -3284
rect 522 -3317 526 -3313
rect 536 -3296 540 -3292
rect 546 -3303 550 -3299
rect 560 -3288 564 -3284
rect 564 -3317 568 -3313
rect 588 -3296 592 -3292
rect 578 -3303 582 -3299
rect 602 -3317 606 -3313
rect 620 -3288 624 -3284
rect 630 -3303 634 -3299
rect 620 -3310 624 -3306
rect 644 -3288 648 -3284
rect 648 -3296 652 -3292
rect 662 -3303 666 -3299
rect 672 -3310 676 -3306
rect 686 -3296 690 -3292
rect 860 -3296 864 -3292
rect 864 -3310 868 -3306
rect 880 -3288 884 -3284
rect 880 -3317 884 -3313
rect 894 -3296 898 -3292
rect 904 -3303 908 -3299
rect 918 -3288 922 -3284
rect 922 -3317 926 -3313
rect 946 -3296 950 -3292
rect 936 -3303 940 -3299
rect 960 -3317 964 -3313
rect 978 -3288 982 -3284
rect 988 -3303 992 -3299
rect 978 -3310 982 -3306
rect 1002 -3288 1006 -3284
rect 1006 -3296 1010 -3292
rect 1020 -3303 1024 -3299
rect 1030 -3310 1034 -3306
rect 1044 -3296 1048 -3292
rect 1218 -3296 1222 -3292
rect 1222 -3310 1226 -3306
rect 1238 -3288 1242 -3284
rect 1238 -3317 1242 -3313
rect 1252 -3296 1256 -3292
rect 1262 -3303 1266 -3299
rect 1276 -3288 1280 -3284
rect 1280 -3317 1284 -3313
rect 1304 -3296 1308 -3292
rect 1294 -3303 1298 -3299
rect 1318 -3317 1322 -3313
rect 1336 -3288 1340 -3284
rect 1346 -3303 1350 -3299
rect 1336 -3310 1340 -3306
rect 1360 -3288 1364 -3284
rect 1364 -3296 1368 -3292
rect 1378 -3303 1382 -3299
rect 1388 -3310 1392 -3306
rect 1402 -3296 1406 -3292
rect -1308 -3383 -1304 -3379
rect -1297 -3391 -1293 -3387
rect -1290 -3413 -1286 -3409
rect -934 -3383 -930 -3379
rect -923 -3391 -919 -3387
rect -916 -3413 -912 -3409
rect -576 -3383 -572 -3379
rect -565 -3391 -561 -3387
rect -558 -3413 -554 -3409
rect -218 -3383 -214 -3379
rect -207 -3391 -203 -3387
rect -200 -3413 -196 -3409
rect 140 -3383 144 -3379
rect 151 -3391 155 -3387
rect 158 -3413 162 -3409
rect 496 -3383 500 -3379
rect 507 -3391 511 -3387
rect 514 -3413 518 -3409
rect 854 -3383 858 -3379
rect 865 -3391 869 -3387
rect 872 -3413 876 -3409
rect 1212 -3383 1216 -3379
rect 1223 -3391 1227 -3387
rect 1230 -3413 1234 -3409
rect -1223 -3566 -1219 -3562
rect -1227 -3573 -1223 -3569
rect -1207 -3553 -1203 -3549
rect -1197 -3573 -1193 -3569
rect -1183 -3566 -1179 -3562
rect -1173 -3559 -1169 -3555
rect -1163 -3566 -1159 -3562
rect -1149 -3573 -1145 -3569
rect -1145 -3587 -1141 -3583
rect -924 -3529 -920 -3525
rect -928 -3550 -924 -3546
rect -924 -3565 -920 -3561
rect -928 -3579 -924 -3575
rect -898 -3550 -894 -3546
rect -902 -3558 -898 -3554
rect -902 -3572 -898 -3568
rect -882 -3536 -878 -3532
rect -872 -3579 -868 -3575
rect -858 -3529 -854 -3525
rect -848 -3543 -844 -3539
rect -838 -3579 -834 -3575
rect -824 -3529 -820 -3525
rect -820 -3587 -816 -3583
rect -804 -3558 -800 -3554
rect -794 -3572 -790 -3568
rect -780 -3529 -776 -3525
rect -780 -3550 -776 -3546
rect -776 -3565 -772 -3561
rect -760 -3572 -756 -3568
rect -746 -3529 -742 -3525
rect -736 -3580 -732 -3576
rect -720 -3587 -716 -3583
rect -706 -3543 -702 -3539
rect -702 -3580 -698 -3576
rect -566 -3529 -562 -3525
rect -570 -3550 -566 -3546
rect -566 -3565 -562 -3561
rect -570 -3579 -566 -3575
rect -540 -3550 -536 -3546
rect -544 -3558 -540 -3554
rect -544 -3572 -540 -3568
rect -524 -3536 -520 -3532
rect -514 -3579 -510 -3575
rect -500 -3529 -496 -3525
rect -490 -3543 -486 -3539
rect -480 -3579 -476 -3575
rect -466 -3529 -462 -3525
rect -462 -3587 -458 -3583
rect -446 -3558 -442 -3554
rect -436 -3572 -432 -3568
rect -422 -3529 -418 -3525
rect -422 -3550 -418 -3546
rect -418 -3565 -414 -3561
rect -402 -3572 -398 -3568
rect -388 -3529 -384 -3525
rect -378 -3580 -374 -3576
rect -362 -3587 -358 -3583
rect -348 -3543 -344 -3539
rect -344 -3580 -340 -3576
rect -208 -3529 -204 -3525
rect -212 -3550 -208 -3546
rect -208 -3565 -204 -3561
rect -212 -3579 -208 -3575
rect -182 -3550 -178 -3546
rect -186 -3558 -182 -3554
rect -186 -3572 -182 -3568
rect -166 -3536 -162 -3532
rect -156 -3579 -152 -3575
rect -142 -3529 -138 -3525
rect -132 -3543 -128 -3539
rect -122 -3579 -118 -3575
rect -108 -3529 -104 -3525
rect -104 -3587 -100 -3583
rect -88 -3558 -84 -3554
rect -78 -3572 -74 -3568
rect -64 -3529 -60 -3525
rect -64 -3550 -60 -3546
rect -60 -3565 -56 -3561
rect -44 -3572 -40 -3568
rect -30 -3529 -26 -3525
rect -20 -3580 -16 -3576
rect -4 -3587 0 -3583
rect 10 -3543 14 -3539
rect 14 -3580 18 -3576
rect 150 -3529 154 -3525
rect 146 -3550 150 -3546
rect 150 -3565 154 -3561
rect 146 -3579 150 -3575
rect 176 -3550 180 -3546
rect 172 -3558 176 -3554
rect 172 -3572 176 -3568
rect 192 -3536 196 -3532
rect 202 -3579 206 -3575
rect 216 -3529 220 -3525
rect 226 -3543 230 -3539
rect 236 -3579 240 -3575
rect 250 -3529 254 -3525
rect 254 -3587 258 -3583
rect 270 -3558 274 -3554
rect 280 -3572 284 -3568
rect 294 -3529 298 -3525
rect 294 -3550 298 -3546
rect 298 -3565 302 -3561
rect 314 -3572 318 -3568
rect 328 -3529 332 -3525
rect 338 -3580 342 -3576
rect 354 -3587 358 -3583
rect 368 -3543 372 -3539
rect 372 -3580 376 -3576
rect 506 -3529 510 -3525
rect 502 -3550 506 -3546
rect 506 -3565 510 -3561
rect 502 -3579 506 -3575
rect 532 -3550 536 -3546
rect 528 -3558 532 -3554
rect 528 -3572 532 -3568
rect 548 -3536 552 -3532
rect 558 -3579 562 -3575
rect 572 -3529 576 -3525
rect 582 -3543 586 -3539
rect 592 -3579 596 -3575
rect 606 -3529 610 -3525
rect 610 -3587 614 -3583
rect 626 -3558 630 -3554
rect 636 -3572 640 -3568
rect 650 -3529 654 -3525
rect 650 -3550 654 -3546
rect 654 -3565 658 -3561
rect 670 -3572 674 -3568
rect 684 -3529 688 -3525
rect 694 -3580 698 -3576
rect 710 -3587 714 -3583
rect 724 -3543 728 -3539
rect 728 -3580 732 -3576
rect 864 -3529 868 -3525
rect 860 -3550 864 -3546
rect 864 -3565 868 -3561
rect 860 -3579 864 -3575
rect 890 -3550 894 -3546
rect 886 -3558 890 -3554
rect 886 -3572 890 -3568
rect 906 -3536 910 -3532
rect 916 -3579 920 -3575
rect 930 -3529 934 -3525
rect 940 -3543 944 -3539
rect 950 -3579 954 -3575
rect 964 -3529 968 -3525
rect 968 -3587 972 -3583
rect 984 -3558 988 -3554
rect 994 -3572 998 -3568
rect 1008 -3529 1012 -3525
rect 1008 -3550 1012 -3546
rect 1012 -3565 1016 -3561
rect 1028 -3572 1032 -3568
rect 1042 -3529 1046 -3525
rect 1052 -3580 1056 -3576
rect 1068 -3587 1072 -3583
rect 1082 -3543 1086 -3539
rect 1086 -3580 1090 -3576
rect 1222 -3529 1226 -3525
rect 1218 -3550 1222 -3546
rect 1222 -3565 1226 -3561
rect 1218 -3579 1222 -3575
rect 1248 -3550 1252 -3546
rect 1244 -3558 1248 -3554
rect 1244 -3572 1248 -3568
rect 1264 -3536 1268 -3532
rect 1274 -3579 1278 -3575
rect 1288 -3529 1292 -3525
rect 1298 -3543 1302 -3539
rect 1308 -3579 1312 -3575
rect 1322 -3529 1326 -3525
rect 1326 -3587 1330 -3583
rect 1342 -3558 1346 -3554
rect 1352 -3572 1356 -3568
rect 1366 -3529 1370 -3525
rect 1366 -3550 1370 -3546
rect 1370 -3565 1374 -3561
rect 1386 -3572 1390 -3568
rect 1400 -3529 1404 -3525
rect 1410 -3580 1414 -3576
rect 1426 -3587 1430 -3583
rect 1440 -3543 1444 -3539
rect 1444 -3580 1448 -3576
rect -1815 -3696 -1811 -3692
rect -1811 -3710 -1807 -3706
rect -1795 -3688 -1791 -3684
rect -1795 -3717 -1791 -3713
rect -1781 -3696 -1777 -3692
rect -1771 -3703 -1767 -3699
rect -1757 -3688 -1753 -3684
rect -1753 -3717 -1749 -3713
rect -1729 -3696 -1725 -3692
rect -1739 -3703 -1735 -3699
rect -1715 -3717 -1711 -3713
rect -1697 -3688 -1693 -3684
rect -1687 -3703 -1683 -3699
rect -1697 -3710 -1693 -3706
rect -1673 -3688 -1669 -3684
rect -1669 -3696 -1665 -3692
rect -1655 -3703 -1651 -3699
rect -1645 -3710 -1641 -3706
rect -1631 -3696 -1627 -3692
rect -1552 -3696 -1548 -3692
rect -1548 -3710 -1544 -3706
rect -1532 -3688 -1528 -3684
rect -1532 -3717 -1528 -3713
rect -1518 -3696 -1514 -3692
rect -1508 -3703 -1504 -3699
rect -1494 -3688 -1490 -3684
rect -1490 -3717 -1486 -3713
rect -1466 -3696 -1462 -3692
rect -1476 -3703 -1472 -3699
rect -1452 -3717 -1448 -3713
rect -1434 -3688 -1430 -3684
rect -1424 -3703 -1420 -3699
rect -1434 -3710 -1430 -3706
rect -1410 -3688 -1406 -3684
rect -1406 -3696 -1402 -3692
rect -1392 -3703 -1388 -3699
rect -1382 -3710 -1378 -3706
rect -1368 -3696 -1364 -3692
rect -1227 -3696 -1223 -3692
rect -1223 -3710 -1219 -3706
rect -1207 -3688 -1203 -3684
rect -1207 -3717 -1203 -3713
rect -1193 -3696 -1189 -3692
rect -1183 -3703 -1179 -3699
rect -1169 -3688 -1165 -3684
rect -1165 -3717 -1161 -3713
rect -1141 -3696 -1137 -3692
rect -1151 -3703 -1147 -3699
rect -1127 -3717 -1123 -3713
rect -1109 -3688 -1105 -3684
rect -1099 -3703 -1095 -3699
rect -1109 -3710 -1105 -3706
rect -1085 -3688 -1081 -3684
rect -1081 -3696 -1077 -3692
rect -1067 -3703 -1063 -3699
rect -1057 -3710 -1053 -3706
rect -1043 -3696 -1039 -3692
rect -927 -3696 -923 -3692
rect -923 -3710 -919 -3706
rect -907 -3688 -903 -3684
rect -907 -3717 -903 -3713
rect -893 -3696 -889 -3692
rect -883 -3703 -879 -3699
rect -869 -3688 -865 -3684
rect -865 -3717 -861 -3713
rect -841 -3696 -837 -3692
rect -851 -3703 -847 -3699
rect -827 -3717 -823 -3713
rect -809 -3688 -805 -3684
rect -799 -3703 -795 -3699
rect -809 -3710 -805 -3706
rect -785 -3688 -781 -3684
rect -781 -3696 -777 -3692
rect -767 -3703 -763 -3699
rect -757 -3710 -753 -3706
rect -743 -3696 -739 -3692
rect -570 -3696 -566 -3692
rect -566 -3710 -562 -3706
rect -550 -3688 -546 -3684
rect -550 -3717 -546 -3713
rect -536 -3696 -532 -3692
rect -526 -3703 -522 -3699
rect -512 -3688 -508 -3684
rect -508 -3717 -504 -3713
rect -484 -3696 -480 -3692
rect -494 -3703 -490 -3699
rect -470 -3717 -466 -3713
rect -452 -3688 -448 -3684
rect -442 -3703 -438 -3699
rect -452 -3710 -448 -3706
rect -428 -3688 -424 -3684
rect -424 -3696 -420 -3692
rect -410 -3703 -406 -3699
rect -400 -3710 -396 -3706
rect -386 -3696 -382 -3692
rect -212 -3696 -208 -3692
rect -208 -3710 -204 -3706
rect -192 -3688 -188 -3684
rect -192 -3717 -188 -3713
rect -178 -3696 -174 -3692
rect -168 -3703 -164 -3699
rect -154 -3688 -150 -3684
rect -150 -3717 -146 -3713
rect -126 -3696 -122 -3692
rect -136 -3703 -132 -3699
rect -112 -3717 -108 -3713
rect -94 -3688 -90 -3684
rect -84 -3703 -80 -3699
rect -94 -3710 -90 -3706
rect -70 -3688 -66 -3684
rect -66 -3696 -62 -3692
rect -52 -3703 -48 -3699
rect -42 -3710 -38 -3706
rect -28 -3696 -24 -3692
rect -1552 -3867 -1548 -3863
rect -1548 -3881 -1544 -3877
rect -1532 -3859 -1528 -3855
rect -1532 -3888 -1528 -3884
rect -1518 -3867 -1514 -3863
rect -1508 -3874 -1504 -3870
rect -1494 -3859 -1490 -3855
rect -1490 -3888 -1486 -3884
rect -1466 -3867 -1462 -3863
rect -1476 -3874 -1472 -3870
rect -1452 -3888 -1448 -3884
rect -1434 -3859 -1430 -3855
rect -1424 -3874 -1420 -3870
rect -1434 -3881 -1430 -3877
rect -1410 -3859 -1406 -3855
rect -1406 -3867 -1402 -3863
rect -1392 -3874 -1388 -3870
rect -1382 -3881 -1378 -3877
rect -1368 -3867 -1364 -3863
rect -1227 -3867 -1223 -3863
rect -1223 -3881 -1219 -3877
rect -1207 -3859 -1203 -3855
rect -1207 -3888 -1203 -3884
rect -1193 -3867 -1189 -3863
rect -1183 -3874 -1179 -3870
rect -1169 -3859 -1165 -3855
rect -1165 -3888 -1161 -3884
rect -1141 -3867 -1137 -3863
rect -1151 -3874 -1147 -3870
rect -1127 -3888 -1123 -3884
rect -1109 -3859 -1105 -3855
rect -1099 -3874 -1095 -3870
rect -1109 -3881 -1105 -3877
rect -1085 -3859 -1081 -3855
rect -1081 -3867 -1077 -3863
rect -1067 -3874 -1063 -3870
rect -1057 -3881 -1053 -3877
rect -1043 -3867 -1039 -3863
rect -927 -3867 -923 -3863
rect -923 -3881 -919 -3877
rect -907 -3859 -903 -3855
rect -907 -3888 -903 -3884
rect -893 -3867 -889 -3863
rect -883 -3874 -879 -3870
rect -869 -3859 -865 -3855
rect -865 -3888 -861 -3884
rect -841 -3867 -837 -3863
rect -851 -3874 -847 -3870
rect -827 -3888 -823 -3884
rect -809 -3859 -805 -3855
rect -799 -3874 -795 -3870
rect -809 -3881 -805 -3877
rect -785 -3859 -781 -3855
rect -781 -3867 -777 -3863
rect -767 -3874 -763 -3870
rect -757 -3881 -753 -3877
rect -743 -3867 -739 -3863
rect -570 -3867 -566 -3863
rect -566 -3881 -562 -3877
rect -550 -3859 -546 -3855
rect -550 -3888 -546 -3884
rect -536 -3867 -532 -3863
rect -526 -3874 -522 -3870
rect -512 -3859 -508 -3855
rect -508 -3888 -504 -3884
rect -484 -3867 -480 -3863
rect -494 -3874 -490 -3870
rect -470 -3888 -466 -3884
rect -452 -3859 -448 -3855
rect -442 -3874 -438 -3870
rect -452 -3881 -448 -3877
rect -428 -3859 -424 -3855
rect -424 -3867 -420 -3863
rect -410 -3874 -406 -3870
rect -400 -3881 -396 -3877
rect -386 -3867 -382 -3863
rect -212 -3867 -208 -3863
rect -208 -3881 -204 -3877
rect -192 -3859 -188 -3855
rect -192 -3888 -188 -3884
rect -178 -3867 -174 -3863
rect -168 -3874 -164 -3870
rect -154 -3859 -150 -3855
rect -150 -3888 -146 -3884
rect -126 -3867 -122 -3863
rect -136 -3874 -132 -3870
rect -112 -3888 -108 -3884
rect -94 -3859 -90 -3855
rect -84 -3874 -80 -3870
rect -94 -3881 -90 -3877
rect -70 -3859 -66 -3855
rect -66 -3867 -62 -3863
rect -52 -3874 -48 -3870
rect -42 -3881 -38 -3877
rect -28 -3867 -24 -3863
rect 146 -3867 150 -3863
rect 150 -3881 154 -3877
rect 166 -3859 170 -3855
rect 166 -3888 170 -3884
rect 180 -3867 184 -3863
rect 190 -3874 194 -3870
rect 204 -3859 208 -3855
rect 208 -3888 212 -3884
rect 232 -3867 236 -3863
rect 222 -3874 226 -3870
rect 246 -3888 250 -3884
rect 264 -3859 268 -3855
rect 274 -3874 278 -3870
rect 264 -3881 268 -3877
rect 288 -3859 292 -3855
rect 292 -3867 296 -3863
rect 306 -3874 310 -3870
rect 316 -3881 320 -3877
rect 330 -3867 334 -3863
rect 502 -3867 506 -3863
rect 506 -3881 510 -3877
rect 522 -3859 526 -3855
rect 522 -3888 526 -3884
rect 536 -3867 540 -3863
rect 546 -3874 550 -3870
rect 560 -3859 564 -3855
rect 564 -3888 568 -3884
rect 588 -3867 592 -3863
rect 578 -3874 582 -3870
rect 602 -3888 606 -3884
rect 620 -3859 624 -3855
rect 630 -3874 634 -3870
rect 620 -3881 624 -3877
rect 644 -3859 648 -3855
rect 648 -3867 652 -3863
rect 662 -3874 666 -3870
rect 672 -3881 676 -3877
rect 686 -3867 690 -3863
rect 860 -3867 864 -3863
rect 864 -3881 868 -3877
rect 880 -3859 884 -3855
rect 880 -3888 884 -3884
rect 894 -3867 898 -3863
rect 904 -3874 908 -3870
rect 918 -3859 922 -3855
rect 922 -3888 926 -3884
rect 946 -3867 950 -3863
rect 936 -3874 940 -3870
rect 960 -3888 964 -3884
rect 978 -3859 982 -3855
rect 988 -3874 992 -3870
rect 978 -3881 982 -3877
rect 1002 -3859 1006 -3855
rect 1006 -3867 1010 -3863
rect 1020 -3874 1024 -3870
rect 1030 -3881 1034 -3877
rect 1044 -3867 1048 -3863
rect 1218 -3867 1222 -3863
rect 1222 -3881 1226 -3877
rect 1238 -3859 1242 -3855
rect 1238 -3888 1242 -3884
rect 1252 -3867 1256 -3863
rect 1262 -3874 1266 -3870
rect 1276 -3859 1280 -3855
rect 1280 -3888 1284 -3884
rect 1304 -3867 1308 -3863
rect 1294 -3874 1298 -3870
rect 1318 -3888 1322 -3884
rect 1336 -3859 1340 -3855
rect 1346 -3874 1350 -3870
rect 1336 -3881 1340 -3877
rect 1360 -3859 1364 -3855
rect 1364 -3867 1368 -3863
rect 1378 -3874 1382 -3870
rect 1388 -3881 1392 -3877
rect 1402 -3867 1406 -3863
rect -1552 -4042 -1548 -4038
rect -1548 -4056 -1544 -4052
rect -1532 -4034 -1528 -4030
rect -1532 -4063 -1528 -4059
rect -1518 -4042 -1514 -4038
rect -1508 -4049 -1504 -4045
rect -1494 -4034 -1490 -4030
rect -1490 -4063 -1486 -4059
rect -1466 -4042 -1462 -4038
rect -1476 -4049 -1472 -4045
rect -1452 -4063 -1448 -4059
rect -1434 -4034 -1430 -4030
rect -1424 -4049 -1420 -4045
rect -1434 -4056 -1430 -4052
rect -1410 -4034 -1406 -4030
rect -1406 -4042 -1402 -4038
rect -1392 -4049 -1388 -4045
rect -1382 -4056 -1378 -4052
rect -1368 -4042 -1364 -4038
rect -1227 -4042 -1223 -4038
rect -1223 -4056 -1219 -4052
rect -1207 -4034 -1203 -4030
rect -1207 -4063 -1203 -4059
rect -1193 -4042 -1189 -4038
rect -1183 -4049 -1179 -4045
rect -1169 -4034 -1165 -4030
rect -1165 -4063 -1161 -4059
rect -1141 -4042 -1137 -4038
rect -1151 -4049 -1147 -4045
rect -1127 -4063 -1123 -4059
rect -1109 -4034 -1105 -4030
rect -1099 -4049 -1095 -4045
rect -1109 -4056 -1105 -4052
rect -1085 -4034 -1081 -4030
rect -1081 -4042 -1077 -4038
rect -1067 -4049 -1063 -4045
rect -1057 -4056 -1053 -4052
rect -1043 -4042 -1039 -4038
rect -928 -4042 -924 -4038
rect -924 -4056 -920 -4052
rect -908 -4034 -904 -4030
rect -908 -4063 -904 -4059
rect -894 -4042 -890 -4038
rect -884 -4049 -880 -4045
rect -870 -4034 -866 -4030
rect -866 -4063 -862 -4059
rect -842 -4042 -838 -4038
rect -852 -4049 -848 -4045
rect -828 -4063 -824 -4059
rect -810 -4034 -806 -4030
rect -800 -4049 -796 -4045
rect -810 -4056 -806 -4052
rect -786 -4034 -782 -4030
rect -782 -4042 -778 -4038
rect -768 -4049 -764 -4045
rect -758 -4056 -754 -4052
rect -744 -4042 -740 -4038
rect -570 -4042 -566 -4038
rect -566 -4056 -562 -4052
rect -550 -4034 -546 -4030
rect -550 -4063 -546 -4059
rect -536 -4042 -532 -4038
rect -526 -4049 -522 -4045
rect -512 -4034 -508 -4030
rect -508 -4063 -504 -4059
rect -484 -4042 -480 -4038
rect -494 -4049 -490 -4045
rect -470 -4063 -466 -4059
rect -452 -4034 -448 -4030
rect -442 -4049 -438 -4045
rect -452 -4056 -448 -4052
rect -428 -4034 -424 -4030
rect -424 -4042 -420 -4038
rect -410 -4049 -406 -4045
rect -400 -4056 -396 -4052
rect -386 -4042 -382 -4038
rect -212 -4042 -208 -4038
rect -208 -4056 -204 -4052
rect -192 -4034 -188 -4030
rect -192 -4063 -188 -4059
rect -178 -4042 -174 -4038
rect -168 -4049 -164 -4045
rect -154 -4034 -150 -4030
rect -150 -4063 -146 -4059
rect -126 -4042 -122 -4038
rect -136 -4049 -132 -4045
rect -112 -4063 -108 -4059
rect -94 -4034 -90 -4030
rect -84 -4049 -80 -4045
rect -94 -4056 -90 -4052
rect -70 -4034 -66 -4030
rect -66 -4042 -62 -4038
rect -52 -4049 -48 -4045
rect -42 -4056 -38 -4052
rect -28 -4042 -24 -4038
rect 146 -4042 150 -4038
rect 150 -4056 154 -4052
rect 166 -4034 170 -4030
rect 166 -4063 170 -4059
rect 180 -4042 184 -4038
rect 190 -4049 194 -4045
rect 204 -4034 208 -4030
rect 208 -4063 212 -4059
rect 232 -4042 236 -4038
rect 222 -4049 226 -4045
rect 246 -4063 250 -4059
rect 264 -4034 268 -4030
rect 274 -4049 278 -4045
rect 264 -4056 268 -4052
rect 288 -4034 292 -4030
rect 292 -4042 296 -4038
rect 306 -4049 310 -4045
rect 316 -4056 320 -4052
rect 330 -4042 334 -4038
rect 502 -4042 506 -4038
rect 506 -4056 510 -4052
rect 522 -4034 526 -4030
rect 522 -4063 526 -4059
rect 536 -4042 540 -4038
rect 546 -4049 550 -4045
rect 560 -4034 564 -4030
rect 564 -4063 568 -4059
rect 588 -4042 592 -4038
rect 578 -4049 582 -4045
rect 602 -4063 606 -4059
rect 620 -4034 624 -4030
rect 630 -4049 634 -4045
rect 620 -4056 624 -4052
rect 644 -4034 648 -4030
rect 648 -4042 652 -4038
rect 662 -4049 666 -4045
rect 672 -4056 676 -4052
rect 686 -4042 690 -4038
rect 860 -4042 864 -4038
rect 864 -4056 868 -4052
rect 880 -4034 884 -4030
rect 880 -4063 884 -4059
rect 894 -4042 898 -4038
rect 904 -4049 908 -4045
rect 918 -4034 922 -4030
rect 922 -4063 926 -4059
rect 946 -4042 950 -4038
rect 936 -4049 940 -4045
rect 960 -4063 964 -4059
rect 978 -4034 982 -4030
rect 988 -4049 992 -4045
rect 978 -4056 982 -4052
rect 1002 -4034 1006 -4030
rect 1006 -4042 1010 -4038
rect 1020 -4049 1024 -4045
rect 1030 -4056 1034 -4052
rect 1044 -4042 1048 -4038
rect 1218 -4042 1222 -4038
rect 1222 -4056 1226 -4052
rect 1238 -4034 1242 -4030
rect 1238 -4063 1242 -4059
rect 1252 -4042 1256 -4038
rect 1262 -4049 1266 -4045
rect 1276 -4034 1280 -4030
rect 1280 -4063 1284 -4059
rect 1304 -4042 1308 -4038
rect 1294 -4049 1298 -4045
rect 1318 -4063 1322 -4059
rect 1336 -4034 1340 -4030
rect 1346 -4049 1350 -4045
rect 1336 -4056 1340 -4052
rect 1360 -4034 1364 -4030
rect 1364 -4042 1368 -4038
rect 1378 -4049 1382 -4045
rect 1388 -4056 1392 -4052
rect 1402 -4042 1406 -4038
rect -1308 -4133 -1304 -4129
rect -1297 -4141 -1293 -4137
rect -1290 -4163 -1286 -4159
rect -934 -4133 -930 -4129
rect -923 -4141 -919 -4137
rect -916 -4163 -912 -4159
rect -576 -4133 -572 -4129
rect -565 -4141 -561 -4137
rect -558 -4163 -554 -4159
rect -218 -4133 -214 -4129
rect -207 -4141 -203 -4137
rect -200 -4163 -196 -4159
rect 140 -4133 144 -4129
rect 151 -4141 155 -4137
rect 158 -4163 162 -4159
rect 496 -4133 500 -4129
rect 507 -4141 511 -4137
rect 514 -4163 518 -4159
rect 854 -4133 858 -4129
rect 865 -4141 869 -4137
rect 872 -4163 876 -4159
rect 1212 -4133 1216 -4129
rect 1223 -4141 1227 -4137
rect 1230 -4163 1234 -4159
rect -1223 -4316 -1219 -4312
rect -1227 -4323 -1223 -4319
rect -1207 -4303 -1203 -4299
rect -1197 -4323 -1193 -4319
rect -1183 -4316 -1179 -4312
rect -1173 -4309 -1169 -4305
rect -1163 -4316 -1159 -4312
rect -1149 -4323 -1145 -4319
rect -1145 -4337 -1141 -4333
rect -924 -4279 -920 -4275
rect -928 -4300 -924 -4296
rect -924 -4315 -920 -4311
rect -928 -4329 -924 -4325
rect -898 -4300 -894 -4296
rect -902 -4308 -898 -4304
rect -902 -4322 -898 -4318
rect -882 -4286 -878 -4282
rect -872 -4329 -868 -4325
rect -858 -4279 -854 -4275
rect -848 -4293 -844 -4289
rect -838 -4329 -834 -4325
rect -824 -4279 -820 -4275
rect -820 -4337 -816 -4333
rect -804 -4308 -800 -4304
rect -794 -4322 -790 -4318
rect -780 -4279 -776 -4275
rect -780 -4300 -776 -4296
rect -776 -4315 -772 -4311
rect -760 -4322 -756 -4318
rect -746 -4279 -742 -4275
rect -736 -4330 -732 -4326
rect -720 -4337 -716 -4333
rect -706 -4293 -702 -4289
rect -702 -4330 -698 -4326
rect -566 -4279 -562 -4275
rect -570 -4300 -566 -4296
rect -566 -4315 -562 -4311
rect -570 -4329 -566 -4325
rect -540 -4300 -536 -4296
rect -544 -4308 -540 -4304
rect -544 -4322 -540 -4318
rect -524 -4286 -520 -4282
rect -514 -4329 -510 -4325
rect -500 -4279 -496 -4275
rect -490 -4293 -486 -4289
rect -480 -4329 -476 -4325
rect -466 -4279 -462 -4275
rect -462 -4337 -458 -4333
rect -446 -4308 -442 -4304
rect -436 -4322 -432 -4318
rect -422 -4279 -418 -4275
rect -422 -4300 -418 -4296
rect -418 -4315 -414 -4311
rect -402 -4322 -398 -4318
rect -388 -4279 -384 -4275
rect -378 -4330 -374 -4326
rect -362 -4337 -358 -4333
rect -348 -4293 -344 -4289
rect -344 -4330 -340 -4326
rect -208 -4279 -204 -4275
rect -212 -4300 -208 -4296
rect -208 -4315 -204 -4311
rect -212 -4329 -208 -4325
rect -182 -4300 -178 -4296
rect -186 -4308 -182 -4304
rect -186 -4322 -182 -4318
rect -166 -4286 -162 -4282
rect -156 -4329 -152 -4325
rect -142 -4279 -138 -4275
rect -132 -4293 -128 -4289
rect -122 -4329 -118 -4325
rect -108 -4279 -104 -4275
rect -104 -4337 -100 -4333
rect -88 -4308 -84 -4304
rect -78 -4322 -74 -4318
rect -64 -4279 -60 -4275
rect -64 -4300 -60 -4296
rect -60 -4315 -56 -4311
rect -44 -4322 -40 -4318
rect -30 -4279 -26 -4275
rect -20 -4330 -16 -4326
rect -4 -4337 0 -4333
rect 10 -4293 14 -4289
rect 14 -4330 18 -4326
rect 150 -4279 154 -4275
rect 146 -4300 150 -4296
rect 150 -4315 154 -4311
rect 146 -4329 150 -4325
rect 176 -4300 180 -4296
rect 172 -4308 176 -4304
rect 172 -4322 176 -4318
rect 192 -4286 196 -4282
rect 202 -4329 206 -4325
rect 216 -4279 220 -4275
rect 226 -4293 230 -4289
rect 236 -4329 240 -4325
rect 250 -4279 254 -4275
rect 254 -4337 258 -4333
rect 270 -4308 274 -4304
rect 280 -4322 284 -4318
rect 294 -4279 298 -4275
rect 294 -4300 298 -4296
rect 298 -4315 302 -4311
rect 314 -4322 318 -4318
rect 328 -4279 332 -4275
rect 338 -4330 342 -4326
rect 354 -4337 358 -4333
rect 368 -4293 372 -4289
rect 372 -4330 376 -4326
rect 506 -4279 510 -4275
rect 502 -4300 506 -4296
rect 506 -4315 510 -4311
rect 502 -4329 506 -4325
rect 532 -4300 536 -4296
rect 528 -4308 532 -4304
rect 528 -4322 532 -4318
rect 548 -4286 552 -4282
rect 558 -4329 562 -4325
rect 572 -4279 576 -4275
rect 582 -4293 586 -4289
rect 592 -4329 596 -4325
rect 606 -4279 610 -4275
rect 610 -4337 614 -4333
rect 626 -4308 630 -4304
rect 636 -4322 640 -4318
rect 650 -4279 654 -4275
rect 650 -4300 654 -4296
rect 654 -4315 658 -4311
rect 670 -4322 674 -4318
rect 684 -4279 688 -4275
rect 694 -4330 698 -4326
rect 710 -4337 714 -4333
rect 724 -4293 728 -4289
rect 728 -4330 732 -4326
rect 864 -4279 868 -4275
rect 860 -4300 864 -4296
rect 864 -4315 868 -4311
rect 860 -4329 864 -4325
rect 890 -4300 894 -4296
rect 886 -4308 890 -4304
rect 886 -4322 890 -4318
rect 906 -4286 910 -4282
rect 916 -4329 920 -4325
rect 930 -4279 934 -4275
rect 940 -4293 944 -4289
rect 950 -4329 954 -4325
rect 964 -4279 968 -4275
rect 968 -4337 972 -4333
rect 984 -4308 988 -4304
rect 994 -4322 998 -4318
rect 1008 -4279 1012 -4275
rect 1008 -4300 1012 -4296
rect 1012 -4315 1016 -4311
rect 1028 -4322 1032 -4318
rect 1042 -4279 1046 -4275
rect 1052 -4330 1056 -4326
rect 1068 -4337 1072 -4333
rect 1082 -4293 1086 -4289
rect 1086 -4330 1090 -4326
rect 1222 -4279 1226 -4275
rect 1218 -4300 1222 -4296
rect 1222 -4315 1226 -4311
rect 1218 -4329 1222 -4325
rect 1248 -4300 1252 -4296
rect 1244 -4308 1248 -4304
rect 1244 -4322 1248 -4318
rect 1264 -4286 1268 -4282
rect 1274 -4329 1278 -4325
rect 1288 -4279 1292 -4275
rect 1298 -4293 1302 -4289
rect 1308 -4329 1312 -4325
rect 1322 -4279 1326 -4275
rect 1326 -4337 1330 -4333
rect 1342 -4308 1346 -4304
rect 1352 -4322 1356 -4318
rect 1366 -4279 1370 -4275
rect 1366 -4300 1370 -4296
rect 1370 -4315 1374 -4311
rect 1386 -4322 1390 -4318
rect 1400 -4279 1404 -4275
rect 1410 -4330 1414 -4326
rect 1426 -4337 1430 -4333
rect 1440 -4293 1444 -4289
rect 1444 -4330 1448 -4326
rect -1807 -4439 -1803 -4435
rect -1803 -4453 -1799 -4449
rect -1787 -4431 -1783 -4427
rect -1787 -4460 -1783 -4456
rect -1773 -4439 -1769 -4435
rect -1763 -4446 -1759 -4442
rect -1749 -4431 -1745 -4427
rect -1745 -4460 -1741 -4456
rect -1721 -4439 -1717 -4435
rect -1731 -4446 -1727 -4442
rect -1707 -4460 -1703 -4456
rect -1689 -4431 -1685 -4427
rect -1679 -4446 -1675 -4442
rect -1689 -4453 -1685 -4449
rect -1665 -4431 -1661 -4427
rect -1661 -4439 -1657 -4435
rect -1647 -4446 -1643 -4442
rect -1637 -4453 -1633 -4449
rect -1623 -4439 -1619 -4435
rect -1544 -4439 -1540 -4435
rect -1540 -4453 -1536 -4449
rect -1524 -4431 -1520 -4427
rect -1524 -4460 -1520 -4456
rect -1510 -4439 -1506 -4435
rect -1500 -4446 -1496 -4442
rect -1486 -4431 -1482 -4427
rect -1482 -4460 -1478 -4456
rect -1458 -4439 -1454 -4435
rect -1468 -4446 -1464 -4442
rect -1444 -4460 -1440 -4456
rect -1426 -4431 -1422 -4427
rect -1416 -4446 -1412 -4442
rect -1426 -4453 -1422 -4449
rect -1402 -4431 -1398 -4427
rect -1398 -4439 -1394 -4435
rect -1384 -4446 -1380 -4442
rect -1374 -4453 -1370 -4449
rect -1360 -4439 -1356 -4435
rect -1227 -4439 -1223 -4435
rect -1223 -4453 -1219 -4449
rect -1207 -4431 -1203 -4427
rect -1207 -4460 -1203 -4456
rect -1193 -4439 -1189 -4435
rect -1183 -4446 -1179 -4442
rect -1169 -4431 -1165 -4427
rect -1165 -4460 -1161 -4456
rect -1141 -4439 -1137 -4435
rect -1151 -4446 -1147 -4442
rect -1127 -4460 -1123 -4456
rect -1109 -4431 -1105 -4427
rect -1099 -4446 -1095 -4442
rect -1109 -4453 -1105 -4449
rect -1085 -4431 -1081 -4427
rect -1081 -4439 -1077 -4435
rect -1067 -4446 -1063 -4442
rect -1057 -4453 -1053 -4449
rect -1043 -4439 -1039 -4435
rect -928 -4439 -924 -4435
rect -924 -4453 -920 -4449
rect -908 -4431 -904 -4427
rect -908 -4460 -904 -4456
rect -894 -4439 -890 -4435
rect -884 -4446 -880 -4442
rect -870 -4431 -866 -4427
rect -866 -4460 -862 -4456
rect -842 -4439 -838 -4435
rect -852 -4446 -848 -4442
rect -828 -4460 -824 -4456
rect -810 -4431 -806 -4427
rect -800 -4446 -796 -4442
rect -810 -4453 -806 -4449
rect -786 -4431 -782 -4427
rect -782 -4439 -778 -4435
rect -768 -4446 -764 -4442
rect -758 -4453 -754 -4449
rect -744 -4439 -740 -4435
rect -570 -4439 -566 -4435
rect -566 -4453 -562 -4449
rect -550 -4431 -546 -4427
rect -550 -4460 -546 -4456
rect -536 -4439 -532 -4435
rect -526 -4446 -522 -4442
rect -512 -4431 -508 -4427
rect -508 -4460 -504 -4456
rect -484 -4439 -480 -4435
rect -494 -4446 -490 -4442
rect -470 -4460 -466 -4456
rect -452 -4431 -448 -4427
rect -442 -4446 -438 -4442
rect -452 -4453 -448 -4449
rect -428 -4431 -424 -4427
rect -424 -4439 -420 -4435
rect -410 -4446 -406 -4442
rect -400 -4453 -396 -4449
rect -386 -4439 -382 -4435
rect -1807 -4610 -1803 -4606
rect -1803 -4624 -1799 -4620
rect -1787 -4602 -1783 -4598
rect -1787 -4631 -1783 -4627
rect -1773 -4610 -1769 -4606
rect -1763 -4617 -1759 -4613
rect -1749 -4602 -1745 -4598
rect -1745 -4631 -1741 -4627
rect -1721 -4610 -1717 -4606
rect -1731 -4617 -1727 -4613
rect -1707 -4631 -1703 -4627
rect -1689 -4602 -1685 -4598
rect -1679 -4617 -1675 -4613
rect -1689 -4624 -1685 -4620
rect -1665 -4602 -1661 -4598
rect -1661 -4610 -1657 -4606
rect -1647 -4617 -1643 -4613
rect -1637 -4624 -1633 -4620
rect -1623 -4610 -1619 -4606
rect -1544 -4610 -1540 -4606
rect -1540 -4624 -1536 -4620
rect -1524 -4602 -1520 -4598
rect -1524 -4631 -1520 -4627
rect -1510 -4610 -1506 -4606
rect -1500 -4617 -1496 -4613
rect -1486 -4602 -1482 -4598
rect -1482 -4631 -1478 -4627
rect -1458 -4610 -1454 -4606
rect -1468 -4617 -1464 -4613
rect -1444 -4631 -1440 -4627
rect -1426 -4602 -1422 -4598
rect -1416 -4617 -1412 -4613
rect -1426 -4624 -1422 -4620
rect -1402 -4602 -1398 -4598
rect -1398 -4610 -1394 -4606
rect -1384 -4617 -1380 -4613
rect -1374 -4624 -1370 -4620
rect -1360 -4610 -1356 -4606
rect -1227 -4610 -1223 -4606
rect -1223 -4624 -1219 -4620
rect -1207 -4602 -1203 -4598
rect -1207 -4631 -1203 -4627
rect -1193 -4610 -1189 -4606
rect -1183 -4617 -1179 -4613
rect -1169 -4602 -1165 -4598
rect -1165 -4631 -1161 -4627
rect -1141 -4610 -1137 -4606
rect -1151 -4617 -1147 -4613
rect -1127 -4631 -1123 -4627
rect -1109 -4602 -1105 -4598
rect -1099 -4617 -1095 -4613
rect -1109 -4624 -1105 -4620
rect -1085 -4602 -1081 -4598
rect -1081 -4610 -1077 -4606
rect -1067 -4617 -1063 -4613
rect -1057 -4624 -1053 -4620
rect -1043 -4610 -1039 -4606
rect -928 -4610 -924 -4606
rect -924 -4624 -920 -4620
rect -908 -4602 -904 -4598
rect -908 -4631 -904 -4627
rect -894 -4610 -890 -4606
rect -884 -4617 -880 -4613
rect -870 -4602 -866 -4598
rect -866 -4631 -862 -4627
rect -842 -4610 -838 -4606
rect -852 -4617 -848 -4613
rect -828 -4631 -824 -4627
rect -810 -4602 -806 -4598
rect -800 -4617 -796 -4613
rect -810 -4624 -806 -4620
rect -786 -4602 -782 -4598
rect -782 -4610 -778 -4606
rect -768 -4617 -764 -4613
rect -758 -4624 -754 -4620
rect -744 -4610 -740 -4606
rect -570 -4610 -566 -4606
rect -566 -4624 -562 -4620
rect -550 -4602 -546 -4598
rect -550 -4631 -546 -4627
rect -536 -4610 -532 -4606
rect -526 -4617 -522 -4613
rect -512 -4602 -508 -4598
rect -508 -4631 -504 -4627
rect -484 -4610 -480 -4606
rect -494 -4617 -490 -4613
rect -470 -4631 -466 -4627
rect -452 -4602 -448 -4598
rect -442 -4617 -438 -4613
rect -452 -4624 -448 -4620
rect -428 -4602 -424 -4598
rect -424 -4610 -420 -4606
rect -410 -4617 -406 -4613
rect -400 -4624 -396 -4620
rect -386 -4610 -382 -4606
rect -212 -4610 -208 -4606
rect -208 -4624 -204 -4620
rect -192 -4602 -188 -4598
rect -192 -4631 -188 -4627
rect -178 -4610 -174 -4606
rect -168 -4617 -164 -4613
rect -154 -4602 -150 -4598
rect -150 -4631 -146 -4627
rect -126 -4610 -122 -4606
rect -136 -4617 -132 -4613
rect -112 -4631 -108 -4627
rect -94 -4602 -90 -4598
rect -84 -4617 -80 -4613
rect -94 -4624 -90 -4620
rect -70 -4602 -66 -4598
rect -66 -4610 -62 -4606
rect -52 -4617 -48 -4613
rect -42 -4624 -38 -4620
rect -28 -4610 -24 -4606
rect 146 -4610 150 -4606
rect 150 -4624 154 -4620
rect 166 -4602 170 -4598
rect 166 -4631 170 -4627
rect 180 -4610 184 -4606
rect 190 -4617 194 -4613
rect 204 -4602 208 -4598
rect 208 -4631 212 -4627
rect 232 -4610 236 -4606
rect 222 -4617 226 -4613
rect 246 -4631 250 -4627
rect 264 -4602 268 -4598
rect 274 -4617 278 -4613
rect 264 -4624 268 -4620
rect 288 -4602 292 -4598
rect 292 -4610 296 -4606
rect 306 -4617 310 -4613
rect 316 -4624 320 -4620
rect 330 -4610 334 -4606
rect 502 -4610 506 -4606
rect 506 -4624 510 -4620
rect 522 -4602 526 -4598
rect 522 -4631 526 -4627
rect 536 -4610 540 -4606
rect 546 -4617 550 -4613
rect 560 -4602 564 -4598
rect 564 -4631 568 -4627
rect 588 -4610 592 -4606
rect 578 -4617 582 -4613
rect 602 -4631 606 -4627
rect 620 -4602 624 -4598
rect 630 -4617 634 -4613
rect 620 -4624 624 -4620
rect 644 -4602 648 -4598
rect 648 -4610 652 -4606
rect 662 -4617 666 -4613
rect 672 -4624 676 -4620
rect 686 -4610 690 -4606
rect 860 -4610 864 -4606
rect 864 -4624 868 -4620
rect 880 -4602 884 -4598
rect 880 -4631 884 -4627
rect 894 -4610 898 -4606
rect 904 -4617 908 -4613
rect 918 -4602 922 -4598
rect 922 -4631 926 -4627
rect 946 -4610 950 -4606
rect 936 -4617 940 -4613
rect 960 -4631 964 -4627
rect 978 -4602 982 -4598
rect 988 -4617 992 -4613
rect 978 -4624 982 -4620
rect 1002 -4602 1006 -4598
rect 1006 -4610 1010 -4606
rect 1020 -4617 1024 -4613
rect 1030 -4624 1034 -4620
rect 1044 -4610 1048 -4606
rect 1218 -4610 1222 -4606
rect 1222 -4624 1226 -4620
rect 1238 -4602 1242 -4598
rect 1238 -4631 1242 -4627
rect 1252 -4610 1256 -4606
rect 1262 -4617 1266 -4613
rect 1276 -4602 1280 -4598
rect 1280 -4631 1284 -4627
rect 1304 -4610 1308 -4606
rect 1294 -4617 1298 -4613
rect 1318 -4631 1322 -4627
rect 1336 -4602 1340 -4598
rect 1346 -4617 1350 -4613
rect 1336 -4624 1340 -4620
rect 1360 -4602 1364 -4598
rect 1364 -4610 1368 -4606
rect 1378 -4617 1382 -4613
rect 1388 -4624 1392 -4620
rect 1402 -4610 1406 -4606
rect -1544 -4781 -1540 -4777
rect -1540 -4795 -1536 -4791
rect -1524 -4773 -1520 -4769
rect -1524 -4802 -1520 -4798
rect -1510 -4781 -1506 -4777
rect -1500 -4788 -1496 -4784
rect -1486 -4773 -1482 -4769
rect -1482 -4802 -1478 -4798
rect -1458 -4781 -1454 -4777
rect -1468 -4788 -1464 -4784
rect -1444 -4802 -1440 -4798
rect -1426 -4773 -1422 -4769
rect -1416 -4788 -1412 -4784
rect -1426 -4795 -1422 -4791
rect -1402 -4773 -1398 -4769
rect -1398 -4781 -1394 -4777
rect -1384 -4788 -1380 -4784
rect -1374 -4795 -1370 -4791
rect -1360 -4781 -1356 -4777
rect -1227 -4781 -1223 -4777
rect -1223 -4795 -1219 -4791
rect -1207 -4773 -1203 -4769
rect -1207 -4802 -1203 -4798
rect -1193 -4781 -1189 -4777
rect -1183 -4788 -1179 -4784
rect -1169 -4773 -1165 -4769
rect -1165 -4802 -1161 -4798
rect -1141 -4781 -1137 -4777
rect -1151 -4788 -1147 -4784
rect -1127 -4802 -1123 -4798
rect -1109 -4773 -1105 -4769
rect -1099 -4788 -1095 -4784
rect -1109 -4795 -1105 -4791
rect -1085 -4773 -1081 -4769
rect -1081 -4781 -1077 -4777
rect -1067 -4788 -1063 -4784
rect -1057 -4795 -1053 -4791
rect -1043 -4781 -1039 -4777
rect -928 -4781 -924 -4777
rect -924 -4795 -920 -4791
rect -908 -4773 -904 -4769
rect -908 -4802 -904 -4798
rect -894 -4781 -890 -4777
rect -884 -4788 -880 -4784
rect -870 -4773 -866 -4769
rect -866 -4802 -862 -4798
rect -842 -4781 -838 -4777
rect -852 -4788 -848 -4784
rect -828 -4802 -824 -4798
rect -810 -4773 -806 -4769
rect -800 -4788 -796 -4784
rect -810 -4795 -806 -4791
rect -786 -4773 -782 -4769
rect -782 -4781 -778 -4777
rect -768 -4788 -764 -4784
rect -758 -4795 -754 -4791
rect -744 -4781 -740 -4777
rect -570 -4781 -566 -4777
rect -566 -4795 -562 -4791
rect -550 -4773 -546 -4769
rect -550 -4802 -546 -4798
rect -536 -4781 -532 -4777
rect -526 -4788 -522 -4784
rect -512 -4773 -508 -4769
rect -508 -4802 -504 -4798
rect -484 -4781 -480 -4777
rect -494 -4788 -490 -4784
rect -470 -4802 -466 -4798
rect -452 -4773 -448 -4769
rect -442 -4788 -438 -4784
rect -452 -4795 -448 -4791
rect -428 -4773 -424 -4769
rect -424 -4781 -420 -4777
rect -410 -4788 -406 -4784
rect -400 -4795 -396 -4791
rect -386 -4781 -382 -4777
rect -212 -4781 -208 -4777
rect -208 -4795 -204 -4791
rect -192 -4773 -188 -4769
rect -192 -4802 -188 -4798
rect -178 -4781 -174 -4777
rect -168 -4788 -164 -4784
rect -154 -4773 -150 -4769
rect -150 -4802 -146 -4798
rect -126 -4781 -122 -4777
rect -136 -4788 -132 -4784
rect -112 -4802 -108 -4798
rect -94 -4773 -90 -4769
rect -84 -4788 -80 -4784
rect -94 -4795 -90 -4791
rect -70 -4773 -66 -4769
rect -66 -4781 -62 -4777
rect -52 -4788 -48 -4784
rect -42 -4795 -38 -4791
rect -28 -4781 -24 -4777
rect 146 -4781 150 -4777
rect 150 -4795 154 -4791
rect 166 -4773 170 -4769
rect 166 -4802 170 -4798
rect 180 -4781 184 -4777
rect 190 -4788 194 -4784
rect 204 -4773 208 -4769
rect 208 -4802 212 -4798
rect 232 -4781 236 -4777
rect 222 -4788 226 -4784
rect 246 -4802 250 -4798
rect 264 -4773 268 -4769
rect 274 -4788 278 -4784
rect 264 -4795 268 -4791
rect 288 -4773 292 -4769
rect 292 -4781 296 -4777
rect 306 -4788 310 -4784
rect 316 -4795 320 -4791
rect 330 -4781 334 -4777
rect 502 -4781 506 -4777
rect 506 -4795 510 -4791
rect 522 -4773 526 -4769
rect 522 -4802 526 -4798
rect 536 -4781 540 -4777
rect 546 -4788 550 -4784
rect 560 -4773 564 -4769
rect 564 -4802 568 -4798
rect 588 -4781 592 -4777
rect 578 -4788 582 -4784
rect 602 -4802 606 -4798
rect 620 -4773 624 -4769
rect 630 -4788 634 -4784
rect 620 -4795 624 -4791
rect 644 -4773 648 -4769
rect 648 -4781 652 -4777
rect 662 -4788 666 -4784
rect 672 -4795 676 -4791
rect 686 -4781 690 -4777
rect 860 -4781 864 -4777
rect 864 -4795 868 -4791
rect 880 -4773 884 -4769
rect 880 -4802 884 -4798
rect 894 -4781 898 -4777
rect 904 -4788 908 -4784
rect 918 -4773 922 -4769
rect 922 -4802 926 -4798
rect 946 -4781 950 -4777
rect 936 -4788 940 -4784
rect 960 -4802 964 -4798
rect 978 -4773 982 -4769
rect 988 -4788 992 -4784
rect 978 -4795 982 -4791
rect 1002 -4773 1006 -4769
rect 1006 -4781 1010 -4777
rect 1020 -4788 1024 -4784
rect 1030 -4795 1034 -4791
rect 1044 -4781 1048 -4777
rect 1218 -4781 1222 -4777
rect 1222 -4795 1226 -4791
rect 1238 -4773 1242 -4769
rect 1238 -4802 1242 -4798
rect 1252 -4781 1256 -4777
rect 1262 -4788 1266 -4784
rect 1276 -4773 1280 -4769
rect 1280 -4802 1284 -4798
rect 1304 -4781 1308 -4777
rect 1294 -4788 1298 -4784
rect 1318 -4802 1322 -4798
rect 1336 -4773 1340 -4769
rect 1346 -4788 1350 -4784
rect 1336 -4795 1340 -4791
rect 1360 -4773 1364 -4769
rect 1364 -4781 1368 -4777
rect 1378 -4788 1382 -4784
rect 1388 -4795 1392 -4791
rect 1402 -4781 1406 -4777
rect -1308 -4872 -1304 -4868
rect -1297 -4880 -1293 -4876
rect -1290 -4902 -1286 -4898
rect -934 -4872 -930 -4868
rect -923 -4880 -919 -4876
rect -916 -4902 -912 -4898
rect -576 -4872 -572 -4868
rect -565 -4880 -561 -4876
rect -558 -4902 -554 -4898
rect -218 -4872 -214 -4868
rect -207 -4880 -203 -4876
rect -200 -4902 -196 -4898
rect 140 -4872 144 -4868
rect 151 -4880 155 -4876
rect 158 -4902 162 -4898
rect 496 -4872 500 -4868
rect 507 -4880 511 -4876
rect 514 -4902 518 -4898
rect 854 -4872 858 -4868
rect 865 -4880 869 -4876
rect 872 -4902 876 -4898
rect 1212 -4872 1216 -4868
rect 1223 -4880 1227 -4876
rect 1230 -4902 1234 -4898
rect -1223 -5055 -1219 -5051
rect -1227 -5062 -1223 -5058
rect -1207 -5042 -1203 -5038
rect -1197 -5062 -1193 -5058
rect -1183 -5055 -1179 -5051
rect -1173 -5048 -1169 -5044
rect -1163 -5055 -1159 -5051
rect -1149 -5062 -1145 -5058
rect -1145 -5076 -1141 -5072
rect -924 -5018 -920 -5014
rect -928 -5039 -924 -5035
rect -924 -5054 -920 -5050
rect -928 -5068 -924 -5064
rect -898 -5039 -894 -5035
rect -902 -5047 -898 -5043
rect -902 -5061 -898 -5057
rect -882 -5025 -878 -5021
rect -872 -5068 -868 -5064
rect -858 -5018 -854 -5014
rect -848 -5032 -844 -5028
rect -838 -5068 -834 -5064
rect -824 -5018 -820 -5014
rect -820 -5076 -816 -5072
rect -804 -5047 -800 -5043
rect -794 -5061 -790 -5057
rect -780 -5018 -776 -5014
rect -780 -5039 -776 -5035
rect -776 -5054 -772 -5050
rect -760 -5061 -756 -5057
rect -746 -5018 -742 -5014
rect -736 -5069 -732 -5065
rect -720 -5076 -716 -5072
rect -706 -5032 -702 -5028
rect -702 -5069 -698 -5065
rect -566 -5018 -562 -5014
rect -570 -5039 -566 -5035
rect -566 -5054 -562 -5050
rect -570 -5068 -566 -5064
rect -540 -5039 -536 -5035
rect -544 -5047 -540 -5043
rect -544 -5061 -540 -5057
rect -524 -5025 -520 -5021
rect -514 -5068 -510 -5064
rect -500 -5018 -496 -5014
rect -490 -5032 -486 -5028
rect -480 -5068 -476 -5064
rect -466 -5018 -462 -5014
rect -462 -5076 -458 -5072
rect -446 -5047 -442 -5043
rect -436 -5061 -432 -5057
rect -422 -5018 -418 -5014
rect -422 -5039 -418 -5035
rect -418 -5054 -414 -5050
rect -402 -5061 -398 -5057
rect -388 -5018 -384 -5014
rect -378 -5069 -374 -5065
rect -362 -5076 -358 -5072
rect -348 -5032 -344 -5028
rect -344 -5069 -340 -5065
rect -208 -5018 -204 -5014
rect -212 -5039 -208 -5035
rect -208 -5054 -204 -5050
rect -212 -5068 -208 -5064
rect -182 -5039 -178 -5035
rect -186 -5047 -182 -5043
rect -186 -5061 -182 -5057
rect -166 -5025 -162 -5021
rect -156 -5068 -152 -5064
rect -142 -5018 -138 -5014
rect -132 -5032 -128 -5028
rect -122 -5068 -118 -5064
rect -108 -5018 -104 -5014
rect -104 -5076 -100 -5072
rect -88 -5047 -84 -5043
rect -78 -5061 -74 -5057
rect -64 -5018 -60 -5014
rect -64 -5039 -60 -5035
rect -60 -5054 -56 -5050
rect -44 -5061 -40 -5057
rect -30 -5018 -26 -5014
rect -20 -5069 -16 -5065
rect -4 -5076 0 -5072
rect 10 -5032 14 -5028
rect 14 -5069 18 -5065
rect 150 -5018 154 -5014
rect 146 -5039 150 -5035
rect 150 -5054 154 -5050
rect 146 -5068 150 -5064
rect 176 -5039 180 -5035
rect 172 -5047 176 -5043
rect 172 -5061 176 -5057
rect 192 -5025 196 -5021
rect 202 -5068 206 -5064
rect 216 -5018 220 -5014
rect 226 -5032 230 -5028
rect 236 -5068 240 -5064
rect 250 -5018 254 -5014
rect 254 -5076 258 -5072
rect 270 -5047 274 -5043
rect 280 -5061 284 -5057
rect 294 -5018 298 -5014
rect 294 -5039 298 -5035
rect 298 -5054 302 -5050
rect 314 -5061 318 -5057
rect 328 -5018 332 -5014
rect 338 -5069 342 -5065
rect 354 -5076 358 -5072
rect 368 -5032 372 -5028
rect 372 -5069 376 -5065
rect 506 -5018 510 -5014
rect 502 -5039 506 -5035
rect 506 -5054 510 -5050
rect 502 -5068 506 -5064
rect 532 -5039 536 -5035
rect 528 -5047 532 -5043
rect 528 -5061 532 -5057
rect 548 -5025 552 -5021
rect 558 -5068 562 -5064
rect 572 -5018 576 -5014
rect 582 -5032 586 -5028
rect 592 -5068 596 -5064
rect 606 -5018 610 -5014
rect 610 -5076 614 -5072
rect 626 -5047 630 -5043
rect 636 -5061 640 -5057
rect 650 -5018 654 -5014
rect 650 -5039 654 -5035
rect 654 -5054 658 -5050
rect 670 -5061 674 -5057
rect 684 -5018 688 -5014
rect 694 -5069 698 -5065
rect 710 -5076 714 -5072
rect 724 -5032 728 -5028
rect 728 -5069 732 -5065
rect 864 -5018 868 -5014
rect 860 -5039 864 -5035
rect 864 -5054 868 -5050
rect 860 -5068 864 -5064
rect 890 -5039 894 -5035
rect 886 -5047 890 -5043
rect 886 -5061 890 -5057
rect 906 -5025 910 -5021
rect 916 -5068 920 -5064
rect 930 -5018 934 -5014
rect 940 -5032 944 -5028
rect 950 -5068 954 -5064
rect 964 -5018 968 -5014
rect 968 -5076 972 -5072
rect 984 -5047 988 -5043
rect 994 -5061 998 -5057
rect 1008 -5018 1012 -5014
rect 1008 -5039 1012 -5035
rect 1012 -5054 1016 -5050
rect 1028 -5061 1032 -5057
rect 1042 -5018 1046 -5014
rect 1052 -5069 1056 -5065
rect 1068 -5076 1072 -5072
rect 1082 -5032 1086 -5028
rect 1086 -5069 1090 -5065
rect 1222 -5018 1226 -5014
rect 1218 -5039 1222 -5035
rect 1222 -5054 1226 -5050
rect 1218 -5068 1222 -5064
rect 1248 -5039 1252 -5035
rect 1244 -5047 1248 -5043
rect 1244 -5061 1248 -5057
rect 1264 -5025 1268 -5021
rect 1274 -5068 1278 -5064
rect 1288 -5018 1292 -5014
rect 1298 -5032 1302 -5028
rect 1308 -5068 1312 -5064
rect 1322 -5018 1326 -5014
rect 1326 -5076 1330 -5072
rect 1342 -5047 1346 -5043
rect 1352 -5061 1356 -5057
rect 1366 -5018 1370 -5014
rect 1366 -5039 1370 -5035
rect 1370 -5054 1374 -5050
rect 1386 -5061 1390 -5057
rect 1400 -5018 1404 -5014
rect 1410 -5069 1414 -5065
rect 1426 -5076 1430 -5072
rect 1440 -5032 1444 -5028
rect 1444 -5069 1448 -5065
rect -1803 -5174 -1799 -5170
rect -1799 -5188 -1795 -5184
rect -1783 -5166 -1779 -5162
rect -1783 -5195 -1779 -5191
rect -1769 -5174 -1765 -5170
rect -1759 -5181 -1755 -5177
rect -1745 -5166 -1741 -5162
rect -1741 -5195 -1737 -5191
rect -1717 -5174 -1713 -5170
rect -1727 -5181 -1723 -5177
rect -1703 -5195 -1699 -5191
rect -1685 -5166 -1681 -5162
rect -1675 -5181 -1671 -5177
rect -1685 -5188 -1681 -5184
rect -1661 -5166 -1657 -5162
rect -1657 -5174 -1653 -5170
rect -1643 -5181 -1639 -5177
rect -1633 -5188 -1629 -5184
rect -1619 -5174 -1615 -5170
rect -1540 -5174 -1536 -5170
rect -1536 -5188 -1532 -5184
rect -1520 -5166 -1516 -5162
rect -1520 -5195 -1516 -5191
rect -1506 -5174 -1502 -5170
rect -1496 -5181 -1492 -5177
rect -1482 -5166 -1478 -5162
rect -1478 -5195 -1474 -5191
rect -1454 -5174 -1450 -5170
rect -1464 -5181 -1460 -5177
rect -1440 -5195 -1436 -5191
rect -1422 -5166 -1418 -5162
rect -1412 -5181 -1408 -5177
rect -1422 -5188 -1418 -5184
rect -1398 -5166 -1394 -5162
rect -1394 -5174 -1390 -5170
rect -1380 -5181 -1376 -5177
rect -1370 -5188 -1366 -5184
rect -1356 -5174 -1352 -5170
rect -1227 -5174 -1223 -5170
rect -1223 -5188 -1219 -5184
rect -1207 -5166 -1203 -5162
rect -1207 -5195 -1203 -5191
rect -1193 -5174 -1189 -5170
rect -1183 -5181 -1179 -5177
rect -1169 -5166 -1165 -5162
rect -1165 -5195 -1161 -5191
rect -1141 -5174 -1137 -5170
rect -1151 -5181 -1147 -5177
rect -1127 -5195 -1123 -5191
rect -1109 -5166 -1105 -5162
rect -1099 -5181 -1095 -5177
rect -1109 -5188 -1105 -5184
rect -1085 -5166 -1081 -5162
rect -1081 -5174 -1077 -5170
rect -1067 -5181 -1063 -5177
rect -1057 -5188 -1053 -5184
rect -1043 -5174 -1039 -5170
rect -928 -5174 -924 -5170
rect -924 -5188 -920 -5184
rect -908 -5166 -904 -5162
rect -908 -5195 -904 -5191
rect -894 -5174 -890 -5170
rect -884 -5181 -880 -5177
rect -870 -5166 -866 -5162
rect -866 -5195 -862 -5191
rect -842 -5174 -838 -5170
rect -852 -5181 -848 -5177
rect -828 -5195 -824 -5191
rect -810 -5166 -806 -5162
rect -800 -5181 -796 -5177
rect -810 -5188 -806 -5184
rect -786 -5166 -782 -5162
rect -782 -5174 -778 -5170
rect -768 -5181 -764 -5177
rect -758 -5188 -754 -5184
rect -744 -5174 -740 -5170
rect -1803 -5345 -1799 -5341
rect -1799 -5359 -1795 -5355
rect -1783 -5337 -1779 -5333
rect -1783 -5366 -1779 -5362
rect -1769 -5345 -1765 -5341
rect -1759 -5352 -1755 -5348
rect -1745 -5337 -1741 -5333
rect -1741 -5366 -1737 -5362
rect -1717 -5345 -1713 -5341
rect -1727 -5352 -1723 -5348
rect -1703 -5366 -1699 -5362
rect -1685 -5337 -1681 -5333
rect -1675 -5352 -1671 -5348
rect -1685 -5359 -1681 -5355
rect -1661 -5337 -1657 -5333
rect -1657 -5345 -1653 -5341
rect -1643 -5352 -1639 -5348
rect -1633 -5359 -1629 -5355
rect -1619 -5345 -1615 -5341
rect -1540 -5345 -1536 -5341
rect -1536 -5359 -1532 -5355
rect -1520 -5337 -1516 -5333
rect -1520 -5366 -1516 -5362
rect -1506 -5345 -1502 -5341
rect -1496 -5352 -1492 -5348
rect -1482 -5337 -1478 -5333
rect -1478 -5366 -1474 -5362
rect -1454 -5345 -1450 -5341
rect -1464 -5352 -1460 -5348
rect -1440 -5366 -1436 -5362
rect -1422 -5337 -1418 -5333
rect -1412 -5352 -1408 -5348
rect -1422 -5359 -1418 -5355
rect -1398 -5337 -1394 -5333
rect -1394 -5345 -1390 -5341
rect -1380 -5352 -1376 -5348
rect -1370 -5359 -1366 -5355
rect -1356 -5345 -1352 -5341
rect -1227 -5345 -1223 -5341
rect -1223 -5359 -1219 -5355
rect -1207 -5337 -1203 -5333
rect -1207 -5366 -1203 -5362
rect -1193 -5345 -1189 -5341
rect -1183 -5352 -1179 -5348
rect -1169 -5337 -1165 -5333
rect -1165 -5366 -1161 -5362
rect -1141 -5345 -1137 -5341
rect -1151 -5352 -1147 -5348
rect -1127 -5366 -1123 -5362
rect -1109 -5337 -1105 -5333
rect -1099 -5352 -1095 -5348
rect -1109 -5359 -1105 -5355
rect -1085 -5337 -1081 -5333
rect -1081 -5345 -1077 -5341
rect -1067 -5352 -1063 -5348
rect -1057 -5359 -1053 -5355
rect -1043 -5345 -1039 -5341
rect -928 -5345 -924 -5341
rect -924 -5359 -920 -5355
rect -908 -5337 -904 -5333
rect -908 -5366 -904 -5362
rect -894 -5345 -890 -5341
rect -884 -5352 -880 -5348
rect -870 -5337 -866 -5333
rect -866 -5366 -862 -5362
rect -842 -5345 -838 -5341
rect -852 -5352 -848 -5348
rect -828 -5366 -824 -5362
rect -810 -5337 -806 -5333
rect -800 -5352 -796 -5348
rect -810 -5359 -806 -5355
rect -786 -5337 -782 -5333
rect -782 -5345 -778 -5341
rect -768 -5352 -764 -5348
rect -758 -5359 -754 -5355
rect -744 -5345 -740 -5341
rect -570 -5345 -566 -5341
rect -566 -5359 -562 -5355
rect -550 -5337 -546 -5333
rect -550 -5366 -546 -5362
rect -536 -5345 -532 -5341
rect -526 -5352 -522 -5348
rect -512 -5337 -508 -5333
rect -508 -5366 -504 -5362
rect -484 -5345 -480 -5341
rect -494 -5352 -490 -5348
rect -470 -5366 -466 -5362
rect -452 -5337 -448 -5333
rect -442 -5352 -438 -5348
rect -452 -5359 -448 -5355
rect -428 -5337 -424 -5333
rect -424 -5345 -420 -5341
rect -410 -5352 -406 -5348
rect -400 -5359 -396 -5355
rect -386 -5345 -382 -5341
rect -212 -5345 -208 -5341
rect -208 -5359 -204 -5355
rect -192 -5337 -188 -5333
rect -192 -5366 -188 -5362
rect -178 -5345 -174 -5341
rect -168 -5352 -164 -5348
rect -154 -5337 -150 -5333
rect -150 -5366 -146 -5362
rect -126 -5345 -122 -5341
rect -136 -5352 -132 -5348
rect -112 -5366 -108 -5362
rect -94 -5337 -90 -5333
rect -84 -5352 -80 -5348
rect -94 -5359 -90 -5355
rect -70 -5337 -66 -5333
rect -66 -5345 -62 -5341
rect -52 -5352 -48 -5348
rect -42 -5359 -38 -5355
rect -28 -5345 -24 -5341
rect 146 -5345 150 -5341
rect 150 -5359 154 -5355
rect 166 -5337 170 -5333
rect 166 -5366 170 -5362
rect 180 -5345 184 -5341
rect 190 -5352 194 -5348
rect 204 -5337 208 -5333
rect 208 -5366 212 -5362
rect 232 -5345 236 -5341
rect 222 -5352 226 -5348
rect 246 -5366 250 -5362
rect 264 -5337 268 -5333
rect 274 -5352 278 -5348
rect 264 -5359 268 -5355
rect 288 -5337 292 -5333
rect 292 -5345 296 -5341
rect 306 -5352 310 -5348
rect 316 -5359 320 -5355
rect 330 -5345 334 -5341
rect 502 -5345 506 -5341
rect 506 -5359 510 -5355
rect 522 -5337 526 -5333
rect 522 -5366 526 -5362
rect 536 -5345 540 -5341
rect 546 -5352 550 -5348
rect 560 -5337 564 -5333
rect 564 -5366 568 -5362
rect 588 -5345 592 -5341
rect 578 -5352 582 -5348
rect 602 -5366 606 -5362
rect 620 -5337 624 -5333
rect 630 -5352 634 -5348
rect 620 -5359 624 -5355
rect 644 -5337 648 -5333
rect 648 -5345 652 -5341
rect 662 -5352 666 -5348
rect 672 -5359 676 -5355
rect 686 -5345 690 -5341
rect 860 -5345 864 -5341
rect 864 -5359 868 -5355
rect 880 -5337 884 -5333
rect 880 -5366 884 -5362
rect 894 -5345 898 -5341
rect 904 -5352 908 -5348
rect 918 -5337 922 -5333
rect 922 -5366 926 -5362
rect 946 -5345 950 -5341
rect 936 -5352 940 -5348
rect 960 -5366 964 -5362
rect 978 -5337 982 -5333
rect 988 -5352 992 -5348
rect 978 -5359 982 -5355
rect 1002 -5337 1006 -5333
rect 1006 -5345 1010 -5341
rect 1020 -5352 1024 -5348
rect 1030 -5359 1034 -5355
rect 1044 -5345 1048 -5341
rect 1218 -5345 1222 -5341
rect 1222 -5359 1226 -5355
rect 1238 -5337 1242 -5333
rect 1238 -5366 1242 -5362
rect 1252 -5345 1256 -5341
rect 1262 -5352 1266 -5348
rect 1276 -5337 1280 -5333
rect 1280 -5366 1284 -5362
rect 1304 -5345 1308 -5341
rect 1294 -5352 1298 -5348
rect 1318 -5366 1322 -5362
rect 1336 -5337 1340 -5333
rect 1346 -5352 1350 -5348
rect 1336 -5359 1340 -5355
rect 1360 -5337 1364 -5333
rect 1364 -5345 1368 -5341
rect 1378 -5352 1382 -5348
rect 1388 -5359 1392 -5355
rect 1402 -5345 1406 -5341
rect -1803 -5505 -1799 -5501
rect -1799 -5519 -1795 -5515
rect -1783 -5497 -1779 -5493
rect -1783 -5526 -1779 -5522
rect -1769 -5505 -1765 -5501
rect -1759 -5512 -1755 -5508
rect -1745 -5497 -1741 -5493
rect -1741 -5526 -1737 -5522
rect -1717 -5505 -1713 -5501
rect -1727 -5512 -1723 -5508
rect -1703 -5526 -1699 -5522
rect -1685 -5497 -1681 -5493
rect -1675 -5512 -1671 -5508
rect -1685 -5519 -1681 -5515
rect -1661 -5497 -1657 -5493
rect -1657 -5505 -1653 -5501
rect -1643 -5512 -1639 -5508
rect -1633 -5519 -1629 -5515
rect -1619 -5505 -1615 -5501
rect -1540 -5505 -1536 -5501
rect -1536 -5519 -1532 -5515
rect -1520 -5497 -1516 -5493
rect -1520 -5526 -1516 -5522
rect -1506 -5505 -1502 -5501
rect -1496 -5512 -1492 -5508
rect -1482 -5497 -1478 -5493
rect -1478 -5526 -1474 -5522
rect -1454 -5505 -1450 -5501
rect -1464 -5512 -1460 -5508
rect -1440 -5526 -1436 -5522
rect -1422 -5497 -1418 -5493
rect -1412 -5512 -1408 -5508
rect -1422 -5519 -1418 -5515
rect -1398 -5497 -1394 -5493
rect -1394 -5505 -1390 -5501
rect -1380 -5512 -1376 -5508
rect -1370 -5519 -1366 -5515
rect -1356 -5505 -1352 -5501
rect -1227 -5505 -1223 -5501
rect -1223 -5519 -1219 -5515
rect -1207 -5497 -1203 -5493
rect -1207 -5526 -1203 -5522
rect -1193 -5505 -1189 -5501
rect -1183 -5512 -1179 -5508
rect -1169 -5497 -1165 -5493
rect -1165 -5526 -1161 -5522
rect -1141 -5505 -1137 -5501
rect -1151 -5512 -1147 -5508
rect -1127 -5526 -1123 -5522
rect -1109 -5497 -1105 -5493
rect -1099 -5512 -1095 -5508
rect -1109 -5519 -1105 -5515
rect -1085 -5497 -1081 -5493
rect -1081 -5505 -1077 -5501
rect -1067 -5512 -1063 -5508
rect -1057 -5519 -1053 -5515
rect -1043 -5505 -1039 -5501
rect -928 -5505 -924 -5501
rect -924 -5519 -920 -5515
rect -908 -5497 -904 -5493
rect -908 -5526 -904 -5522
rect -894 -5505 -890 -5501
rect -884 -5512 -880 -5508
rect -870 -5497 -866 -5493
rect -866 -5526 -862 -5522
rect -842 -5505 -838 -5501
rect -852 -5512 -848 -5508
rect -828 -5526 -824 -5522
rect -810 -5497 -806 -5493
rect -800 -5512 -796 -5508
rect -810 -5519 -806 -5515
rect -786 -5497 -782 -5493
rect -782 -5505 -778 -5501
rect -768 -5512 -764 -5508
rect -758 -5519 -754 -5515
rect -744 -5505 -740 -5501
rect -570 -5505 -566 -5501
rect -566 -5519 -562 -5515
rect -550 -5497 -546 -5493
rect -550 -5526 -546 -5522
rect -536 -5505 -532 -5501
rect -526 -5512 -522 -5508
rect -512 -5497 -508 -5493
rect -508 -5526 -504 -5522
rect -484 -5505 -480 -5501
rect -494 -5512 -490 -5508
rect -470 -5526 -466 -5522
rect -452 -5497 -448 -5493
rect -442 -5512 -438 -5508
rect -452 -5519 -448 -5515
rect -428 -5497 -424 -5493
rect -424 -5505 -420 -5501
rect -410 -5512 -406 -5508
rect -400 -5519 -396 -5515
rect -386 -5505 -382 -5501
rect -212 -5505 -208 -5501
rect -208 -5519 -204 -5515
rect -192 -5497 -188 -5493
rect -192 -5526 -188 -5522
rect -178 -5505 -174 -5501
rect -168 -5512 -164 -5508
rect -154 -5497 -150 -5493
rect -150 -5526 -146 -5522
rect -126 -5505 -122 -5501
rect -136 -5512 -132 -5508
rect -112 -5526 -108 -5522
rect -94 -5497 -90 -5493
rect -84 -5512 -80 -5508
rect -94 -5519 -90 -5515
rect -70 -5497 -66 -5493
rect -66 -5505 -62 -5501
rect -52 -5512 -48 -5508
rect -42 -5519 -38 -5515
rect -28 -5505 -24 -5501
rect 146 -5505 150 -5501
rect 150 -5519 154 -5515
rect 166 -5497 170 -5493
rect 166 -5526 170 -5522
rect 180 -5505 184 -5501
rect 190 -5512 194 -5508
rect 204 -5497 208 -5493
rect 208 -5526 212 -5522
rect 232 -5505 236 -5501
rect 222 -5512 226 -5508
rect 246 -5526 250 -5522
rect 264 -5497 268 -5493
rect 274 -5512 278 -5508
rect 264 -5519 268 -5515
rect 288 -5497 292 -5493
rect 292 -5505 296 -5501
rect 306 -5512 310 -5508
rect 316 -5519 320 -5515
rect 330 -5505 334 -5501
rect 502 -5505 506 -5501
rect 506 -5519 510 -5515
rect 522 -5497 526 -5493
rect 522 -5526 526 -5522
rect 536 -5505 540 -5501
rect 546 -5512 550 -5508
rect 560 -5497 564 -5493
rect 564 -5526 568 -5522
rect 588 -5505 592 -5501
rect 578 -5512 582 -5508
rect 602 -5526 606 -5522
rect 620 -5497 624 -5493
rect 630 -5512 634 -5508
rect 620 -5519 624 -5515
rect 644 -5497 648 -5493
rect 648 -5505 652 -5501
rect 662 -5512 666 -5508
rect 672 -5519 676 -5515
rect 686 -5505 690 -5501
rect 860 -5505 864 -5501
rect 864 -5519 868 -5515
rect 880 -5497 884 -5493
rect 880 -5526 884 -5522
rect 894 -5505 898 -5501
rect 904 -5512 908 -5508
rect 918 -5497 922 -5493
rect 922 -5526 926 -5522
rect 946 -5505 950 -5501
rect 936 -5512 940 -5508
rect 960 -5526 964 -5522
rect 978 -5497 982 -5493
rect 988 -5512 992 -5508
rect 978 -5519 982 -5515
rect 1002 -5497 1006 -5493
rect 1006 -5505 1010 -5501
rect 1020 -5512 1024 -5508
rect 1030 -5519 1034 -5515
rect 1044 -5505 1048 -5501
rect 1218 -5505 1222 -5501
rect 1222 -5519 1226 -5515
rect 1238 -5497 1242 -5493
rect 1238 -5526 1242 -5522
rect 1252 -5505 1256 -5501
rect 1262 -5512 1266 -5508
rect 1276 -5497 1280 -5493
rect 1280 -5526 1284 -5522
rect 1304 -5505 1308 -5501
rect 1294 -5512 1298 -5508
rect 1318 -5526 1322 -5522
rect 1336 -5497 1340 -5493
rect 1346 -5512 1350 -5508
rect 1336 -5519 1340 -5515
rect 1360 -5497 1364 -5493
rect 1364 -5505 1368 -5501
rect 1378 -5512 1382 -5508
rect 1388 -5519 1392 -5515
rect 1402 -5505 1406 -5501
rect -1308 -5595 -1304 -5591
rect -1297 -5603 -1293 -5599
rect -1290 -5625 -1286 -5621
rect -934 -5595 -930 -5591
rect -923 -5603 -919 -5599
rect -916 -5625 -912 -5621
rect -576 -5595 -572 -5591
rect -565 -5603 -561 -5599
rect -558 -5625 -554 -5621
rect -218 -5595 -214 -5591
rect -207 -5603 -203 -5599
rect -200 -5625 -196 -5621
rect 140 -5595 144 -5591
rect 151 -5603 155 -5599
rect 158 -5625 162 -5621
rect 496 -5595 500 -5591
rect 507 -5603 511 -5599
rect 514 -5625 518 -5621
rect 854 -5595 858 -5591
rect 865 -5603 869 -5599
rect 872 -5625 876 -5621
rect 1212 -5595 1216 -5591
rect 1223 -5603 1227 -5599
rect 1230 -5625 1234 -5621
rect -1223 -5778 -1219 -5774
rect -1227 -5785 -1223 -5781
rect -1207 -5765 -1203 -5761
rect -1197 -5785 -1193 -5781
rect -1183 -5778 -1179 -5774
rect -1173 -5771 -1169 -5767
rect -1163 -5778 -1159 -5774
rect -1149 -5785 -1145 -5781
rect -1145 -5799 -1141 -5795
rect -924 -5741 -920 -5737
rect -928 -5762 -924 -5758
rect -924 -5777 -920 -5773
rect -928 -5791 -924 -5787
rect -898 -5762 -894 -5758
rect -902 -5770 -898 -5766
rect -902 -5784 -898 -5780
rect -882 -5748 -878 -5744
rect -872 -5791 -868 -5787
rect -858 -5741 -854 -5737
rect -848 -5755 -844 -5751
rect -838 -5791 -834 -5787
rect -824 -5741 -820 -5737
rect -820 -5799 -816 -5795
rect -804 -5770 -800 -5766
rect -794 -5784 -790 -5780
rect -780 -5741 -776 -5737
rect -780 -5762 -776 -5758
rect -776 -5777 -772 -5773
rect -760 -5784 -756 -5780
rect -746 -5741 -742 -5737
rect -736 -5792 -732 -5788
rect -720 -5799 -716 -5795
rect -706 -5755 -702 -5751
rect -702 -5792 -698 -5788
rect -566 -5741 -562 -5737
rect -570 -5762 -566 -5758
rect -566 -5777 -562 -5773
rect -570 -5791 -566 -5787
rect -540 -5762 -536 -5758
rect -544 -5770 -540 -5766
rect -544 -5784 -540 -5780
rect -524 -5748 -520 -5744
rect -514 -5791 -510 -5787
rect -500 -5741 -496 -5737
rect -490 -5755 -486 -5751
rect -480 -5791 -476 -5787
rect -466 -5741 -462 -5737
rect -462 -5799 -458 -5795
rect -446 -5770 -442 -5766
rect -436 -5784 -432 -5780
rect -422 -5741 -418 -5737
rect -422 -5762 -418 -5758
rect -418 -5777 -414 -5773
rect -402 -5784 -398 -5780
rect -388 -5741 -384 -5737
rect -378 -5792 -374 -5788
rect -362 -5799 -358 -5795
rect -348 -5755 -344 -5751
rect -344 -5792 -340 -5788
rect -208 -5741 -204 -5737
rect -212 -5762 -208 -5758
rect -208 -5777 -204 -5773
rect -212 -5791 -208 -5787
rect -182 -5762 -178 -5758
rect -186 -5770 -182 -5766
rect -186 -5784 -182 -5780
rect -166 -5748 -162 -5744
rect -156 -5791 -152 -5787
rect -142 -5741 -138 -5737
rect -132 -5755 -128 -5751
rect -122 -5791 -118 -5787
rect -108 -5741 -104 -5737
rect -104 -5799 -100 -5795
rect -88 -5770 -84 -5766
rect -78 -5784 -74 -5780
rect -64 -5741 -60 -5737
rect -64 -5762 -60 -5758
rect -60 -5777 -56 -5773
rect -44 -5784 -40 -5780
rect -30 -5741 -26 -5737
rect -20 -5792 -16 -5788
rect -4 -5799 0 -5795
rect 10 -5755 14 -5751
rect 14 -5792 18 -5788
rect 150 -5741 154 -5737
rect 146 -5762 150 -5758
rect 150 -5777 154 -5773
rect 146 -5791 150 -5787
rect 176 -5762 180 -5758
rect 172 -5770 176 -5766
rect 172 -5784 176 -5780
rect 192 -5748 196 -5744
rect 202 -5791 206 -5787
rect 216 -5741 220 -5737
rect 226 -5755 230 -5751
rect 236 -5791 240 -5787
rect 250 -5741 254 -5737
rect 254 -5799 258 -5795
rect 270 -5770 274 -5766
rect 280 -5784 284 -5780
rect 294 -5741 298 -5737
rect 294 -5762 298 -5758
rect 298 -5777 302 -5773
rect 314 -5784 318 -5780
rect 328 -5741 332 -5737
rect 338 -5792 342 -5788
rect 354 -5799 358 -5795
rect 368 -5755 372 -5751
rect 372 -5792 376 -5788
rect 506 -5741 510 -5737
rect 502 -5762 506 -5758
rect 506 -5777 510 -5773
rect 502 -5791 506 -5787
rect 532 -5762 536 -5758
rect 528 -5770 532 -5766
rect 528 -5784 532 -5780
rect 548 -5748 552 -5744
rect 558 -5791 562 -5787
rect 572 -5741 576 -5737
rect 582 -5755 586 -5751
rect 592 -5791 596 -5787
rect 606 -5741 610 -5737
rect 610 -5799 614 -5795
rect 626 -5770 630 -5766
rect 636 -5784 640 -5780
rect 650 -5741 654 -5737
rect 650 -5762 654 -5758
rect 654 -5777 658 -5773
rect 670 -5784 674 -5780
rect 684 -5741 688 -5737
rect 694 -5792 698 -5788
rect 710 -5799 714 -5795
rect 724 -5755 728 -5751
rect 728 -5792 732 -5788
rect 864 -5741 868 -5737
rect 860 -5762 864 -5758
rect 864 -5777 868 -5773
rect 860 -5791 864 -5787
rect 890 -5762 894 -5758
rect 886 -5770 890 -5766
rect 886 -5784 890 -5780
rect 906 -5748 910 -5744
rect 916 -5791 920 -5787
rect 930 -5741 934 -5737
rect 940 -5755 944 -5751
rect 950 -5791 954 -5787
rect 964 -5741 968 -5737
rect 968 -5799 972 -5795
rect 984 -5770 988 -5766
rect 994 -5784 998 -5780
rect 1008 -5741 1012 -5737
rect 1008 -5762 1012 -5758
rect 1012 -5777 1016 -5773
rect 1028 -5784 1032 -5780
rect 1042 -5741 1046 -5737
rect 1052 -5792 1056 -5788
rect 1068 -5799 1072 -5795
rect 1082 -5755 1086 -5751
rect 1086 -5792 1090 -5788
rect 1222 -5741 1226 -5737
rect 1218 -5762 1222 -5758
rect 1222 -5777 1226 -5773
rect 1218 -5791 1222 -5787
rect 1248 -5762 1252 -5758
rect 1244 -5770 1248 -5766
rect 1244 -5784 1248 -5780
rect 1264 -5748 1268 -5744
rect 1274 -5791 1278 -5787
rect 1288 -5741 1292 -5737
rect 1298 -5755 1302 -5751
rect 1308 -5791 1312 -5787
rect 1322 -5741 1326 -5737
rect 1326 -5799 1330 -5795
rect 1342 -5770 1346 -5766
rect 1352 -5784 1356 -5780
rect 1366 -5741 1370 -5737
rect 1366 -5762 1370 -5758
rect 1370 -5777 1374 -5773
rect 1386 -5784 1390 -5780
rect 1400 -5741 1404 -5737
rect 1410 -5792 1414 -5788
rect 1426 -5799 1430 -5795
rect 1440 -5755 1444 -5751
rect 1444 -5792 1448 -5788
rect -1227 -5901 -1223 -5897
rect -1223 -5915 -1219 -5911
rect -1207 -5893 -1203 -5889
rect -1207 -5922 -1203 -5918
rect -1193 -5901 -1189 -5897
rect -1183 -5908 -1179 -5904
rect -1169 -5893 -1165 -5889
rect -1165 -5922 -1161 -5918
rect -1141 -5901 -1137 -5897
rect -1151 -5908 -1147 -5904
rect -1127 -5922 -1123 -5918
rect -1109 -5893 -1105 -5889
rect -1099 -5908 -1095 -5904
rect -1109 -5915 -1105 -5911
rect -1085 -5893 -1081 -5889
rect -1081 -5901 -1077 -5897
rect -1067 -5908 -1063 -5904
rect -1057 -5915 -1053 -5911
rect -1043 -5901 -1039 -5897
rect -928 -5901 -924 -5897
rect -924 -5915 -920 -5911
rect -908 -5893 -904 -5889
rect -908 -5922 -904 -5918
rect -894 -5901 -890 -5897
rect -884 -5908 -880 -5904
rect -870 -5893 -866 -5889
rect -866 -5922 -862 -5918
rect -842 -5901 -838 -5897
rect -852 -5908 -848 -5904
rect -828 -5922 -824 -5918
rect -810 -5893 -806 -5889
rect -800 -5908 -796 -5904
rect -810 -5915 -806 -5911
rect -786 -5893 -782 -5889
rect -782 -5901 -778 -5897
rect -768 -5908 -764 -5904
rect -758 -5915 -754 -5911
rect -744 -5901 -740 -5897
rect -570 -5901 -566 -5897
rect -566 -5915 -562 -5911
rect -550 -5893 -546 -5889
rect -550 -5922 -546 -5918
rect -536 -5901 -532 -5897
rect -526 -5908 -522 -5904
rect -512 -5893 -508 -5889
rect -508 -5922 -504 -5918
rect -484 -5901 -480 -5897
rect -494 -5908 -490 -5904
rect -470 -5922 -466 -5918
rect -452 -5893 -448 -5889
rect -442 -5908 -438 -5904
rect -452 -5915 -448 -5911
rect -428 -5893 -424 -5889
rect -424 -5901 -420 -5897
rect -410 -5908 -406 -5904
rect -400 -5915 -396 -5911
rect -386 -5901 -382 -5897
rect -212 -5901 -208 -5897
rect -208 -5915 -204 -5911
rect -192 -5893 -188 -5889
rect -192 -5922 -188 -5918
rect -178 -5901 -174 -5897
rect -168 -5908 -164 -5904
rect -154 -5893 -150 -5889
rect -150 -5922 -146 -5918
rect -126 -5901 -122 -5897
rect -136 -5908 -132 -5904
rect -112 -5922 -108 -5918
rect -94 -5893 -90 -5889
rect -84 -5908 -80 -5904
rect -94 -5915 -90 -5911
rect -70 -5893 -66 -5889
rect -66 -5901 -62 -5897
rect -52 -5908 -48 -5904
rect -42 -5915 -38 -5911
rect -28 -5901 -24 -5897
rect 146 -5901 150 -5897
rect 150 -5915 154 -5911
rect 166 -5893 170 -5889
rect 166 -5922 170 -5918
rect 180 -5901 184 -5897
rect 190 -5908 194 -5904
rect 204 -5893 208 -5889
rect 208 -5922 212 -5918
rect 232 -5901 236 -5897
rect 222 -5908 226 -5904
rect 246 -5922 250 -5918
rect 264 -5893 268 -5889
rect 274 -5908 278 -5904
rect 264 -5915 268 -5911
rect 288 -5893 292 -5889
rect 292 -5901 296 -5897
rect 306 -5908 310 -5904
rect 316 -5915 320 -5911
rect 330 -5901 334 -5897
rect 502 -5901 506 -5897
rect 506 -5915 510 -5911
rect 522 -5893 526 -5889
rect 522 -5922 526 -5918
rect 536 -5901 540 -5897
rect 546 -5908 550 -5904
rect 560 -5893 564 -5889
rect 564 -5922 568 -5918
rect 588 -5901 592 -5897
rect 578 -5908 582 -5904
rect 602 -5922 606 -5918
rect 620 -5893 624 -5889
rect 630 -5908 634 -5904
rect 620 -5915 624 -5911
rect 644 -5893 648 -5889
rect 648 -5901 652 -5897
rect 662 -5908 666 -5904
rect 672 -5915 676 -5911
rect 686 -5901 690 -5897
rect 860 -5901 864 -5897
rect 864 -5915 868 -5911
rect 880 -5893 884 -5889
rect 880 -5922 884 -5918
rect 894 -5901 898 -5897
rect 904 -5908 908 -5904
rect 918 -5893 922 -5889
rect 922 -5922 926 -5918
rect 946 -5901 950 -5897
rect 936 -5908 940 -5904
rect 960 -5922 964 -5918
rect 978 -5893 982 -5889
rect 988 -5908 992 -5904
rect 978 -5915 982 -5911
rect 1002 -5893 1006 -5889
rect 1006 -5901 1010 -5897
rect 1020 -5908 1024 -5904
rect 1030 -5915 1034 -5911
rect 1044 -5901 1048 -5897
rect 1218 -5901 1222 -5897
rect 1222 -5915 1226 -5911
rect 1238 -5893 1242 -5889
rect 1238 -5922 1242 -5918
rect 1252 -5901 1256 -5897
rect 1262 -5908 1266 -5904
rect 1276 -5893 1280 -5889
rect 1280 -5922 1284 -5918
rect 1304 -5901 1308 -5897
rect 1294 -5908 1298 -5904
rect 1318 -5922 1322 -5918
rect 1336 -5893 1340 -5889
rect 1346 -5908 1350 -5904
rect 1336 -5915 1340 -5911
rect 1360 -5893 1364 -5889
rect 1364 -5901 1368 -5897
rect 1378 -5908 1382 -5904
rect 1388 -5915 1392 -5911
rect 1402 -5901 1406 -5897
rect 1562 -5901 1566 -5897
rect 1566 -5915 1570 -5911
rect 1582 -5893 1586 -5889
rect 1582 -5922 1586 -5918
rect 1596 -5901 1600 -5897
rect 1606 -5908 1610 -5904
rect 1620 -5893 1624 -5889
rect 1624 -5922 1628 -5918
rect 1648 -5901 1652 -5897
rect 1638 -5908 1642 -5904
rect 1662 -5922 1666 -5918
rect 1680 -5893 1684 -5889
rect 1690 -5908 1694 -5904
rect 1680 -5915 1684 -5911
rect 1704 -5893 1708 -5889
rect 1708 -5901 1712 -5897
rect 1722 -5908 1726 -5904
rect 1732 -5915 1736 -5911
rect 1746 -5901 1750 -5897
<< ndcontact >>
rect -1307 -868 -1303 -864
rect -1290 -868 -1286 -864
rect -1281 -868 -1277 -864
rect -936 -868 -932 -864
rect -919 -868 -915 -864
rect -910 -868 -906 -864
rect -577 -868 -573 -864
rect -560 -868 -556 -864
rect -551 -868 -547 -864
rect -219 -868 -215 -864
rect -202 -868 -198 -864
rect -193 -868 -189 -864
rect 138 -868 142 -864
rect 155 -868 159 -864
rect 164 -868 168 -864
rect 495 -868 499 -864
rect 512 -868 516 -864
rect 521 -868 525 -864
rect 853 -868 857 -864
rect 870 -868 874 -864
rect 879 -868 883 -864
rect 1211 -868 1215 -864
rect 1228 -868 1232 -864
rect 1237 -868 1241 -864
rect -1230 -1102 -1226 -1098
rect -1221 -1102 -1217 -1098
rect -1212 -1102 -1208 -1098
rect -1204 -1102 -1200 -1098
rect -1188 -1102 -1184 -1098
rect -1180 -1102 -1176 -1098
rect -1163 -1102 -1159 -1098
rect -1146 -1102 -1142 -1098
rect -1138 -1102 -1134 -1098
rect -1121 -1102 -1117 -1098
rect -1104 -1102 -1100 -1098
rect -1096 -1102 -1092 -1098
rect -1079 -1102 -1075 -1098
rect -1062 -1102 -1058 -1098
rect -1054 -1102 -1050 -1098
rect -1038 -1102 -1034 -1098
rect -935 -1102 -931 -1098
rect -926 -1102 -922 -1098
rect -917 -1102 -913 -1098
rect -909 -1102 -905 -1098
rect -893 -1102 -889 -1098
rect -885 -1102 -881 -1098
rect -868 -1102 -864 -1098
rect -851 -1102 -847 -1098
rect -843 -1102 -839 -1098
rect -826 -1102 -822 -1098
rect -809 -1102 -805 -1098
rect -801 -1102 -797 -1098
rect -784 -1102 -780 -1098
rect -767 -1102 -763 -1098
rect -759 -1102 -755 -1098
rect -743 -1102 -739 -1098
rect -577 -1102 -573 -1098
rect -568 -1102 -564 -1098
rect -559 -1102 -555 -1098
rect -551 -1102 -547 -1098
rect -535 -1102 -531 -1098
rect -527 -1102 -523 -1098
rect -510 -1102 -506 -1098
rect -493 -1102 -489 -1098
rect -485 -1102 -481 -1098
rect -468 -1102 -464 -1098
rect -451 -1102 -447 -1098
rect -443 -1102 -439 -1098
rect -426 -1102 -422 -1098
rect -409 -1102 -405 -1098
rect -401 -1102 -397 -1098
rect -385 -1102 -381 -1098
rect -219 -1102 -215 -1098
rect -210 -1102 -206 -1098
rect -201 -1102 -197 -1098
rect -193 -1102 -189 -1098
rect -177 -1102 -173 -1098
rect -169 -1102 -165 -1098
rect -152 -1102 -148 -1098
rect -135 -1102 -131 -1098
rect -127 -1102 -123 -1098
rect -110 -1102 -106 -1098
rect -93 -1102 -89 -1098
rect -85 -1102 -81 -1098
rect -68 -1102 -64 -1098
rect -51 -1102 -47 -1098
rect -43 -1102 -39 -1098
rect -27 -1102 -23 -1098
rect 139 -1102 143 -1098
rect 148 -1102 152 -1098
rect 157 -1102 161 -1098
rect 165 -1102 169 -1098
rect 181 -1102 185 -1098
rect 189 -1102 193 -1098
rect 206 -1102 210 -1098
rect 223 -1102 227 -1098
rect 231 -1102 235 -1098
rect 248 -1102 252 -1098
rect 265 -1102 269 -1098
rect 273 -1102 277 -1098
rect 290 -1102 294 -1098
rect 307 -1102 311 -1098
rect 315 -1102 319 -1098
rect 331 -1102 335 -1098
rect 495 -1102 499 -1098
rect 504 -1102 508 -1098
rect 513 -1102 517 -1098
rect 521 -1102 525 -1098
rect 537 -1102 541 -1098
rect 545 -1102 549 -1098
rect 562 -1102 566 -1098
rect 579 -1102 583 -1098
rect 587 -1102 591 -1098
rect 604 -1102 608 -1098
rect 621 -1102 625 -1098
rect 629 -1102 633 -1098
rect 646 -1102 650 -1098
rect 663 -1102 667 -1098
rect 671 -1102 675 -1098
rect 687 -1102 691 -1098
rect 853 -1102 857 -1098
rect 862 -1102 866 -1098
rect 871 -1102 875 -1098
rect 879 -1102 883 -1098
rect 895 -1102 899 -1098
rect 903 -1102 907 -1098
rect 920 -1102 924 -1098
rect 937 -1102 941 -1098
rect 945 -1102 949 -1098
rect 962 -1102 966 -1098
rect 979 -1102 983 -1098
rect 987 -1102 991 -1098
rect 1004 -1102 1008 -1098
rect 1021 -1102 1025 -1098
rect 1029 -1102 1033 -1098
rect 1045 -1102 1049 -1098
rect -1309 -1218 -1305 -1214
rect -1292 -1218 -1288 -1214
rect -1283 -1218 -1279 -1214
rect -935 -1218 -931 -1214
rect -918 -1218 -914 -1214
rect -909 -1218 -905 -1214
rect -577 -1218 -573 -1214
rect -560 -1218 -556 -1214
rect -551 -1218 -547 -1214
rect -219 -1218 -215 -1214
rect -202 -1218 -198 -1214
rect -193 -1218 -189 -1214
rect 139 -1218 143 -1214
rect 156 -1218 160 -1214
rect 165 -1218 169 -1214
rect 495 -1218 499 -1214
rect 512 -1218 516 -1214
rect 521 -1218 525 -1214
rect 853 -1218 857 -1214
rect 870 -1218 874 -1214
rect 879 -1218 883 -1214
rect 1211 -1218 1215 -1214
rect 1228 -1218 1232 -1214
rect 1237 -1218 1241 -1214
rect -1230 -1382 -1226 -1378
rect -1221 -1382 -1217 -1378
rect -1212 -1382 -1208 -1378
rect -1204 -1382 -1200 -1378
rect -1195 -1382 -1191 -1378
rect -1177 -1382 -1173 -1378
rect -1168 -1382 -1164 -1378
rect -1160 -1382 -1156 -1378
rect -1143 -1382 -1139 -1378
rect -1134 -1382 -1130 -1378
rect -935 -1382 -931 -1378
rect -926 -1382 -922 -1378
rect -917 -1382 -913 -1378
rect -909 -1382 -905 -1378
rect -900 -1382 -896 -1378
rect -891 -1382 -887 -1378
rect -883 -1382 -879 -1378
rect -875 -1382 -871 -1378
rect -857 -1382 -853 -1378
rect -847 -1382 -843 -1378
rect -839 -1382 -835 -1378
rect -822 -1382 -818 -1378
rect -813 -1382 -809 -1378
rect -805 -1382 -801 -1378
rect -796 -1382 -792 -1378
rect -778 -1382 -774 -1378
rect -769 -1382 -765 -1378
rect -761 -1382 -757 -1378
rect -745 -1382 -741 -1378
rect -737 -1382 -733 -1378
rect -725 -1382 -721 -1378
rect -713 -1382 -709 -1378
rect -704 -1382 -700 -1378
rect -695 -1382 -691 -1378
rect -577 -1382 -573 -1378
rect -568 -1382 -564 -1378
rect -559 -1382 -555 -1378
rect -551 -1382 -547 -1378
rect -542 -1382 -538 -1378
rect -533 -1382 -529 -1378
rect -525 -1382 -521 -1378
rect -517 -1382 -513 -1378
rect -499 -1382 -495 -1378
rect -489 -1382 -485 -1378
rect -481 -1382 -477 -1378
rect -464 -1382 -460 -1378
rect -455 -1382 -451 -1378
rect -447 -1382 -443 -1378
rect -438 -1382 -434 -1378
rect -420 -1382 -416 -1378
rect -411 -1382 -407 -1378
rect -403 -1382 -399 -1378
rect -387 -1382 -383 -1378
rect -379 -1382 -375 -1378
rect -367 -1382 -363 -1378
rect -355 -1382 -351 -1378
rect -346 -1382 -342 -1378
rect -337 -1382 -333 -1378
rect -219 -1382 -215 -1378
rect -210 -1382 -206 -1378
rect -201 -1382 -197 -1378
rect -193 -1382 -189 -1378
rect -184 -1382 -180 -1378
rect -175 -1382 -171 -1378
rect -167 -1382 -163 -1378
rect -159 -1382 -155 -1378
rect -141 -1382 -137 -1378
rect -131 -1382 -127 -1378
rect -123 -1382 -119 -1378
rect -106 -1382 -102 -1378
rect -97 -1382 -93 -1378
rect -89 -1382 -85 -1378
rect -80 -1382 -76 -1378
rect -62 -1382 -58 -1378
rect -53 -1382 -49 -1378
rect -45 -1382 -41 -1378
rect -29 -1382 -25 -1378
rect -21 -1382 -17 -1378
rect -9 -1382 -5 -1378
rect 3 -1382 7 -1378
rect 12 -1382 16 -1378
rect 21 -1382 25 -1378
rect 139 -1382 143 -1378
rect 148 -1382 152 -1378
rect 157 -1382 161 -1378
rect 165 -1382 169 -1378
rect 174 -1382 178 -1378
rect 183 -1382 187 -1378
rect 191 -1382 195 -1378
rect 199 -1382 203 -1378
rect 217 -1382 221 -1378
rect 227 -1382 231 -1378
rect 235 -1382 239 -1378
rect 252 -1382 256 -1378
rect 261 -1382 265 -1378
rect 269 -1382 273 -1378
rect 278 -1382 282 -1378
rect 296 -1382 300 -1378
rect 305 -1382 309 -1378
rect 313 -1382 317 -1378
rect 329 -1382 333 -1378
rect 337 -1382 341 -1378
rect 349 -1382 353 -1378
rect 361 -1382 365 -1378
rect 370 -1382 374 -1378
rect 379 -1382 383 -1378
rect 495 -1382 499 -1378
rect 504 -1382 508 -1378
rect 513 -1382 517 -1378
rect 521 -1382 525 -1378
rect 530 -1382 534 -1378
rect 539 -1382 543 -1378
rect 547 -1382 551 -1378
rect 555 -1382 559 -1378
rect 573 -1382 577 -1378
rect 583 -1382 587 -1378
rect 591 -1382 595 -1378
rect 608 -1382 612 -1378
rect 617 -1382 621 -1378
rect 625 -1382 629 -1378
rect 634 -1382 638 -1378
rect 652 -1382 656 -1378
rect 661 -1382 665 -1378
rect 669 -1382 673 -1378
rect 685 -1382 689 -1378
rect 693 -1382 697 -1378
rect 705 -1382 709 -1378
rect 717 -1382 721 -1378
rect 726 -1382 730 -1378
rect 735 -1382 739 -1378
rect 853 -1382 857 -1378
rect 862 -1382 866 -1378
rect 871 -1382 875 -1378
rect 879 -1382 883 -1378
rect 888 -1382 892 -1378
rect 897 -1382 901 -1378
rect 905 -1382 909 -1378
rect 913 -1382 917 -1378
rect 931 -1382 935 -1378
rect 941 -1382 945 -1378
rect 949 -1382 953 -1378
rect 966 -1382 970 -1378
rect 975 -1382 979 -1378
rect 983 -1382 987 -1378
rect 992 -1382 996 -1378
rect 1010 -1382 1014 -1378
rect 1019 -1382 1023 -1378
rect 1027 -1382 1031 -1378
rect 1043 -1382 1047 -1378
rect 1051 -1382 1055 -1378
rect 1063 -1382 1067 -1378
rect 1075 -1382 1079 -1378
rect 1084 -1382 1088 -1378
rect 1093 -1382 1097 -1378
rect 1211 -1382 1215 -1378
rect 1220 -1382 1224 -1378
rect 1229 -1382 1233 -1378
rect 1237 -1382 1241 -1378
rect 1246 -1382 1250 -1378
rect 1264 -1382 1268 -1378
rect 1273 -1382 1277 -1378
rect 1281 -1382 1285 -1378
rect 1298 -1382 1302 -1378
rect 1307 -1382 1311 -1378
rect -1230 -1505 -1226 -1501
rect -1221 -1505 -1217 -1501
rect -1212 -1505 -1208 -1501
rect -1204 -1505 -1200 -1501
rect -1188 -1505 -1184 -1501
rect -1180 -1505 -1176 -1501
rect -1163 -1505 -1159 -1501
rect -1146 -1505 -1142 -1501
rect -1138 -1505 -1134 -1501
rect -1121 -1505 -1117 -1501
rect -1104 -1505 -1100 -1501
rect -1096 -1505 -1092 -1501
rect -1079 -1505 -1075 -1501
rect -1062 -1505 -1058 -1501
rect -1054 -1505 -1050 -1501
rect -1038 -1505 -1034 -1501
rect -935 -1505 -931 -1501
rect -926 -1505 -922 -1501
rect -917 -1505 -913 -1501
rect -909 -1505 -905 -1501
rect -893 -1505 -889 -1501
rect -885 -1505 -881 -1501
rect -868 -1505 -864 -1501
rect -851 -1505 -847 -1501
rect -843 -1505 -839 -1501
rect -826 -1505 -822 -1501
rect -809 -1505 -805 -1501
rect -801 -1505 -797 -1501
rect -784 -1505 -780 -1501
rect -767 -1505 -763 -1501
rect -759 -1505 -755 -1501
rect -743 -1505 -739 -1501
rect -577 -1505 -573 -1501
rect -568 -1505 -564 -1501
rect -559 -1505 -555 -1501
rect -551 -1505 -547 -1501
rect -535 -1505 -531 -1501
rect -527 -1505 -523 -1501
rect -510 -1505 -506 -1501
rect -493 -1505 -489 -1501
rect -485 -1505 -481 -1501
rect -468 -1505 -464 -1501
rect -451 -1505 -447 -1501
rect -443 -1505 -439 -1501
rect -426 -1505 -422 -1501
rect -409 -1505 -405 -1501
rect -401 -1505 -397 -1501
rect -385 -1505 -381 -1501
rect -219 -1505 -215 -1501
rect -210 -1505 -206 -1501
rect -201 -1505 -197 -1501
rect -193 -1505 -189 -1501
rect -177 -1505 -173 -1501
rect -169 -1505 -165 -1501
rect -152 -1505 -148 -1501
rect -135 -1505 -131 -1501
rect -127 -1505 -123 -1501
rect -110 -1505 -106 -1501
rect -93 -1505 -89 -1501
rect -85 -1505 -81 -1501
rect -68 -1505 -64 -1501
rect -51 -1505 -47 -1501
rect -43 -1505 -39 -1501
rect -27 -1505 -23 -1501
rect 139 -1505 143 -1501
rect 148 -1505 152 -1501
rect 157 -1505 161 -1501
rect 165 -1505 169 -1501
rect 181 -1505 185 -1501
rect 189 -1505 193 -1501
rect 206 -1505 210 -1501
rect 223 -1505 227 -1501
rect 231 -1505 235 -1501
rect 248 -1505 252 -1501
rect 265 -1505 269 -1501
rect 273 -1505 277 -1501
rect 290 -1505 294 -1501
rect 307 -1505 311 -1501
rect 315 -1505 319 -1501
rect 331 -1505 335 -1501
rect 495 -1505 499 -1501
rect 504 -1505 508 -1501
rect 513 -1505 517 -1501
rect 521 -1505 525 -1501
rect 537 -1505 541 -1501
rect 545 -1505 549 -1501
rect 562 -1505 566 -1501
rect 579 -1505 583 -1501
rect 587 -1505 591 -1501
rect 604 -1505 608 -1501
rect 621 -1505 625 -1501
rect 629 -1505 633 -1501
rect 646 -1505 650 -1501
rect 663 -1505 667 -1501
rect 671 -1505 675 -1501
rect 687 -1505 691 -1501
rect 853 -1505 857 -1501
rect 862 -1505 866 -1501
rect 871 -1505 875 -1501
rect 879 -1505 883 -1501
rect 895 -1505 899 -1501
rect 903 -1505 907 -1501
rect 920 -1505 924 -1501
rect 937 -1505 941 -1501
rect 945 -1505 949 -1501
rect 962 -1505 966 -1501
rect 979 -1505 983 -1501
rect 987 -1505 991 -1501
rect 1004 -1505 1008 -1501
rect 1021 -1505 1025 -1501
rect 1029 -1505 1033 -1501
rect 1045 -1505 1049 -1501
rect -1230 -1676 -1226 -1672
rect -1221 -1676 -1217 -1672
rect -1212 -1676 -1208 -1672
rect -1204 -1676 -1200 -1672
rect -1188 -1676 -1184 -1672
rect -1180 -1676 -1176 -1672
rect -1163 -1676 -1159 -1672
rect -1146 -1676 -1142 -1672
rect -1138 -1676 -1134 -1672
rect -1121 -1676 -1117 -1672
rect -1104 -1676 -1100 -1672
rect -1096 -1676 -1092 -1672
rect -1079 -1676 -1075 -1672
rect -1062 -1676 -1058 -1672
rect -1054 -1676 -1050 -1672
rect -1038 -1676 -1034 -1672
rect -935 -1676 -931 -1672
rect -926 -1676 -922 -1672
rect -917 -1676 -913 -1672
rect -909 -1676 -905 -1672
rect -893 -1676 -889 -1672
rect -885 -1676 -881 -1672
rect -868 -1676 -864 -1672
rect -851 -1676 -847 -1672
rect -843 -1676 -839 -1672
rect -826 -1676 -822 -1672
rect -809 -1676 -805 -1672
rect -801 -1676 -797 -1672
rect -784 -1676 -780 -1672
rect -767 -1676 -763 -1672
rect -759 -1676 -755 -1672
rect -743 -1676 -739 -1672
rect -577 -1676 -573 -1672
rect -568 -1676 -564 -1672
rect -559 -1676 -555 -1672
rect -551 -1676 -547 -1672
rect -535 -1676 -531 -1672
rect -527 -1676 -523 -1672
rect -510 -1676 -506 -1672
rect -493 -1676 -489 -1672
rect -485 -1676 -481 -1672
rect -468 -1676 -464 -1672
rect -451 -1676 -447 -1672
rect -443 -1676 -439 -1672
rect -426 -1676 -422 -1672
rect -409 -1676 -405 -1672
rect -401 -1676 -397 -1672
rect -385 -1676 -381 -1672
rect -219 -1676 -215 -1672
rect -210 -1676 -206 -1672
rect -201 -1676 -197 -1672
rect -193 -1676 -189 -1672
rect -177 -1676 -173 -1672
rect -169 -1676 -165 -1672
rect -152 -1676 -148 -1672
rect -135 -1676 -131 -1672
rect -127 -1676 -123 -1672
rect -110 -1676 -106 -1672
rect -93 -1676 -89 -1672
rect -85 -1676 -81 -1672
rect -68 -1676 -64 -1672
rect -51 -1676 -47 -1672
rect -43 -1676 -39 -1672
rect -27 -1676 -23 -1672
rect 139 -1676 143 -1672
rect 148 -1676 152 -1672
rect 157 -1676 161 -1672
rect 165 -1676 169 -1672
rect 181 -1676 185 -1672
rect 189 -1676 193 -1672
rect 206 -1676 210 -1672
rect 223 -1676 227 -1672
rect 231 -1676 235 -1672
rect 248 -1676 252 -1672
rect 265 -1676 269 -1672
rect 273 -1676 277 -1672
rect 290 -1676 294 -1672
rect 307 -1676 311 -1672
rect 315 -1676 319 -1672
rect 331 -1676 335 -1672
rect 495 -1676 499 -1672
rect 504 -1676 508 -1672
rect 513 -1676 517 -1672
rect 521 -1676 525 -1672
rect 537 -1676 541 -1672
rect 545 -1676 549 -1672
rect 562 -1676 566 -1672
rect 579 -1676 583 -1672
rect 587 -1676 591 -1672
rect 604 -1676 608 -1672
rect 621 -1676 625 -1672
rect 629 -1676 633 -1672
rect 646 -1676 650 -1672
rect 663 -1676 667 -1672
rect 671 -1676 675 -1672
rect 687 -1676 691 -1672
rect 853 -1676 857 -1672
rect 862 -1676 866 -1672
rect 871 -1676 875 -1672
rect 879 -1676 883 -1672
rect 895 -1676 899 -1672
rect 903 -1676 907 -1672
rect 920 -1676 924 -1672
rect 937 -1676 941 -1672
rect 945 -1676 949 -1672
rect 962 -1676 966 -1672
rect 979 -1676 983 -1672
rect 987 -1676 991 -1672
rect 1004 -1676 1008 -1672
rect 1021 -1676 1025 -1672
rect 1029 -1676 1033 -1672
rect 1045 -1676 1049 -1672
rect 1211 -1676 1215 -1672
rect 1220 -1676 1224 -1672
rect 1229 -1676 1233 -1672
rect 1237 -1676 1241 -1672
rect 1253 -1676 1257 -1672
rect 1261 -1676 1265 -1672
rect 1278 -1676 1282 -1672
rect 1295 -1676 1299 -1672
rect 1303 -1676 1307 -1672
rect 1320 -1676 1324 -1672
rect 1337 -1676 1341 -1672
rect 1345 -1676 1349 -1672
rect 1362 -1676 1366 -1672
rect 1379 -1676 1383 -1672
rect 1387 -1676 1391 -1672
rect 1403 -1676 1407 -1672
rect -1559 -1847 -1555 -1843
rect -1550 -1847 -1546 -1843
rect -1541 -1847 -1537 -1843
rect -1533 -1847 -1529 -1843
rect -1517 -1847 -1513 -1843
rect -1509 -1847 -1505 -1843
rect -1492 -1847 -1488 -1843
rect -1475 -1847 -1471 -1843
rect -1467 -1847 -1463 -1843
rect -1450 -1847 -1446 -1843
rect -1433 -1847 -1429 -1843
rect -1425 -1847 -1421 -1843
rect -1408 -1847 -1404 -1843
rect -1391 -1847 -1387 -1843
rect -1383 -1847 -1379 -1843
rect -1367 -1847 -1363 -1843
rect -1230 -1847 -1226 -1843
rect -1221 -1847 -1217 -1843
rect -1212 -1847 -1208 -1843
rect -1204 -1847 -1200 -1843
rect -1188 -1847 -1184 -1843
rect -1180 -1847 -1176 -1843
rect -1163 -1847 -1159 -1843
rect -1146 -1847 -1142 -1843
rect -1138 -1847 -1134 -1843
rect -1121 -1847 -1117 -1843
rect -1104 -1847 -1100 -1843
rect -1096 -1847 -1092 -1843
rect -1079 -1847 -1075 -1843
rect -1062 -1847 -1058 -1843
rect -1054 -1847 -1050 -1843
rect -1038 -1847 -1034 -1843
rect -935 -1847 -931 -1843
rect -926 -1847 -922 -1843
rect -917 -1847 -913 -1843
rect -909 -1847 -905 -1843
rect -893 -1847 -889 -1843
rect -885 -1847 -881 -1843
rect -868 -1847 -864 -1843
rect -851 -1847 -847 -1843
rect -843 -1847 -839 -1843
rect -826 -1847 -822 -1843
rect -809 -1847 -805 -1843
rect -801 -1847 -797 -1843
rect -784 -1847 -780 -1843
rect -767 -1847 -763 -1843
rect -759 -1847 -755 -1843
rect -743 -1847 -739 -1843
rect -577 -1847 -573 -1843
rect -568 -1847 -564 -1843
rect -559 -1847 -555 -1843
rect -551 -1847 -547 -1843
rect -535 -1847 -531 -1843
rect -527 -1847 -523 -1843
rect -510 -1847 -506 -1843
rect -493 -1847 -489 -1843
rect -485 -1847 -481 -1843
rect -468 -1847 -464 -1843
rect -451 -1847 -447 -1843
rect -443 -1847 -439 -1843
rect -426 -1847 -422 -1843
rect -409 -1847 -405 -1843
rect -401 -1847 -397 -1843
rect -385 -1847 -381 -1843
rect -219 -1847 -215 -1843
rect -210 -1847 -206 -1843
rect -201 -1847 -197 -1843
rect -193 -1847 -189 -1843
rect -177 -1847 -173 -1843
rect -169 -1847 -165 -1843
rect -152 -1847 -148 -1843
rect -135 -1847 -131 -1843
rect -127 -1847 -123 -1843
rect -110 -1847 -106 -1843
rect -93 -1847 -89 -1843
rect -85 -1847 -81 -1843
rect -68 -1847 -64 -1843
rect -51 -1847 -47 -1843
rect -43 -1847 -39 -1843
rect -27 -1847 -23 -1843
rect 139 -1847 143 -1843
rect 148 -1847 152 -1843
rect 157 -1847 161 -1843
rect 165 -1847 169 -1843
rect 181 -1847 185 -1843
rect 189 -1847 193 -1843
rect 206 -1847 210 -1843
rect 223 -1847 227 -1843
rect 231 -1847 235 -1843
rect 248 -1847 252 -1843
rect 265 -1847 269 -1843
rect 273 -1847 277 -1843
rect 290 -1847 294 -1843
rect 307 -1847 311 -1843
rect 315 -1847 319 -1843
rect 331 -1847 335 -1843
rect 495 -1847 499 -1843
rect 504 -1847 508 -1843
rect 513 -1847 517 -1843
rect 521 -1847 525 -1843
rect 537 -1847 541 -1843
rect 545 -1847 549 -1843
rect 562 -1847 566 -1843
rect 579 -1847 583 -1843
rect 587 -1847 591 -1843
rect 604 -1847 608 -1843
rect 621 -1847 625 -1843
rect 629 -1847 633 -1843
rect 646 -1847 650 -1843
rect 663 -1847 667 -1843
rect 671 -1847 675 -1843
rect 687 -1847 691 -1843
rect 853 -1847 857 -1843
rect 862 -1847 866 -1843
rect 871 -1847 875 -1843
rect 879 -1847 883 -1843
rect 895 -1847 899 -1843
rect 903 -1847 907 -1843
rect 920 -1847 924 -1843
rect 937 -1847 941 -1843
rect 945 -1847 949 -1843
rect 962 -1847 966 -1843
rect 979 -1847 983 -1843
rect 987 -1847 991 -1843
rect 1004 -1847 1008 -1843
rect 1021 -1847 1025 -1843
rect 1029 -1847 1033 -1843
rect 1045 -1847 1049 -1843
rect 1211 -1847 1215 -1843
rect 1220 -1847 1224 -1843
rect 1229 -1847 1233 -1843
rect 1237 -1847 1241 -1843
rect 1253 -1847 1257 -1843
rect 1261 -1847 1265 -1843
rect 1278 -1847 1282 -1843
rect 1295 -1847 1299 -1843
rect 1303 -1847 1307 -1843
rect 1320 -1847 1324 -1843
rect 1337 -1847 1341 -1843
rect 1345 -1847 1349 -1843
rect 1362 -1847 1366 -1843
rect 1379 -1847 1383 -1843
rect 1387 -1847 1391 -1843
rect 1403 -1847 1407 -1843
rect -1309 -1954 -1305 -1950
rect -1292 -1954 -1288 -1950
rect -1283 -1954 -1279 -1950
rect -935 -1954 -931 -1950
rect -918 -1954 -914 -1950
rect -909 -1954 -905 -1950
rect -577 -1954 -573 -1950
rect -560 -1954 -556 -1950
rect -551 -1954 -547 -1950
rect -219 -1954 -215 -1950
rect -202 -1954 -198 -1950
rect -193 -1954 -189 -1950
rect 139 -1954 143 -1950
rect 156 -1954 160 -1950
rect 165 -1954 169 -1950
rect 495 -1954 499 -1950
rect 512 -1954 516 -1950
rect 521 -1954 525 -1950
rect 853 -1954 857 -1950
rect 870 -1954 874 -1950
rect 879 -1954 883 -1950
rect 1211 -1954 1215 -1950
rect 1228 -1954 1232 -1950
rect 1237 -1954 1241 -1950
rect -1234 -2113 -1230 -2109
rect -1225 -2113 -1221 -2109
rect -1216 -2113 -1212 -2109
rect -1208 -2113 -1204 -2109
rect -1199 -2113 -1195 -2109
rect -1181 -2113 -1177 -2109
rect -1172 -2113 -1168 -2109
rect -1164 -2113 -1160 -2109
rect -1147 -2113 -1143 -2109
rect -1138 -2113 -1134 -2109
rect -935 -2113 -931 -2109
rect -926 -2113 -922 -2109
rect -917 -2113 -913 -2109
rect -909 -2113 -905 -2109
rect -900 -2113 -896 -2109
rect -891 -2113 -887 -2109
rect -883 -2113 -879 -2109
rect -875 -2113 -871 -2109
rect -857 -2113 -853 -2109
rect -847 -2113 -843 -2109
rect -839 -2113 -835 -2109
rect -822 -2113 -818 -2109
rect -813 -2113 -809 -2109
rect -805 -2113 -801 -2109
rect -796 -2113 -792 -2109
rect -778 -2113 -774 -2109
rect -769 -2113 -765 -2109
rect -761 -2113 -757 -2109
rect -745 -2113 -741 -2109
rect -737 -2113 -733 -2109
rect -725 -2113 -721 -2109
rect -713 -2113 -709 -2109
rect -704 -2113 -700 -2109
rect -695 -2113 -691 -2109
rect -577 -2113 -573 -2109
rect -568 -2113 -564 -2109
rect -559 -2113 -555 -2109
rect -551 -2113 -547 -2109
rect -542 -2113 -538 -2109
rect -533 -2113 -529 -2109
rect -525 -2113 -521 -2109
rect -517 -2113 -513 -2109
rect -499 -2113 -495 -2109
rect -489 -2113 -485 -2109
rect -481 -2113 -477 -2109
rect -464 -2113 -460 -2109
rect -455 -2113 -451 -2109
rect -447 -2113 -443 -2109
rect -438 -2113 -434 -2109
rect -420 -2113 -416 -2109
rect -411 -2113 -407 -2109
rect -403 -2113 -399 -2109
rect -387 -2113 -383 -2109
rect -379 -2113 -375 -2109
rect -367 -2113 -363 -2109
rect -355 -2113 -351 -2109
rect -346 -2113 -342 -2109
rect -337 -2113 -333 -2109
rect -219 -2113 -215 -2109
rect -210 -2113 -206 -2109
rect -201 -2113 -197 -2109
rect -193 -2113 -189 -2109
rect -184 -2113 -180 -2109
rect -175 -2113 -171 -2109
rect -167 -2113 -163 -2109
rect -159 -2113 -155 -2109
rect -141 -2113 -137 -2109
rect -131 -2113 -127 -2109
rect -123 -2113 -119 -2109
rect -106 -2113 -102 -2109
rect -97 -2113 -93 -2109
rect -89 -2113 -85 -2109
rect -80 -2113 -76 -2109
rect -62 -2113 -58 -2109
rect -53 -2113 -49 -2109
rect -45 -2113 -41 -2109
rect -29 -2113 -25 -2109
rect -21 -2113 -17 -2109
rect -9 -2113 -5 -2109
rect 3 -2113 7 -2109
rect 12 -2113 16 -2109
rect 21 -2113 25 -2109
rect 139 -2113 143 -2109
rect 148 -2113 152 -2109
rect 157 -2113 161 -2109
rect 165 -2113 169 -2109
rect 174 -2113 178 -2109
rect 183 -2113 187 -2109
rect 191 -2113 195 -2109
rect 199 -2113 203 -2109
rect 217 -2113 221 -2109
rect 227 -2113 231 -2109
rect 235 -2113 239 -2109
rect 252 -2113 256 -2109
rect 261 -2113 265 -2109
rect 269 -2113 273 -2109
rect 278 -2113 282 -2109
rect 296 -2113 300 -2109
rect 305 -2113 309 -2109
rect 313 -2113 317 -2109
rect 329 -2113 333 -2109
rect 337 -2113 341 -2109
rect 349 -2113 353 -2109
rect 361 -2113 365 -2109
rect 370 -2113 374 -2109
rect 379 -2113 383 -2109
rect 495 -2113 499 -2109
rect 504 -2113 508 -2109
rect 513 -2113 517 -2109
rect 521 -2113 525 -2109
rect 530 -2113 534 -2109
rect 539 -2113 543 -2109
rect 547 -2113 551 -2109
rect 555 -2113 559 -2109
rect 573 -2113 577 -2109
rect 583 -2113 587 -2109
rect 591 -2113 595 -2109
rect 608 -2113 612 -2109
rect 617 -2113 621 -2109
rect 625 -2113 629 -2109
rect 634 -2113 638 -2109
rect 652 -2113 656 -2109
rect 661 -2113 665 -2109
rect 669 -2113 673 -2109
rect 685 -2113 689 -2109
rect 693 -2113 697 -2109
rect 705 -2113 709 -2109
rect 717 -2113 721 -2109
rect 726 -2113 730 -2109
rect 735 -2113 739 -2109
rect 853 -2113 857 -2109
rect 862 -2113 866 -2109
rect 871 -2113 875 -2109
rect 879 -2113 883 -2109
rect 888 -2113 892 -2109
rect 897 -2113 901 -2109
rect 905 -2113 909 -2109
rect 913 -2113 917 -2109
rect 931 -2113 935 -2109
rect 941 -2113 945 -2109
rect 949 -2113 953 -2109
rect 966 -2113 970 -2109
rect 975 -2113 979 -2109
rect 983 -2113 987 -2109
rect 992 -2113 996 -2109
rect 1010 -2113 1014 -2109
rect 1019 -2113 1023 -2109
rect 1027 -2113 1031 -2109
rect 1043 -2113 1047 -2109
rect 1051 -2113 1055 -2109
rect 1063 -2113 1067 -2109
rect 1075 -2113 1079 -2109
rect 1084 -2113 1088 -2109
rect 1093 -2113 1097 -2109
rect 1211 -2113 1215 -2109
rect 1220 -2113 1224 -2109
rect 1229 -2113 1233 -2109
rect 1237 -2113 1241 -2109
rect 1246 -2113 1250 -2109
rect 1255 -2113 1259 -2109
rect 1263 -2113 1267 -2109
rect 1271 -2113 1275 -2109
rect 1289 -2113 1293 -2109
rect 1299 -2113 1303 -2109
rect 1307 -2113 1311 -2109
rect 1324 -2113 1328 -2109
rect 1333 -2113 1337 -2109
rect 1341 -2113 1345 -2109
rect 1350 -2113 1354 -2109
rect 1368 -2113 1372 -2109
rect 1377 -2113 1381 -2109
rect 1385 -2113 1389 -2109
rect 1401 -2113 1405 -2109
rect 1409 -2113 1413 -2109
rect 1421 -2113 1425 -2109
rect 1433 -2113 1437 -2109
rect 1442 -2113 1446 -2109
rect 1451 -2113 1455 -2109
rect -1234 -2257 -1230 -2253
rect -1225 -2257 -1221 -2253
rect -1216 -2257 -1212 -2253
rect -1208 -2257 -1204 -2253
rect -1192 -2257 -1188 -2253
rect -1184 -2257 -1180 -2253
rect -1167 -2257 -1163 -2253
rect -1150 -2257 -1146 -2253
rect -1142 -2257 -1138 -2253
rect -1125 -2257 -1121 -2253
rect -1108 -2257 -1104 -2253
rect -1100 -2257 -1096 -2253
rect -1083 -2257 -1079 -2253
rect -1066 -2257 -1062 -2253
rect -1058 -2257 -1054 -2253
rect -1042 -2257 -1038 -2253
rect -935 -2257 -931 -2253
rect -926 -2257 -922 -2253
rect -917 -2257 -913 -2253
rect -909 -2257 -905 -2253
rect -893 -2257 -889 -2253
rect -885 -2257 -881 -2253
rect -868 -2257 -864 -2253
rect -851 -2257 -847 -2253
rect -843 -2257 -839 -2253
rect -826 -2257 -822 -2253
rect -809 -2257 -805 -2253
rect -801 -2257 -797 -2253
rect -784 -2257 -780 -2253
rect -767 -2257 -763 -2253
rect -759 -2257 -755 -2253
rect -743 -2257 -739 -2253
rect -577 -2257 -573 -2253
rect -568 -2257 -564 -2253
rect -559 -2257 -555 -2253
rect -551 -2257 -547 -2253
rect -535 -2257 -531 -2253
rect -527 -2257 -523 -2253
rect -510 -2257 -506 -2253
rect -493 -2257 -489 -2253
rect -485 -2257 -481 -2253
rect -468 -2257 -464 -2253
rect -451 -2257 -447 -2253
rect -443 -2257 -439 -2253
rect -426 -2257 -422 -2253
rect -409 -2257 -405 -2253
rect -401 -2257 -397 -2253
rect -385 -2257 -381 -2253
rect -219 -2257 -215 -2253
rect -210 -2257 -206 -2253
rect -201 -2257 -197 -2253
rect -193 -2257 -189 -2253
rect -177 -2257 -173 -2253
rect -169 -2257 -165 -2253
rect -152 -2257 -148 -2253
rect -135 -2257 -131 -2253
rect -127 -2257 -123 -2253
rect -110 -2257 -106 -2253
rect -93 -2257 -89 -2253
rect -85 -2257 -81 -2253
rect -68 -2257 -64 -2253
rect -51 -2257 -47 -2253
rect -43 -2257 -39 -2253
rect -27 -2257 -23 -2253
rect 139 -2257 143 -2253
rect 148 -2257 152 -2253
rect 157 -2257 161 -2253
rect 165 -2257 169 -2253
rect 181 -2257 185 -2253
rect 189 -2257 193 -2253
rect 206 -2257 210 -2253
rect 223 -2257 227 -2253
rect 231 -2257 235 -2253
rect 248 -2257 252 -2253
rect 265 -2257 269 -2253
rect 273 -2257 277 -2253
rect 290 -2257 294 -2253
rect 307 -2257 311 -2253
rect 315 -2257 319 -2253
rect 331 -2257 335 -2253
rect 495 -2257 499 -2253
rect 504 -2257 508 -2253
rect 513 -2257 517 -2253
rect 521 -2257 525 -2253
rect 537 -2257 541 -2253
rect 545 -2257 549 -2253
rect 562 -2257 566 -2253
rect 579 -2257 583 -2253
rect 587 -2257 591 -2253
rect 604 -2257 608 -2253
rect 621 -2257 625 -2253
rect 629 -2257 633 -2253
rect 646 -2257 650 -2253
rect 663 -2257 667 -2253
rect 671 -2257 675 -2253
rect 687 -2257 691 -2253
rect -1559 -2428 -1555 -2424
rect -1550 -2428 -1546 -2424
rect -1541 -2428 -1537 -2424
rect -1533 -2428 -1529 -2424
rect -1517 -2428 -1513 -2424
rect -1509 -2428 -1505 -2424
rect -1492 -2428 -1488 -2424
rect -1475 -2428 -1471 -2424
rect -1467 -2428 -1463 -2424
rect -1450 -2428 -1446 -2424
rect -1433 -2428 -1429 -2424
rect -1425 -2428 -1421 -2424
rect -1408 -2428 -1404 -2424
rect -1391 -2428 -1387 -2424
rect -1383 -2428 -1379 -2424
rect -1367 -2428 -1363 -2424
rect -1234 -2428 -1230 -2424
rect -1225 -2428 -1221 -2424
rect -1216 -2428 -1212 -2424
rect -1208 -2428 -1204 -2424
rect -1192 -2428 -1188 -2424
rect -1184 -2428 -1180 -2424
rect -1167 -2428 -1163 -2424
rect -1150 -2428 -1146 -2424
rect -1142 -2428 -1138 -2424
rect -1125 -2428 -1121 -2424
rect -1108 -2428 -1104 -2424
rect -1100 -2428 -1096 -2424
rect -1083 -2428 -1079 -2424
rect -1066 -2428 -1062 -2424
rect -1058 -2428 -1054 -2424
rect -1042 -2428 -1038 -2424
rect -935 -2428 -931 -2424
rect -926 -2428 -922 -2424
rect -917 -2428 -913 -2424
rect -909 -2428 -905 -2424
rect -893 -2428 -889 -2424
rect -885 -2428 -881 -2424
rect -868 -2428 -864 -2424
rect -851 -2428 -847 -2424
rect -843 -2428 -839 -2424
rect -826 -2428 -822 -2424
rect -809 -2428 -805 -2424
rect -801 -2428 -797 -2424
rect -784 -2428 -780 -2424
rect -767 -2428 -763 -2424
rect -759 -2428 -755 -2424
rect -743 -2428 -739 -2424
rect -577 -2428 -573 -2424
rect -568 -2428 -564 -2424
rect -559 -2428 -555 -2424
rect -551 -2428 -547 -2424
rect -535 -2428 -531 -2424
rect -527 -2428 -523 -2424
rect -510 -2428 -506 -2424
rect -493 -2428 -489 -2424
rect -485 -2428 -481 -2424
rect -468 -2428 -464 -2424
rect -451 -2428 -447 -2424
rect -443 -2428 -439 -2424
rect -426 -2428 -422 -2424
rect -409 -2428 -405 -2424
rect -401 -2428 -397 -2424
rect -385 -2428 -381 -2424
rect -219 -2428 -215 -2424
rect -210 -2428 -206 -2424
rect -201 -2428 -197 -2424
rect -193 -2428 -189 -2424
rect -177 -2428 -173 -2424
rect -169 -2428 -165 -2424
rect -152 -2428 -148 -2424
rect -135 -2428 -131 -2424
rect -127 -2428 -123 -2424
rect -110 -2428 -106 -2424
rect -93 -2428 -89 -2424
rect -85 -2428 -81 -2424
rect -68 -2428 -64 -2424
rect -51 -2428 -47 -2424
rect -43 -2428 -39 -2424
rect -27 -2428 -23 -2424
rect 139 -2428 143 -2424
rect 148 -2428 152 -2424
rect 157 -2428 161 -2424
rect 165 -2428 169 -2424
rect 181 -2428 185 -2424
rect 189 -2428 193 -2424
rect 206 -2428 210 -2424
rect 223 -2428 227 -2424
rect 231 -2428 235 -2424
rect 248 -2428 252 -2424
rect 265 -2428 269 -2424
rect 273 -2428 277 -2424
rect 290 -2428 294 -2424
rect 307 -2428 311 -2424
rect 315 -2428 319 -2424
rect 331 -2428 335 -2424
rect 495 -2428 499 -2424
rect 504 -2428 508 -2424
rect 513 -2428 517 -2424
rect 521 -2428 525 -2424
rect 537 -2428 541 -2424
rect 545 -2428 549 -2424
rect 562 -2428 566 -2424
rect 579 -2428 583 -2424
rect 587 -2428 591 -2424
rect 604 -2428 608 -2424
rect 621 -2428 625 -2424
rect 629 -2428 633 -2424
rect 646 -2428 650 -2424
rect 663 -2428 667 -2424
rect 671 -2428 675 -2424
rect 687 -2428 691 -2424
rect 853 -2428 857 -2424
rect 862 -2428 866 -2424
rect 871 -2428 875 -2424
rect 879 -2428 883 -2424
rect 895 -2428 899 -2424
rect 903 -2428 907 -2424
rect 920 -2428 924 -2424
rect 937 -2428 941 -2424
rect 945 -2428 949 -2424
rect 962 -2428 966 -2424
rect 979 -2428 983 -2424
rect 987 -2428 991 -2424
rect 1004 -2428 1008 -2424
rect 1021 -2428 1025 -2424
rect 1029 -2428 1033 -2424
rect 1045 -2428 1049 -2424
rect 1211 -2428 1215 -2424
rect 1220 -2428 1224 -2424
rect 1229 -2428 1233 -2424
rect 1237 -2428 1241 -2424
rect 1253 -2428 1257 -2424
rect 1261 -2428 1265 -2424
rect 1278 -2428 1282 -2424
rect 1295 -2428 1299 -2424
rect 1303 -2428 1307 -2424
rect 1320 -2428 1324 -2424
rect 1337 -2428 1341 -2424
rect 1345 -2428 1349 -2424
rect 1362 -2428 1366 -2424
rect 1379 -2428 1383 -2424
rect 1387 -2428 1391 -2424
rect 1403 -2428 1407 -2424
rect -1559 -2599 -1555 -2595
rect -1550 -2599 -1546 -2595
rect -1541 -2599 -1537 -2595
rect -1533 -2599 -1529 -2595
rect -1517 -2599 -1513 -2595
rect -1509 -2599 -1505 -2595
rect -1492 -2599 -1488 -2595
rect -1475 -2599 -1471 -2595
rect -1467 -2599 -1463 -2595
rect -1450 -2599 -1446 -2595
rect -1433 -2599 -1429 -2595
rect -1425 -2599 -1421 -2595
rect -1408 -2599 -1404 -2595
rect -1391 -2599 -1387 -2595
rect -1383 -2599 -1379 -2595
rect -1367 -2599 -1363 -2595
rect -1234 -2599 -1230 -2595
rect -1225 -2599 -1221 -2595
rect -1216 -2599 -1212 -2595
rect -1208 -2599 -1204 -2595
rect -1192 -2599 -1188 -2595
rect -1184 -2599 -1180 -2595
rect -1167 -2599 -1163 -2595
rect -1150 -2599 -1146 -2595
rect -1142 -2599 -1138 -2595
rect -1125 -2599 -1121 -2595
rect -1108 -2599 -1104 -2595
rect -1100 -2599 -1096 -2595
rect -1083 -2599 -1079 -2595
rect -1066 -2599 -1062 -2595
rect -1058 -2599 -1054 -2595
rect -1042 -2599 -1038 -2595
rect -935 -2599 -931 -2595
rect -926 -2599 -922 -2595
rect -917 -2599 -913 -2595
rect -909 -2599 -905 -2595
rect -893 -2599 -889 -2595
rect -885 -2599 -881 -2595
rect -868 -2599 -864 -2595
rect -851 -2599 -847 -2595
rect -843 -2599 -839 -2595
rect -826 -2599 -822 -2595
rect -809 -2599 -805 -2595
rect -801 -2599 -797 -2595
rect -784 -2599 -780 -2595
rect -767 -2599 -763 -2595
rect -759 -2599 -755 -2595
rect -743 -2599 -739 -2595
rect -577 -2599 -573 -2595
rect -568 -2599 -564 -2595
rect -559 -2599 -555 -2595
rect -551 -2599 -547 -2595
rect -535 -2599 -531 -2595
rect -527 -2599 -523 -2595
rect -510 -2599 -506 -2595
rect -493 -2599 -489 -2595
rect -485 -2599 -481 -2595
rect -468 -2599 -464 -2595
rect -451 -2599 -447 -2595
rect -443 -2599 -439 -2595
rect -426 -2599 -422 -2595
rect -409 -2599 -405 -2595
rect -401 -2599 -397 -2595
rect -385 -2599 -381 -2595
rect -220 -2599 -216 -2595
rect -211 -2599 -207 -2595
rect -202 -2599 -198 -2595
rect -194 -2599 -190 -2595
rect -178 -2599 -174 -2595
rect -170 -2599 -166 -2595
rect -153 -2599 -149 -2595
rect -136 -2599 -132 -2595
rect -128 -2599 -124 -2595
rect -111 -2599 -107 -2595
rect -94 -2599 -90 -2595
rect -86 -2599 -82 -2595
rect -69 -2599 -65 -2595
rect -52 -2599 -48 -2595
rect -44 -2599 -40 -2595
rect -28 -2599 -24 -2595
rect 139 -2599 143 -2595
rect 148 -2599 152 -2595
rect 157 -2599 161 -2595
rect 165 -2599 169 -2595
rect 181 -2599 185 -2595
rect 189 -2599 193 -2595
rect 206 -2599 210 -2595
rect 223 -2599 227 -2595
rect 231 -2599 235 -2595
rect 248 -2599 252 -2595
rect 265 -2599 269 -2595
rect 273 -2599 277 -2595
rect 290 -2599 294 -2595
rect 307 -2599 311 -2595
rect 315 -2599 319 -2595
rect 331 -2599 335 -2595
rect 495 -2599 499 -2595
rect 504 -2599 508 -2595
rect 513 -2599 517 -2595
rect 521 -2599 525 -2595
rect 537 -2599 541 -2595
rect 545 -2599 549 -2595
rect 562 -2599 566 -2595
rect 579 -2599 583 -2595
rect 587 -2599 591 -2595
rect 604 -2599 608 -2595
rect 621 -2599 625 -2595
rect 629 -2599 633 -2595
rect 646 -2599 650 -2595
rect 663 -2599 667 -2595
rect 671 -2599 675 -2595
rect 687 -2599 691 -2595
rect 853 -2599 857 -2595
rect 862 -2599 866 -2595
rect 871 -2599 875 -2595
rect 879 -2599 883 -2595
rect 895 -2599 899 -2595
rect 903 -2599 907 -2595
rect 920 -2599 924 -2595
rect 937 -2599 941 -2595
rect 945 -2599 949 -2595
rect 962 -2599 966 -2595
rect 979 -2599 983 -2595
rect 987 -2599 991 -2595
rect 1004 -2599 1008 -2595
rect 1021 -2599 1025 -2595
rect 1029 -2599 1033 -2595
rect 1045 -2599 1049 -2595
rect 1211 -2599 1215 -2595
rect 1220 -2599 1224 -2595
rect 1229 -2599 1233 -2595
rect 1237 -2599 1241 -2595
rect 1253 -2599 1257 -2595
rect 1261 -2599 1265 -2595
rect 1278 -2599 1282 -2595
rect 1295 -2599 1299 -2595
rect 1303 -2599 1307 -2595
rect 1320 -2599 1324 -2595
rect 1337 -2599 1341 -2595
rect 1345 -2599 1349 -2595
rect 1362 -2599 1366 -2595
rect 1379 -2599 1383 -2595
rect 1387 -2599 1391 -2595
rect 1403 -2599 1407 -2595
rect -1309 -2704 -1305 -2700
rect -1292 -2704 -1288 -2700
rect -1283 -2704 -1279 -2700
rect -935 -2704 -931 -2700
rect -918 -2704 -914 -2700
rect -909 -2704 -905 -2700
rect -577 -2704 -573 -2700
rect -560 -2704 -556 -2700
rect -551 -2704 -547 -2700
rect -219 -2704 -215 -2700
rect -202 -2704 -198 -2700
rect -193 -2704 -189 -2700
rect 139 -2704 143 -2700
rect 156 -2704 160 -2700
rect 165 -2704 169 -2700
rect 495 -2704 499 -2700
rect 512 -2704 516 -2700
rect 521 -2704 525 -2700
rect 853 -2704 857 -2700
rect 870 -2704 874 -2700
rect 879 -2704 883 -2700
rect 1211 -2704 1215 -2700
rect 1228 -2704 1232 -2700
rect 1237 -2704 1241 -2700
rect -1234 -2863 -1230 -2859
rect -1225 -2863 -1221 -2859
rect -1216 -2863 -1212 -2859
rect -1208 -2863 -1204 -2859
rect -1199 -2863 -1195 -2859
rect -1181 -2863 -1177 -2859
rect -1172 -2863 -1168 -2859
rect -1164 -2863 -1160 -2859
rect -1147 -2863 -1143 -2859
rect -1138 -2863 -1134 -2859
rect -935 -2863 -931 -2859
rect -926 -2863 -922 -2859
rect -917 -2863 -913 -2859
rect -909 -2863 -905 -2859
rect -900 -2863 -896 -2859
rect -891 -2863 -887 -2859
rect -883 -2863 -879 -2859
rect -875 -2863 -871 -2859
rect -857 -2863 -853 -2859
rect -847 -2863 -843 -2859
rect -839 -2863 -835 -2859
rect -822 -2863 -818 -2859
rect -813 -2863 -809 -2859
rect -805 -2863 -801 -2859
rect -796 -2863 -792 -2859
rect -778 -2863 -774 -2859
rect -769 -2863 -765 -2859
rect -761 -2863 -757 -2859
rect -745 -2863 -741 -2859
rect -737 -2863 -733 -2859
rect -725 -2863 -721 -2859
rect -713 -2863 -709 -2859
rect -704 -2863 -700 -2859
rect -695 -2863 -691 -2859
rect -577 -2863 -573 -2859
rect -568 -2863 -564 -2859
rect -559 -2863 -555 -2859
rect -551 -2863 -547 -2859
rect -542 -2863 -538 -2859
rect -533 -2863 -529 -2859
rect -525 -2863 -521 -2859
rect -517 -2863 -513 -2859
rect -499 -2863 -495 -2859
rect -489 -2863 -485 -2859
rect -481 -2863 -477 -2859
rect -464 -2863 -460 -2859
rect -455 -2863 -451 -2859
rect -447 -2863 -443 -2859
rect -438 -2863 -434 -2859
rect -420 -2863 -416 -2859
rect -411 -2863 -407 -2859
rect -403 -2863 -399 -2859
rect -387 -2863 -383 -2859
rect -379 -2863 -375 -2859
rect -367 -2863 -363 -2859
rect -355 -2863 -351 -2859
rect -346 -2863 -342 -2859
rect -337 -2863 -333 -2859
rect -219 -2863 -215 -2859
rect -210 -2863 -206 -2859
rect -201 -2863 -197 -2859
rect -193 -2863 -189 -2859
rect -184 -2863 -180 -2859
rect -175 -2863 -171 -2859
rect -167 -2863 -163 -2859
rect -159 -2863 -155 -2859
rect -141 -2863 -137 -2859
rect -131 -2863 -127 -2859
rect -123 -2863 -119 -2859
rect -106 -2863 -102 -2859
rect -97 -2863 -93 -2859
rect -89 -2863 -85 -2859
rect -80 -2863 -76 -2859
rect -62 -2863 -58 -2859
rect -53 -2863 -49 -2859
rect -45 -2863 -41 -2859
rect -29 -2863 -25 -2859
rect -21 -2863 -17 -2859
rect -9 -2863 -5 -2859
rect 3 -2863 7 -2859
rect 12 -2863 16 -2859
rect 21 -2863 25 -2859
rect 139 -2863 143 -2859
rect 148 -2863 152 -2859
rect 157 -2863 161 -2859
rect 165 -2863 169 -2859
rect 174 -2863 178 -2859
rect 183 -2863 187 -2859
rect 191 -2863 195 -2859
rect 199 -2863 203 -2859
rect 217 -2863 221 -2859
rect 227 -2863 231 -2859
rect 235 -2863 239 -2859
rect 252 -2863 256 -2859
rect 261 -2863 265 -2859
rect 269 -2863 273 -2859
rect 278 -2863 282 -2859
rect 296 -2863 300 -2859
rect 305 -2863 309 -2859
rect 313 -2863 317 -2859
rect 329 -2863 333 -2859
rect 337 -2863 341 -2859
rect 349 -2863 353 -2859
rect 361 -2863 365 -2859
rect 370 -2863 374 -2859
rect 379 -2863 383 -2859
rect 495 -2863 499 -2859
rect 504 -2863 508 -2859
rect 513 -2863 517 -2859
rect 521 -2863 525 -2859
rect 530 -2863 534 -2859
rect 539 -2863 543 -2859
rect 547 -2863 551 -2859
rect 555 -2863 559 -2859
rect 573 -2863 577 -2859
rect 583 -2863 587 -2859
rect 591 -2863 595 -2859
rect 608 -2863 612 -2859
rect 617 -2863 621 -2859
rect 625 -2863 629 -2859
rect 634 -2863 638 -2859
rect 652 -2863 656 -2859
rect 661 -2863 665 -2859
rect 669 -2863 673 -2859
rect 685 -2863 689 -2859
rect 693 -2863 697 -2859
rect 705 -2863 709 -2859
rect 717 -2863 721 -2859
rect 726 -2863 730 -2859
rect 735 -2863 739 -2859
rect 853 -2863 857 -2859
rect 862 -2863 866 -2859
rect 871 -2863 875 -2859
rect 879 -2863 883 -2859
rect 888 -2863 892 -2859
rect 897 -2863 901 -2859
rect 905 -2863 909 -2859
rect 913 -2863 917 -2859
rect 931 -2863 935 -2859
rect 941 -2863 945 -2859
rect 949 -2863 953 -2859
rect 966 -2863 970 -2859
rect 975 -2863 979 -2859
rect 983 -2863 987 -2859
rect 992 -2863 996 -2859
rect 1010 -2863 1014 -2859
rect 1019 -2863 1023 -2859
rect 1027 -2863 1031 -2859
rect 1043 -2863 1047 -2859
rect 1051 -2863 1055 -2859
rect 1063 -2863 1067 -2859
rect 1075 -2863 1079 -2859
rect 1084 -2863 1088 -2859
rect 1093 -2863 1097 -2859
rect 1211 -2863 1215 -2859
rect 1220 -2863 1224 -2859
rect 1229 -2863 1233 -2859
rect 1237 -2863 1241 -2859
rect 1246 -2863 1250 -2859
rect 1255 -2863 1259 -2859
rect 1263 -2863 1267 -2859
rect 1271 -2863 1275 -2859
rect 1289 -2863 1293 -2859
rect 1299 -2863 1303 -2859
rect 1307 -2863 1311 -2859
rect 1324 -2863 1328 -2859
rect 1333 -2863 1337 -2859
rect 1341 -2863 1345 -2859
rect 1350 -2863 1354 -2859
rect 1368 -2863 1372 -2859
rect 1377 -2863 1381 -2859
rect 1385 -2863 1389 -2859
rect 1401 -2863 1405 -2859
rect 1409 -2863 1413 -2859
rect 1421 -2863 1425 -2859
rect 1433 -2863 1437 -2859
rect 1442 -2863 1446 -2859
rect 1451 -2863 1455 -2859
rect -1559 -2982 -1555 -2978
rect -1550 -2982 -1546 -2978
rect -1541 -2982 -1537 -2978
rect -1533 -2982 -1529 -2978
rect -1517 -2982 -1513 -2978
rect -1509 -2982 -1505 -2978
rect -1492 -2982 -1488 -2978
rect -1475 -2982 -1471 -2978
rect -1467 -2982 -1463 -2978
rect -1450 -2982 -1446 -2978
rect -1433 -2982 -1429 -2978
rect -1425 -2982 -1421 -2978
rect -1408 -2982 -1404 -2978
rect -1391 -2982 -1387 -2978
rect -1383 -2982 -1379 -2978
rect -1367 -2982 -1363 -2978
rect -1234 -2982 -1230 -2978
rect -1225 -2982 -1221 -2978
rect -1216 -2982 -1212 -2978
rect -1208 -2982 -1204 -2978
rect -1192 -2982 -1188 -2978
rect -1184 -2982 -1180 -2978
rect -1167 -2982 -1163 -2978
rect -1150 -2982 -1146 -2978
rect -1142 -2982 -1138 -2978
rect -1125 -2982 -1121 -2978
rect -1108 -2982 -1104 -2978
rect -1100 -2982 -1096 -2978
rect -1083 -2982 -1079 -2978
rect -1066 -2982 -1062 -2978
rect -1058 -2982 -1054 -2978
rect -1042 -2982 -1038 -2978
rect -935 -2982 -931 -2978
rect -926 -2982 -922 -2978
rect -917 -2982 -913 -2978
rect -909 -2982 -905 -2978
rect -893 -2982 -889 -2978
rect -885 -2982 -881 -2978
rect -868 -2982 -864 -2978
rect -851 -2982 -847 -2978
rect -843 -2982 -839 -2978
rect -826 -2982 -822 -2978
rect -809 -2982 -805 -2978
rect -801 -2982 -797 -2978
rect -784 -2982 -780 -2978
rect -767 -2982 -763 -2978
rect -759 -2982 -755 -2978
rect -743 -2982 -739 -2978
rect -577 -2982 -573 -2978
rect -568 -2982 -564 -2978
rect -559 -2982 -555 -2978
rect -551 -2982 -547 -2978
rect -535 -2982 -531 -2978
rect -527 -2982 -523 -2978
rect -510 -2982 -506 -2978
rect -493 -2982 -489 -2978
rect -485 -2982 -481 -2978
rect -468 -2982 -464 -2978
rect -451 -2982 -447 -2978
rect -443 -2982 -439 -2978
rect -426 -2982 -422 -2978
rect -409 -2982 -405 -2978
rect -401 -2982 -397 -2978
rect -385 -2982 -381 -2978
rect -219 -2982 -215 -2978
rect -210 -2982 -206 -2978
rect -201 -2982 -197 -2978
rect -193 -2982 -189 -2978
rect -177 -2982 -173 -2978
rect -169 -2982 -165 -2978
rect -152 -2982 -148 -2978
rect -135 -2982 -131 -2978
rect -127 -2982 -123 -2978
rect -110 -2982 -106 -2978
rect -93 -2982 -89 -2978
rect -85 -2982 -81 -2978
rect -68 -2982 -64 -2978
rect -51 -2982 -47 -2978
rect -43 -2982 -39 -2978
rect -27 -2982 -23 -2978
rect 139 -2982 143 -2978
rect 148 -2982 152 -2978
rect 157 -2982 161 -2978
rect 165 -2982 169 -2978
rect 181 -2982 185 -2978
rect 189 -2982 193 -2978
rect 206 -2982 210 -2978
rect 223 -2982 227 -2978
rect 231 -2982 235 -2978
rect 248 -2982 252 -2978
rect 265 -2982 269 -2978
rect 273 -2982 277 -2978
rect 290 -2982 294 -2978
rect 307 -2982 311 -2978
rect 315 -2982 319 -2978
rect 331 -2982 335 -2978
rect -1559 -3153 -1555 -3149
rect -1550 -3153 -1546 -3149
rect -1541 -3153 -1537 -3149
rect -1533 -3153 -1529 -3149
rect -1517 -3153 -1513 -3149
rect -1509 -3153 -1505 -3149
rect -1492 -3153 -1488 -3149
rect -1475 -3153 -1471 -3149
rect -1467 -3153 -1463 -3149
rect -1450 -3153 -1446 -3149
rect -1433 -3153 -1429 -3149
rect -1425 -3153 -1421 -3149
rect -1408 -3153 -1404 -3149
rect -1391 -3153 -1387 -3149
rect -1383 -3153 -1379 -3149
rect -1367 -3153 -1363 -3149
rect -1234 -3153 -1230 -3149
rect -1225 -3153 -1221 -3149
rect -1216 -3153 -1212 -3149
rect -1208 -3153 -1204 -3149
rect -1192 -3153 -1188 -3149
rect -1184 -3153 -1180 -3149
rect -1167 -3153 -1163 -3149
rect -1150 -3153 -1146 -3149
rect -1142 -3153 -1138 -3149
rect -1125 -3153 -1121 -3149
rect -1108 -3153 -1104 -3149
rect -1100 -3153 -1096 -3149
rect -1083 -3153 -1079 -3149
rect -1066 -3153 -1062 -3149
rect -1058 -3153 -1054 -3149
rect -1042 -3153 -1038 -3149
rect -935 -3153 -931 -3149
rect -926 -3153 -922 -3149
rect -917 -3153 -913 -3149
rect -909 -3153 -905 -3149
rect -893 -3153 -889 -3149
rect -885 -3153 -881 -3149
rect -868 -3153 -864 -3149
rect -851 -3153 -847 -3149
rect -843 -3153 -839 -3149
rect -826 -3153 -822 -3149
rect -809 -3153 -805 -3149
rect -801 -3153 -797 -3149
rect -784 -3153 -780 -3149
rect -767 -3153 -763 -3149
rect -759 -3153 -755 -3149
rect -743 -3153 -739 -3149
rect -577 -3153 -573 -3149
rect -568 -3153 -564 -3149
rect -559 -3153 -555 -3149
rect -551 -3153 -547 -3149
rect -535 -3153 -531 -3149
rect -527 -3153 -523 -3149
rect -510 -3153 -506 -3149
rect -493 -3153 -489 -3149
rect -485 -3153 -481 -3149
rect -468 -3153 -464 -3149
rect -451 -3153 -447 -3149
rect -443 -3153 -439 -3149
rect -426 -3153 -422 -3149
rect -409 -3153 -405 -3149
rect -401 -3153 -397 -3149
rect -385 -3153 -381 -3149
rect -219 -3153 -215 -3149
rect -210 -3153 -206 -3149
rect -201 -3153 -197 -3149
rect -193 -3153 -189 -3149
rect -177 -3153 -173 -3149
rect -169 -3153 -165 -3149
rect -152 -3153 -148 -3149
rect -135 -3153 -131 -3149
rect -127 -3153 -123 -3149
rect -110 -3153 -106 -3149
rect -93 -3153 -89 -3149
rect -85 -3153 -81 -3149
rect -68 -3153 -64 -3149
rect -51 -3153 -47 -3149
rect -43 -3153 -39 -3149
rect -27 -3153 -23 -3149
rect 139 -3153 143 -3149
rect 148 -3153 152 -3149
rect 157 -3153 161 -3149
rect 165 -3153 169 -3149
rect 181 -3153 185 -3149
rect 189 -3153 193 -3149
rect 206 -3153 210 -3149
rect 223 -3153 227 -3149
rect 231 -3153 235 -3149
rect 248 -3153 252 -3149
rect 265 -3153 269 -3149
rect 273 -3153 277 -3149
rect 290 -3153 294 -3149
rect 307 -3153 311 -3149
rect 315 -3153 319 -3149
rect 331 -3153 335 -3149
rect 495 -3153 499 -3149
rect 504 -3153 508 -3149
rect 513 -3153 517 -3149
rect 521 -3153 525 -3149
rect 537 -3153 541 -3149
rect 545 -3153 549 -3149
rect 562 -3153 566 -3149
rect 579 -3153 583 -3149
rect 587 -3153 591 -3149
rect 604 -3153 608 -3149
rect 621 -3153 625 -3149
rect 629 -3153 633 -3149
rect 646 -3153 650 -3149
rect 663 -3153 667 -3149
rect 671 -3153 675 -3149
rect 687 -3153 691 -3149
rect 853 -3153 857 -3149
rect 862 -3153 866 -3149
rect 871 -3153 875 -3149
rect 879 -3153 883 -3149
rect 895 -3153 899 -3149
rect 903 -3153 907 -3149
rect 920 -3153 924 -3149
rect 937 -3153 941 -3149
rect 945 -3153 949 -3149
rect 962 -3153 966 -3149
rect 979 -3153 983 -3149
rect 987 -3153 991 -3149
rect 1004 -3153 1008 -3149
rect 1021 -3153 1025 -3149
rect 1029 -3153 1033 -3149
rect 1045 -3153 1049 -3149
rect 1211 -3153 1215 -3149
rect 1220 -3153 1224 -3149
rect 1229 -3153 1233 -3149
rect 1237 -3153 1241 -3149
rect 1253 -3153 1257 -3149
rect 1261 -3153 1265 -3149
rect 1278 -3153 1282 -3149
rect 1295 -3153 1299 -3149
rect 1303 -3153 1307 -3149
rect 1320 -3153 1324 -3149
rect 1337 -3153 1341 -3149
rect 1345 -3153 1349 -3149
rect 1362 -3153 1366 -3149
rect 1379 -3153 1383 -3149
rect 1387 -3153 1391 -3149
rect 1403 -3153 1407 -3149
rect -1559 -3324 -1555 -3320
rect -1550 -3324 -1546 -3320
rect -1541 -3324 -1537 -3320
rect -1533 -3324 -1529 -3320
rect -1517 -3324 -1513 -3320
rect -1509 -3324 -1505 -3320
rect -1492 -3324 -1488 -3320
rect -1475 -3324 -1471 -3320
rect -1467 -3324 -1463 -3320
rect -1450 -3324 -1446 -3320
rect -1433 -3324 -1429 -3320
rect -1425 -3324 -1421 -3320
rect -1408 -3324 -1404 -3320
rect -1391 -3324 -1387 -3320
rect -1383 -3324 -1379 -3320
rect -1367 -3324 -1363 -3320
rect -1234 -3324 -1230 -3320
rect -1225 -3324 -1221 -3320
rect -1216 -3324 -1212 -3320
rect -1208 -3324 -1204 -3320
rect -1192 -3324 -1188 -3320
rect -1184 -3324 -1180 -3320
rect -1167 -3324 -1163 -3320
rect -1150 -3324 -1146 -3320
rect -1142 -3324 -1138 -3320
rect -1125 -3324 -1121 -3320
rect -1108 -3324 -1104 -3320
rect -1100 -3324 -1096 -3320
rect -1083 -3324 -1079 -3320
rect -1066 -3324 -1062 -3320
rect -1058 -3324 -1054 -3320
rect -1042 -3324 -1038 -3320
rect -935 -3324 -931 -3320
rect -926 -3324 -922 -3320
rect -917 -3324 -913 -3320
rect -909 -3324 -905 -3320
rect -893 -3324 -889 -3320
rect -885 -3324 -881 -3320
rect -868 -3324 -864 -3320
rect -851 -3324 -847 -3320
rect -843 -3324 -839 -3320
rect -826 -3324 -822 -3320
rect -809 -3324 -805 -3320
rect -801 -3324 -797 -3320
rect -784 -3324 -780 -3320
rect -767 -3324 -763 -3320
rect -759 -3324 -755 -3320
rect -743 -3324 -739 -3320
rect -577 -3324 -573 -3320
rect -568 -3324 -564 -3320
rect -559 -3324 -555 -3320
rect -551 -3324 -547 -3320
rect -535 -3324 -531 -3320
rect -527 -3324 -523 -3320
rect -510 -3324 -506 -3320
rect -493 -3324 -489 -3320
rect -485 -3324 -481 -3320
rect -468 -3324 -464 -3320
rect -451 -3324 -447 -3320
rect -443 -3324 -439 -3320
rect -426 -3324 -422 -3320
rect -409 -3324 -405 -3320
rect -401 -3324 -397 -3320
rect -385 -3324 -381 -3320
rect -219 -3324 -215 -3320
rect -210 -3324 -206 -3320
rect -201 -3324 -197 -3320
rect -193 -3324 -189 -3320
rect -177 -3324 -173 -3320
rect -169 -3324 -165 -3320
rect -152 -3324 -148 -3320
rect -135 -3324 -131 -3320
rect -127 -3324 -123 -3320
rect -110 -3324 -106 -3320
rect -93 -3324 -89 -3320
rect -85 -3324 -81 -3320
rect -68 -3324 -64 -3320
rect -51 -3324 -47 -3320
rect -43 -3324 -39 -3320
rect -27 -3324 -23 -3320
rect 139 -3324 143 -3320
rect 148 -3324 152 -3320
rect 157 -3324 161 -3320
rect 165 -3324 169 -3320
rect 181 -3324 185 -3320
rect 189 -3324 193 -3320
rect 206 -3324 210 -3320
rect 223 -3324 227 -3320
rect 231 -3324 235 -3320
rect 248 -3324 252 -3320
rect 265 -3324 269 -3320
rect 273 -3324 277 -3320
rect 290 -3324 294 -3320
rect 307 -3324 311 -3320
rect 315 -3324 319 -3320
rect 331 -3324 335 -3320
rect 495 -3324 499 -3320
rect 504 -3324 508 -3320
rect 513 -3324 517 -3320
rect 521 -3324 525 -3320
rect 537 -3324 541 -3320
rect 545 -3324 549 -3320
rect 562 -3324 566 -3320
rect 579 -3324 583 -3320
rect 587 -3324 591 -3320
rect 604 -3324 608 -3320
rect 621 -3324 625 -3320
rect 629 -3324 633 -3320
rect 646 -3324 650 -3320
rect 663 -3324 667 -3320
rect 671 -3324 675 -3320
rect 687 -3324 691 -3320
rect 853 -3324 857 -3320
rect 862 -3324 866 -3320
rect 871 -3324 875 -3320
rect 879 -3324 883 -3320
rect 895 -3324 899 -3320
rect 903 -3324 907 -3320
rect 920 -3324 924 -3320
rect 937 -3324 941 -3320
rect 945 -3324 949 -3320
rect 962 -3324 966 -3320
rect 979 -3324 983 -3320
rect 987 -3324 991 -3320
rect 1004 -3324 1008 -3320
rect 1021 -3324 1025 -3320
rect 1029 -3324 1033 -3320
rect 1045 -3324 1049 -3320
rect 1211 -3324 1215 -3320
rect 1220 -3324 1224 -3320
rect 1229 -3324 1233 -3320
rect 1237 -3324 1241 -3320
rect 1253 -3324 1257 -3320
rect 1261 -3324 1265 -3320
rect 1278 -3324 1282 -3320
rect 1295 -3324 1299 -3320
rect 1303 -3324 1307 -3320
rect 1320 -3324 1324 -3320
rect 1337 -3324 1341 -3320
rect 1345 -3324 1349 -3320
rect 1362 -3324 1366 -3320
rect 1379 -3324 1383 -3320
rect 1387 -3324 1391 -3320
rect 1403 -3324 1407 -3320
rect -1309 -3435 -1305 -3431
rect -1292 -3435 -1288 -3431
rect -1283 -3435 -1279 -3431
rect -935 -3435 -931 -3431
rect -918 -3435 -914 -3431
rect -909 -3435 -905 -3431
rect -577 -3435 -573 -3431
rect -560 -3435 -556 -3431
rect -551 -3435 -547 -3431
rect -219 -3435 -215 -3431
rect -202 -3435 -198 -3431
rect -193 -3435 -189 -3431
rect 139 -3435 143 -3431
rect 156 -3435 160 -3431
rect 165 -3435 169 -3431
rect 495 -3435 499 -3431
rect 512 -3435 516 -3431
rect 521 -3435 525 -3431
rect 853 -3435 857 -3431
rect 870 -3435 874 -3431
rect 879 -3435 883 -3431
rect 1211 -3435 1215 -3431
rect 1228 -3435 1232 -3431
rect 1237 -3435 1241 -3431
rect -1234 -3594 -1230 -3590
rect -1225 -3594 -1221 -3590
rect -1216 -3594 -1212 -3590
rect -1208 -3594 -1204 -3590
rect -1199 -3594 -1195 -3590
rect -1181 -3594 -1177 -3590
rect -1172 -3594 -1168 -3590
rect -1164 -3594 -1160 -3590
rect -1147 -3594 -1143 -3590
rect -1138 -3594 -1134 -3590
rect -935 -3594 -931 -3590
rect -926 -3594 -922 -3590
rect -917 -3594 -913 -3590
rect -909 -3594 -905 -3590
rect -900 -3594 -896 -3590
rect -891 -3594 -887 -3590
rect -883 -3594 -879 -3590
rect -875 -3594 -871 -3590
rect -857 -3594 -853 -3590
rect -847 -3594 -843 -3590
rect -839 -3594 -835 -3590
rect -822 -3594 -818 -3590
rect -813 -3594 -809 -3590
rect -805 -3594 -801 -3590
rect -796 -3594 -792 -3590
rect -778 -3594 -774 -3590
rect -769 -3594 -765 -3590
rect -761 -3594 -757 -3590
rect -745 -3594 -741 -3590
rect -737 -3594 -733 -3590
rect -725 -3594 -721 -3590
rect -713 -3594 -709 -3590
rect -704 -3594 -700 -3590
rect -695 -3594 -691 -3590
rect -577 -3594 -573 -3590
rect -568 -3594 -564 -3590
rect -559 -3594 -555 -3590
rect -551 -3594 -547 -3590
rect -542 -3594 -538 -3590
rect -533 -3594 -529 -3590
rect -525 -3594 -521 -3590
rect -517 -3594 -513 -3590
rect -499 -3594 -495 -3590
rect -489 -3594 -485 -3590
rect -481 -3594 -477 -3590
rect -464 -3594 -460 -3590
rect -455 -3594 -451 -3590
rect -447 -3594 -443 -3590
rect -438 -3594 -434 -3590
rect -420 -3594 -416 -3590
rect -411 -3594 -407 -3590
rect -403 -3594 -399 -3590
rect -387 -3594 -383 -3590
rect -379 -3594 -375 -3590
rect -367 -3594 -363 -3590
rect -355 -3594 -351 -3590
rect -346 -3594 -342 -3590
rect -337 -3594 -333 -3590
rect -219 -3594 -215 -3590
rect -210 -3594 -206 -3590
rect -201 -3594 -197 -3590
rect -193 -3594 -189 -3590
rect -184 -3594 -180 -3590
rect -175 -3594 -171 -3590
rect -167 -3594 -163 -3590
rect -159 -3594 -155 -3590
rect -141 -3594 -137 -3590
rect -131 -3594 -127 -3590
rect -123 -3594 -119 -3590
rect -106 -3594 -102 -3590
rect -97 -3594 -93 -3590
rect -89 -3594 -85 -3590
rect -80 -3594 -76 -3590
rect -62 -3594 -58 -3590
rect -53 -3594 -49 -3590
rect -45 -3594 -41 -3590
rect -29 -3594 -25 -3590
rect -21 -3594 -17 -3590
rect -9 -3594 -5 -3590
rect 3 -3594 7 -3590
rect 12 -3594 16 -3590
rect 21 -3594 25 -3590
rect 139 -3594 143 -3590
rect 148 -3594 152 -3590
rect 157 -3594 161 -3590
rect 165 -3594 169 -3590
rect 174 -3594 178 -3590
rect 183 -3594 187 -3590
rect 191 -3594 195 -3590
rect 199 -3594 203 -3590
rect 217 -3594 221 -3590
rect 227 -3594 231 -3590
rect 235 -3594 239 -3590
rect 252 -3594 256 -3590
rect 261 -3594 265 -3590
rect 269 -3594 273 -3590
rect 278 -3594 282 -3590
rect 296 -3594 300 -3590
rect 305 -3594 309 -3590
rect 313 -3594 317 -3590
rect 329 -3594 333 -3590
rect 337 -3594 341 -3590
rect 349 -3594 353 -3590
rect 361 -3594 365 -3590
rect 370 -3594 374 -3590
rect 379 -3594 383 -3590
rect 495 -3594 499 -3590
rect 504 -3594 508 -3590
rect 513 -3594 517 -3590
rect 521 -3594 525 -3590
rect 530 -3594 534 -3590
rect 539 -3594 543 -3590
rect 547 -3594 551 -3590
rect 555 -3594 559 -3590
rect 573 -3594 577 -3590
rect 583 -3594 587 -3590
rect 591 -3594 595 -3590
rect 608 -3594 612 -3590
rect 617 -3594 621 -3590
rect 625 -3594 629 -3590
rect 634 -3594 638 -3590
rect 652 -3594 656 -3590
rect 661 -3594 665 -3590
rect 669 -3594 673 -3590
rect 685 -3594 689 -3590
rect 693 -3594 697 -3590
rect 705 -3594 709 -3590
rect 717 -3594 721 -3590
rect 726 -3594 730 -3590
rect 735 -3594 739 -3590
rect 853 -3594 857 -3590
rect 862 -3594 866 -3590
rect 871 -3594 875 -3590
rect 879 -3594 883 -3590
rect 888 -3594 892 -3590
rect 897 -3594 901 -3590
rect 905 -3594 909 -3590
rect 913 -3594 917 -3590
rect 931 -3594 935 -3590
rect 941 -3594 945 -3590
rect 949 -3594 953 -3590
rect 966 -3594 970 -3590
rect 975 -3594 979 -3590
rect 983 -3594 987 -3590
rect 992 -3594 996 -3590
rect 1010 -3594 1014 -3590
rect 1019 -3594 1023 -3590
rect 1027 -3594 1031 -3590
rect 1043 -3594 1047 -3590
rect 1051 -3594 1055 -3590
rect 1063 -3594 1067 -3590
rect 1075 -3594 1079 -3590
rect 1084 -3594 1088 -3590
rect 1093 -3594 1097 -3590
rect 1211 -3594 1215 -3590
rect 1220 -3594 1224 -3590
rect 1229 -3594 1233 -3590
rect 1237 -3594 1241 -3590
rect 1246 -3594 1250 -3590
rect 1255 -3594 1259 -3590
rect 1263 -3594 1267 -3590
rect 1271 -3594 1275 -3590
rect 1289 -3594 1293 -3590
rect 1299 -3594 1303 -3590
rect 1307 -3594 1311 -3590
rect 1324 -3594 1328 -3590
rect 1333 -3594 1337 -3590
rect 1341 -3594 1345 -3590
rect 1350 -3594 1354 -3590
rect 1368 -3594 1372 -3590
rect 1377 -3594 1381 -3590
rect 1385 -3594 1389 -3590
rect 1401 -3594 1405 -3590
rect 1409 -3594 1413 -3590
rect 1421 -3594 1425 -3590
rect 1433 -3594 1437 -3590
rect 1442 -3594 1446 -3590
rect 1451 -3594 1455 -3590
rect -1822 -3724 -1818 -3720
rect -1813 -3724 -1809 -3720
rect -1804 -3724 -1800 -3720
rect -1796 -3724 -1792 -3720
rect -1780 -3724 -1776 -3720
rect -1772 -3724 -1768 -3720
rect -1755 -3724 -1751 -3720
rect -1738 -3724 -1734 -3720
rect -1730 -3724 -1726 -3720
rect -1713 -3724 -1709 -3720
rect -1696 -3724 -1692 -3720
rect -1688 -3724 -1684 -3720
rect -1671 -3724 -1667 -3720
rect -1654 -3724 -1650 -3720
rect -1646 -3724 -1642 -3720
rect -1630 -3724 -1626 -3720
rect -1559 -3724 -1555 -3720
rect -1550 -3724 -1546 -3720
rect -1541 -3724 -1537 -3720
rect -1533 -3724 -1529 -3720
rect -1517 -3724 -1513 -3720
rect -1509 -3724 -1505 -3720
rect -1492 -3724 -1488 -3720
rect -1475 -3724 -1471 -3720
rect -1467 -3724 -1463 -3720
rect -1450 -3724 -1446 -3720
rect -1433 -3724 -1429 -3720
rect -1425 -3724 -1421 -3720
rect -1408 -3724 -1404 -3720
rect -1391 -3724 -1387 -3720
rect -1383 -3724 -1379 -3720
rect -1367 -3724 -1363 -3720
rect -1234 -3724 -1230 -3720
rect -1225 -3724 -1221 -3720
rect -1216 -3724 -1212 -3720
rect -1208 -3724 -1204 -3720
rect -1192 -3724 -1188 -3720
rect -1184 -3724 -1180 -3720
rect -1167 -3724 -1163 -3720
rect -1150 -3724 -1146 -3720
rect -1142 -3724 -1138 -3720
rect -1125 -3724 -1121 -3720
rect -1108 -3724 -1104 -3720
rect -1100 -3724 -1096 -3720
rect -1083 -3724 -1079 -3720
rect -1066 -3724 -1062 -3720
rect -1058 -3724 -1054 -3720
rect -1042 -3724 -1038 -3720
rect -934 -3724 -930 -3720
rect -925 -3724 -921 -3720
rect -916 -3724 -912 -3720
rect -908 -3724 -904 -3720
rect -892 -3724 -888 -3720
rect -884 -3724 -880 -3720
rect -867 -3724 -863 -3720
rect -850 -3724 -846 -3720
rect -842 -3724 -838 -3720
rect -825 -3724 -821 -3720
rect -808 -3724 -804 -3720
rect -800 -3724 -796 -3720
rect -783 -3724 -779 -3720
rect -766 -3724 -762 -3720
rect -758 -3724 -754 -3720
rect -742 -3724 -738 -3720
rect -577 -3724 -573 -3720
rect -568 -3724 -564 -3720
rect -559 -3724 -555 -3720
rect -551 -3724 -547 -3720
rect -535 -3724 -531 -3720
rect -527 -3724 -523 -3720
rect -510 -3724 -506 -3720
rect -493 -3724 -489 -3720
rect -485 -3724 -481 -3720
rect -468 -3724 -464 -3720
rect -451 -3724 -447 -3720
rect -443 -3724 -439 -3720
rect -426 -3724 -422 -3720
rect -409 -3724 -405 -3720
rect -401 -3724 -397 -3720
rect -385 -3724 -381 -3720
rect -219 -3724 -215 -3720
rect -210 -3724 -206 -3720
rect -201 -3724 -197 -3720
rect -193 -3724 -189 -3720
rect -177 -3724 -173 -3720
rect -169 -3724 -165 -3720
rect -152 -3724 -148 -3720
rect -135 -3724 -131 -3720
rect -127 -3724 -123 -3720
rect -110 -3724 -106 -3720
rect -93 -3724 -89 -3720
rect -85 -3724 -81 -3720
rect -68 -3724 -64 -3720
rect -51 -3724 -47 -3720
rect -43 -3724 -39 -3720
rect -27 -3724 -23 -3720
rect -1559 -3895 -1555 -3891
rect -1550 -3895 -1546 -3891
rect -1541 -3895 -1537 -3891
rect -1533 -3895 -1529 -3891
rect -1517 -3895 -1513 -3891
rect -1509 -3895 -1505 -3891
rect -1492 -3895 -1488 -3891
rect -1475 -3895 -1471 -3891
rect -1467 -3895 -1463 -3891
rect -1450 -3895 -1446 -3891
rect -1433 -3895 -1429 -3891
rect -1425 -3895 -1421 -3891
rect -1408 -3895 -1404 -3891
rect -1391 -3895 -1387 -3891
rect -1383 -3895 -1379 -3891
rect -1367 -3895 -1363 -3891
rect -1234 -3895 -1230 -3891
rect -1225 -3895 -1221 -3891
rect -1216 -3895 -1212 -3891
rect -1208 -3895 -1204 -3891
rect -1192 -3895 -1188 -3891
rect -1184 -3895 -1180 -3891
rect -1167 -3895 -1163 -3891
rect -1150 -3895 -1146 -3891
rect -1142 -3895 -1138 -3891
rect -1125 -3895 -1121 -3891
rect -1108 -3895 -1104 -3891
rect -1100 -3895 -1096 -3891
rect -1083 -3895 -1079 -3891
rect -1066 -3895 -1062 -3891
rect -1058 -3895 -1054 -3891
rect -1042 -3895 -1038 -3891
rect -934 -3895 -930 -3891
rect -925 -3895 -921 -3891
rect -916 -3895 -912 -3891
rect -908 -3895 -904 -3891
rect -892 -3895 -888 -3891
rect -884 -3895 -880 -3891
rect -867 -3895 -863 -3891
rect -850 -3895 -846 -3891
rect -842 -3895 -838 -3891
rect -825 -3895 -821 -3891
rect -808 -3895 -804 -3891
rect -800 -3895 -796 -3891
rect -783 -3895 -779 -3891
rect -766 -3895 -762 -3891
rect -758 -3895 -754 -3891
rect -742 -3895 -738 -3891
rect -577 -3895 -573 -3891
rect -568 -3895 -564 -3891
rect -559 -3895 -555 -3891
rect -551 -3895 -547 -3891
rect -535 -3895 -531 -3891
rect -527 -3895 -523 -3891
rect -510 -3895 -506 -3891
rect -493 -3895 -489 -3891
rect -485 -3895 -481 -3891
rect -468 -3895 -464 -3891
rect -451 -3895 -447 -3891
rect -443 -3895 -439 -3891
rect -426 -3895 -422 -3891
rect -409 -3895 -405 -3891
rect -401 -3895 -397 -3891
rect -385 -3895 -381 -3891
rect -219 -3895 -215 -3891
rect -210 -3895 -206 -3891
rect -201 -3895 -197 -3891
rect -193 -3895 -189 -3891
rect -177 -3895 -173 -3891
rect -169 -3895 -165 -3891
rect -152 -3895 -148 -3891
rect -135 -3895 -131 -3891
rect -127 -3895 -123 -3891
rect -110 -3895 -106 -3891
rect -93 -3895 -89 -3891
rect -85 -3895 -81 -3891
rect -68 -3895 -64 -3891
rect -51 -3895 -47 -3891
rect -43 -3895 -39 -3891
rect -27 -3895 -23 -3891
rect 139 -3895 143 -3891
rect 148 -3895 152 -3891
rect 157 -3895 161 -3891
rect 165 -3895 169 -3891
rect 181 -3895 185 -3891
rect 189 -3895 193 -3891
rect 206 -3895 210 -3891
rect 223 -3895 227 -3891
rect 231 -3895 235 -3891
rect 248 -3895 252 -3891
rect 265 -3895 269 -3891
rect 273 -3895 277 -3891
rect 290 -3895 294 -3891
rect 307 -3895 311 -3891
rect 315 -3895 319 -3891
rect 331 -3895 335 -3891
rect 495 -3895 499 -3891
rect 504 -3895 508 -3891
rect 513 -3895 517 -3891
rect 521 -3895 525 -3891
rect 537 -3895 541 -3891
rect 545 -3895 549 -3891
rect 562 -3895 566 -3891
rect 579 -3895 583 -3891
rect 587 -3895 591 -3891
rect 604 -3895 608 -3891
rect 621 -3895 625 -3891
rect 629 -3895 633 -3891
rect 646 -3895 650 -3891
rect 663 -3895 667 -3891
rect 671 -3895 675 -3891
rect 687 -3895 691 -3891
rect 853 -3895 857 -3891
rect 862 -3895 866 -3891
rect 871 -3895 875 -3891
rect 879 -3895 883 -3891
rect 895 -3895 899 -3891
rect 903 -3895 907 -3891
rect 920 -3895 924 -3891
rect 937 -3895 941 -3891
rect 945 -3895 949 -3891
rect 962 -3895 966 -3891
rect 979 -3895 983 -3891
rect 987 -3895 991 -3891
rect 1004 -3895 1008 -3891
rect 1021 -3895 1025 -3891
rect 1029 -3895 1033 -3891
rect 1045 -3895 1049 -3891
rect 1211 -3895 1215 -3891
rect 1220 -3895 1224 -3891
rect 1229 -3895 1233 -3891
rect 1237 -3895 1241 -3891
rect 1253 -3895 1257 -3891
rect 1261 -3895 1265 -3891
rect 1278 -3895 1282 -3891
rect 1295 -3895 1299 -3891
rect 1303 -3895 1307 -3891
rect 1320 -3895 1324 -3891
rect 1337 -3895 1341 -3891
rect 1345 -3895 1349 -3891
rect 1362 -3895 1366 -3891
rect 1379 -3895 1383 -3891
rect 1387 -3895 1391 -3891
rect 1403 -3895 1407 -3891
rect -1559 -4070 -1555 -4066
rect -1550 -4070 -1546 -4066
rect -1541 -4070 -1537 -4066
rect -1533 -4070 -1529 -4066
rect -1517 -4070 -1513 -4066
rect -1509 -4070 -1505 -4066
rect -1492 -4070 -1488 -4066
rect -1475 -4070 -1471 -4066
rect -1467 -4070 -1463 -4066
rect -1450 -4070 -1446 -4066
rect -1433 -4070 -1429 -4066
rect -1425 -4070 -1421 -4066
rect -1408 -4070 -1404 -4066
rect -1391 -4070 -1387 -4066
rect -1383 -4070 -1379 -4066
rect -1367 -4070 -1363 -4066
rect -1234 -4070 -1230 -4066
rect -1225 -4070 -1221 -4066
rect -1216 -4070 -1212 -4066
rect -1208 -4070 -1204 -4066
rect -1192 -4070 -1188 -4066
rect -1184 -4070 -1180 -4066
rect -1167 -4070 -1163 -4066
rect -1150 -4070 -1146 -4066
rect -1142 -4070 -1138 -4066
rect -1125 -4070 -1121 -4066
rect -1108 -4070 -1104 -4066
rect -1100 -4070 -1096 -4066
rect -1083 -4070 -1079 -4066
rect -1066 -4070 -1062 -4066
rect -1058 -4070 -1054 -4066
rect -1042 -4070 -1038 -4066
rect -935 -4070 -931 -4066
rect -926 -4070 -922 -4066
rect -917 -4070 -913 -4066
rect -909 -4070 -905 -4066
rect -893 -4070 -889 -4066
rect -885 -4070 -881 -4066
rect -868 -4070 -864 -4066
rect -851 -4070 -847 -4066
rect -843 -4070 -839 -4066
rect -826 -4070 -822 -4066
rect -809 -4070 -805 -4066
rect -801 -4070 -797 -4066
rect -784 -4070 -780 -4066
rect -767 -4070 -763 -4066
rect -759 -4070 -755 -4066
rect -743 -4070 -739 -4066
rect -577 -4070 -573 -4066
rect -568 -4070 -564 -4066
rect -559 -4070 -555 -4066
rect -551 -4070 -547 -4066
rect -535 -4070 -531 -4066
rect -527 -4070 -523 -4066
rect -510 -4070 -506 -4066
rect -493 -4070 -489 -4066
rect -485 -4070 -481 -4066
rect -468 -4070 -464 -4066
rect -451 -4070 -447 -4066
rect -443 -4070 -439 -4066
rect -426 -4070 -422 -4066
rect -409 -4070 -405 -4066
rect -401 -4070 -397 -4066
rect -385 -4070 -381 -4066
rect -219 -4070 -215 -4066
rect -210 -4070 -206 -4066
rect -201 -4070 -197 -4066
rect -193 -4070 -189 -4066
rect -177 -4070 -173 -4066
rect -169 -4070 -165 -4066
rect -152 -4070 -148 -4066
rect -135 -4070 -131 -4066
rect -127 -4070 -123 -4066
rect -110 -4070 -106 -4066
rect -93 -4070 -89 -4066
rect -85 -4070 -81 -4066
rect -68 -4070 -64 -4066
rect -51 -4070 -47 -4066
rect -43 -4070 -39 -4066
rect -27 -4070 -23 -4066
rect 139 -4070 143 -4066
rect 148 -4070 152 -4066
rect 157 -4070 161 -4066
rect 165 -4070 169 -4066
rect 181 -4070 185 -4066
rect 189 -4070 193 -4066
rect 206 -4070 210 -4066
rect 223 -4070 227 -4066
rect 231 -4070 235 -4066
rect 248 -4070 252 -4066
rect 265 -4070 269 -4066
rect 273 -4070 277 -4066
rect 290 -4070 294 -4066
rect 307 -4070 311 -4066
rect 315 -4070 319 -4066
rect 331 -4070 335 -4066
rect 495 -4070 499 -4066
rect 504 -4070 508 -4066
rect 513 -4070 517 -4066
rect 521 -4070 525 -4066
rect 537 -4070 541 -4066
rect 545 -4070 549 -4066
rect 562 -4070 566 -4066
rect 579 -4070 583 -4066
rect 587 -4070 591 -4066
rect 604 -4070 608 -4066
rect 621 -4070 625 -4066
rect 629 -4070 633 -4066
rect 646 -4070 650 -4066
rect 663 -4070 667 -4066
rect 671 -4070 675 -4066
rect 687 -4070 691 -4066
rect 853 -4070 857 -4066
rect 862 -4070 866 -4066
rect 871 -4070 875 -4066
rect 879 -4070 883 -4066
rect 895 -4070 899 -4066
rect 903 -4070 907 -4066
rect 920 -4070 924 -4066
rect 937 -4070 941 -4066
rect 945 -4070 949 -4066
rect 962 -4070 966 -4066
rect 979 -4070 983 -4066
rect 987 -4070 991 -4066
rect 1004 -4070 1008 -4066
rect 1021 -4070 1025 -4066
rect 1029 -4070 1033 -4066
rect 1045 -4070 1049 -4066
rect 1211 -4070 1215 -4066
rect 1220 -4070 1224 -4066
rect 1229 -4070 1233 -4066
rect 1237 -4070 1241 -4066
rect 1253 -4070 1257 -4066
rect 1261 -4070 1265 -4066
rect 1278 -4070 1282 -4066
rect 1295 -4070 1299 -4066
rect 1303 -4070 1307 -4066
rect 1320 -4070 1324 -4066
rect 1337 -4070 1341 -4066
rect 1345 -4070 1349 -4066
rect 1362 -4070 1366 -4066
rect 1379 -4070 1383 -4066
rect 1387 -4070 1391 -4066
rect 1403 -4070 1407 -4066
rect -1309 -4185 -1305 -4181
rect -1292 -4185 -1288 -4181
rect -1283 -4185 -1279 -4181
rect -935 -4185 -931 -4181
rect -918 -4185 -914 -4181
rect -909 -4185 -905 -4181
rect -577 -4185 -573 -4181
rect -560 -4185 -556 -4181
rect -551 -4185 -547 -4181
rect -219 -4185 -215 -4181
rect -202 -4185 -198 -4181
rect -193 -4185 -189 -4181
rect 139 -4185 143 -4181
rect 156 -4185 160 -4181
rect 165 -4185 169 -4181
rect 495 -4185 499 -4181
rect 512 -4185 516 -4181
rect 521 -4185 525 -4181
rect 853 -4185 857 -4181
rect 870 -4185 874 -4181
rect 879 -4185 883 -4181
rect 1211 -4185 1215 -4181
rect 1228 -4185 1232 -4181
rect 1237 -4185 1241 -4181
rect -1234 -4344 -1230 -4340
rect -1225 -4344 -1221 -4340
rect -1216 -4344 -1212 -4340
rect -1208 -4344 -1204 -4340
rect -1199 -4344 -1195 -4340
rect -1181 -4344 -1177 -4340
rect -1172 -4344 -1168 -4340
rect -1164 -4344 -1160 -4340
rect -1147 -4344 -1143 -4340
rect -1138 -4344 -1134 -4340
rect -935 -4344 -931 -4340
rect -926 -4344 -922 -4340
rect -917 -4344 -913 -4340
rect -909 -4344 -905 -4340
rect -900 -4344 -896 -4340
rect -891 -4344 -887 -4340
rect -883 -4344 -879 -4340
rect -875 -4344 -871 -4340
rect -857 -4344 -853 -4340
rect -847 -4344 -843 -4340
rect -839 -4344 -835 -4340
rect -822 -4344 -818 -4340
rect -813 -4344 -809 -4340
rect -805 -4344 -801 -4340
rect -796 -4344 -792 -4340
rect -778 -4344 -774 -4340
rect -769 -4344 -765 -4340
rect -761 -4344 -757 -4340
rect -745 -4344 -741 -4340
rect -737 -4344 -733 -4340
rect -725 -4344 -721 -4340
rect -713 -4344 -709 -4340
rect -704 -4344 -700 -4340
rect -695 -4344 -691 -4340
rect -577 -4344 -573 -4340
rect -568 -4344 -564 -4340
rect -559 -4344 -555 -4340
rect -551 -4344 -547 -4340
rect -542 -4344 -538 -4340
rect -533 -4344 -529 -4340
rect -525 -4344 -521 -4340
rect -517 -4344 -513 -4340
rect -499 -4344 -495 -4340
rect -489 -4344 -485 -4340
rect -481 -4344 -477 -4340
rect -464 -4344 -460 -4340
rect -455 -4344 -451 -4340
rect -447 -4344 -443 -4340
rect -438 -4344 -434 -4340
rect -420 -4344 -416 -4340
rect -411 -4344 -407 -4340
rect -403 -4344 -399 -4340
rect -387 -4344 -383 -4340
rect -379 -4344 -375 -4340
rect -367 -4344 -363 -4340
rect -355 -4344 -351 -4340
rect -346 -4344 -342 -4340
rect -337 -4344 -333 -4340
rect -219 -4344 -215 -4340
rect -210 -4344 -206 -4340
rect -201 -4344 -197 -4340
rect -193 -4344 -189 -4340
rect -184 -4344 -180 -4340
rect -175 -4344 -171 -4340
rect -167 -4344 -163 -4340
rect -159 -4344 -155 -4340
rect -141 -4344 -137 -4340
rect -131 -4344 -127 -4340
rect -123 -4344 -119 -4340
rect -106 -4344 -102 -4340
rect -97 -4344 -93 -4340
rect -89 -4344 -85 -4340
rect -80 -4344 -76 -4340
rect -62 -4344 -58 -4340
rect -53 -4344 -49 -4340
rect -45 -4344 -41 -4340
rect -29 -4344 -25 -4340
rect -21 -4344 -17 -4340
rect -9 -4344 -5 -4340
rect 3 -4344 7 -4340
rect 12 -4344 16 -4340
rect 21 -4344 25 -4340
rect 139 -4344 143 -4340
rect 148 -4344 152 -4340
rect 157 -4344 161 -4340
rect 165 -4344 169 -4340
rect 174 -4344 178 -4340
rect 183 -4344 187 -4340
rect 191 -4344 195 -4340
rect 199 -4344 203 -4340
rect 217 -4344 221 -4340
rect 227 -4344 231 -4340
rect 235 -4344 239 -4340
rect 252 -4344 256 -4340
rect 261 -4344 265 -4340
rect 269 -4344 273 -4340
rect 278 -4344 282 -4340
rect 296 -4344 300 -4340
rect 305 -4344 309 -4340
rect 313 -4344 317 -4340
rect 329 -4344 333 -4340
rect 337 -4344 341 -4340
rect 349 -4344 353 -4340
rect 361 -4344 365 -4340
rect 370 -4344 374 -4340
rect 379 -4344 383 -4340
rect 495 -4344 499 -4340
rect 504 -4344 508 -4340
rect 513 -4344 517 -4340
rect 521 -4344 525 -4340
rect 530 -4344 534 -4340
rect 539 -4344 543 -4340
rect 547 -4344 551 -4340
rect 555 -4344 559 -4340
rect 573 -4344 577 -4340
rect 583 -4344 587 -4340
rect 591 -4344 595 -4340
rect 608 -4344 612 -4340
rect 617 -4344 621 -4340
rect 625 -4344 629 -4340
rect 634 -4344 638 -4340
rect 652 -4344 656 -4340
rect 661 -4344 665 -4340
rect 669 -4344 673 -4340
rect 685 -4344 689 -4340
rect 693 -4344 697 -4340
rect 705 -4344 709 -4340
rect 717 -4344 721 -4340
rect 726 -4344 730 -4340
rect 735 -4344 739 -4340
rect 853 -4344 857 -4340
rect 862 -4344 866 -4340
rect 871 -4344 875 -4340
rect 879 -4344 883 -4340
rect 888 -4344 892 -4340
rect 897 -4344 901 -4340
rect 905 -4344 909 -4340
rect 913 -4344 917 -4340
rect 931 -4344 935 -4340
rect 941 -4344 945 -4340
rect 949 -4344 953 -4340
rect 966 -4344 970 -4340
rect 975 -4344 979 -4340
rect 983 -4344 987 -4340
rect 992 -4344 996 -4340
rect 1010 -4344 1014 -4340
rect 1019 -4344 1023 -4340
rect 1027 -4344 1031 -4340
rect 1043 -4344 1047 -4340
rect 1051 -4344 1055 -4340
rect 1063 -4344 1067 -4340
rect 1075 -4344 1079 -4340
rect 1084 -4344 1088 -4340
rect 1093 -4344 1097 -4340
rect 1211 -4344 1215 -4340
rect 1220 -4344 1224 -4340
rect 1229 -4344 1233 -4340
rect 1237 -4344 1241 -4340
rect 1246 -4344 1250 -4340
rect 1255 -4344 1259 -4340
rect 1263 -4344 1267 -4340
rect 1271 -4344 1275 -4340
rect 1289 -4344 1293 -4340
rect 1299 -4344 1303 -4340
rect 1307 -4344 1311 -4340
rect 1324 -4344 1328 -4340
rect 1333 -4344 1337 -4340
rect 1341 -4344 1345 -4340
rect 1350 -4344 1354 -4340
rect 1368 -4344 1372 -4340
rect 1377 -4344 1381 -4340
rect 1385 -4344 1389 -4340
rect 1401 -4344 1405 -4340
rect 1409 -4344 1413 -4340
rect 1421 -4344 1425 -4340
rect 1433 -4344 1437 -4340
rect 1442 -4344 1446 -4340
rect 1451 -4344 1455 -4340
rect -1814 -4467 -1810 -4463
rect -1805 -4467 -1801 -4463
rect -1796 -4467 -1792 -4463
rect -1788 -4467 -1784 -4463
rect -1772 -4467 -1768 -4463
rect -1764 -4467 -1760 -4463
rect -1747 -4467 -1743 -4463
rect -1730 -4467 -1726 -4463
rect -1722 -4467 -1718 -4463
rect -1705 -4467 -1701 -4463
rect -1688 -4467 -1684 -4463
rect -1680 -4467 -1676 -4463
rect -1663 -4467 -1659 -4463
rect -1646 -4467 -1642 -4463
rect -1638 -4467 -1634 -4463
rect -1622 -4467 -1618 -4463
rect -1551 -4467 -1547 -4463
rect -1542 -4467 -1538 -4463
rect -1533 -4467 -1529 -4463
rect -1525 -4467 -1521 -4463
rect -1509 -4467 -1505 -4463
rect -1501 -4467 -1497 -4463
rect -1484 -4467 -1480 -4463
rect -1467 -4467 -1463 -4463
rect -1459 -4467 -1455 -4463
rect -1442 -4467 -1438 -4463
rect -1425 -4467 -1421 -4463
rect -1417 -4467 -1413 -4463
rect -1400 -4467 -1396 -4463
rect -1383 -4467 -1379 -4463
rect -1375 -4467 -1371 -4463
rect -1359 -4467 -1355 -4463
rect -1234 -4467 -1230 -4463
rect -1225 -4467 -1221 -4463
rect -1216 -4467 -1212 -4463
rect -1208 -4467 -1204 -4463
rect -1192 -4467 -1188 -4463
rect -1184 -4467 -1180 -4463
rect -1167 -4467 -1163 -4463
rect -1150 -4467 -1146 -4463
rect -1142 -4467 -1138 -4463
rect -1125 -4467 -1121 -4463
rect -1108 -4467 -1104 -4463
rect -1100 -4467 -1096 -4463
rect -1083 -4467 -1079 -4463
rect -1066 -4467 -1062 -4463
rect -1058 -4467 -1054 -4463
rect -1042 -4467 -1038 -4463
rect -935 -4467 -931 -4463
rect -926 -4467 -922 -4463
rect -917 -4467 -913 -4463
rect -909 -4467 -905 -4463
rect -893 -4467 -889 -4463
rect -885 -4467 -881 -4463
rect -868 -4467 -864 -4463
rect -851 -4467 -847 -4463
rect -843 -4467 -839 -4463
rect -826 -4467 -822 -4463
rect -809 -4467 -805 -4463
rect -801 -4467 -797 -4463
rect -784 -4467 -780 -4463
rect -767 -4467 -763 -4463
rect -759 -4467 -755 -4463
rect -743 -4467 -739 -4463
rect -577 -4467 -573 -4463
rect -568 -4467 -564 -4463
rect -559 -4467 -555 -4463
rect -551 -4467 -547 -4463
rect -535 -4467 -531 -4463
rect -527 -4467 -523 -4463
rect -510 -4467 -506 -4463
rect -493 -4467 -489 -4463
rect -485 -4467 -481 -4463
rect -468 -4467 -464 -4463
rect -451 -4467 -447 -4463
rect -443 -4467 -439 -4463
rect -426 -4467 -422 -4463
rect -409 -4467 -405 -4463
rect -401 -4467 -397 -4463
rect -385 -4467 -381 -4463
rect -1814 -4638 -1810 -4634
rect -1805 -4638 -1801 -4634
rect -1796 -4638 -1792 -4634
rect -1788 -4638 -1784 -4634
rect -1772 -4638 -1768 -4634
rect -1764 -4638 -1760 -4634
rect -1747 -4638 -1743 -4634
rect -1730 -4638 -1726 -4634
rect -1722 -4638 -1718 -4634
rect -1705 -4638 -1701 -4634
rect -1688 -4638 -1684 -4634
rect -1680 -4638 -1676 -4634
rect -1663 -4638 -1659 -4634
rect -1646 -4638 -1642 -4634
rect -1638 -4638 -1634 -4634
rect -1622 -4638 -1618 -4634
rect -1551 -4638 -1547 -4634
rect -1542 -4638 -1538 -4634
rect -1533 -4638 -1529 -4634
rect -1525 -4638 -1521 -4634
rect -1509 -4638 -1505 -4634
rect -1501 -4638 -1497 -4634
rect -1484 -4638 -1480 -4634
rect -1467 -4638 -1463 -4634
rect -1459 -4638 -1455 -4634
rect -1442 -4638 -1438 -4634
rect -1425 -4638 -1421 -4634
rect -1417 -4638 -1413 -4634
rect -1400 -4638 -1396 -4634
rect -1383 -4638 -1379 -4634
rect -1375 -4638 -1371 -4634
rect -1359 -4638 -1355 -4634
rect -1234 -4638 -1230 -4634
rect -1225 -4638 -1221 -4634
rect -1216 -4638 -1212 -4634
rect -1208 -4638 -1204 -4634
rect -1192 -4638 -1188 -4634
rect -1184 -4638 -1180 -4634
rect -1167 -4638 -1163 -4634
rect -1150 -4638 -1146 -4634
rect -1142 -4638 -1138 -4634
rect -1125 -4638 -1121 -4634
rect -1108 -4638 -1104 -4634
rect -1100 -4638 -1096 -4634
rect -1083 -4638 -1079 -4634
rect -1066 -4638 -1062 -4634
rect -1058 -4638 -1054 -4634
rect -1042 -4638 -1038 -4634
rect -935 -4638 -931 -4634
rect -926 -4638 -922 -4634
rect -917 -4638 -913 -4634
rect -909 -4638 -905 -4634
rect -893 -4638 -889 -4634
rect -885 -4638 -881 -4634
rect -868 -4638 -864 -4634
rect -851 -4638 -847 -4634
rect -843 -4638 -839 -4634
rect -826 -4638 -822 -4634
rect -809 -4638 -805 -4634
rect -801 -4638 -797 -4634
rect -784 -4638 -780 -4634
rect -767 -4638 -763 -4634
rect -759 -4638 -755 -4634
rect -743 -4638 -739 -4634
rect -577 -4638 -573 -4634
rect -568 -4638 -564 -4634
rect -559 -4638 -555 -4634
rect -551 -4638 -547 -4634
rect -535 -4638 -531 -4634
rect -527 -4638 -523 -4634
rect -510 -4638 -506 -4634
rect -493 -4638 -489 -4634
rect -485 -4638 -481 -4634
rect -468 -4638 -464 -4634
rect -451 -4638 -447 -4634
rect -443 -4638 -439 -4634
rect -426 -4638 -422 -4634
rect -409 -4638 -405 -4634
rect -401 -4638 -397 -4634
rect -385 -4638 -381 -4634
rect -219 -4638 -215 -4634
rect -210 -4638 -206 -4634
rect -201 -4638 -197 -4634
rect -193 -4638 -189 -4634
rect -177 -4638 -173 -4634
rect -169 -4638 -165 -4634
rect -152 -4638 -148 -4634
rect -135 -4638 -131 -4634
rect -127 -4638 -123 -4634
rect -110 -4638 -106 -4634
rect -93 -4638 -89 -4634
rect -85 -4638 -81 -4634
rect -68 -4638 -64 -4634
rect -51 -4638 -47 -4634
rect -43 -4638 -39 -4634
rect -27 -4638 -23 -4634
rect 139 -4638 143 -4634
rect 148 -4638 152 -4634
rect 157 -4638 161 -4634
rect 165 -4638 169 -4634
rect 181 -4638 185 -4634
rect 189 -4638 193 -4634
rect 206 -4638 210 -4634
rect 223 -4638 227 -4634
rect 231 -4638 235 -4634
rect 248 -4638 252 -4634
rect 265 -4638 269 -4634
rect 273 -4638 277 -4634
rect 290 -4638 294 -4634
rect 307 -4638 311 -4634
rect 315 -4638 319 -4634
rect 331 -4638 335 -4634
rect 495 -4638 499 -4634
rect 504 -4638 508 -4634
rect 513 -4638 517 -4634
rect 521 -4638 525 -4634
rect 537 -4638 541 -4634
rect 545 -4638 549 -4634
rect 562 -4638 566 -4634
rect 579 -4638 583 -4634
rect 587 -4638 591 -4634
rect 604 -4638 608 -4634
rect 621 -4638 625 -4634
rect 629 -4638 633 -4634
rect 646 -4638 650 -4634
rect 663 -4638 667 -4634
rect 671 -4638 675 -4634
rect 687 -4638 691 -4634
rect 853 -4638 857 -4634
rect 862 -4638 866 -4634
rect 871 -4638 875 -4634
rect 879 -4638 883 -4634
rect 895 -4638 899 -4634
rect 903 -4638 907 -4634
rect 920 -4638 924 -4634
rect 937 -4638 941 -4634
rect 945 -4638 949 -4634
rect 962 -4638 966 -4634
rect 979 -4638 983 -4634
rect 987 -4638 991 -4634
rect 1004 -4638 1008 -4634
rect 1021 -4638 1025 -4634
rect 1029 -4638 1033 -4634
rect 1045 -4638 1049 -4634
rect 1211 -4638 1215 -4634
rect 1220 -4638 1224 -4634
rect 1229 -4638 1233 -4634
rect 1237 -4638 1241 -4634
rect 1253 -4638 1257 -4634
rect 1261 -4638 1265 -4634
rect 1278 -4638 1282 -4634
rect 1295 -4638 1299 -4634
rect 1303 -4638 1307 -4634
rect 1320 -4638 1324 -4634
rect 1337 -4638 1341 -4634
rect 1345 -4638 1349 -4634
rect 1362 -4638 1366 -4634
rect 1379 -4638 1383 -4634
rect 1387 -4638 1391 -4634
rect 1403 -4638 1407 -4634
rect -1551 -4809 -1547 -4805
rect -1542 -4809 -1538 -4805
rect -1533 -4809 -1529 -4805
rect -1525 -4809 -1521 -4805
rect -1509 -4809 -1505 -4805
rect -1501 -4809 -1497 -4805
rect -1484 -4809 -1480 -4805
rect -1467 -4809 -1463 -4805
rect -1459 -4809 -1455 -4805
rect -1442 -4809 -1438 -4805
rect -1425 -4809 -1421 -4805
rect -1417 -4809 -1413 -4805
rect -1400 -4809 -1396 -4805
rect -1383 -4809 -1379 -4805
rect -1375 -4809 -1371 -4805
rect -1359 -4809 -1355 -4805
rect -1234 -4809 -1230 -4805
rect -1225 -4809 -1221 -4805
rect -1216 -4809 -1212 -4805
rect -1208 -4809 -1204 -4805
rect -1192 -4809 -1188 -4805
rect -1184 -4809 -1180 -4805
rect -1167 -4809 -1163 -4805
rect -1150 -4809 -1146 -4805
rect -1142 -4809 -1138 -4805
rect -1125 -4809 -1121 -4805
rect -1108 -4809 -1104 -4805
rect -1100 -4809 -1096 -4805
rect -1083 -4809 -1079 -4805
rect -1066 -4809 -1062 -4805
rect -1058 -4809 -1054 -4805
rect -1042 -4809 -1038 -4805
rect -935 -4809 -931 -4805
rect -926 -4809 -922 -4805
rect -917 -4809 -913 -4805
rect -909 -4809 -905 -4805
rect -893 -4809 -889 -4805
rect -885 -4809 -881 -4805
rect -868 -4809 -864 -4805
rect -851 -4809 -847 -4805
rect -843 -4809 -839 -4805
rect -826 -4809 -822 -4805
rect -809 -4809 -805 -4805
rect -801 -4809 -797 -4805
rect -784 -4809 -780 -4805
rect -767 -4809 -763 -4805
rect -759 -4809 -755 -4805
rect -743 -4809 -739 -4805
rect -577 -4809 -573 -4805
rect -568 -4809 -564 -4805
rect -559 -4809 -555 -4805
rect -551 -4809 -547 -4805
rect -535 -4809 -531 -4805
rect -527 -4809 -523 -4805
rect -510 -4809 -506 -4805
rect -493 -4809 -489 -4805
rect -485 -4809 -481 -4805
rect -468 -4809 -464 -4805
rect -451 -4809 -447 -4805
rect -443 -4809 -439 -4805
rect -426 -4809 -422 -4805
rect -409 -4809 -405 -4805
rect -401 -4809 -397 -4805
rect -385 -4809 -381 -4805
rect -219 -4809 -215 -4805
rect -210 -4809 -206 -4805
rect -201 -4809 -197 -4805
rect -193 -4809 -189 -4805
rect -177 -4809 -173 -4805
rect -169 -4809 -165 -4805
rect -152 -4809 -148 -4805
rect -135 -4809 -131 -4805
rect -127 -4809 -123 -4805
rect -110 -4809 -106 -4805
rect -93 -4809 -89 -4805
rect -85 -4809 -81 -4805
rect -68 -4809 -64 -4805
rect -51 -4809 -47 -4805
rect -43 -4809 -39 -4805
rect -27 -4809 -23 -4805
rect 139 -4809 143 -4805
rect 148 -4809 152 -4805
rect 157 -4809 161 -4805
rect 165 -4809 169 -4805
rect 181 -4809 185 -4805
rect 189 -4809 193 -4805
rect 206 -4809 210 -4805
rect 223 -4809 227 -4805
rect 231 -4809 235 -4805
rect 248 -4809 252 -4805
rect 265 -4809 269 -4805
rect 273 -4809 277 -4805
rect 290 -4809 294 -4805
rect 307 -4809 311 -4805
rect 315 -4809 319 -4805
rect 331 -4809 335 -4805
rect 495 -4809 499 -4805
rect 504 -4809 508 -4805
rect 513 -4809 517 -4805
rect 521 -4809 525 -4805
rect 537 -4809 541 -4805
rect 545 -4809 549 -4805
rect 562 -4809 566 -4805
rect 579 -4809 583 -4805
rect 587 -4809 591 -4805
rect 604 -4809 608 -4805
rect 621 -4809 625 -4805
rect 629 -4809 633 -4805
rect 646 -4809 650 -4805
rect 663 -4809 667 -4805
rect 671 -4809 675 -4805
rect 687 -4809 691 -4805
rect 853 -4809 857 -4805
rect 862 -4809 866 -4805
rect 871 -4809 875 -4805
rect 879 -4809 883 -4805
rect 895 -4809 899 -4805
rect 903 -4809 907 -4805
rect 920 -4809 924 -4805
rect 937 -4809 941 -4805
rect 945 -4809 949 -4805
rect 962 -4809 966 -4805
rect 979 -4809 983 -4805
rect 987 -4809 991 -4805
rect 1004 -4809 1008 -4805
rect 1021 -4809 1025 -4805
rect 1029 -4809 1033 -4805
rect 1045 -4809 1049 -4805
rect 1211 -4809 1215 -4805
rect 1220 -4809 1224 -4805
rect 1229 -4809 1233 -4805
rect 1237 -4809 1241 -4805
rect 1253 -4809 1257 -4805
rect 1261 -4809 1265 -4805
rect 1278 -4809 1282 -4805
rect 1295 -4809 1299 -4805
rect 1303 -4809 1307 -4805
rect 1320 -4809 1324 -4805
rect 1337 -4809 1341 -4805
rect 1345 -4809 1349 -4805
rect 1362 -4809 1366 -4805
rect 1379 -4809 1383 -4805
rect 1387 -4809 1391 -4805
rect 1403 -4809 1407 -4805
rect -1309 -4924 -1305 -4920
rect -1292 -4924 -1288 -4920
rect -1283 -4924 -1279 -4920
rect -935 -4924 -931 -4920
rect -918 -4924 -914 -4920
rect -909 -4924 -905 -4920
rect -577 -4924 -573 -4920
rect -560 -4924 -556 -4920
rect -551 -4924 -547 -4920
rect -219 -4924 -215 -4920
rect -202 -4924 -198 -4920
rect -193 -4924 -189 -4920
rect 139 -4924 143 -4920
rect 156 -4924 160 -4920
rect 165 -4924 169 -4920
rect 495 -4924 499 -4920
rect 512 -4924 516 -4920
rect 521 -4924 525 -4920
rect 853 -4924 857 -4920
rect 870 -4924 874 -4920
rect 879 -4924 883 -4920
rect 1211 -4924 1215 -4920
rect 1228 -4924 1232 -4920
rect 1237 -4924 1241 -4920
rect -1234 -5083 -1230 -5079
rect -1225 -5083 -1221 -5079
rect -1216 -5083 -1212 -5079
rect -1208 -5083 -1204 -5079
rect -1199 -5083 -1195 -5079
rect -1181 -5083 -1177 -5079
rect -1172 -5083 -1168 -5079
rect -1164 -5083 -1160 -5079
rect -1147 -5083 -1143 -5079
rect -1138 -5083 -1134 -5079
rect -935 -5083 -931 -5079
rect -926 -5083 -922 -5079
rect -917 -5083 -913 -5079
rect -909 -5083 -905 -5079
rect -900 -5083 -896 -5079
rect -891 -5083 -887 -5079
rect -883 -5083 -879 -5079
rect -875 -5083 -871 -5079
rect -857 -5083 -853 -5079
rect -847 -5083 -843 -5079
rect -839 -5083 -835 -5079
rect -822 -5083 -818 -5079
rect -813 -5083 -809 -5079
rect -805 -5083 -801 -5079
rect -796 -5083 -792 -5079
rect -778 -5083 -774 -5079
rect -769 -5083 -765 -5079
rect -761 -5083 -757 -5079
rect -745 -5083 -741 -5079
rect -737 -5083 -733 -5079
rect -725 -5083 -721 -5079
rect -713 -5083 -709 -5079
rect -704 -5083 -700 -5079
rect -695 -5083 -691 -5079
rect -577 -5083 -573 -5079
rect -568 -5083 -564 -5079
rect -559 -5083 -555 -5079
rect -551 -5083 -547 -5079
rect -542 -5083 -538 -5079
rect -533 -5083 -529 -5079
rect -525 -5083 -521 -5079
rect -517 -5083 -513 -5079
rect -499 -5083 -495 -5079
rect -489 -5083 -485 -5079
rect -481 -5083 -477 -5079
rect -464 -5083 -460 -5079
rect -455 -5083 -451 -5079
rect -447 -5083 -443 -5079
rect -438 -5083 -434 -5079
rect -420 -5083 -416 -5079
rect -411 -5083 -407 -5079
rect -403 -5083 -399 -5079
rect -387 -5083 -383 -5079
rect -379 -5083 -375 -5079
rect -367 -5083 -363 -5079
rect -355 -5083 -351 -5079
rect -346 -5083 -342 -5079
rect -337 -5083 -333 -5079
rect -219 -5083 -215 -5079
rect -210 -5083 -206 -5079
rect -201 -5083 -197 -5079
rect -193 -5083 -189 -5079
rect -184 -5083 -180 -5079
rect -175 -5083 -171 -5079
rect -167 -5083 -163 -5079
rect -159 -5083 -155 -5079
rect -141 -5083 -137 -5079
rect -131 -5083 -127 -5079
rect -123 -5083 -119 -5079
rect -106 -5083 -102 -5079
rect -97 -5083 -93 -5079
rect -89 -5083 -85 -5079
rect -80 -5083 -76 -5079
rect -62 -5083 -58 -5079
rect -53 -5083 -49 -5079
rect -45 -5083 -41 -5079
rect -29 -5083 -25 -5079
rect -21 -5083 -17 -5079
rect -9 -5083 -5 -5079
rect 3 -5083 7 -5079
rect 12 -5083 16 -5079
rect 21 -5083 25 -5079
rect 139 -5083 143 -5079
rect 148 -5083 152 -5079
rect 157 -5083 161 -5079
rect 165 -5083 169 -5079
rect 174 -5083 178 -5079
rect 183 -5083 187 -5079
rect 191 -5083 195 -5079
rect 199 -5083 203 -5079
rect 217 -5083 221 -5079
rect 227 -5083 231 -5079
rect 235 -5083 239 -5079
rect 252 -5083 256 -5079
rect 261 -5083 265 -5079
rect 269 -5083 273 -5079
rect 278 -5083 282 -5079
rect 296 -5083 300 -5079
rect 305 -5083 309 -5079
rect 313 -5083 317 -5079
rect 329 -5083 333 -5079
rect 337 -5083 341 -5079
rect 349 -5083 353 -5079
rect 361 -5083 365 -5079
rect 370 -5083 374 -5079
rect 379 -5083 383 -5079
rect 495 -5083 499 -5079
rect 504 -5083 508 -5079
rect 513 -5083 517 -5079
rect 521 -5083 525 -5079
rect 530 -5083 534 -5079
rect 539 -5083 543 -5079
rect 547 -5083 551 -5079
rect 555 -5083 559 -5079
rect 573 -5083 577 -5079
rect 583 -5083 587 -5079
rect 591 -5083 595 -5079
rect 608 -5083 612 -5079
rect 617 -5083 621 -5079
rect 625 -5083 629 -5079
rect 634 -5083 638 -5079
rect 652 -5083 656 -5079
rect 661 -5083 665 -5079
rect 669 -5083 673 -5079
rect 685 -5083 689 -5079
rect 693 -5083 697 -5079
rect 705 -5083 709 -5079
rect 717 -5083 721 -5079
rect 726 -5083 730 -5079
rect 735 -5083 739 -5079
rect 853 -5083 857 -5079
rect 862 -5083 866 -5079
rect 871 -5083 875 -5079
rect 879 -5083 883 -5079
rect 888 -5083 892 -5079
rect 897 -5083 901 -5079
rect 905 -5083 909 -5079
rect 913 -5083 917 -5079
rect 931 -5083 935 -5079
rect 941 -5083 945 -5079
rect 949 -5083 953 -5079
rect 966 -5083 970 -5079
rect 975 -5083 979 -5079
rect 983 -5083 987 -5079
rect 992 -5083 996 -5079
rect 1010 -5083 1014 -5079
rect 1019 -5083 1023 -5079
rect 1027 -5083 1031 -5079
rect 1043 -5083 1047 -5079
rect 1051 -5083 1055 -5079
rect 1063 -5083 1067 -5079
rect 1075 -5083 1079 -5079
rect 1084 -5083 1088 -5079
rect 1093 -5083 1097 -5079
rect 1211 -5083 1215 -5079
rect 1220 -5083 1224 -5079
rect 1229 -5083 1233 -5079
rect 1237 -5083 1241 -5079
rect 1246 -5083 1250 -5079
rect 1255 -5083 1259 -5079
rect 1263 -5083 1267 -5079
rect 1271 -5083 1275 -5079
rect 1289 -5083 1293 -5079
rect 1299 -5083 1303 -5079
rect 1307 -5083 1311 -5079
rect 1324 -5083 1328 -5079
rect 1333 -5083 1337 -5079
rect 1341 -5083 1345 -5079
rect 1350 -5083 1354 -5079
rect 1368 -5083 1372 -5079
rect 1377 -5083 1381 -5079
rect 1385 -5083 1389 -5079
rect 1401 -5083 1405 -5079
rect 1409 -5083 1413 -5079
rect 1421 -5083 1425 -5079
rect 1433 -5083 1437 -5079
rect 1442 -5083 1446 -5079
rect 1451 -5083 1455 -5079
rect -1810 -5202 -1806 -5198
rect -1801 -5202 -1797 -5198
rect -1792 -5202 -1788 -5198
rect -1784 -5202 -1780 -5198
rect -1768 -5202 -1764 -5198
rect -1760 -5202 -1756 -5198
rect -1743 -5202 -1739 -5198
rect -1726 -5202 -1722 -5198
rect -1718 -5202 -1714 -5198
rect -1701 -5202 -1697 -5198
rect -1684 -5202 -1680 -5198
rect -1676 -5202 -1672 -5198
rect -1659 -5202 -1655 -5198
rect -1642 -5202 -1638 -5198
rect -1634 -5202 -1630 -5198
rect -1618 -5202 -1614 -5198
rect -1547 -5202 -1543 -5198
rect -1538 -5202 -1534 -5198
rect -1529 -5202 -1525 -5198
rect -1521 -5202 -1517 -5198
rect -1505 -5202 -1501 -5198
rect -1497 -5202 -1493 -5198
rect -1480 -5202 -1476 -5198
rect -1463 -5202 -1459 -5198
rect -1455 -5202 -1451 -5198
rect -1438 -5202 -1434 -5198
rect -1421 -5202 -1417 -5198
rect -1413 -5202 -1409 -5198
rect -1396 -5202 -1392 -5198
rect -1379 -5202 -1375 -5198
rect -1371 -5202 -1367 -5198
rect -1355 -5202 -1351 -5198
rect -1234 -5202 -1230 -5198
rect -1225 -5202 -1221 -5198
rect -1216 -5202 -1212 -5198
rect -1208 -5202 -1204 -5198
rect -1192 -5202 -1188 -5198
rect -1184 -5202 -1180 -5198
rect -1167 -5202 -1163 -5198
rect -1150 -5202 -1146 -5198
rect -1142 -5202 -1138 -5198
rect -1125 -5202 -1121 -5198
rect -1108 -5202 -1104 -5198
rect -1100 -5202 -1096 -5198
rect -1083 -5202 -1079 -5198
rect -1066 -5202 -1062 -5198
rect -1058 -5202 -1054 -5198
rect -1042 -5202 -1038 -5198
rect -935 -5202 -931 -5198
rect -926 -5202 -922 -5198
rect -917 -5202 -913 -5198
rect -909 -5202 -905 -5198
rect -893 -5202 -889 -5198
rect -885 -5202 -881 -5198
rect -868 -5202 -864 -5198
rect -851 -5202 -847 -5198
rect -843 -5202 -839 -5198
rect -826 -5202 -822 -5198
rect -809 -5202 -805 -5198
rect -801 -5202 -797 -5198
rect -784 -5202 -780 -5198
rect -767 -5202 -763 -5198
rect -759 -5202 -755 -5198
rect -743 -5202 -739 -5198
rect -1810 -5373 -1806 -5369
rect -1801 -5373 -1797 -5369
rect -1792 -5373 -1788 -5369
rect -1784 -5373 -1780 -5369
rect -1768 -5373 -1764 -5369
rect -1760 -5373 -1756 -5369
rect -1743 -5373 -1739 -5369
rect -1726 -5373 -1722 -5369
rect -1718 -5373 -1714 -5369
rect -1701 -5373 -1697 -5369
rect -1684 -5373 -1680 -5369
rect -1676 -5373 -1672 -5369
rect -1659 -5373 -1655 -5369
rect -1642 -5373 -1638 -5369
rect -1634 -5373 -1630 -5369
rect -1618 -5373 -1614 -5369
rect -1547 -5373 -1543 -5369
rect -1538 -5373 -1534 -5369
rect -1529 -5373 -1525 -5369
rect -1521 -5373 -1517 -5369
rect -1505 -5373 -1501 -5369
rect -1497 -5373 -1493 -5369
rect -1480 -5373 -1476 -5369
rect -1463 -5373 -1459 -5369
rect -1455 -5373 -1451 -5369
rect -1438 -5373 -1434 -5369
rect -1421 -5373 -1417 -5369
rect -1413 -5373 -1409 -5369
rect -1396 -5373 -1392 -5369
rect -1379 -5373 -1375 -5369
rect -1371 -5373 -1367 -5369
rect -1355 -5373 -1351 -5369
rect -1234 -5373 -1230 -5369
rect -1225 -5373 -1221 -5369
rect -1216 -5373 -1212 -5369
rect -1208 -5373 -1204 -5369
rect -1192 -5373 -1188 -5369
rect -1184 -5373 -1180 -5369
rect -1167 -5373 -1163 -5369
rect -1150 -5373 -1146 -5369
rect -1142 -5373 -1138 -5369
rect -1125 -5373 -1121 -5369
rect -1108 -5373 -1104 -5369
rect -1100 -5373 -1096 -5369
rect -1083 -5373 -1079 -5369
rect -1066 -5373 -1062 -5369
rect -1058 -5373 -1054 -5369
rect -1042 -5373 -1038 -5369
rect -935 -5373 -931 -5369
rect -926 -5373 -922 -5369
rect -917 -5373 -913 -5369
rect -909 -5373 -905 -5369
rect -893 -5373 -889 -5369
rect -885 -5373 -881 -5369
rect -868 -5373 -864 -5369
rect -851 -5373 -847 -5369
rect -843 -5373 -839 -5369
rect -826 -5373 -822 -5369
rect -809 -5373 -805 -5369
rect -801 -5373 -797 -5369
rect -784 -5373 -780 -5369
rect -767 -5373 -763 -5369
rect -759 -5373 -755 -5369
rect -743 -5373 -739 -5369
rect -577 -5373 -573 -5369
rect -568 -5373 -564 -5369
rect -559 -5373 -555 -5369
rect -551 -5373 -547 -5369
rect -535 -5373 -531 -5369
rect -527 -5373 -523 -5369
rect -510 -5373 -506 -5369
rect -493 -5373 -489 -5369
rect -485 -5373 -481 -5369
rect -468 -5373 -464 -5369
rect -451 -5373 -447 -5369
rect -443 -5373 -439 -5369
rect -426 -5373 -422 -5369
rect -409 -5373 -405 -5369
rect -401 -5373 -397 -5369
rect -385 -5373 -381 -5369
rect -219 -5373 -215 -5369
rect -210 -5373 -206 -5369
rect -201 -5373 -197 -5369
rect -193 -5373 -189 -5369
rect -177 -5373 -173 -5369
rect -169 -5373 -165 -5369
rect -152 -5373 -148 -5369
rect -135 -5373 -131 -5369
rect -127 -5373 -123 -5369
rect -110 -5373 -106 -5369
rect -93 -5373 -89 -5369
rect -85 -5373 -81 -5369
rect -68 -5373 -64 -5369
rect -51 -5373 -47 -5369
rect -43 -5373 -39 -5369
rect -27 -5373 -23 -5369
rect 139 -5373 143 -5369
rect 148 -5373 152 -5369
rect 157 -5373 161 -5369
rect 165 -5373 169 -5369
rect 181 -5373 185 -5369
rect 189 -5373 193 -5369
rect 206 -5373 210 -5369
rect 223 -5373 227 -5369
rect 231 -5373 235 -5369
rect 248 -5373 252 -5369
rect 265 -5373 269 -5369
rect 273 -5373 277 -5369
rect 290 -5373 294 -5369
rect 307 -5373 311 -5369
rect 315 -5373 319 -5369
rect 331 -5373 335 -5369
rect 495 -5373 499 -5369
rect 504 -5373 508 -5369
rect 513 -5373 517 -5369
rect 521 -5373 525 -5369
rect 537 -5373 541 -5369
rect 545 -5373 549 -5369
rect 562 -5373 566 -5369
rect 579 -5373 583 -5369
rect 587 -5373 591 -5369
rect 604 -5373 608 -5369
rect 621 -5373 625 -5369
rect 629 -5373 633 -5369
rect 646 -5373 650 -5369
rect 663 -5373 667 -5369
rect 671 -5373 675 -5369
rect 687 -5373 691 -5369
rect 853 -5373 857 -5369
rect 862 -5373 866 -5369
rect 871 -5373 875 -5369
rect 879 -5373 883 -5369
rect 895 -5373 899 -5369
rect 903 -5373 907 -5369
rect 920 -5373 924 -5369
rect 937 -5373 941 -5369
rect 945 -5373 949 -5369
rect 962 -5373 966 -5369
rect 979 -5373 983 -5369
rect 987 -5373 991 -5369
rect 1004 -5373 1008 -5369
rect 1021 -5373 1025 -5369
rect 1029 -5373 1033 -5369
rect 1045 -5373 1049 -5369
rect 1211 -5373 1215 -5369
rect 1220 -5373 1224 -5369
rect 1229 -5373 1233 -5369
rect 1237 -5373 1241 -5369
rect 1253 -5373 1257 -5369
rect 1261 -5373 1265 -5369
rect 1278 -5373 1282 -5369
rect 1295 -5373 1299 -5369
rect 1303 -5373 1307 -5369
rect 1320 -5373 1324 -5369
rect 1337 -5373 1341 -5369
rect 1345 -5373 1349 -5369
rect 1362 -5373 1366 -5369
rect 1379 -5373 1383 -5369
rect 1387 -5373 1391 -5369
rect 1403 -5373 1407 -5369
rect -1810 -5533 -1806 -5529
rect -1801 -5533 -1797 -5529
rect -1792 -5533 -1788 -5529
rect -1784 -5533 -1780 -5529
rect -1768 -5533 -1764 -5529
rect -1760 -5533 -1756 -5529
rect -1743 -5533 -1739 -5529
rect -1726 -5533 -1722 -5529
rect -1718 -5533 -1714 -5529
rect -1701 -5533 -1697 -5529
rect -1684 -5533 -1680 -5529
rect -1676 -5533 -1672 -5529
rect -1659 -5533 -1655 -5529
rect -1642 -5533 -1638 -5529
rect -1634 -5533 -1630 -5529
rect -1618 -5533 -1614 -5529
rect -1547 -5533 -1543 -5529
rect -1538 -5533 -1534 -5529
rect -1529 -5533 -1525 -5529
rect -1521 -5533 -1517 -5529
rect -1505 -5533 -1501 -5529
rect -1497 -5533 -1493 -5529
rect -1480 -5533 -1476 -5529
rect -1463 -5533 -1459 -5529
rect -1455 -5533 -1451 -5529
rect -1438 -5533 -1434 -5529
rect -1421 -5533 -1417 -5529
rect -1413 -5533 -1409 -5529
rect -1396 -5533 -1392 -5529
rect -1379 -5533 -1375 -5529
rect -1371 -5533 -1367 -5529
rect -1355 -5533 -1351 -5529
rect -1234 -5533 -1230 -5529
rect -1225 -5533 -1221 -5529
rect -1216 -5533 -1212 -5529
rect -1208 -5533 -1204 -5529
rect -1192 -5533 -1188 -5529
rect -1184 -5533 -1180 -5529
rect -1167 -5533 -1163 -5529
rect -1150 -5533 -1146 -5529
rect -1142 -5533 -1138 -5529
rect -1125 -5533 -1121 -5529
rect -1108 -5533 -1104 -5529
rect -1100 -5533 -1096 -5529
rect -1083 -5533 -1079 -5529
rect -1066 -5533 -1062 -5529
rect -1058 -5533 -1054 -5529
rect -1042 -5533 -1038 -5529
rect -935 -5533 -931 -5529
rect -926 -5533 -922 -5529
rect -917 -5533 -913 -5529
rect -909 -5533 -905 -5529
rect -893 -5533 -889 -5529
rect -885 -5533 -881 -5529
rect -868 -5533 -864 -5529
rect -851 -5533 -847 -5529
rect -843 -5533 -839 -5529
rect -826 -5533 -822 -5529
rect -809 -5533 -805 -5529
rect -801 -5533 -797 -5529
rect -784 -5533 -780 -5529
rect -767 -5533 -763 -5529
rect -759 -5533 -755 -5529
rect -743 -5533 -739 -5529
rect -577 -5533 -573 -5529
rect -568 -5533 -564 -5529
rect -559 -5533 -555 -5529
rect -551 -5533 -547 -5529
rect -535 -5533 -531 -5529
rect -527 -5533 -523 -5529
rect -510 -5533 -506 -5529
rect -493 -5533 -489 -5529
rect -485 -5533 -481 -5529
rect -468 -5533 -464 -5529
rect -451 -5533 -447 -5529
rect -443 -5533 -439 -5529
rect -426 -5533 -422 -5529
rect -409 -5533 -405 -5529
rect -401 -5533 -397 -5529
rect -385 -5533 -381 -5529
rect -219 -5533 -215 -5529
rect -210 -5533 -206 -5529
rect -201 -5533 -197 -5529
rect -193 -5533 -189 -5529
rect -177 -5533 -173 -5529
rect -169 -5533 -165 -5529
rect -152 -5533 -148 -5529
rect -135 -5533 -131 -5529
rect -127 -5533 -123 -5529
rect -110 -5533 -106 -5529
rect -93 -5533 -89 -5529
rect -85 -5533 -81 -5529
rect -68 -5533 -64 -5529
rect -51 -5533 -47 -5529
rect -43 -5533 -39 -5529
rect -27 -5533 -23 -5529
rect 139 -5533 143 -5529
rect 148 -5533 152 -5529
rect 157 -5533 161 -5529
rect 165 -5533 169 -5529
rect 181 -5533 185 -5529
rect 189 -5533 193 -5529
rect 206 -5533 210 -5529
rect 223 -5533 227 -5529
rect 231 -5533 235 -5529
rect 248 -5533 252 -5529
rect 265 -5533 269 -5529
rect 273 -5533 277 -5529
rect 290 -5533 294 -5529
rect 307 -5533 311 -5529
rect 315 -5533 319 -5529
rect 331 -5533 335 -5529
rect 495 -5533 499 -5529
rect 504 -5533 508 -5529
rect 513 -5533 517 -5529
rect 521 -5533 525 -5529
rect 537 -5533 541 -5529
rect 545 -5533 549 -5529
rect 562 -5533 566 -5529
rect 579 -5533 583 -5529
rect 587 -5533 591 -5529
rect 604 -5533 608 -5529
rect 621 -5533 625 -5529
rect 629 -5533 633 -5529
rect 646 -5533 650 -5529
rect 663 -5533 667 -5529
rect 671 -5533 675 -5529
rect 687 -5533 691 -5529
rect 853 -5533 857 -5529
rect 862 -5533 866 -5529
rect 871 -5533 875 -5529
rect 879 -5533 883 -5529
rect 895 -5533 899 -5529
rect 903 -5533 907 -5529
rect 920 -5533 924 -5529
rect 937 -5533 941 -5529
rect 945 -5533 949 -5529
rect 962 -5533 966 -5529
rect 979 -5533 983 -5529
rect 987 -5533 991 -5529
rect 1004 -5533 1008 -5529
rect 1021 -5533 1025 -5529
rect 1029 -5533 1033 -5529
rect 1045 -5533 1049 -5529
rect 1211 -5533 1215 -5529
rect 1220 -5533 1224 -5529
rect 1229 -5533 1233 -5529
rect 1237 -5533 1241 -5529
rect 1253 -5533 1257 -5529
rect 1261 -5533 1265 -5529
rect 1278 -5533 1282 -5529
rect 1295 -5533 1299 -5529
rect 1303 -5533 1307 -5529
rect 1320 -5533 1324 -5529
rect 1337 -5533 1341 -5529
rect 1345 -5533 1349 -5529
rect 1362 -5533 1366 -5529
rect 1379 -5533 1383 -5529
rect 1387 -5533 1391 -5529
rect 1403 -5533 1407 -5529
rect -1309 -5647 -1305 -5643
rect -1292 -5647 -1288 -5643
rect -1283 -5647 -1279 -5643
rect -935 -5647 -931 -5643
rect -918 -5647 -914 -5643
rect -909 -5647 -905 -5643
rect -577 -5647 -573 -5643
rect -560 -5647 -556 -5643
rect -551 -5647 -547 -5643
rect -219 -5647 -215 -5643
rect -202 -5647 -198 -5643
rect -193 -5647 -189 -5643
rect 139 -5647 143 -5643
rect 156 -5647 160 -5643
rect 165 -5647 169 -5643
rect 495 -5647 499 -5643
rect 512 -5647 516 -5643
rect 521 -5647 525 -5643
rect 853 -5647 857 -5643
rect 870 -5647 874 -5643
rect 879 -5647 883 -5643
rect 1211 -5647 1215 -5643
rect 1228 -5647 1232 -5643
rect 1237 -5647 1241 -5643
rect -1234 -5806 -1230 -5802
rect -1225 -5806 -1221 -5802
rect -1216 -5806 -1212 -5802
rect -1208 -5806 -1204 -5802
rect -1199 -5806 -1195 -5802
rect -1181 -5806 -1177 -5802
rect -1172 -5806 -1168 -5802
rect -1164 -5806 -1160 -5802
rect -1147 -5806 -1143 -5802
rect -1138 -5806 -1134 -5802
rect -935 -5806 -931 -5802
rect -926 -5806 -922 -5802
rect -917 -5806 -913 -5802
rect -909 -5806 -905 -5802
rect -900 -5806 -896 -5802
rect -891 -5806 -887 -5802
rect -883 -5806 -879 -5802
rect -875 -5806 -871 -5802
rect -857 -5806 -853 -5802
rect -847 -5806 -843 -5802
rect -839 -5806 -835 -5802
rect -822 -5806 -818 -5802
rect -813 -5806 -809 -5802
rect -805 -5806 -801 -5802
rect -796 -5806 -792 -5802
rect -778 -5806 -774 -5802
rect -769 -5806 -765 -5802
rect -761 -5806 -757 -5802
rect -745 -5806 -741 -5802
rect -737 -5806 -733 -5802
rect -725 -5806 -721 -5802
rect -713 -5806 -709 -5802
rect -704 -5806 -700 -5802
rect -695 -5806 -691 -5802
rect -577 -5806 -573 -5802
rect -568 -5806 -564 -5802
rect -559 -5806 -555 -5802
rect -551 -5806 -547 -5802
rect -542 -5806 -538 -5802
rect -533 -5806 -529 -5802
rect -525 -5806 -521 -5802
rect -517 -5806 -513 -5802
rect -499 -5806 -495 -5802
rect -489 -5806 -485 -5802
rect -481 -5806 -477 -5802
rect -464 -5806 -460 -5802
rect -455 -5806 -451 -5802
rect -447 -5806 -443 -5802
rect -438 -5806 -434 -5802
rect -420 -5806 -416 -5802
rect -411 -5806 -407 -5802
rect -403 -5806 -399 -5802
rect -387 -5806 -383 -5802
rect -379 -5806 -375 -5802
rect -367 -5806 -363 -5802
rect -355 -5806 -351 -5802
rect -346 -5806 -342 -5802
rect -337 -5806 -333 -5802
rect -219 -5806 -215 -5802
rect -210 -5806 -206 -5802
rect -201 -5806 -197 -5802
rect -193 -5806 -189 -5802
rect -184 -5806 -180 -5802
rect -175 -5806 -171 -5802
rect -167 -5806 -163 -5802
rect -159 -5806 -155 -5802
rect -141 -5806 -137 -5802
rect -131 -5806 -127 -5802
rect -123 -5806 -119 -5802
rect -106 -5806 -102 -5802
rect -97 -5806 -93 -5802
rect -89 -5806 -85 -5802
rect -80 -5806 -76 -5802
rect -62 -5806 -58 -5802
rect -53 -5806 -49 -5802
rect -45 -5806 -41 -5802
rect -29 -5806 -25 -5802
rect -21 -5806 -17 -5802
rect -9 -5806 -5 -5802
rect 3 -5806 7 -5802
rect 12 -5806 16 -5802
rect 21 -5806 25 -5802
rect 139 -5806 143 -5802
rect 148 -5806 152 -5802
rect 157 -5806 161 -5802
rect 165 -5806 169 -5802
rect 174 -5806 178 -5802
rect 183 -5806 187 -5802
rect 191 -5806 195 -5802
rect 199 -5806 203 -5802
rect 217 -5806 221 -5802
rect 227 -5806 231 -5802
rect 235 -5806 239 -5802
rect 252 -5806 256 -5802
rect 261 -5806 265 -5802
rect 269 -5806 273 -5802
rect 278 -5806 282 -5802
rect 296 -5806 300 -5802
rect 305 -5806 309 -5802
rect 313 -5806 317 -5802
rect 329 -5806 333 -5802
rect 337 -5806 341 -5802
rect 349 -5806 353 -5802
rect 361 -5806 365 -5802
rect 370 -5806 374 -5802
rect 379 -5806 383 -5802
rect 495 -5806 499 -5802
rect 504 -5806 508 -5802
rect 513 -5806 517 -5802
rect 521 -5806 525 -5802
rect 530 -5806 534 -5802
rect 539 -5806 543 -5802
rect 547 -5806 551 -5802
rect 555 -5806 559 -5802
rect 573 -5806 577 -5802
rect 583 -5806 587 -5802
rect 591 -5806 595 -5802
rect 608 -5806 612 -5802
rect 617 -5806 621 -5802
rect 625 -5806 629 -5802
rect 634 -5806 638 -5802
rect 652 -5806 656 -5802
rect 661 -5806 665 -5802
rect 669 -5806 673 -5802
rect 685 -5806 689 -5802
rect 693 -5806 697 -5802
rect 705 -5806 709 -5802
rect 717 -5806 721 -5802
rect 726 -5806 730 -5802
rect 735 -5806 739 -5802
rect 853 -5806 857 -5802
rect 862 -5806 866 -5802
rect 871 -5806 875 -5802
rect 879 -5806 883 -5802
rect 888 -5806 892 -5802
rect 897 -5806 901 -5802
rect 905 -5806 909 -5802
rect 913 -5806 917 -5802
rect 931 -5806 935 -5802
rect 941 -5806 945 -5802
rect 949 -5806 953 -5802
rect 966 -5806 970 -5802
rect 975 -5806 979 -5802
rect 983 -5806 987 -5802
rect 992 -5806 996 -5802
rect 1010 -5806 1014 -5802
rect 1019 -5806 1023 -5802
rect 1027 -5806 1031 -5802
rect 1043 -5806 1047 -5802
rect 1051 -5806 1055 -5802
rect 1063 -5806 1067 -5802
rect 1075 -5806 1079 -5802
rect 1084 -5806 1088 -5802
rect 1093 -5806 1097 -5802
rect 1211 -5806 1215 -5802
rect 1220 -5806 1224 -5802
rect 1229 -5806 1233 -5802
rect 1237 -5806 1241 -5802
rect 1246 -5806 1250 -5802
rect 1255 -5806 1259 -5802
rect 1263 -5806 1267 -5802
rect 1271 -5806 1275 -5802
rect 1289 -5806 1293 -5802
rect 1299 -5806 1303 -5802
rect 1307 -5806 1311 -5802
rect 1324 -5806 1328 -5802
rect 1333 -5806 1337 -5802
rect 1341 -5806 1345 -5802
rect 1350 -5806 1354 -5802
rect 1368 -5806 1372 -5802
rect 1377 -5806 1381 -5802
rect 1385 -5806 1389 -5802
rect 1401 -5806 1405 -5802
rect 1409 -5806 1413 -5802
rect 1421 -5806 1425 -5802
rect 1433 -5806 1437 -5802
rect 1442 -5806 1446 -5802
rect 1451 -5806 1455 -5802
rect -1234 -5929 -1230 -5925
rect -1225 -5929 -1221 -5925
rect -1216 -5929 -1212 -5925
rect -1208 -5929 -1204 -5925
rect -1192 -5929 -1188 -5925
rect -1184 -5929 -1180 -5925
rect -1167 -5929 -1163 -5925
rect -1150 -5929 -1146 -5925
rect -1142 -5929 -1138 -5925
rect -1125 -5929 -1121 -5925
rect -1108 -5929 -1104 -5925
rect -1100 -5929 -1096 -5925
rect -1083 -5929 -1079 -5925
rect -1066 -5929 -1062 -5925
rect -1058 -5929 -1054 -5925
rect -1042 -5929 -1038 -5925
rect -935 -5929 -931 -5925
rect -926 -5929 -922 -5925
rect -917 -5929 -913 -5925
rect -909 -5929 -905 -5925
rect -893 -5929 -889 -5925
rect -885 -5929 -881 -5925
rect -868 -5929 -864 -5925
rect -851 -5929 -847 -5925
rect -843 -5929 -839 -5925
rect -826 -5929 -822 -5925
rect -809 -5929 -805 -5925
rect -801 -5929 -797 -5925
rect -784 -5929 -780 -5925
rect -767 -5929 -763 -5925
rect -759 -5929 -755 -5925
rect -743 -5929 -739 -5925
rect -577 -5929 -573 -5925
rect -568 -5929 -564 -5925
rect -559 -5929 -555 -5925
rect -551 -5929 -547 -5925
rect -535 -5929 -531 -5925
rect -527 -5929 -523 -5925
rect -510 -5929 -506 -5925
rect -493 -5929 -489 -5925
rect -485 -5929 -481 -5925
rect -468 -5929 -464 -5925
rect -451 -5929 -447 -5925
rect -443 -5929 -439 -5925
rect -426 -5929 -422 -5925
rect -409 -5929 -405 -5925
rect -401 -5929 -397 -5925
rect -385 -5929 -381 -5925
rect -219 -5929 -215 -5925
rect -210 -5929 -206 -5925
rect -201 -5929 -197 -5925
rect -193 -5929 -189 -5925
rect -177 -5929 -173 -5925
rect -169 -5929 -165 -5925
rect -152 -5929 -148 -5925
rect -135 -5929 -131 -5925
rect -127 -5929 -123 -5925
rect -110 -5929 -106 -5925
rect -93 -5929 -89 -5925
rect -85 -5929 -81 -5925
rect -68 -5929 -64 -5925
rect -51 -5929 -47 -5925
rect -43 -5929 -39 -5925
rect -27 -5929 -23 -5925
rect 139 -5929 143 -5925
rect 148 -5929 152 -5925
rect 157 -5929 161 -5925
rect 165 -5929 169 -5925
rect 181 -5929 185 -5925
rect 189 -5929 193 -5925
rect 206 -5929 210 -5925
rect 223 -5929 227 -5925
rect 231 -5929 235 -5925
rect 248 -5929 252 -5925
rect 265 -5929 269 -5925
rect 273 -5929 277 -5925
rect 290 -5929 294 -5925
rect 307 -5929 311 -5925
rect 315 -5929 319 -5925
rect 331 -5929 335 -5925
rect 495 -5929 499 -5925
rect 504 -5929 508 -5925
rect 513 -5929 517 -5925
rect 521 -5929 525 -5925
rect 537 -5929 541 -5925
rect 545 -5929 549 -5925
rect 562 -5929 566 -5925
rect 579 -5929 583 -5925
rect 587 -5929 591 -5925
rect 604 -5929 608 -5925
rect 621 -5929 625 -5925
rect 629 -5929 633 -5925
rect 646 -5929 650 -5925
rect 663 -5929 667 -5925
rect 671 -5929 675 -5925
rect 687 -5929 691 -5925
rect 853 -5929 857 -5925
rect 862 -5929 866 -5925
rect 871 -5929 875 -5925
rect 879 -5929 883 -5925
rect 895 -5929 899 -5925
rect 903 -5929 907 -5925
rect 920 -5929 924 -5925
rect 937 -5929 941 -5925
rect 945 -5929 949 -5925
rect 962 -5929 966 -5925
rect 979 -5929 983 -5925
rect 987 -5929 991 -5925
rect 1004 -5929 1008 -5925
rect 1021 -5929 1025 -5925
rect 1029 -5929 1033 -5925
rect 1045 -5929 1049 -5925
rect 1211 -5929 1215 -5925
rect 1220 -5929 1224 -5925
rect 1229 -5929 1233 -5925
rect 1237 -5929 1241 -5925
rect 1253 -5929 1257 -5925
rect 1261 -5929 1265 -5925
rect 1278 -5929 1282 -5925
rect 1295 -5929 1299 -5925
rect 1303 -5929 1307 -5925
rect 1320 -5929 1324 -5925
rect 1337 -5929 1341 -5925
rect 1345 -5929 1349 -5925
rect 1362 -5929 1366 -5925
rect 1379 -5929 1383 -5925
rect 1387 -5929 1391 -5925
rect 1403 -5929 1407 -5925
rect 1555 -5929 1559 -5925
rect 1564 -5929 1568 -5925
rect 1573 -5929 1577 -5925
rect 1581 -5929 1585 -5925
rect 1597 -5929 1601 -5925
rect 1605 -5929 1609 -5925
rect 1622 -5929 1626 -5925
rect 1639 -5929 1643 -5925
rect 1647 -5929 1651 -5925
rect 1664 -5929 1668 -5925
rect 1681 -5929 1685 -5925
rect 1689 -5929 1693 -5925
rect 1706 -5929 1710 -5925
rect 1723 -5929 1727 -5925
rect 1731 -5929 1735 -5925
rect 1747 -5929 1751 -5925
<< pdcontact >>
rect -1307 -796 -1303 -788
rect -1299 -796 -1295 -788
rect -1290 -796 -1286 -788
rect -1281 -796 -1277 -788
rect -936 -796 -932 -788
rect -928 -796 -924 -788
rect -919 -796 -915 -788
rect -910 -796 -906 -788
rect -577 -796 -573 -788
rect -569 -796 -565 -788
rect -560 -796 -556 -788
rect -551 -796 -547 -788
rect -219 -796 -215 -788
rect -211 -796 -207 -788
rect -202 -796 -198 -788
rect -193 -796 -189 -788
rect 138 -796 142 -788
rect 146 -796 150 -788
rect 155 -796 159 -788
rect 164 -796 168 -788
rect 495 -796 499 -788
rect 503 -796 507 -788
rect 512 -796 516 -788
rect 521 -796 525 -788
rect 853 -796 857 -788
rect 861 -796 865 -788
rect 870 -796 874 -788
rect 879 -796 883 -788
rect 1211 -796 1215 -788
rect 1219 -796 1223 -788
rect 1228 -796 1232 -788
rect 1237 -796 1241 -788
rect -1230 -1030 -1226 -1022
rect -1221 -1030 -1217 -1022
rect -1212 -1030 -1208 -1022
rect -1204 -1030 -1200 -1022
rect -1196 -1030 -1192 -1022
rect -1184 -1030 -1180 -1022
rect -1172 -1030 -1168 -1022
rect -1163 -1030 -1159 -1022
rect -1154 -1030 -1150 -1022
rect -1142 -1030 -1138 -1022
rect -1130 -1030 -1126 -1022
rect -1121 -1030 -1117 -1022
rect -1112 -1030 -1108 -1022
rect -1100 -1030 -1096 -1022
rect -1088 -1030 -1084 -1022
rect -1079 -1030 -1075 -1022
rect -1070 -1030 -1066 -1022
rect -1058 -1030 -1054 -1022
rect -1046 -1030 -1042 -1022
rect -1038 -1030 -1034 -1022
rect -935 -1030 -931 -1022
rect -926 -1030 -922 -1022
rect -917 -1030 -913 -1022
rect -909 -1030 -905 -1022
rect -901 -1030 -897 -1022
rect -889 -1030 -885 -1022
rect -877 -1030 -873 -1022
rect -868 -1030 -864 -1022
rect -859 -1030 -855 -1022
rect -847 -1030 -843 -1022
rect -835 -1030 -831 -1022
rect -826 -1030 -822 -1022
rect -817 -1030 -813 -1022
rect -805 -1030 -801 -1022
rect -793 -1030 -789 -1022
rect -784 -1030 -780 -1022
rect -775 -1030 -771 -1022
rect -763 -1030 -759 -1022
rect -751 -1030 -747 -1022
rect -743 -1030 -739 -1022
rect -577 -1030 -573 -1022
rect -568 -1030 -564 -1022
rect -559 -1030 -555 -1022
rect -551 -1030 -547 -1022
rect -543 -1030 -539 -1022
rect -531 -1030 -527 -1022
rect -519 -1030 -515 -1022
rect -510 -1030 -506 -1022
rect -501 -1030 -497 -1022
rect -489 -1030 -485 -1022
rect -477 -1030 -473 -1022
rect -468 -1030 -464 -1022
rect -459 -1030 -455 -1022
rect -447 -1030 -443 -1022
rect -435 -1030 -431 -1022
rect -426 -1030 -422 -1022
rect -417 -1030 -413 -1022
rect -405 -1030 -401 -1022
rect -393 -1030 -389 -1022
rect -385 -1030 -381 -1022
rect -219 -1030 -215 -1022
rect -210 -1030 -206 -1022
rect -201 -1030 -197 -1022
rect -193 -1030 -189 -1022
rect -185 -1030 -181 -1022
rect -173 -1030 -169 -1022
rect -161 -1030 -157 -1022
rect -152 -1030 -148 -1022
rect -143 -1030 -139 -1022
rect -131 -1030 -127 -1022
rect -119 -1030 -115 -1022
rect -110 -1030 -106 -1022
rect -101 -1030 -97 -1022
rect -89 -1030 -85 -1022
rect -77 -1030 -73 -1022
rect -68 -1030 -64 -1022
rect -59 -1030 -55 -1022
rect -47 -1030 -43 -1022
rect -35 -1030 -31 -1022
rect -27 -1030 -23 -1022
rect 139 -1030 143 -1022
rect 148 -1030 152 -1022
rect 157 -1030 161 -1022
rect 165 -1030 169 -1022
rect 173 -1030 177 -1022
rect 185 -1030 189 -1022
rect 197 -1030 201 -1022
rect 206 -1030 210 -1022
rect 215 -1030 219 -1022
rect 227 -1030 231 -1022
rect 239 -1030 243 -1022
rect 248 -1030 252 -1022
rect 257 -1030 261 -1022
rect 269 -1030 273 -1022
rect 281 -1030 285 -1022
rect 290 -1030 294 -1022
rect 299 -1030 303 -1022
rect 311 -1030 315 -1022
rect 323 -1030 327 -1022
rect 331 -1030 335 -1022
rect 495 -1030 499 -1022
rect 504 -1030 508 -1022
rect 513 -1030 517 -1022
rect 521 -1030 525 -1022
rect 529 -1030 533 -1022
rect 541 -1030 545 -1022
rect 553 -1030 557 -1022
rect 562 -1030 566 -1022
rect 571 -1030 575 -1022
rect 583 -1030 587 -1022
rect 595 -1030 599 -1022
rect 604 -1030 608 -1022
rect 613 -1030 617 -1022
rect 625 -1030 629 -1022
rect 637 -1030 641 -1022
rect 646 -1030 650 -1022
rect 655 -1030 659 -1022
rect 667 -1030 671 -1022
rect 679 -1030 683 -1022
rect 687 -1030 691 -1022
rect 853 -1030 857 -1022
rect 862 -1030 866 -1022
rect 871 -1030 875 -1022
rect 879 -1030 883 -1022
rect 887 -1030 891 -1022
rect 899 -1030 903 -1022
rect 911 -1030 915 -1022
rect 920 -1030 924 -1022
rect 929 -1030 933 -1022
rect 941 -1030 945 -1022
rect 953 -1030 957 -1022
rect 962 -1030 966 -1022
rect 971 -1030 975 -1022
rect 983 -1030 987 -1022
rect 995 -1030 999 -1022
rect 1004 -1030 1008 -1022
rect 1013 -1030 1017 -1022
rect 1025 -1030 1029 -1022
rect 1037 -1030 1041 -1022
rect 1045 -1030 1049 -1022
rect -1309 -1146 -1305 -1138
rect -1301 -1146 -1297 -1138
rect -1292 -1146 -1288 -1138
rect -1283 -1146 -1279 -1138
rect -935 -1146 -931 -1138
rect -927 -1146 -923 -1138
rect -918 -1146 -914 -1138
rect -909 -1146 -905 -1138
rect -577 -1146 -573 -1138
rect -569 -1146 -565 -1138
rect -560 -1146 -556 -1138
rect -551 -1146 -547 -1138
rect -219 -1146 -215 -1138
rect -211 -1146 -207 -1138
rect -202 -1146 -198 -1138
rect -193 -1146 -189 -1138
rect 139 -1146 143 -1138
rect 147 -1146 151 -1138
rect 156 -1146 160 -1138
rect 165 -1146 169 -1138
rect 495 -1146 499 -1138
rect 503 -1146 507 -1138
rect 512 -1146 516 -1138
rect 521 -1146 525 -1138
rect 853 -1146 857 -1138
rect 861 -1146 865 -1138
rect 870 -1146 874 -1138
rect 879 -1146 883 -1138
rect 1211 -1146 1215 -1138
rect 1219 -1146 1223 -1138
rect 1228 -1146 1232 -1138
rect 1237 -1146 1241 -1138
rect -1230 -1310 -1226 -1302
rect -1221 -1310 -1217 -1302
rect -1212 -1310 -1208 -1302
rect -1204 -1310 -1200 -1302
rect -1186 -1310 -1182 -1302
rect -1164 -1310 -1160 -1302
rect -1152 -1310 -1148 -1302
rect -1143 -1310 -1139 -1302
rect -1134 -1310 -1130 -1302
rect -935 -1310 -931 -1302
rect -926 -1310 -922 -1302
rect -917 -1310 -913 -1302
rect -909 -1310 -905 -1302
rect -900 -1310 -896 -1302
rect -891 -1310 -887 -1302
rect -883 -1310 -879 -1302
rect -865 -1310 -861 -1302
rect -843 -1310 -839 -1302
rect -831 -1310 -827 -1302
rect -822 -1310 -818 -1302
rect -813 -1310 -809 -1302
rect -805 -1310 -801 -1302
rect -787 -1310 -783 -1302
rect -765 -1310 -761 -1302
rect -753 -1310 -749 -1302
rect -741 -1310 -737 -1302
rect -729 -1310 -725 -1302
rect -721 -1310 -717 -1302
rect -704 -1310 -700 -1302
rect -695 -1310 -691 -1302
rect -577 -1310 -573 -1302
rect -568 -1310 -564 -1302
rect -559 -1310 -555 -1302
rect -551 -1310 -547 -1302
rect -542 -1310 -538 -1302
rect -533 -1310 -529 -1302
rect -525 -1310 -521 -1302
rect -507 -1310 -503 -1302
rect -485 -1310 -481 -1302
rect -473 -1310 -469 -1302
rect -464 -1310 -460 -1302
rect -455 -1310 -451 -1302
rect -447 -1310 -443 -1302
rect -429 -1310 -425 -1302
rect -407 -1310 -403 -1302
rect -395 -1310 -391 -1302
rect -383 -1310 -379 -1302
rect -371 -1310 -367 -1302
rect -363 -1310 -359 -1302
rect -346 -1310 -342 -1302
rect -337 -1310 -333 -1302
rect -219 -1310 -215 -1302
rect -210 -1310 -206 -1302
rect -201 -1310 -197 -1302
rect -193 -1310 -189 -1302
rect -184 -1310 -180 -1302
rect -175 -1310 -171 -1302
rect -167 -1310 -163 -1302
rect -149 -1310 -145 -1302
rect -127 -1310 -123 -1302
rect -115 -1310 -111 -1302
rect -106 -1310 -102 -1302
rect -97 -1310 -93 -1302
rect -89 -1310 -85 -1302
rect -71 -1310 -67 -1302
rect -49 -1310 -45 -1302
rect -37 -1310 -33 -1302
rect -25 -1310 -21 -1302
rect -13 -1310 -9 -1302
rect -5 -1310 -1 -1302
rect 12 -1310 16 -1302
rect 21 -1310 25 -1302
rect 139 -1310 143 -1302
rect 148 -1310 152 -1302
rect 157 -1310 161 -1302
rect 165 -1310 169 -1302
rect 174 -1310 178 -1302
rect 183 -1310 187 -1302
rect 191 -1310 195 -1302
rect 209 -1310 213 -1302
rect 231 -1310 235 -1302
rect 243 -1310 247 -1302
rect 252 -1310 256 -1302
rect 261 -1310 265 -1302
rect 269 -1310 273 -1302
rect 287 -1310 291 -1302
rect 309 -1310 313 -1302
rect 321 -1310 325 -1302
rect 333 -1310 337 -1302
rect 345 -1310 349 -1302
rect 353 -1310 357 -1302
rect 370 -1310 374 -1302
rect 379 -1310 383 -1302
rect 495 -1310 499 -1302
rect 504 -1310 508 -1302
rect 513 -1310 517 -1302
rect 521 -1310 525 -1302
rect 530 -1310 534 -1302
rect 539 -1310 543 -1302
rect 547 -1310 551 -1302
rect 565 -1310 569 -1302
rect 587 -1310 591 -1302
rect 599 -1310 603 -1302
rect 608 -1310 612 -1302
rect 617 -1310 621 -1302
rect 625 -1310 629 -1302
rect 643 -1310 647 -1302
rect 665 -1310 669 -1302
rect 677 -1310 681 -1302
rect 689 -1310 693 -1302
rect 701 -1310 705 -1302
rect 709 -1310 713 -1302
rect 726 -1310 730 -1302
rect 735 -1310 739 -1302
rect 853 -1310 857 -1302
rect 862 -1310 866 -1302
rect 871 -1310 875 -1302
rect 879 -1310 883 -1302
rect 888 -1310 892 -1302
rect 897 -1310 901 -1302
rect 905 -1310 909 -1302
rect 923 -1310 927 -1302
rect 945 -1310 949 -1302
rect 957 -1310 961 -1302
rect 966 -1310 970 -1302
rect 975 -1310 979 -1302
rect 983 -1310 987 -1302
rect 1001 -1310 1005 -1302
rect 1023 -1310 1027 -1302
rect 1035 -1310 1039 -1302
rect 1047 -1310 1051 -1302
rect 1059 -1310 1063 -1302
rect 1067 -1310 1071 -1302
rect 1084 -1310 1088 -1302
rect 1093 -1310 1097 -1302
rect 1211 -1310 1215 -1302
rect 1220 -1310 1224 -1302
rect 1229 -1310 1233 -1302
rect 1237 -1310 1241 -1302
rect 1255 -1310 1259 -1302
rect 1277 -1310 1281 -1302
rect 1289 -1310 1293 -1302
rect 1298 -1310 1302 -1302
rect 1307 -1310 1311 -1302
rect -1230 -1433 -1226 -1425
rect -1221 -1433 -1217 -1425
rect -1212 -1433 -1208 -1425
rect -1204 -1433 -1200 -1425
rect -1196 -1433 -1192 -1425
rect -1184 -1433 -1180 -1425
rect -1172 -1433 -1168 -1425
rect -1163 -1433 -1159 -1425
rect -1154 -1433 -1150 -1425
rect -1142 -1433 -1138 -1425
rect -1130 -1433 -1126 -1425
rect -1121 -1433 -1117 -1425
rect -1112 -1433 -1108 -1425
rect -1100 -1433 -1096 -1425
rect -1088 -1433 -1084 -1425
rect -1079 -1433 -1075 -1425
rect -1070 -1433 -1066 -1425
rect -1058 -1433 -1054 -1425
rect -1046 -1433 -1042 -1425
rect -1038 -1433 -1034 -1425
rect -935 -1433 -931 -1425
rect -926 -1433 -922 -1425
rect -917 -1433 -913 -1425
rect -909 -1433 -905 -1425
rect -901 -1433 -897 -1425
rect -889 -1433 -885 -1425
rect -877 -1433 -873 -1425
rect -868 -1433 -864 -1425
rect -859 -1433 -855 -1425
rect -847 -1433 -843 -1425
rect -835 -1433 -831 -1425
rect -826 -1433 -822 -1425
rect -817 -1433 -813 -1425
rect -805 -1433 -801 -1425
rect -793 -1433 -789 -1425
rect -784 -1433 -780 -1425
rect -775 -1433 -771 -1425
rect -763 -1433 -759 -1425
rect -751 -1433 -747 -1425
rect -743 -1433 -739 -1425
rect -577 -1433 -573 -1425
rect -568 -1433 -564 -1425
rect -559 -1433 -555 -1425
rect -551 -1433 -547 -1425
rect -543 -1433 -539 -1425
rect -531 -1433 -527 -1425
rect -519 -1433 -515 -1425
rect -510 -1433 -506 -1425
rect -501 -1433 -497 -1425
rect -489 -1433 -485 -1425
rect -477 -1433 -473 -1425
rect -468 -1433 -464 -1425
rect -459 -1433 -455 -1425
rect -447 -1433 -443 -1425
rect -435 -1433 -431 -1425
rect -426 -1433 -422 -1425
rect -417 -1433 -413 -1425
rect -405 -1433 -401 -1425
rect -393 -1433 -389 -1425
rect -385 -1433 -381 -1425
rect -219 -1433 -215 -1425
rect -210 -1433 -206 -1425
rect -201 -1433 -197 -1425
rect -193 -1433 -189 -1425
rect -185 -1433 -181 -1425
rect -173 -1433 -169 -1425
rect -161 -1433 -157 -1425
rect -152 -1433 -148 -1425
rect -143 -1433 -139 -1425
rect -131 -1433 -127 -1425
rect -119 -1433 -115 -1425
rect -110 -1433 -106 -1425
rect -101 -1433 -97 -1425
rect -89 -1433 -85 -1425
rect -77 -1433 -73 -1425
rect -68 -1433 -64 -1425
rect -59 -1433 -55 -1425
rect -47 -1433 -43 -1425
rect -35 -1433 -31 -1425
rect -27 -1433 -23 -1425
rect 139 -1433 143 -1425
rect 148 -1433 152 -1425
rect 157 -1433 161 -1425
rect 165 -1433 169 -1425
rect 173 -1433 177 -1425
rect 185 -1433 189 -1425
rect 197 -1433 201 -1425
rect 206 -1433 210 -1425
rect 215 -1433 219 -1425
rect 227 -1433 231 -1425
rect 239 -1433 243 -1425
rect 248 -1433 252 -1425
rect 257 -1433 261 -1425
rect 269 -1433 273 -1425
rect 281 -1433 285 -1425
rect 290 -1433 294 -1425
rect 299 -1433 303 -1425
rect 311 -1433 315 -1425
rect 323 -1433 327 -1425
rect 331 -1433 335 -1425
rect 495 -1433 499 -1425
rect 504 -1433 508 -1425
rect 513 -1433 517 -1425
rect 521 -1433 525 -1425
rect 529 -1433 533 -1425
rect 541 -1433 545 -1425
rect 553 -1433 557 -1425
rect 562 -1433 566 -1425
rect 571 -1433 575 -1425
rect 583 -1433 587 -1425
rect 595 -1433 599 -1425
rect 604 -1433 608 -1425
rect 613 -1433 617 -1425
rect 625 -1433 629 -1425
rect 637 -1433 641 -1425
rect 646 -1433 650 -1425
rect 655 -1433 659 -1425
rect 667 -1433 671 -1425
rect 679 -1433 683 -1425
rect 687 -1433 691 -1425
rect 853 -1433 857 -1425
rect 862 -1433 866 -1425
rect 871 -1433 875 -1425
rect 879 -1433 883 -1425
rect 887 -1433 891 -1425
rect 899 -1433 903 -1425
rect 911 -1433 915 -1425
rect 920 -1433 924 -1425
rect 929 -1433 933 -1425
rect 941 -1433 945 -1425
rect 953 -1433 957 -1425
rect 962 -1433 966 -1425
rect 971 -1433 975 -1425
rect 983 -1433 987 -1425
rect 995 -1433 999 -1425
rect 1004 -1433 1008 -1425
rect 1013 -1433 1017 -1425
rect 1025 -1433 1029 -1425
rect 1037 -1433 1041 -1425
rect 1045 -1433 1049 -1425
rect -1230 -1604 -1226 -1596
rect -1221 -1604 -1217 -1596
rect -1212 -1604 -1208 -1596
rect -1204 -1604 -1200 -1596
rect -1196 -1604 -1192 -1596
rect -1184 -1604 -1180 -1596
rect -1172 -1604 -1168 -1596
rect -1163 -1604 -1159 -1596
rect -1154 -1604 -1150 -1596
rect -1142 -1604 -1138 -1596
rect -1130 -1604 -1126 -1596
rect -1121 -1604 -1117 -1596
rect -1112 -1604 -1108 -1596
rect -1100 -1604 -1096 -1596
rect -1088 -1604 -1084 -1596
rect -1079 -1604 -1075 -1596
rect -1070 -1604 -1066 -1596
rect -1058 -1604 -1054 -1596
rect -1046 -1604 -1042 -1596
rect -1038 -1604 -1034 -1596
rect -935 -1604 -931 -1596
rect -926 -1604 -922 -1596
rect -917 -1604 -913 -1596
rect -909 -1604 -905 -1596
rect -901 -1604 -897 -1596
rect -889 -1604 -885 -1596
rect -877 -1604 -873 -1596
rect -868 -1604 -864 -1596
rect -859 -1604 -855 -1596
rect -847 -1604 -843 -1596
rect -835 -1604 -831 -1596
rect -826 -1604 -822 -1596
rect -817 -1604 -813 -1596
rect -805 -1604 -801 -1596
rect -793 -1604 -789 -1596
rect -784 -1604 -780 -1596
rect -775 -1604 -771 -1596
rect -763 -1604 -759 -1596
rect -751 -1604 -747 -1596
rect -743 -1604 -739 -1596
rect -577 -1604 -573 -1596
rect -568 -1604 -564 -1596
rect -559 -1604 -555 -1596
rect -551 -1604 -547 -1596
rect -543 -1604 -539 -1596
rect -531 -1604 -527 -1596
rect -519 -1604 -515 -1596
rect -510 -1604 -506 -1596
rect -501 -1604 -497 -1596
rect -489 -1604 -485 -1596
rect -477 -1604 -473 -1596
rect -468 -1604 -464 -1596
rect -459 -1604 -455 -1596
rect -447 -1604 -443 -1596
rect -435 -1604 -431 -1596
rect -426 -1604 -422 -1596
rect -417 -1604 -413 -1596
rect -405 -1604 -401 -1596
rect -393 -1604 -389 -1596
rect -385 -1604 -381 -1596
rect -219 -1604 -215 -1596
rect -210 -1604 -206 -1596
rect -201 -1604 -197 -1596
rect -193 -1604 -189 -1596
rect -185 -1604 -181 -1596
rect -173 -1604 -169 -1596
rect -161 -1604 -157 -1596
rect -152 -1604 -148 -1596
rect -143 -1604 -139 -1596
rect -131 -1604 -127 -1596
rect -119 -1604 -115 -1596
rect -110 -1604 -106 -1596
rect -101 -1604 -97 -1596
rect -89 -1604 -85 -1596
rect -77 -1604 -73 -1596
rect -68 -1604 -64 -1596
rect -59 -1604 -55 -1596
rect -47 -1604 -43 -1596
rect -35 -1604 -31 -1596
rect -27 -1604 -23 -1596
rect 139 -1604 143 -1596
rect 148 -1604 152 -1596
rect 157 -1604 161 -1596
rect 165 -1604 169 -1596
rect 173 -1604 177 -1596
rect 185 -1604 189 -1596
rect 197 -1604 201 -1596
rect 206 -1604 210 -1596
rect 215 -1604 219 -1596
rect 227 -1604 231 -1596
rect 239 -1604 243 -1596
rect 248 -1604 252 -1596
rect 257 -1604 261 -1596
rect 269 -1604 273 -1596
rect 281 -1604 285 -1596
rect 290 -1604 294 -1596
rect 299 -1604 303 -1596
rect 311 -1604 315 -1596
rect 323 -1604 327 -1596
rect 331 -1604 335 -1596
rect 495 -1604 499 -1596
rect 504 -1604 508 -1596
rect 513 -1604 517 -1596
rect 521 -1604 525 -1596
rect 529 -1604 533 -1596
rect 541 -1604 545 -1596
rect 553 -1604 557 -1596
rect 562 -1604 566 -1596
rect 571 -1604 575 -1596
rect 583 -1604 587 -1596
rect 595 -1604 599 -1596
rect 604 -1604 608 -1596
rect 613 -1604 617 -1596
rect 625 -1604 629 -1596
rect 637 -1604 641 -1596
rect 646 -1604 650 -1596
rect 655 -1604 659 -1596
rect 667 -1604 671 -1596
rect 679 -1604 683 -1596
rect 687 -1604 691 -1596
rect 853 -1604 857 -1596
rect 862 -1604 866 -1596
rect 871 -1604 875 -1596
rect 879 -1604 883 -1596
rect 887 -1604 891 -1596
rect 899 -1604 903 -1596
rect 911 -1604 915 -1596
rect 920 -1604 924 -1596
rect 929 -1604 933 -1596
rect 941 -1604 945 -1596
rect 953 -1604 957 -1596
rect 962 -1604 966 -1596
rect 971 -1604 975 -1596
rect 983 -1604 987 -1596
rect 995 -1604 999 -1596
rect 1004 -1604 1008 -1596
rect 1013 -1604 1017 -1596
rect 1025 -1604 1029 -1596
rect 1037 -1604 1041 -1596
rect 1045 -1604 1049 -1596
rect 1211 -1604 1215 -1596
rect 1220 -1604 1224 -1596
rect 1229 -1604 1233 -1596
rect 1237 -1604 1241 -1596
rect 1245 -1604 1249 -1596
rect 1257 -1604 1261 -1596
rect 1269 -1604 1273 -1596
rect 1278 -1604 1282 -1596
rect 1287 -1604 1291 -1596
rect 1299 -1604 1303 -1596
rect 1311 -1604 1315 -1596
rect 1320 -1604 1324 -1596
rect 1329 -1604 1333 -1596
rect 1341 -1604 1345 -1596
rect 1353 -1604 1357 -1596
rect 1362 -1604 1366 -1596
rect 1371 -1604 1375 -1596
rect 1383 -1604 1387 -1596
rect 1395 -1604 1399 -1596
rect 1403 -1604 1407 -1596
rect -1559 -1775 -1555 -1767
rect -1550 -1775 -1546 -1767
rect -1541 -1775 -1537 -1767
rect -1533 -1775 -1529 -1767
rect -1525 -1775 -1521 -1767
rect -1513 -1775 -1509 -1767
rect -1501 -1775 -1497 -1767
rect -1492 -1775 -1488 -1767
rect -1483 -1775 -1479 -1767
rect -1471 -1775 -1467 -1767
rect -1459 -1775 -1455 -1767
rect -1450 -1775 -1446 -1767
rect -1441 -1775 -1437 -1767
rect -1429 -1775 -1425 -1767
rect -1417 -1775 -1413 -1767
rect -1408 -1775 -1404 -1767
rect -1399 -1775 -1395 -1767
rect -1387 -1775 -1383 -1767
rect -1375 -1775 -1371 -1767
rect -1367 -1775 -1363 -1767
rect -1230 -1775 -1226 -1767
rect -1221 -1775 -1217 -1767
rect -1212 -1775 -1208 -1767
rect -1204 -1775 -1200 -1767
rect -1196 -1775 -1192 -1767
rect -1184 -1775 -1180 -1767
rect -1172 -1775 -1168 -1767
rect -1163 -1775 -1159 -1767
rect -1154 -1775 -1150 -1767
rect -1142 -1775 -1138 -1767
rect -1130 -1775 -1126 -1767
rect -1121 -1775 -1117 -1767
rect -1112 -1775 -1108 -1767
rect -1100 -1775 -1096 -1767
rect -1088 -1775 -1084 -1767
rect -1079 -1775 -1075 -1767
rect -1070 -1775 -1066 -1767
rect -1058 -1775 -1054 -1767
rect -1046 -1775 -1042 -1767
rect -1038 -1775 -1034 -1767
rect -935 -1775 -931 -1767
rect -926 -1775 -922 -1767
rect -917 -1775 -913 -1767
rect -909 -1775 -905 -1767
rect -901 -1775 -897 -1767
rect -889 -1775 -885 -1767
rect -877 -1775 -873 -1767
rect -868 -1775 -864 -1767
rect -859 -1775 -855 -1767
rect -847 -1775 -843 -1767
rect -835 -1775 -831 -1767
rect -826 -1775 -822 -1767
rect -817 -1775 -813 -1767
rect -805 -1775 -801 -1767
rect -793 -1775 -789 -1767
rect -784 -1775 -780 -1767
rect -775 -1775 -771 -1767
rect -763 -1775 -759 -1767
rect -751 -1775 -747 -1767
rect -743 -1775 -739 -1767
rect -577 -1775 -573 -1767
rect -568 -1775 -564 -1767
rect -559 -1775 -555 -1767
rect -551 -1775 -547 -1767
rect -543 -1775 -539 -1767
rect -531 -1775 -527 -1767
rect -519 -1775 -515 -1767
rect -510 -1775 -506 -1767
rect -501 -1775 -497 -1767
rect -489 -1775 -485 -1767
rect -477 -1775 -473 -1767
rect -468 -1775 -464 -1767
rect -459 -1775 -455 -1767
rect -447 -1775 -443 -1767
rect -435 -1775 -431 -1767
rect -426 -1775 -422 -1767
rect -417 -1775 -413 -1767
rect -405 -1775 -401 -1767
rect -393 -1775 -389 -1767
rect -385 -1775 -381 -1767
rect -219 -1775 -215 -1767
rect -210 -1775 -206 -1767
rect -201 -1775 -197 -1767
rect -193 -1775 -189 -1767
rect -185 -1775 -181 -1767
rect -173 -1775 -169 -1767
rect -161 -1775 -157 -1767
rect -152 -1775 -148 -1767
rect -143 -1775 -139 -1767
rect -131 -1775 -127 -1767
rect -119 -1775 -115 -1767
rect -110 -1775 -106 -1767
rect -101 -1775 -97 -1767
rect -89 -1775 -85 -1767
rect -77 -1775 -73 -1767
rect -68 -1775 -64 -1767
rect -59 -1775 -55 -1767
rect -47 -1775 -43 -1767
rect -35 -1775 -31 -1767
rect -27 -1775 -23 -1767
rect 139 -1775 143 -1767
rect 148 -1775 152 -1767
rect 157 -1775 161 -1767
rect 165 -1775 169 -1767
rect 173 -1775 177 -1767
rect 185 -1775 189 -1767
rect 197 -1775 201 -1767
rect 206 -1775 210 -1767
rect 215 -1775 219 -1767
rect 227 -1775 231 -1767
rect 239 -1775 243 -1767
rect 248 -1775 252 -1767
rect 257 -1775 261 -1767
rect 269 -1775 273 -1767
rect 281 -1775 285 -1767
rect 290 -1775 294 -1767
rect 299 -1775 303 -1767
rect 311 -1775 315 -1767
rect 323 -1775 327 -1767
rect 331 -1775 335 -1767
rect 495 -1775 499 -1767
rect 504 -1775 508 -1767
rect 513 -1775 517 -1767
rect 521 -1775 525 -1767
rect 529 -1775 533 -1767
rect 541 -1775 545 -1767
rect 553 -1775 557 -1767
rect 562 -1775 566 -1767
rect 571 -1775 575 -1767
rect 583 -1775 587 -1767
rect 595 -1775 599 -1767
rect 604 -1775 608 -1767
rect 613 -1775 617 -1767
rect 625 -1775 629 -1767
rect 637 -1775 641 -1767
rect 646 -1775 650 -1767
rect 655 -1775 659 -1767
rect 667 -1775 671 -1767
rect 679 -1775 683 -1767
rect 687 -1775 691 -1767
rect 853 -1775 857 -1767
rect 862 -1775 866 -1767
rect 871 -1775 875 -1767
rect 879 -1775 883 -1767
rect 887 -1775 891 -1767
rect 899 -1775 903 -1767
rect 911 -1775 915 -1767
rect 920 -1775 924 -1767
rect 929 -1775 933 -1767
rect 941 -1775 945 -1767
rect 953 -1775 957 -1767
rect 962 -1775 966 -1767
rect 971 -1775 975 -1767
rect 983 -1775 987 -1767
rect 995 -1775 999 -1767
rect 1004 -1775 1008 -1767
rect 1013 -1775 1017 -1767
rect 1025 -1775 1029 -1767
rect 1037 -1775 1041 -1767
rect 1045 -1775 1049 -1767
rect 1211 -1775 1215 -1767
rect 1220 -1775 1224 -1767
rect 1229 -1775 1233 -1767
rect 1237 -1775 1241 -1767
rect 1245 -1775 1249 -1767
rect 1257 -1775 1261 -1767
rect 1269 -1775 1273 -1767
rect 1278 -1775 1282 -1767
rect 1287 -1775 1291 -1767
rect 1299 -1775 1303 -1767
rect 1311 -1775 1315 -1767
rect 1320 -1775 1324 -1767
rect 1329 -1775 1333 -1767
rect 1341 -1775 1345 -1767
rect 1353 -1775 1357 -1767
rect 1362 -1775 1366 -1767
rect 1371 -1775 1375 -1767
rect 1383 -1775 1387 -1767
rect 1395 -1775 1399 -1767
rect 1403 -1775 1407 -1767
rect -1309 -1882 -1305 -1874
rect -1301 -1882 -1297 -1874
rect -1292 -1882 -1288 -1874
rect -1283 -1882 -1279 -1874
rect -935 -1882 -931 -1874
rect -927 -1882 -923 -1874
rect -918 -1882 -914 -1874
rect -909 -1882 -905 -1874
rect -577 -1882 -573 -1874
rect -569 -1882 -565 -1874
rect -560 -1882 -556 -1874
rect -551 -1882 -547 -1874
rect -219 -1882 -215 -1874
rect -211 -1882 -207 -1874
rect -202 -1882 -198 -1874
rect -193 -1882 -189 -1874
rect 139 -1882 143 -1874
rect 147 -1882 151 -1874
rect 156 -1882 160 -1874
rect 165 -1882 169 -1874
rect 495 -1882 499 -1874
rect 503 -1882 507 -1874
rect 512 -1882 516 -1874
rect 521 -1882 525 -1874
rect 853 -1882 857 -1874
rect 861 -1882 865 -1874
rect 870 -1882 874 -1874
rect 879 -1882 883 -1874
rect 1211 -1882 1215 -1874
rect 1219 -1882 1223 -1874
rect 1228 -1882 1232 -1874
rect 1237 -1882 1241 -1874
rect -1234 -2041 -1230 -2033
rect -1225 -2041 -1221 -2033
rect -1216 -2041 -1212 -2033
rect -1208 -2041 -1204 -2033
rect -1190 -2041 -1186 -2033
rect -1168 -2041 -1164 -2033
rect -1156 -2041 -1152 -2033
rect -1147 -2041 -1143 -2033
rect -1138 -2041 -1134 -2033
rect -935 -2041 -931 -2033
rect -926 -2041 -922 -2033
rect -917 -2041 -913 -2033
rect -909 -2041 -905 -2033
rect -900 -2041 -896 -2033
rect -891 -2041 -887 -2033
rect -883 -2041 -879 -2033
rect -865 -2041 -861 -2033
rect -843 -2041 -839 -2033
rect -831 -2041 -827 -2033
rect -822 -2041 -818 -2033
rect -813 -2041 -809 -2033
rect -805 -2041 -801 -2033
rect -787 -2041 -783 -2033
rect -765 -2041 -761 -2033
rect -753 -2041 -749 -2033
rect -741 -2041 -737 -2033
rect -729 -2041 -725 -2033
rect -721 -2041 -717 -2033
rect -704 -2041 -700 -2033
rect -695 -2041 -691 -2033
rect -577 -2041 -573 -2033
rect -568 -2041 -564 -2033
rect -559 -2041 -555 -2033
rect -551 -2041 -547 -2033
rect -542 -2041 -538 -2033
rect -533 -2041 -529 -2033
rect -525 -2041 -521 -2033
rect -507 -2041 -503 -2033
rect -485 -2041 -481 -2033
rect -473 -2041 -469 -2033
rect -464 -2041 -460 -2033
rect -455 -2041 -451 -2033
rect -447 -2041 -443 -2033
rect -429 -2041 -425 -2033
rect -407 -2041 -403 -2033
rect -395 -2041 -391 -2033
rect -383 -2041 -379 -2033
rect -371 -2041 -367 -2033
rect -363 -2041 -359 -2033
rect -346 -2041 -342 -2033
rect -337 -2041 -333 -2033
rect -219 -2041 -215 -2033
rect -210 -2041 -206 -2033
rect -201 -2041 -197 -2033
rect -193 -2041 -189 -2033
rect -184 -2041 -180 -2033
rect -175 -2041 -171 -2033
rect -167 -2041 -163 -2033
rect -149 -2041 -145 -2033
rect -127 -2041 -123 -2033
rect -115 -2041 -111 -2033
rect -106 -2041 -102 -2033
rect -97 -2041 -93 -2033
rect -89 -2041 -85 -2033
rect -71 -2041 -67 -2033
rect -49 -2041 -45 -2033
rect -37 -2041 -33 -2033
rect -25 -2041 -21 -2033
rect -13 -2041 -9 -2033
rect -5 -2041 -1 -2033
rect 12 -2041 16 -2033
rect 21 -2041 25 -2033
rect 139 -2041 143 -2033
rect 148 -2041 152 -2033
rect 157 -2041 161 -2033
rect 165 -2041 169 -2033
rect 174 -2041 178 -2033
rect 183 -2041 187 -2033
rect 191 -2041 195 -2033
rect 209 -2041 213 -2033
rect 231 -2041 235 -2033
rect 243 -2041 247 -2033
rect 252 -2041 256 -2033
rect 261 -2041 265 -2033
rect 269 -2041 273 -2033
rect 287 -2041 291 -2033
rect 309 -2041 313 -2033
rect 321 -2041 325 -2033
rect 333 -2041 337 -2033
rect 345 -2041 349 -2033
rect 353 -2041 357 -2033
rect 370 -2041 374 -2033
rect 379 -2041 383 -2033
rect 495 -2041 499 -2033
rect 504 -2041 508 -2033
rect 513 -2041 517 -2033
rect 521 -2041 525 -2033
rect 530 -2041 534 -2033
rect 539 -2041 543 -2033
rect 547 -2041 551 -2033
rect 565 -2041 569 -2033
rect 587 -2041 591 -2033
rect 599 -2041 603 -2033
rect 608 -2041 612 -2033
rect 617 -2041 621 -2033
rect 625 -2041 629 -2033
rect 643 -2041 647 -2033
rect 665 -2041 669 -2033
rect 677 -2041 681 -2033
rect 689 -2041 693 -2033
rect 701 -2041 705 -2033
rect 709 -2041 713 -2033
rect 726 -2041 730 -2033
rect 735 -2041 739 -2033
rect 853 -2041 857 -2033
rect 862 -2041 866 -2033
rect 871 -2041 875 -2033
rect 879 -2041 883 -2033
rect 888 -2041 892 -2033
rect 897 -2041 901 -2033
rect 905 -2041 909 -2033
rect 923 -2041 927 -2033
rect 945 -2041 949 -2033
rect 957 -2041 961 -2033
rect 966 -2041 970 -2033
rect 975 -2041 979 -2033
rect 983 -2041 987 -2033
rect 1001 -2041 1005 -2033
rect 1023 -2041 1027 -2033
rect 1035 -2041 1039 -2033
rect 1047 -2041 1051 -2033
rect 1059 -2041 1063 -2033
rect 1067 -2041 1071 -2033
rect 1084 -2041 1088 -2033
rect 1093 -2041 1097 -2033
rect 1211 -2041 1215 -2033
rect 1220 -2041 1224 -2033
rect 1229 -2041 1233 -2033
rect 1237 -2041 1241 -2033
rect 1246 -2041 1250 -2033
rect 1255 -2041 1259 -2033
rect 1263 -2041 1267 -2033
rect 1281 -2041 1285 -2033
rect 1303 -2041 1307 -2033
rect 1315 -2041 1319 -2033
rect 1324 -2041 1328 -2033
rect 1333 -2041 1337 -2033
rect 1341 -2041 1345 -2033
rect 1359 -2041 1363 -2033
rect 1381 -2041 1385 -2033
rect 1393 -2041 1397 -2033
rect 1405 -2041 1409 -2033
rect 1417 -2041 1421 -2033
rect 1425 -2041 1429 -2033
rect 1442 -2041 1446 -2033
rect 1451 -2041 1455 -2033
rect -1234 -2185 -1230 -2177
rect -1225 -2185 -1221 -2177
rect -1216 -2185 -1212 -2177
rect -1208 -2185 -1204 -2177
rect -1200 -2185 -1196 -2177
rect -1188 -2185 -1184 -2177
rect -1176 -2185 -1172 -2177
rect -1167 -2185 -1163 -2177
rect -1158 -2185 -1154 -2177
rect -1146 -2185 -1142 -2177
rect -1134 -2185 -1130 -2177
rect -1125 -2185 -1121 -2177
rect -1116 -2185 -1112 -2177
rect -1104 -2185 -1100 -2177
rect -1092 -2185 -1088 -2177
rect -1083 -2185 -1079 -2177
rect -1074 -2185 -1070 -2177
rect -1062 -2185 -1058 -2177
rect -1050 -2185 -1046 -2177
rect -1042 -2185 -1038 -2177
rect -935 -2185 -931 -2177
rect -926 -2185 -922 -2177
rect -917 -2185 -913 -2177
rect -909 -2185 -905 -2177
rect -901 -2185 -897 -2177
rect -889 -2185 -885 -2177
rect -877 -2185 -873 -2177
rect -868 -2185 -864 -2177
rect -859 -2185 -855 -2177
rect -847 -2185 -843 -2177
rect -835 -2185 -831 -2177
rect -826 -2185 -822 -2177
rect -817 -2185 -813 -2177
rect -805 -2185 -801 -2177
rect -793 -2185 -789 -2177
rect -784 -2185 -780 -2177
rect -775 -2185 -771 -2177
rect -763 -2185 -759 -2177
rect -751 -2185 -747 -2177
rect -743 -2185 -739 -2177
rect -577 -2185 -573 -2177
rect -568 -2185 -564 -2177
rect -559 -2185 -555 -2177
rect -551 -2185 -547 -2177
rect -543 -2185 -539 -2177
rect -531 -2185 -527 -2177
rect -519 -2185 -515 -2177
rect -510 -2185 -506 -2177
rect -501 -2185 -497 -2177
rect -489 -2185 -485 -2177
rect -477 -2185 -473 -2177
rect -468 -2185 -464 -2177
rect -459 -2185 -455 -2177
rect -447 -2185 -443 -2177
rect -435 -2185 -431 -2177
rect -426 -2185 -422 -2177
rect -417 -2185 -413 -2177
rect -405 -2185 -401 -2177
rect -393 -2185 -389 -2177
rect -385 -2185 -381 -2177
rect -219 -2185 -215 -2177
rect -210 -2185 -206 -2177
rect -201 -2185 -197 -2177
rect -193 -2185 -189 -2177
rect -185 -2185 -181 -2177
rect -173 -2185 -169 -2177
rect -161 -2185 -157 -2177
rect -152 -2185 -148 -2177
rect -143 -2185 -139 -2177
rect -131 -2185 -127 -2177
rect -119 -2185 -115 -2177
rect -110 -2185 -106 -2177
rect -101 -2185 -97 -2177
rect -89 -2185 -85 -2177
rect -77 -2185 -73 -2177
rect -68 -2185 -64 -2177
rect -59 -2185 -55 -2177
rect -47 -2185 -43 -2177
rect -35 -2185 -31 -2177
rect -27 -2185 -23 -2177
rect 139 -2185 143 -2177
rect 148 -2185 152 -2177
rect 157 -2185 161 -2177
rect 165 -2185 169 -2177
rect 173 -2185 177 -2177
rect 185 -2185 189 -2177
rect 197 -2185 201 -2177
rect 206 -2185 210 -2177
rect 215 -2185 219 -2177
rect 227 -2185 231 -2177
rect 239 -2185 243 -2177
rect 248 -2185 252 -2177
rect 257 -2185 261 -2177
rect 269 -2185 273 -2177
rect 281 -2185 285 -2177
rect 290 -2185 294 -2177
rect 299 -2185 303 -2177
rect 311 -2185 315 -2177
rect 323 -2185 327 -2177
rect 331 -2185 335 -2177
rect 495 -2185 499 -2177
rect 504 -2185 508 -2177
rect 513 -2185 517 -2177
rect 521 -2185 525 -2177
rect 529 -2185 533 -2177
rect 541 -2185 545 -2177
rect 553 -2185 557 -2177
rect 562 -2185 566 -2177
rect 571 -2185 575 -2177
rect 583 -2185 587 -2177
rect 595 -2185 599 -2177
rect 604 -2185 608 -2177
rect 613 -2185 617 -2177
rect 625 -2185 629 -2177
rect 637 -2185 641 -2177
rect 646 -2185 650 -2177
rect 655 -2185 659 -2177
rect 667 -2185 671 -2177
rect 679 -2185 683 -2177
rect 687 -2185 691 -2177
rect -1559 -2356 -1555 -2348
rect -1550 -2356 -1546 -2348
rect -1541 -2356 -1537 -2348
rect -1533 -2356 -1529 -2348
rect -1525 -2356 -1521 -2348
rect -1513 -2356 -1509 -2348
rect -1501 -2356 -1497 -2348
rect -1492 -2356 -1488 -2348
rect -1483 -2356 -1479 -2348
rect -1471 -2356 -1467 -2348
rect -1459 -2356 -1455 -2348
rect -1450 -2356 -1446 -2348
rect -1441 -2356 -1437 -2348
rect -1429 -2356 -1425 -2348
rect -1417 -2356 -1413 -2348
rect -1408 -2356 -1404 -2348
rect -1399 -2356 -1395 -2348
rect -1387 -2356 -1383 -2348
rect -1375 -2356 -1371 -2348
rect -1367 -2356 -1363 -2348
rect -1234 -2356 -1230 -2348
rect -1225 -2356 -1221 -2348
rect -1216 -2356 -1212 -2348
rect -1208 -2356 -1204 -2348
rect -1200 -2356 -1196 -2348
rect -1188 -2356 -1184 -2348
rect -1176 -2356 -1172 -2348
rect -1167 -2356 -1163 -2348
rect -1158 -2356 -1154 -2348
rect -1146 -2356 -1142 -2348
rect -1134 -2356 -1130 -2348
rect -1125 -2356 -1121 -2348
rect -1116 -2356 -1112 -2348
rect -1104 -2356 -1100 -2348
rect -1092 -2356 -1088 -2348
rect -1083 -2356 -1079 -2348
rect -1074 -2356 -1070 -2348
rect -1062 -2356 -1058 -2348
rect -1050 -2356 -1046 -2348
rect -1042 -2356 -1038 -2348
rect -935 -2356 -931 -2348
rect -926 -2356 -922 -2348
rect -917 -2356 -913 -2348
rect -909 -2356 -905 -2348
rect -901 -2356 -897 -2348
rect -889 -2356 -885 -2348
rect -877 -2356 -873 -2348
rect -868 -2356 -864 -2348
rect -859 -2356 -855 -2348
rect -847 -2356 -843 -2348
rect -835 -2356 -831 -2348
rect -826 -2356 -822 -2348
rect -817 -2356 -813 -2348
rect -805 -2356 -801 -2348
rect -793 -2356 -789 -2348
rect -784 -2356 -780 -2348
rect -775 -2356 -771 -2348
rect -763 -2356 -759 -2348
rect -751 -2356 -747 -2348
rect -743 -2356 -739 -2348
rect -577 -2356 -573 -2348
rect -568 -2356 -564 -2348
rect -559 -2356 -555 -2348
rect -551 -2356 -547 -2348
rect -543 -2356 -539 -2348
rect -531 -2356 -527 -2348
rect -519 -2356 -515 -2348
rect -510 -2356 -506 -2348
rect -501 -2356 -497 -2348
rect -489 -2356 -485 -2348
rect -477 -2356 -473 -2348
rect -468 -2356 -464 -2348
rect -459 -2356 -455 -2348
rect -447 -2356 -443 -2348
rect -435 -2356 -431 -2348
rect -426 -2356 -422 -2348
rect -417 -2356 -413 -2348
rect -405 -2356 -401 -2348
rect -393 -2356 -389 -2348
rect -385 -2356 -381 -2348
rect -219 -2356 -215 -2348
rect -210 -2356 -206 -2348
rect -201 -2356 -197 -2348
rect -193 -2356 -189 -2348
rect -185 -2356 -181 -2348
rect -173 -2356 -169 -2348
rect -161 -2356 -157 -2348
rect -152 -2356 -148 -2348
rect -143 -2356 -139 -2348
rect -131 -2356 -127 -2348
rect -119 -2356 -115 -2348
rect -110 -2356 -106 -2348
rect -101 -2356 -97 -2348
rect -89 -2356 -85 -2348
rect -77 -2356 -73 -2348
rect -68 -2356 -64 -2348
rect -59 -2356 -55 -2348
rect -47 -2356 -43 -2348
rect -35 -2356 -31 -2348
rect -27 -2356 -23 -2348
rect 139 -2356 143 -2348
rect 148 -2356 152 -2348
rect 157 -2356 161 -2348
rect 165 -2356 169 -2348
rect 173 -2356 177 -2348
rect 185 -2356 189 -2348
rect 197 -2356 201 -2348
rect 206 -2356 210 -2348
rect 215 -2356 219 -2348
rect 227 -2356 231 -2348
rect 239 -2356 243 -2348
rect 248 -2356 252 -2348
rect 257 -2356 261 -2348
rect 269 -2356 273 -2348
rect 281 -2356 285 -2348
rect 290 -2356 294 -2348
rect 299 -2356 303 -2348
rect 311 -2356 315 -2348
rect 323 -2356 327 -2348
rect 331 -2356 335 -2348
rect 495 -2356 499 -2348
rect 504 -2356 508 -2348
rect 513 -2356 517 -2348
rect 521 -2356 525 -2348
rect 529 -2356 533 -2348
rect 541 -2356 545 -2348
rect 553 -2356 557 -2348
rect 562 -2356 566 -2348
rect 571 -2356 575 -2348
rect 583 -2356 587 -2348
rect 595 -2356 599 -2348
rect 604 -2356 608 -2348
rect 613 -2356 617 -2348
rect 625 -2356 629 -2348
rect 637 -2356 641 -2348
rect 646 -2356 650 -2348
rect 655 -2356 659 -2348
rect 667 -2356 671 -2348
rect 679 -2356 683 -2348
rect 687 -2356 691 -2348
rect 853 -2356 857 -2348
rect 862 -2356 866 -2348
rect 871 -2356 875 -2348
rect 879 -2356 883 -2348
rect 887 -2356 891 -2348
rect 899 -2356 903 -2348
rect 911 -2356 915 -2348
rect 920 -2356 924 -2348
rect 929 -2356 933 -2348
rect 941 -2356 945 -2348
rect 953 -2356 957 -2348
rect 962 -2356 966 -2348
rect 971 -2356 975 -2348
rect 983 -2356 987 -2348
rect 995 -2356 999 -2348
rect 1004 -2356 1008 -2348
rect 1013 -2356 1017 -2348
rect 1025 -2356 1029 -2348
rect 1037 -2356 1041 -2348
rect 1045 -2356 1049 -2348
rect 1211 -2356 1215 -2348
rect 1220 -2356 1224 -2348
rect 1229 -2356 1233 -2348
rect 1237 -2356 1241 -2348
rect 1245 -2356 1249 -2348
rect 1257 -2356 1261 -2348
rect 1269 -2356 1273 -2348
rect 1278 -2356 1282 -2348
rect 1287 -2356 1291 -2348
rect 1299 -2356 1303 -2348
rect 1311 -2356 1315 -2348
rect 1320 -2356 1324 -2348
rect 1329 -2356 1333 -2348
rect 1341 -2356 1345 -2348
rect 1353 -2356 1357 -2348
rect 1362 -2356 1366 -2348
rect 1371 -2356 1375 -2348
rect 1383 -2356 1387 -2348
rect 1395 -2356 1399 -2348
rect 1403 -2356 1407 -2348
rect -1559 -2527 -1555 -2519
rect -1550 -2527 -1546 -2519
rect -1541 -2527 -1537 -2519
rect -1533 -2527 -1529 -2519
rect -1525 -2527 -1521 -2519
rect -1513 -2527 -1509 -2519
rect -1501 -2527 -1497 -2519
rect -1492 -2527 -1488 -2519
rect -1483 -2527 -1479 -2519
rect -1471 -2527 -1467 -2519
rect -1459 -2527 -1455 -2519
rect -1450 -2527 -1446 -2519
rect -1441 -2527 -1437 -2519
rect -1429 -2527 -1425 -2519
rect -1417 -2527 -1413 -2519
rect -1408 -2527 -1404 -2519
rect -1399 -2527 -1395 -2519
rect -1387 -2527 -1383 -2519
rect -1375 -2527 -1371 -2519
rect -1367 -2527 -1363 -2519
rect -1234 -2527 -1230 -2519
rect -1225 -2527 -1221 -2519
rect -1216 -2527 -1212 -2519
rect -1208 -2527 -1204 -2519
rect -1200 -2527 -1196 -2519
rect -1188 -2527 -1184 -2519
rect -1176 -2527 -1172 -2519
rect -1167 -2527 -1163 -2519
rect -1158 -2527 -1154 -2519
rect -1146 -2527 -1142 -2519
rect -1134 -2527 -1130 -2519
rect -1125 -2527 -1121 -2519
rect -1116 -2527 -1112 -2519
rect -1104 -2527 -1100 -2519
rect -1092 -2527 -1088 -2519
rect -1083 -2527 -1079 -2519
rect -1074 -2527 -1070 -2519
rect -1062 -2527 -1058 -2519
rect -1050 -2527 -1046 -2519
rect -1042 -2527 -1038 -2519
rect -935 -2527 -931 -2519
rect -926 -2527 -922 -2519
rect -917 -2527 -913 -2519
rect -909 -2527 -905 -2519
rect -901 -2527 -897 -2519
rect -889 -2527 -885 -2519
rect -877 -2527 -873 -2519
rect -868 -2527 -864 -2519
rect -859 -2527 -855 -2519
rect -847 -2527 -843 -2519
rect -835 -2527 -831 -2519
rect -826 -2527 -822 -2519
rect -817 -2527 -813 -2519
rect -805 -2527 -801 -2519
rect -793 -2527 -789 -2519
rect -784 -2527 -780 -2519
rect -775 -2527 -771 -2519
rect -763 -2527 -759 -2519
rect -751 -2527 -747 -2519
rect -743 -2527 -739 -2519
rect -577 -2527 -573 -2519
rect -568 -2527 -564 -2519
rect -559 -2527 -555 -2519
rect -551 -2527 -547 -2519
rect -543 -2527 -539 -2519
rect -531 -2527 -527 -2519
rect -519 -2527 -515 -2519
rect -510 -2527 -506 -2519
rect -501 -2527 -497 -2519
rect -489 -2527 -485 -2519
rect -477 -2527 -473 -2519
rect -468 -2527 -464 -2519
rect -459 -2527 -455 -2519
rect -447 -2527 -443 -2519
rect -435 -2527 -431 -2519
rect -426 -2527 -422 -2519
rect -417 -2527 -413 -2519
rect -405 -2527 -401 -2519
rect -393 -2527 -389 -2519
rect -385 -2527 -381 -2519
rect -220 -2527 -216 -2519
rect -211 -2527 -207 -2519
rect -202 -2527 -198 -2519
rect -194 -2527 -190 -2519
rect -186 -2527 -182 -2519
rect -174 -2527 -170 -2519
rect -162 -2527 -158 -2519
rect -153 -2527 -149 -2519
rect -144 -2527 -140 -2519
rect -132 -2527 -128 -2519
rect -120 -2527 -116 -2519
rect -111 -2527 -107 -2519
rect -102 -2527 -98 -2519
rect -90 -2527 -86 -2519
rect -78 -2527 -74 -2519
rect -69 -2527 -65 -2519
rect -60 -2527 -56 -2519
rect -48 -2527 -44 -2519
rect -36 -2527 -32 -2519
rect -28 -2527 -24 -2519
rect 139 -2527 143 -2519
rect 148 -2527 152 -2519
rect 157 -2527 161 -2519
rect 165 -2527 169 -2519
rect 173 -2527 177 -2519
rect 185 -2527 189 -2519
rect 197 -2527 201 -2519
rect 206 -2527 210 -2519
rect 215 -2527 219 -2519
rect 227 -2527 231 -2519
rect 239 -2527 243 -2519
rect 248 -2527 252 -2519
rect 257 -2527 261 -2519
rect 269 -2527 273 -2519
rect 281 -2527 285 -2519
rect 290 -2527 294 -2519
rect 299 -2527 303 -2519
rect 311 -2527 315 -2519
rect 323 -2527 327 -2519
rect 331 -2527 335 -2519
rect 495 -2527 499 -2519
rect 504 -2527 508 -2519
rect 513 -2527 517 -2519
rect 521 -2527 525 -2519
rect 529 -2527 533 -2519
rect 541 -2527 545 -2519
rect 553 -2527 557 -2519
rect 562 -2527 566 -2519
rect 571 -2527 575 -2519
rect 583 -2527 587 -2519
rect 595 -2527 599 -2519
rect 604 -2527 608 -2519
rect 613 -2527 617 -2519
rect 625 -2527 629 -2519
rect 637 -2527 641 -2519
rect 646 -2527 650 -2519
rect 655 -2527 659 -2519
rect 667 -2527 671 -2519
rect 679 -2527 683 -2519
rect 687 -2527 691 -2519
rect 853 -2527 857 -2519
rect 862 -2527 866 -2519
rect 871 -2527 875 -2519
rect 879 -2527 883 -2519
rect 887 -2527 891 -2519
rect 899 -2527 903 -2519
rect 911 -2527 915 -2519
rect 920 -2527 924 -2519
rect 929 -2527 933 -2519
rect 941 -2527 945 -2519
rect 953 -2527 957 -2519
rect 962 -2527 966 -2519
rect 971 -2527 975 -2519
rect 983 -2527 987 -2519
rect 995 -2527 999 -2519
rect 1004 -2527 1008 -2519
rect 1013 -2527 1017 -2519
rect 1025 -2527 1029 -2519
rect 1037 -2527 1041 -2519
rect 1045 -2527 1049 -2519
rect 1211 -2527 1215 -2519
rect 1220 -2527 1224 -2519
rect 1229 -2527 1233 -2519
rect 1237 -2527 1241 -2519
rect 1245 -2527 1249 -2519
rect 1257 -2527 1261 -2519
rect 1269 -2527 1273 -2519
rect 1278 -2527 1282 -2519
rect 1287 -2527 1291 -2519
rect 1299 -2527 1303 -2519
rect 1311 -2527 1315 -2519
rect 1320 -2527 1324 -2519
rect 1329 -2527 1333 -2519
rect 1341 -2527 1345 -2519
rect 1353 -2527 1357 -2519
rect 1362 -2527 1366 -2519
rect 1371 -2527 1375 -2519
rect 1383 -2527 1387 -2519
rect 1395 -2527 1399 -2519
rect 1403 -2527 1407 -2519
rect -1309 -2632 -1305 -2624
rect -1301 -2632 -1297 -2624
rect -1292 -2632 -1288 -2624
rect -1283 -2632 -1279 -2624
rect -935 -2632 -931 -2624
rect -927 -2632 -923 -2624
rect -918 -2632 -914 -2624
rect -909 -2632 -905 -2624
rect -577 -2632 -573 -2624
rect -569 -2632 -565 -2624
rect -560 -2632 -556 -2624
rect -551 -2632 -547 -2624
rect -219 -2632 -215 -2624
rect -211 -2632 -207 -2624
rect -202 -2632 -198 -2624
rect -193 -2632 -189 -2624
rect 139 -2632 143 -2624
rect 147 -2632 151 -2624
rect 156 -2632 160 -2624
rect 165 -2632 169 -2624
rect 495 -2632 499 -2624
rect 503 -2632 507 -2624
rect 512 -2632 516 -2624
rect 521 -2632 525 -2624
rect 853 -2632 857 -2624
rect 861 -2632 865 -2624
rect 870 -2632 874 -2624
rect 879 -2632 883 -2624
rect 1211 -2632 1215 -2624
rect 1219 -2632 1223 -2624
rect 1228 -2632 1232 -2624
rect 1237 -2632 1241 -2624
rect -1234 -2791 -1230 -2783
rect -1225 -2791 -1221 -2783
rect -1216 -2791 -1212 -2783
rect -1208 -2791 -1204 -2783
rect -1190 -2791 -1186 -2783
rect -1168 -2791 -1164 -2783
rect -1156 -2791 -1152 -2783
rect -1147 -2791 -1143 -2783
rect -1138 -2791 -1134 -2783
rect -935 -2791 -931 -2783
rect -926 -2791 -922 -2783
rect -917 -2791 -913 -2783
rect -909 -2791 -905 -2783
rect -900 -2791 -896 -2783
rect -891 -2791 -887 -2783
rect -883 -2791 -879 -2783
rect -865 -2791 -861 -2783
rect -843 -2791 -839 -2783
rect -831 -2791 -827 -2783
rect -822 -2791 -818 -2783
rect -813 -2791 -809 -2783
rect -805 -2791 -801 -2783
rect -787 -2791 -783 -2783
rect -765 -2791 -761 -2783
rect -753 -2791 -749 -2783
rect -741 -2791 -737 -2783
rect -729 -2791 -725 -2783
rect -721 -2791 -717 -2783
rect -704 -2791 -700 -2783
rect -695 -2791 -691 -2783
rect -577 -2791 -573 -2783
rect -568 -2791 -564 -2783
rect -559 -2791 -555 -2783
rect -551 -2791 -547 -2783
rect -542 -2791 -538 -2783
rect -533 -2791 -529 -2783
rect -525 -2791 -521 -2783
rect -507 -2791 -503 -2783
rect -485 -2791 -481 -2783
rect -473 -2791 -469 -2783
rect -464 -2791 -460 -2783
rect -455 -2791 -451 -2783
rect -447 -2791 -443 -2783
rect -429 -2791 -425 -2783
rect -407 -2791 -403 -2783
rect -395 -2791 -391 -2783
rect -383 -2791 -379 -2783
rect -371 -2791 -367 -2783
rect -363 -2791 -359 -2783
rect -346 -2791 -342 -2783
rect -337 -2791 -333 -2783
rect -219 -2791 -215 -2783
rect -210 -2791 -206 -2783
rect -201 -2791 -197 -2783
rect -193 -2791 -189 -2783
rect -184 -2791 -180 -2783
rect -175 -2791 -171 -2783
rect -167 -2791 -163 -2783
rect -149 -2791 -145 -2783
rect -127 -2791 -123 -2783
rect -115 -2791 -111 -2783
rect -106 -2791 -102 -2783
rect -97 -2791 -93 -2783
rect -89 -2791 -85 -2783
rect -71 -2791 -67 -2783
rect -49 -2791 -45 -2783
rect -37 -2791 -33 -2783
rect -25 -2791 -21 -2783
rect -13 -2791 -9 -2783
rect -5 -2791 -1 -2783
rect 12 -2791 16 -2783
rect 21 -2791 25 -2783
rect 139 -2791 143 -2783
rect 148 -2791 152 -2783
rect 157 -2791 161 -2783
rect 165 -2791 169 -2783
rect 174 -2791 178 -2783
rect 183 -2791 187 -2783
rect 191 -2791 195 -2783
rect 209 -2791 213 -2783
rect 231 -2791 235 -2783
rect 243 -2791 247 -2783
rect 252 -2791 256 -2783
rect 261 -2791 265 -2783
rect 269 -2791 273 -2783
rect 287 -2791 291 -2783
rect 309 -2791 313 -2783
rect 321 -2791 325 -2783
rect 333 -2791 337 -2783
rect 345 -2791 349 -2783
rect 353 -2791 357 -2783
rect 370 -2791 374 -2783
rect 379 -2791 383 -2783
rect 495 -2791 499 -2783
rect 504 -2791 508 -2783
rect 513 -2791 517 -2783
rect 521 -2791 525 -2783
rect 530 -2791 534 -2783
rect 539 -2791 543 -2783
rect 547 -2791 551 -2783
rect 565 -2791 569 -2783
rect 587 -2791 591 -2783
rect 599 -2791 603 -2783
rect 608 -2791 612 -2783
rect 617 -2791 621 -2783
rect 625 -2791 629 -2783
rect 643 -2791 647 -2783
rect 665 -2791 669 -2783
rect 677 -2791 681 -2783
rect 689 -2791 693 -2783
rect 701 -2791 705 -2783
rect 709 -2791 713 -2783
rect 726 -2791 730 -2783
rect 735 -2791 739 -2783
rect 853 -2791 857 -2783
rect 862 -2791 866 -2783
rect 871 -2791 875 -2783
rect 879 -2791 883 -2783
rect 888 -2791 892 -2783
rect 897 -2791 901 -2783
rect 905 -2791 909 -2783
rect 923 -2791 927 -2783
rect 945 -2791 949 -2783
rect 957 -2791 961 -2783
rect 966 -2791 970 -2783
rect 975 -2791 979 -2783
rect 983 -2791 987 -2783
rect 1001 -2791 1005 -2783
rect 1023 -2791 1027 -2783
rect 1035 -2791 1039 -2783
rect 1047 -2791 1051 -2783
rect 1059 -2791 1063 -2783
rect 1067 -2791 1071 -2783
rect 1084 -2791 1088 -2783
rect 1093 -2791 1097 -2783
rect 1211 -2791 1215 -2783
rect 1220 -2791 1224 -2783
rect 1229 -2791 1233 -2783
rect 1237 -2791 1241 -2783
rect 1246 -2791 1250 -2783
rect 1255 -2791 1259 -2783
rect 1263 -2791 1267 -2783
rect 1281 -2791 1285 -2783
rect 1303 -2791 1307 -2783
rect 1315 -2791 1319 -2783
rect 1324 -2791 1328 -2783
rect 1333 -2791 1337 -2783
rect 1341 -2791 1345 -2783
rect 1359 -2791 1363 -2783
rect 1381 -2791 1385 -2783
rect 1393 -2791 1397 -2783
rect 1405 -2791 1409 -2783
rect 1417 -2791 1421 -2783
rect 1425 -2791 1429 -2783
rect 1442 -2791 1446 -2783
rect 1451 -2791 1455 -2783
rect -1559 -2910 -1555 -2902
rect -1550 -2910 -1546 -2902
rect -1541 -2910 -1537 -2902
rect -1533 -2910 -1529 -2902
rect -1525 -2910 -1521 -2902
rect -1513 -2910 -1509 -2902
rect -1501 -2910 -1497 -2902
rect -1492 -2910 -1488 -2902
rect -1483 -2910 -1479 -2902
rect -1471 -2910 -1467 -2902
rect -1459 -2910 -1455 -2902
rect -1450 -2910 -1446 -2902
rect -1441 -2910 -1437 -2902
rect -1429 -2910 -1425 -2902
rect -1417 -2910 -1413 -2902
rect -1408 -2910 -1404 -2902
rect -1399 -2910 -1395 -2902
rect -1387 -2910 -1383 -2902
rect -1375 -2910 -1371 -2902
rect -1367 -2910 -1363 -2902
rect -1234 -2910 -1230 -2902
rect -1225 -2910 -1221 -2902
rect -1216 -2910 -1212 -2902
rect -1208 -2910 -1204 -2902
rect -1200 -2910 -1196 -2902
rect -1188 -2910 -1184 -2902
rect -1176 -2910 -1172 -2902
rect -1167 -2910 -1163 -2902
rect -1158 -2910 -1154 -2902
rect -1146 -2910 -1142 -2902
rect -1134 -2910 -1130 -2902
rect -1125 -2910 -1121 -2902
rect -1116 -2910 -1112 -2902
rect -1104 -2910 -1100 -2902
rect -1092 -2910 -1088 -2902
rect -1083 -2910 -1079 -2902
rect -1074 -2910 -1070 -2902
rect -1062 -2910 -1058 -2902
rect -1050 -2910 -1046 -2902
rect -1042 -2910 -1038 -2902
rect -935 -2910 -931 -2902
rect -926 -2910 -922 -2902
rect -917 -2910 -913 -2902
rect -909 -2910 -905 -2902
rect -901 -2910 -897 -2902
rect -889 -2910 -885 -2902
rect -877 -2910 -873 -2902
rect -868 -2910 -864 -2902
rect -859 -2910 -855 -2902
rect -847 -2910 -843 -2902
rect -835 -2910 -831 -2902
rect -826 -2910 -822 -2902
rect -817 -2910 -813 -2902
rect -805 -2910 -801 -2902
rect -793 -2910 -789 -2902
rect -784 -2910 -780 -2902
rect -775 -2910 -771 -2902
rect -763 -2910 -759 -2902
rect -751 -2910 -747 -2902
rect -743 -2910 -739 -2902
rect -577 -2910 -573 -2902
rect -568 -2910 -564 -2902
rect -559 -2910 -555 -2902
rect -551 -2910 -547 -2902
rect -543 -2910 -539 -2902
rect -531 -2910 -527 -2902
rect -519 -2910 -515 -2902
rect -510 -2910 -506 -2902
rect -501 -2910 -497 -2902
rect -489 -2910 -485 -2902
rect -477 -2910 -473 -2902
rect -468 -2910 -464 -2902
rect -459 -2910 -455 -2902
rect -447 -2910 -443 -2902
rect -435 -2910 -431 -2902
rect -426 -2910 -422 -2902
rect -417 -2910 -413 -2902
rect -405 -2910 -401 -2902
rect -393 -2910 -389 -2902
rect -385 -2910 -381 -2902
rect -219 -2910 -215 -2902
rect -210 -2910 -206 -2902
rect -201 -2910 -197 -2902
rect -193 -2910 -189 -2902
rect -185 -2910 -181 -2902
rect -173 -2910 -169 -2902
rect -161 -2910 -157 -2902
rect -152 -2910 -148 -2902
rect -143 -2910 -139 -2902
rect -131 -2910 -127 -2902
rect -119 -2910 -115 -2902
rect -110 -2910 -106 -2902
rect -101 -2910 -97 -2902
rect -89 -2910 -85 -2902
rect -77 -2910 -73 -2902
rect -68 -2910 -64 -2902
rect -59 -2910 -55 -2902
rect -47 -2910 -43 -2902
rect -35 -2910 -31 -2902
rect -27 -2910 -23 -2902
rect 139 -2910 143 -2902
rect 148 -2910 152 -2902
rect 157 -2910 161 -2902
rect 165 -2910 169 -2902
rect 173 -2910 177 -2902
rect 185 -2910 189 -2902
rect 197 -2910 201 -2902
rect 206 -2910 210 -2902
rect 215 -2910 219 -2902
rect 227 -2910 231 -2902
rect 239 -2910 243 -2902
rect 248 -2910 252 -2902
rect 257 -2910 261 -2902
rect 269 -2910 273 -2902
rect 281 -2910 285 -2902
rect 290 -2910 294 -2902
rect 299 -2910 303 -2902
rect 311 -2910 315 -2902
rect 323 -2910 327 -2902
rect 331 -2910 335 -2902
rect -1559 -3081 -1555 -3073
rect -1550 -3081 -1546 -3073
rect -1541 -3081 -1537 -3073
rect -1533 -3081 -1529 -3073
rect -1525 -3081 -1521 -3073
rect -1513 -3081 -1509 -3073
rect -1501 -3081 -1497 -3073
rect -1492 -3081 -1488 -3073
rect -1483 -3081 -1479 -3073
rect -1471 -3081 -1467 -3073
rect -1459 -3081 -1455 -3073
rect -1450 -3081 -1446 -3073
rect -1441 -3081 -1437 -3073
rect -1429 -3081 -1425 -3073
rect -1417 -3081 -1413 -3073
rect -1408 -3081 -1404 -3073
rect -1399 -3081 -1395 -3073
rect -1387 -3081 -1383 -3073
rect -1375 -3081 -1371 -3073
rect -1367 -3081 -1363 -3073
rect -1234 -3081 -1230 -3073
rect -1225 -3081 -1221 -3073
rect -1216 -3081 -1212 -3073
rect -1208 -3081 -1204 -3073
rect -1200 -3081 -1196 -3073
rect -1188 -3081 -1184 -3073
rect -1176 -3081 -1172 -3073
rect -1167 -3081 -1163 -3073
rect -1158 -3081 -1154 -3073
rect -1146 -3081 -1142 -3073
rect -1134 -3081 -1130 -3073
rect -1125 -3081 -1121 -3073
rect -1116 -3081 -1112 -3073
rect -1104 -3081 -1100 -3073
rect -1092 -3081 -1088 -3073
rect -1083 -3081 -1079 -3073
rect -1074 -3081 -1070 -3073
rect -1062 -3081 -1058 -3073
rect -1050 -3081 -1046 -3073
rect -1042 -3081 -1038 -3073
rect -935 -3081 -931 -3073
rect -926 -3081 -922 -3073
rect -917 -3081 -913 -3073
rect -909 -3081 -905 -3073
rect -901 -3081 -897 -3073
rect -889 -3081 -885 -3073
rect -877 -3081 -873 -3073
rect -868 -3081 -864 -3073
rect -859 -3081 -855 -3073
rect -847 -3081 -843 -3073
rect -835 -3081 -831 -3073
rect -826 -3081 -822 -3073
rect -817 -3081 -813 -3073
rect -805 -3081 -801 -3073
rect -793 -3081 -789 -3073
rect -784 -3081 -780 -3073
rect -775 -3081 -771 -3073
rect -763 -3081 -759 -3073
rect -751 -3081 -747 -3073
rect -743 -3081 -739 -3073
rect -577 -3081 -573 -3073
rect -568 -3081 -564 -3073
rect -559 -3081 -555 -3073
rect -551 -3081 -547 -3073
rect -543 -3081 -539 -3073
rect -531 -3081 -527 -3073
rect -519 -3081 -515 -3073
rect -510 -3081 -506 -3073
rect -501 -3081 -497 -3073
rect -489 -3081 -485 -3073
rect -477 -3081 -473 -3073
rect -468 -3081 -464 -3073
rect -459 -3081 -455 -3073
rect -447 -3081 -443 -3073
rect -435 -3081 -431 -3073
rect -426 -3081 -422 -3073
rect -417 -3081 -413 -3073
rect -405 -3081 -401 -3073
rect -393 -3081 -389 -3073
rect -385 -3081 -381 -3073
rect -219 -3081 -215 -3073
rect -210 -3081 -206 -3073
rect -201 -3081 -197 -3073
rect -193 -3081 -189 -3073
rect -185 -3081 -181 -3073
rect -173 -3081 -169 -3073
rect -161 -3081 -157 -3073
rect -152 -3081 -148 -3073
rect -143 -3081 -139 -3073
rect -131 -3081 -127 -3073
rect -119 -3081 -115 -3073
rect -110 -3081 -106 -3073
rect -101 -3081 -97 -3073
rect -89 -3081 -85 -3073
rect -77 -3081 -73 -3073
rect -68 -3081 -64 -3073
rect -59 -3081 -55 -3073
rect -47 -3081 -43 -3073
rect -35 -3081 -31 -3073
rect -27 -3081 -23 -3073
rect 139 -3081 143 -3073
rect 148 -3081 152 -3073
rect 157 -3081 161 -3073
rect 165 -3081 169 -3073
rect 173 -3081 177 -3073
rect 185 -3081 189 -3073
rect 197 -3081 201 -3073
rect 206 -3081 210 -3073
rect 215 -3081 219 -3073
rect 227 -3081 231 -3073
rect 239 -3081 243 -3073
rect 248 -3081 252 -3073
rect 257 -3081 261 -3073
rect 269 -3081 273 -3073
rect 281 -3081 285 -3073
rect 290 -3081 294 -3073
rect 299 -3081 303 -3073
rect 311 -3081 315 -3073
rect 323 -3081 327 -3073
rect 331 -3081 335 -3073
rect 495 -3081 499 -3073
rect 504 -3081 508 -3073
rect 513 -3081 517 -3073
rect 521 -3081 525 -3073
rect 529 -3081 533 -3073
rect 541 -3081 545 -3073
rect 553 -3081 557 -3073
rect 562 -3081 566 -3073
rect 571 -3081 575 -3073
rect 583 -3081 587 -3073
rect 595 -3081 599 -3073
rect 604 -3081 608 -3073
rect 613 -3081 617 -3073
rect 625 -3081 629 -3073
rect 637 -3081 641 -3073
rect 646 -3081 650 -3073
rect 655 -3081 659 -3073
rect 667 -3081 671 -3073
rect 679 -3081 683 -3073
rect 687 -3081 691 -3073
rect 853 -3081 857 -3073
rect 862 -3081 866 -3073
rect 871 -3081 875 -3073
rect 879 -3081 883 -3073
rect 887 -3081 891 -3073
rect 899 -3081 903 -3073
rect 911 -3081 915 -3073
rect 920 -3081 924 -3073
rect 929 -3081 933 -3073
rect 941 -3081 945 -3073
rect 953 -3081 957 -3073
rect 962 -3081 966 -3073
rect 971 -3081 975 -3073
rect 983 -3081 987 -3073
rect 995 -3081 999 -3073
rect 1004 -3081 1008 -3073
rect 1013 -3081 1017 -3073
rect 1025 -3081 1029 -3073
rect 1037 -3081 1041 -3073
rect 1045 -3081 1049 -3073
rect 1211 -3081 1215 -3073
rect 1220 -3081 1224 -3073
rect 1229 -3081 1233 -3073
rect 1237 -3081 1241 -3073
rect 1245 -3081 1249 -3073
rect 1257 -3081 1261 -3073
rect 1269 -3081 1273 -3073
rect 1278 -3081 1282 -3073
rect 1287 -3081 1291 -3073
rect 1299 -3081 1303 -3073
rect 1311 -3081 1315 -3073
rect 1320 -3081 1324 -3073
rect 1329 -3081 1333 -3073
rect 1341 -3081 1345 -3073
rect 1353 -3081 1357 -3073
rect 1362 -3081 1366 -3073
rect 1371 -3081 1375 -3073
rect 1383 -3081 1387 -3073
rect 1395 -3081 1399 -3073
rect 1403 -3081 1407 -3073
rect -1559 -3252 -1555 -3244
rect -1550 -3252 -1546 -3244
rect -1541 -3252 -1537 -3244
rect -1533 -3252 -1529 -3244
rect -1525 -3252 -1521 -3244
rect -1513 -3252 -1509 -3244
rect -1501 -3252 -1497 -3244
rect -1492 -3252 -1488 -3244
rect -1483 -3252 -1479 -3244
rect -1471 -3252 -1467 -3244
rect -1459 -3252 -1455 -3244
rect -1450 -3252 -1446 -3244
rect -1441 -3252 -1437 -3244
rect -1429 -3252 -1425 -3244
rect -1417 -3252 -1413 -3244
rect -1408 -3252 -1404 -3244
rect -1399 -3252 -1395 -3244
rect -1387 -3252 -1383 -3244
rect -1375 -3252 -1371 -3244
rect -1367 -3252 -1363 -3244
rect -1234 -3252 -1230 -3244
rect -1225 -3252 -1221 -3244
rect -1216 -3252 -1212 -3244
rect -1208 -3252 -1204 -3244
rect -1200 -3252 -1196 -3244
rect -1188 -3252 -1184 -3244
rect -1176 -3252 -1172 -3244
rect -1167 -3252 -1163 -3244
rect -1158 -3252 -1154 -3244
rect -1146 -3252 -1142 -3244
rect -1134 -3252 -1130 -3244
rect -1125 -3252 -1121 -3244
rect -1116 -3252 -1112 -3244
rect -1104 -3252 -1100 -3244
rect -1092 -3252 -1088 -3244
rect -1083 -3252 -1079 -3244
rect -1074 -3252 -1070 -3244
rect -1062 -3252 -1058 -3244
rect -1050 -3252 -1046 -3244
rect -1042 -3252 -1038 -3244
rect -935 -3252 -931 -3244
rect -926 -3252 -922 -3244
rect -917 -3252 -913 -3244
rect -909 -3252 -905 -3244
rect -901 -3252 -897 -3244
rect -889 -3252 -885 -3244
rect -877 -3252 -873 -3244
rect -868 -3252 -864 -3244
rect -859 -3252 -855 -3244
rect -847 -3252 -843 -3244
rect -835 -3252 -831 -3244
rect -826 -3252 -822 -3244
rect -817 -3252 -813 -3244
rect -805 -3252 -801 -3244
rect -793 -3252 -789 -3244
rect -784 -3252 -780 -3244
rect -775 -3252 -771 -3244
rect -763 -3252 -759 -3244
rect -751 -3252 -747 -3244
rect -743 -3252 -739 -3244
rect -577 -3252 -573 -3244
rect -568 -3252 -564 -3244
rect -559 -3252 -555 -3244
rect -551 -3252 -547 -3244
rect -543 -3252 -539 -3244
rect -531 -3252 -527 -3244
rect -519 -3252 -515 -3244
rect -510 -3252 -506 -3244
rect -501 -3252 -497 -3244
rect -489 -3252 -485 -3244
rect -477 -3252 -473 -3244
rect -468 -3252 -464 -3244
rect -459 -3252 -455 -3244
rect -447 -3252 -443 -3244
rect -435 -3252 -431 -3244
rect -426 -3252 -422 -3244
rect -417 -3252 -413 -3244
rect -405 -3252 -401 -3244
rect -393 -3252 -389 -3244
rect -385 -3252 -381 -3244
rect -219 -3252 -215 -3244
rect -210 -3252 -206 -3244
rect -201 -3252 -197 -3244
rect -193 -3252 -189 -3244
rect -185 -3252 -181 -3244
rect -173 -3252 -169 -3244
rect -161 -3252 -157 -3244
rect -152 -3252 -148 -3244
rect -143 -3252 -139 -3244
rect -131 -3252 -127 -3244
rect -119 -3252 -115 -3244
rect -110 -3252 -106 -3244
rect -101 -3252 -97 -3244
rect -89 -3252 -85 -3244
rect -77 -3252 -73 -3244
rect -68 -3252 -64 -3244
rect -59 -3252 -55 -3244
rect -47 -3252 -43 -3244
rect -35 -3252 -31 -3244
rect -27 -3252 -23 -3244
rect 139 -3252 143 -3244
rect 148 -3252 152 -3244
rect 157 -3252 161 -3244
rect 165 -3252 169 -3244
rect 173 -3252 177 -3244
rect 185 -3252 189 -3244
rect 197 -3252 201 -3244
rect 206 -3252 210 -3244
rect 215 -3252 219 -3244
rect 227 -3252 231 -3244
rect 239 -3252 243 -3244
rect 248 -3252 252 -3244
rect 257 -3252 261 -3244
rect 269 -3252 273 -3244
rect 281 -3252 285 -3244
rect 290 -3252 294 -3244
rect 299 -3252 303 -3244
rect 311 -3252 315 -3244
rect 323 -3252 327 -3244
rect 331 -3252 335 -3244
rect 495 -3252 499 -3244
rect 504 -3252 508 -3244
rect 513 -3252 517 -3244
rect 521 -3252 525 -3244
rect 529 -3252 533 -3244
rect 541 -3252 545 -3244
rect 553 -3252 557 -3244
rect 562 -3252 566 -3244
rect 571 -3252 575 -3244
rect 583 -3252 587 -3244
rect 595 -3252 599 -3244
rect 604 -3252 608 -3244
rect 613 -3252 617 -3244
rect 625 -3252 629 -3244
rect 637 -3252 641 -3244
rect 646 -3252 650 -3244
rect 655 -3252 659 -3244
rect 667 -3252 671 -3244
rect 679 -3252 683 -3244
rect 687 -3252 691 -3244
rect 853 -3252 857 -3244
rect 862 -3252 866 -3244
rect 871 -3252 875 -3244
rect 879 -3252 883 -3244
rect 887 -3252 891 -3244
rect 899 -3252 903 -3244
rect 911 -3252 915 -3244
rect 920 -3252 924 -3244
rect 929 -3252 933 -3244
rect 941 -3252 945 -3244
rect 953 -3252 957 -3244
rect 962 -3252 966 -3244
rect 971 -3252 975 -3244
rect 983 -3252 987 -3244
rect 995 -3252 999 -3244
rect 1004 -3252 1008 -3244
rect 1013 -3252 1017 -3244
rect 1025 -3252 1029 -3244
rect 1037 -3252 1041 -3244
rect 1045 -3252 1049 -3244
rect 1211 -3252 1215 -3244
rect 1220 -3252 1224 -3244
rect 1229 -3252 1233 -3244
rect 1237 -3252 1241 -3244
rect 1245 -3252 1249 -3244
rect 1257 -3252 1261 -3244
rect 1269 -3252 1273 -3244
rect 1278 -3252 1282 -3244
rect 1287 -3252 1291 -3244
rect 1299 -3252 1303 -3244
rect 1311 -3252 1315 -3244
rect 1320 -3252 1324 -3244
rect 1329 -3252 1333 -3244
rect 1341 -3252 1345 -3244
rect 1353 -3252 1357 -3244
rect 1362 -3252 1366 -3244
rect 1371 -3252 1375 -3244
rect 1383 -3252 1387 -3244
rect 1395 -3252 1399 -3244
rect 1403 -3252 1407 -3244
rect -1309 -3363 -1305 -3355
rect -1301 -3363 -1297 -3355
rect -1292 -3363 -1288 -3355
rect -1283 -3363 -1279 -3355
rect -935 -3363 -931 -3355
rect -927 -3363 -923 -3355
rect -918 -3363 -914 -3355
rect -909 -3363 -905 -3355
rect -577 -3363 -573 -3355
rect -569 -3363 -565 -3355
rect -560 -3363 -556 -3355
rect -551 -3363 -547 -3355
rect -219 -3363 -215 -3355
rect -211 -3363 -207 -3355
rect -202 -3363 -198 -3355
rect -193 -3363 -189 -3355
rect 139 -3363 143 -3355
rect 147 -3363 151 -3355
rect 156 -3363 160 -3355
rect 165 -3363 169 -3355
rect 495 -3363 499 -3355
rect 503 -3363 507 -3355
rect 512 -3363 516 -3355
rect 521 -3363 525 -3355
rect 853 -3363 857 -3355
rect 861 -3363 865 -3355
rect 870 -3363 874 -3355
rect 879 -3363 883 -3355
rect 1211 -3363 1215 -3355
rect 1219 -3363 1223 -3355
rect 1228 -3363 1232 -3355
rect 1237 -3363 1241 -3355
rect -1234 -3522 -1230 -3514
rect -1225 -3522 -1221 -3514
rect -1216 -3522 -1212 -3514
rect -1208 -3522 -1204 -3514
rect -1190 -3522 -1186 -3514
rect -1168 -3522 -1164 -3514
rect -1156 -3522 -1152 -3514
rect -1147 -3522 -1143 -3514
rect -1138 -3522 -1134 -3514
rect -935 -3522 -931 -3514
rect -926 -3522 -922 -3514
rect -917 -3522 -913 -3514
rect -909 -3522 -905 -3514
rect -900 -3522 -896 -3514
rect -891 -3522 -887 -3514
rect -883 -3522 -879 -3514
rect -865 -3522 -861 -3514
rect -843 -3522 -839 -3514
rect -831 -3522 -827 -3514
rect -822 -3522 -818 -3514
rect -813 -3522 -809 -3514
rect -805 -3522 -801 -3514
rect -787 -3522 -783 -3514
rect -765 -3522 -761 -3514
rect -753 -3522 -749 -3514
rect -741 -3522 -737 -3514
rect -729 -3522 -725 -3514
rect -721 -3522 -717 -3514
rect -704 -3522 -700 -3514
rect -695 -3522 -691 -3514
rect -577 -3522 -573 -3514
rect -568 -3522 -564 -3514
rect -559 -3522 -555 -3514
rect -551 -3522 -547 -3514
rect -542 -3522 -538 -3514
rect -533 -3522 -529 -3514
rect -525 -3522 -521 -3514
rect -507 -3522 -503 -3514
rect -485 -3522 -481 -3514
rect -473 -3522 -469 -3514
rect -464 -3522 -460 -3514
rect -455 -3522 -451 -3514
rect -447 -3522 -443 -3514
rect -429 -3522 -425 -3514
rect -407 -3522 -403 -3514
rect -395 -3522 -391 -3514
rect -383 -3522 -379 -3514
rect -371 -3522 -367 -3514
rect -363 -3522 -359 -3514
rect -346 -3522 -342 -3514
rect -337 -3522 -333 -3514
rect -219 -3522 -215 -3514
rect -210 -3522 -206 -3514
rect -201 -3522 -197 -3514
rect -193 -3522 -189 -3514
rect -184 -3522 -180 -3514
rect -175 -3522 -171 -3514
rect -167 -3522 -163 -3514
rect -149 -3522 -145 -3514
rect -127 -3522 -123 -3514
rect -115 -3522 -111 -3514
rect -106 -3522 -102 -3514
rect -97 -3522 -93 -3514
rect -89 -3522 -85 -3514
rect -71 -3522 -67 -3514
rect -49 -3522 -45 -3514
rect -37 -3522 -33 -3514
rect -25 -3522 -21 -3514
rect -13 -3522 -9 -3514
rect -5 -3522 -1 -3514
rect 12 -3522 16 -3514
rect 21 -3522 25 -3514
rect 139 -3522 143 -3514
rect 148 -3522 152 -3514
rect 157 -3522 161 -3514
rect 165 -3522 169 -3514
rect 174 -3522 178 -3514
rect 183 -3522 187 -3514
rect 191 -3522 195 -3514
rect 209 -3522 213 -3514
rect 231 -3522 235 -3514
rect 243 -3522 247 -3514
rect 252 -3522 256 -3514
rect 261 -3522 265 -3514
rect 269 -3522 273 -3514
rect 287 -3522 291 -3514
rect 309 -3522 313 -3514
rect 321 -3522 325 -3514
rect 333 -3522 337 -3514
rect 345 -3522 349 -3514
rect 353 -3522 357 -3514
rect 370 -3522 374 -3514
rect 379 -3522 383 -3514
rect 495 -3522 499 -3514
rect 504 -3522 508 -3514
rect 513 -3522 517 -3514
rect 521 -3522 525 -3514
rect 530 -3522 534 -3514
rect 539 -3522 543 -3514
rect 547 -3522 551 -3514
rect 565 -3522 569 -3514
rect 587 -3522 591 -3514
rect 599 -3522 603 -3514
rect 608 -3522 612 -3514
rect 617 -3522 621 -3514
rect 625 -3522 629 -3514
rect 643 -3522 647 -3514
rect 665 -3522 669 -3514
rect 677 -3522 681 -3514
rect 689 -3522 693 -3514
rect 701 -3522 705 -3514
rect 709 -3522 713 -3514
rect 726 -3522 730 -3514
rect 735 -3522 739 -3514
rect 853 -3522 857 -3514
rect 862 -3522 866 -3514
rect 871 -3522 875 -3514
rect 879 -3522 883 -3514
rect 888 -3522 892 -3514
rect 897 -3522 901 -3514
rect 905 -3522 909 -3514
rect 923 -3522 927 -3514
rect 945 -3522 949 -3514
rect 957 -3522 961 -3514
rect 966 -3522 970 -3514
rect 975 -3522 979 -3514
rect 983 -3522 987 -3514
rect 1001 -3522 1005 -3514
rect 1023 -3522 1027 -3514
rect 1035 -3522 1039 -3514
rect 1047 -3522 1051 -3514
rect 1059 -3522 1063 -3514
rect 1067 -3522 1071 -3514
rect 1084 -3522 1088 -3514
rect 1093 -3522 1097 -3514
rect 1211 -3522 1215 -3514
rect 1220 -3522 1224 -3514
rect 1229 -3522 1233 -3514
rect 1237 -3522 1241 -3514
rect 1246 -3522 1250 -3514
rect 1255 -3522 1259 -3514
rect 1263 -3522 1267 -3514
rect 1281 -3522 1285 -3514
rect 1303 -3522 1307 -3514
rect 1315 -3522 1319 -3514
rect 1324 -3522 1328 -3514
rect 1333 -3522 1337 -3514
rect 1341 -3522 1345 -3514
rect 1359 -3522 1363 -3514
rect 1381 -3522 1385 -3514
rect 1393 -3522 1397 -3514
rect 1405 -3522 1409 -3514
rect 1417 -3522 1421 -3514
rect 1425 -3522 1429 -3514
rect 1442 -3522 1446 -3514
rect 1451 -3522 1455 -3514
rect -1822 -3652 -1818 -3644
rect -1813 -3652 -1809 -3644
rect -1804 -3652 -1800 -3644
rect -1796 -3652 -1792 -3644
rect -1788 -3652 -1784 -3644
rect -1776 -3652 -1772 -3644
rect -1764 -3652 -1760 -3644
rect -1755 -3652 -1751 -3644
rect -1746 -3652 -1742 -3644
rect -1734 -3652 -1730 -3644
rect -1722 -3652 -1718 -3644
rect -1713 -3652 -1709 -3644
rect -1704 -3652 -1700 -3644
rect -1692 -3652 -1688 -3644
rect -1680 -3652 -1676 -3644
rect -1671 -3652 -1667 -3644
rect -1662 -3652 -1658 -3644
rect -1650 -3652 -1646 -3644
rect -1638 -3652 -1634 -3644
rect -1630 -3652 -1626 -3644
rect -1559 -3652 -1555 -3644
rect -1550 -3652 -1546 -3644
rect -1541 -3652 -1537 -3644
rect -1533 -3652 -1529 -3644
rect -1525 -3652 -1521 -3644
rect -1513 -3652 -1509 -3644
rect -1501 -3652 -1497 -3644
rect -1492 -3652 -1488 -3644
rect -1483 -3652 -1479 -3644
rect -1471 -3652 -1467 -3644
rect -1459 -3652 -1455 -3644
rect -1450 -3652 -1446 -3644
rect -1441 -3652 -1437 -3644
rect -1429 -3652 -1425 -3644
rect -1417 -3652 -1413 -3644
rect -1408 -3652 -1404 -3644
rect -1399 -3652 -1395 -3644
rect -1387 -3652 -1383 -3644
rect -1375 -3652 -1371 -3644
rect -1367 -3652 -1363 -3644
rect -1234 -3652 -1230 -3644
rect -1225 -3652 -1221 -3644
rect -1216 -3652 -1212 -3644
rect -1208 -3652 -1204 -3644
rect -1200 -3652 -1196 -3644
rect -1188 -3652 -1184 -3644
rect -1176 -3652 -1172 -3644
rect -1167 -3652 -1163 -3644
rect -1158 -3652 -1154 -3644
rect -1146 -3652 -1142 -3644
rect -1134 -3652 -1130 -3644
rect -1125 -3652 -1121 -3644
rect -1116 -3652 -1112 -3644
rect -1104 -3652 -1100 -3644
rect -1092 -3652 -1088 -3644
rect -1083 -3652 -1079 -3644
rect -1074 -3652 -1070 -3644
rect -1062 -3652 -1058 -3644
rect -1050 -3652 -1046 -3644
rect -1042 -3652 -1038 -3644
rect -934 -3652 -930 -3644
rect -925 -3652 -921 -3644
rect -916 -3652 -912 -3644
rect -908 -3652 -904 -3644
rect -900 -3652 -896 -3644
rect -888 -3652 -884 -3644
rect -876 -3652 -872 -3644
rect -867 -3652 -863 -3644
rect -858 -3652 -854 -3644
rect -846 -3652 -842 -3644
rect -834 -3652 -830 -3644
rect -825 -3652 -821 -3644
rect -816 -3652 -812 -3644
rect -804 -3652 -800 -3644
rect -792 -3652 -788 -3644
rect -783 -3652 -779 -3644
rect -774 -3652 -770 -3644
rect -762 -3652 -758 -3644
rect -750 -3652 -746 -3644
rect -742 -3652 -738 -3644
rect -577 -3652 -573 -3644
rect -568 -3652 -564 -3644
rect -559 -3652 -555 -3644
rect -551 -3652 -547 -3644
rect -543 -3652 -539 -3644
rect -531 -3652 -527 -3644
rect -519 -3652 -515 -3644
rect -510 -3652 -506 -3644
rect -501 -3652 -497 -3644
rect -489 -3652 -485 -3644
rect -477 -3652 -473 -3644
rect -468 -3652 -464 -3644
rect -459 -3652 -455 -3644
rect -447 -3652 -443 -3644
rect -435 -3652 -431 -3644
rect -426 -3652 -422 -3644
rect -417 -3652 -413 -3644
rect -405 -3652 -401 -3644
rect -393 -3652 -389 -3644
rect -385 -3652 -381 -3644
rect -219 -3652 -215 -3644
rect -210 -3652 -206 -3644
rect -201 -3652 -197 -3644
rect -193 -3652 -189 -3644
rect -185 -3652 -181 -3644
rect -173 -3652 -169 -3644
rect -161 -3652 -157 -3644
rect -152 -3652 -148 -3644
rect -143 -3652 -139 -3644
rect -131 -3652 -127 -3644
rect -119 -3652 -115 -3644
rect -110 -3652 -106 -3644
rect -101 -3652 -97 -3644
rect -89 -3652 -85 -3644
rect -77 -3652 -73 -3644
rect -68 -3652 -64 -3644
rect -59 -3652 -55 -3644
rect -47 -3652 -43 -3644
rect -35 -3652 -31 -3644
rect -27 -3652 -23 -3644
rect -1559 -3823 -1555 -3815
rect -1550 -3823 -1546 -3815
rect -1541 -3823 -1537 -3815
rect -1533 -3823 -1529 -3815
rect -1525 -3823 -1521 -3815
rect -1513 -3823 -1509 -3815
rect -1501 -3823 -1497 -3815
rect -1492 -3823 -1488 -3815
rect -1483 -3823 -1479 -3815
rect -1471 -3823 -1467 -3815
rect -1459 -3823 -1455 -3815
rect -1450 -3823 -1446 -3815
rect -1441 -3823 -1437 -3815
rect -1429 -3823 -1425 -3815
rect -1417 -3823 -1413 -3815
rect -1408 -3823 -1404 -3815
rect -1399 -3823 -1395 -3815
rect -1387 -3823 -1383 -3815
rect -1375 -3823 -1371 -3815
rect -1367 -3823 -1363 -3815
rect -1234 -3823 -1230 -3815
rect -1225 -3823 -1221 -3815
rect -1216 -3823 -1212 -3815
rect -1208 -3823 -1204 -3815
rect -1200 -3823 -1196 -3815
rect -1188 -3823 -1184 -3815
rect -1176 -3823 -1172 -3815
rect -1167 -3823 -1163 -3815
rect -1158 -3823 -1154 -3815
rect -1146 -3823 -1142 -3815
rect -1134 -3823 -1130 -3815
rect -1125 -3823 -1121 -3815
rect -1116 -3823 -1112 -3815
rect -1104 -3823 -1100 -3815
rect -1092 -3823 -1088 -3815
rect -1083 -3823 -1079 -3815
rect -1074 -3823 -1070 -3815
rect -1062 -3823 -1058 -3815
rect -1050 -3823 -1046 -3815
rect -1042 -3823 -1038 -3815
rect -934 -3823 -930 -3815
rect -925 -3823 -921 -3815
rect -916 -3823 -912 -3815
rect -908 -3823 -904 -3815
rect -900 -3823 -896 -3815
rect -888 -3823 -884 -3815
rect -876 -3823 -872 -3815
rect -867 -3823 -863 -3815
rect -858 -3823 -854 -3815
rect -846 -3823 -842 -3815
rect -834 -3823 -830 -3815
rect -825 -3823 -821 -3815
rect -816 -3823 -812 -3815
rect -804 -3823 -800 -3815
rect -792 -3823 -788 -3815
rect -783 -3823 -779 -3815
rect -774 -3823 -770 -3815
rect -762 -3823 -758 -3815
rect -750 -3823 -746 -3815
rect -742 -3823 -738 -3815
rect -577 -3823 -573 -3815
rect -568 -3823 -564 -3815
rect -559 -3823 -555 -3815
rect -551 -3823 -547 -3815
rect -543 -3823 -539 -3815
rect -531 -3823 -527 -3815
rect -519 -3823 -515 -3815
rect -510 -3823 -506 -3815
rect -501 -3823 -497 -3815
rect -489 -3823 -485 -3815
rect -477 -3823 -473 -3815
rect -468 -3823 -464 -3815
rect -459 -3823 -455 -3815
rect -447 -3823 -443 -3815
rect -435 -3823 -431 -3815
rect -426 -3823 -422 -3815
rect -417 -3823 -413 -3815
rect -405 -3823 -401 -3815
rect -393 -3823 -389 -3815
rect -385 -3823 -381 -3815
rect -219 -3823 -215 -3815
rect -210 -3823 -206 -3815
rect -201 -3823 -197 -3815
rect -193 -3823 -189 -3815
rect -185 -3823 -181 -3815
rect -173 -3823 -169 -3815
rect -161 -3823 -157 -3815
rect -152 -3823 -148 -3815
rect -143 -3823 -139 -3815
rect -131 -3823 -127 -3815
rect -119 -3823 -115 -3815
rect -110 -3823 -106 -3815
rect -101 -3823 -97 -3815
rect -89 -3823 -85 -3815
rect -77 -3823 -73 -3815
rect -68 -3823 -64 -3815
rect -59 -3823 -55 -3815
rect -47 -3823 -43 -3815
rect -35 -3823 -31 -3815
rect -27 -3823 -23 -3815
rect 139 -3823 143 -3815
rect 148 -3823 152 -3815
rect 157 -3823 161 -3815
rect 165 -3823 169 -3815
rect 173 -3823 177 -3815
rect 185 -3823 189 -3815
rect 197 -3823 201 -3815
rect 206 -3823 210 -3815
rect 215 -3823 219 -3815
rect 227 -3823 231 -3815
rect 239 -3823 243 -3815
rect 248 -3823 252 -3815
rect 257 -3823 261 -3815
rect 269 -3823 273 -3815
rect 281 -3823 285 -3815
rect 290 -3823 294 -3815
rect 299 -3823 303 -3815
rect 311 -3823 315 -3815
rect 323 -3823 327 -3815
rect 331 -3823 335 -3815
rect 495 -3823 499 -3815
rect 504 -3823 508 -3815
rect 513 -3823 517 -3815
rect 521 -3823 525 -3815
rect 529 -3823 533 -3815
rect 541 -3823 545 -3815
rect 553 -3823 557 -3815
rect 562 -3823 566 -3815
rect 571 -3823 575 -3815
rect 583 -3823 587 -3815
rect 595 -3823 599 -3815
rect 604 -3823 608 -3815
rect 613 -3823 617 -3815
rect 625 -3823 629 -3815
rect 637 -3823 641 -3815
rect 646 -3823 650 -3815
rect 655 -3823 659 -3815
rect 667 -3823 671 -3815
rect 679 -3823 683 -3815
rect 687 -3823 691 -3815
rect 853 -3823 857 -3815
rect 862 -3823 866 -3815
rect 871 -3823 875 -3815
rect 879 -3823 883 -3815
rect 887 -3823 891 -3815
rect 899 -3823 903 -3815
rect 911 -3823 915 -3815
rect 920 -3823 924 -3815
rect 929 -3823 933 -3815
rect 941 -3823 945 -3815
rect 953 -3823 957 -3815
rect 962 -3823 966 -3815
rect 971 -3823 975 -3815
rect 983 -3823 987 -3815
rect 995 -3823 999 -3815
rect 1004 -3823 1008 -3815
rect 1013 -3823 1017 -3815
rect 1025 -3823 1029 -3815
rect 1037 -3823 1041 -3815
rect 1045 -3823 1049 -3815
rect 1211 -3823 1215 -3815
rect 1220 -3823 1224 -3815
rect 1229 -3823 1233 -3815
rect 1237 -3823 1241 -3815
rect 1245 -3823 1249 -3815
rect 1257 -3823 1261 -3815
rect 1269 -3823 1273 -3815
rect 1278 -3823 1282 -3815
rect 1287 -3823 1291 -3815
rect 1299 -3823 1303 -3815
rect 1311 -3823 1315 -3815
rect 1320 -3823 1324 -3815
rect 1329 -3823 1333 -3815
rect 1341 -3823 1345 -3815
rect 1353 -3823 1357 -3815
rect 1362 -3823 1366 -3815
rect 1371 -3823 1375 -3815
rect 1383 -3823 1387 -3815
rect 1395 -3823 1399 -3815
rect 1403 -3823 1407 -3815
rect -1559 -3998 -1555 -3990
rect -1550 -3998 -1546 -3990
rect -1541 -3998 -1537 -3990
rect -1533 -3998 -1529 -3990
rect -1525 -3998 -1521 -3990
rect -1513 -3998 -1509 -3990
rect -1501 -3998 -1497 -3990
rect -1492 -3998 -1488 -3990
rect -1483 -3998 -1479 -3990
rect -1471 -3998 -1467 -3990
rect -1459 -3998 -1455 -3990
rect -1450 -3998 -1446 -3990
rect -1441 -3998 -1437 -3990
rect -1429 -3998 -1425 -3990
rect -1417 -3998 -1413 -3990
rect -1408 -3998 -1404 -3990
rect -1399 -3998 -1395 -3990
rect -1387 -3998 -1383 -3990
rect -1375 -3998 -1371 -3990
rect -1367 -3998 -1363 -3990
rect -1234 -3998 -1230 -3990
rect -1225 -3998 -1221 -3990
rect -1216 -3998 -1212 -3990
rect -1208 -3998 -1204 -3990
rect -1200 -3998 -1196 -3990
rect -1188 -3998 -1184 -3990
rect -1176 -3998 -1172 -3990
rect -1167 -3998 -1163 -3990
rect -1158 -3998 -1154 -3990
rect -1146 -3998 -1142 -3990
rect -1134 -3998 -1130 -3990
rect -1125 -3998 -1121 -3990
rect -1116 -3998 -1112 -3990
rect -1104 -3998 -1100 -3990
rect -1092 -3998 -1088 -3990
rect -1083 -3998 -1079 -3990
rect -1074 -3998 -1070 -3990
rect -1062 -3998 -1058 -3990
rect -1050 -3998 -1046 -3990
rect -1042 -3998 -1038 -3990
rect -935 -3998 -931 -3990
rect -926 -3998 -922 -3990
rect -917 -3998 -913 -3990
rect -909 -3998 -905 -3990
rect -901 -3998 -897 -3990
rect -889 -3998 -885 -3990
rect -877 -3998 -873 -3990
rect -868 -3998 -864 -3990
rect -859 -3998 -855 -3990
rect -847 -3998 -843 -3990
rect -835 -3998 -831 -3990
rect -826 -3998 -822 -3990
rect -817 -3998 -813 -3990
rect -805 -3998 -801 -3990
rect -793 -3998 -789 -3990
rect -784 -3998 -780 -3990
rect -775 -3998 -771 -3990
rect -763 -3998 -759 -3990
rect -751 -3998 -747 -3990
rect -743 -3998 -739 -3990
rect -577 -3998 -573 -3990
rect -568 -3998 -564 -3990
rect -559 -3998 -555 -3990
rect -551 -3998 -547 -3990
rect -543 -3998 -539 -3990
rect -531 -3998 -527 -3990
rect -519 -3998 -515 -3990
rect -510 -3998 -506 -3990
rect -501 -3998 -497 -3990
rect -489 -3998 -485 -3990
rect -477 -3998 -473 -3990
rect -468 -3998 -464 -3990
rect -459 -3998 -455 -3990
rect -447 -3998 -443 -3990
rect -435 -3998 -431 -3990
rect -426 -3998 -422 -3990
rect -417 -3998 -413 -3990
rect -405 -3998 -401 -3990
rect -393 -3998 -389 -3990
rect -385 -3998 -381 -3990
rect -219 -3998 -215 -3990
rect -210 -3998 -206 -3990
rect -201 -3998 -197 -3990
rect -193 -3998 -189 -3990
rect -185 -3998 -181 -3990
rect -173 -3998 -169 -3990
rect -161 -3998 -157 -3990
rect -152 -3998 -148 -3990
rect -143 -3998 -139 -3990
rect -131 -3998 -127 -3990
rect -119 -3998 -115 -3990
rect -110 -3998 -106 -3990
rect -101 -3998 -97 -3990
rect -89 -3998 -85 -3990
rect -77 -3998 -73 -3990
rect -68 -3998 -64 -3990
rect -59 -3998 -55 -3990
rect -47 -3998 -43 -3990
rect -35 -3998 -31 -3990
rect -27 -3998 -23 -3990
rect 139 -3998 143 -3990
rect 148 -3998 152 -3990
rect 157 -3998 161 -3990
rect 165 -3998 169 -3990
rect 173 -3998 177 -3990
rect 185 -3998 189 -3990
rect 197 -3998 201 -3990
rect 206 -3998 210 -3990
rect 215 -3998 219 -3990
rect 227 -3998 231 -3990
rect 239 -3998 243 -3990
rect 248 -3998 252 -3990
rect 257 -3998 261 -3990
rect 269 -3998 273 -3990
rect 281 -3998 285 -3990
rect 290 -3998 294 -3990
rect 299 -3998 303 -3990
rect 311 -3998 315 -3990
rect 323 -3998 327 -3990
rect 331 -3998 335 -3990
rect 495 -3998 499 -3990
rect 504 -3998 508 -3990
rect 513 -3998 517 -3990
rect 521 -3998 525 -3990
rect 529 -3998 533 -3990
rect 541 -3998 545 -3990
rect 553 -3998 557 -3990
rect 562 -3998 566 -3990
rect 571 -3998 575 -3990
rect 583 -3998 587 -3990
rect 595 -3998 599 -3990
rect 604 -3998 608 -3990
rect 613 -3998 617 -3990
rect 625 -3998 629 -3990
rect 637 -3998 641 -3990
rect 646 -3998 650 -3990
rect 655 -3998 659 -3990
rect 667 -3998 671 -3990
rect 679 -3998 683 -3990
rect 687 -3998 691 -3990
rect 853 -3998 857 -3990
rect 862 -3998 866 -3990
rect 871 -3998 875 -3990
rect 879 -3998 883 -3990
rect 887 -3998 891 -3990
rect 899 -3998 903 -3990
rect 911 -3998 915 -3990
rect 920 -3998 924 -3990
rect 929 -3998 933 -3990
rect 941 -3998 945 -3990
rect 953 -3998 957 -3990
rect 962 -3998 966 -3990
rect 971 -3998 975 -3990
rect 983 -3998 987 -3990
rect 995 -3998 999 -3990
rect 1004 -3998 1008 -3990
rect 1013 -3998 1017 -3990
rect 1025 -3998 1029 -3990
rect 1037 -3998 1041 -3990
rect 1045 -3998 1049 -3990
rect 1211 -3998 1215 -3990
rect 1220 -3998 1224 -3990
rect 1229 -3998 1233 -3990
rect 1237 -3998 1241 -3990
rect 1245 -3998 1249 -3990
rect 1257 -3998 1261 -3990
rect 1269 -3998 1273 -3990
rect 1278 -3998 1282 -3990
rect 1287 -3998 1291 -3990
rect 1299 -3998 1303 -3990
rect 1311 -3998 1315 -3990
rect 1320 -3998 1324 -3990
rect 1329 -3998 1333 -3990
rect 1341 -3998 1345 -3990
rect 1353 -3998 1357 -3990
rect 1362 -3998 1366 -3990
rect 1371 -3998 1375 -3990
rect 1383 -3998 1387 -3990
rect 1395 -3998 1399 -3990
rect 1403 -3998 1407 -3990
rect -1309 -4113 -1305 -4105
rect -1301 -4113 -1297 -4105
rect -1292 -4113 -1288 -4105
rect -1283 -4113 -1279 -4105
rect -935 -4113 -931 -4105
rect -927 -4113 -923 -4105
rect -918 -4113 -914 -4105
rect -909 -4113 -905 -4105
rect -577 -4113 -573 -4105
rect -569 -4113 -565 -4105
rect -560 -4113 -556 -4105
rect -551 -4113 -547 -4105
rect -219 -4113 -215 -4105
rect -211 -4113 -207 -4105
rect -202 -4113 -198 -4105
rect -193 -4113 -189 -4105
rect 139 -4113 143 -4105
rect 147 -4113 151 -4105
rect 156 -4113 160 -4105
rect 165 -4113 169 -4105
rect 495 -4113 499 -4105
rect 503 -4113 507 -4105
rect 512 -4113 516 -4105
rect 521 -4113 525 -4105
rect 853 -4113 857 -4105
rect 861 -4113 865 -4105
rect 870 -4113 874 -4105
rect 879 -4113 883 -4105
rect 1211 -4113 1215 -4105
rect 1219 -4113 1223 -4105
rect 1228 -4113 1232 -4105
rect 1237 -4113 1241 -4105
rect -1234 -4272 -1230 -4264
rect -1225 -4272 -1221 -4264
rect -1216 -4272 -1212 -4264
rect -1208 -4272 -1204 -4264
rect -1190 -4272 -1186 -4264
rect -1168 -4272 -1164 -4264
rect -1156 -4272 -1152 -4264
rect -1147 -4272 -1143 -4264
rect -1138 -4272 -1134 -4264
rect -935 -4272 -931 -4264
rect -926 -4272 -922 -4264
rect -917 -4272 -913 -4264
rect -909 -4272 -905 -4264
rect -900 -4272 -896 -4264
rect -891 -4272 -887 -4264
rect -883 -4272 -879 -4264
rect -865 -4272 -861 -4264
rect -843 -4272 -839 -4264
rect -831 -4272 -827 -4264
rect -822 -4272 -818 -4264
rect -813 -4272 -809 -4264
rect -805 -4272 -801 -4264
rect -787 -4272 -783 -4264
rect -765 -4272 -761 -4264
rect -753 -4272 -749 -4264
rect -741 -4272 -737 -4264
rect -729 -4272 -725 -4264
rect -721 -4272 -717 -4264
rect -704 -4272 -700 -4264
rect -695 -4272 -691 -4264
rect -577 -4272 -573 -4264
rect -568 -4272 -564 -4264
rect -559 -4272 -555 -4264
rect -551 -4272 -547 -4264
rect -542 -4272 -538 -4264
rect -533 -4272 -529 -4264
rect -525 -4272 -521 -4264
rect -507 -4272 -503 -4264
rect -485 -4272 -481 -4264
rect -473 -4272 -469 -4264
rect -464 -4272 -460 -4264
rect -455 -4272 -451 -4264
rect -447 -4272 -443 -4264
rect -429 -4272 -425 -4264
rect -407 -4272 -403 -4264
rect -395 -4272 -391 -4264
rect -383 -4272 -379 -4264
rect -371 -4272 -367 -4264
rect -363 -4272 -359 -4264
rect -346 -4272 -342 -4264
rect -337 -4272 -333 -4264
rect -219 -4272 -215 -4264
rect -210 -4272 -206 -4264
rect -201 -4272 -197 -4264
rect -193 -4272 -189 -4264
rect -184 -4272 -180 -4264
rect -175 -4272 -171 -4264
rect -167 -4272 -163 -4264
rect -149 -4272 -145 -4264
rect -127 -4272 -123 -4264
rect -115 -4272 -111 -4264
rect -106 -4272 -102 -4264
rect -97 -4272 -93 -4264
rect -89 -4272 -85 -4264
rect -71 -4272 -67 -4264
rect -49 -4272 -45 -4264
rect -37 -4272 -33 -4264
rect -25 -4272 -21 -4264
rect -13 -4272 -9 -4264
rect -5 -4272 -1 -4264
rect 12 -4272 16 -4264
rect 21 -4272 25 -4264
rect 139 -4272 143 -4264
rect 148 -4272 152 -4264
rect 157 -4272 161 -4264
rect 165 -4272 169 -4264
rect 174 -4272 178 -4264
rect 183 -4272 187 -4264
rect 191 -4272 195 -4264
rect 209 -4272 213 -4264
rect 231 -4272 235 -4264
rect 243 -4272 247 -4264
rect 252 -4272 256 -4264
rect 261 -4272 265 -4264
rect 269 -4272 273 -4264
rect 287 -4272 291 -4264
rect 309 -4272 313 -4264
rect 321 -4272 325 -4264
rect 333 -4272 337 -4264
rect 345 -4272 349 -4264
rect 353 -4272 357 -4264
rect 370 -4272 374 -4264
rect 379 -4272 383 -4264
rect 495 -4272 499 -4264
rect 504 -4272 508 -4264
rect 513 -4272 517 -4264
rect 521 -4272 525 -4264
rect 530 -4272 534 -4264
rect 539 -4272 543 -4264
rect 547 -4272 551 -4264
rect 565 -4272 569 -4264
rect 587 -4272 591 -4264
rect 599 -4272 603 -4264
rect 608 -4272 612 -4264
rect 617 -4272 621 -4264
rect 625 -4272 629 -4264
rect 643 -4272 647 -4264
rect 665 -4272 669 -4264
rect 677 -4272 681 -4264
rect 689 -4272 693 -4264
rect 701 -4272 705 -4264
rect 709 -4272 713 -4264
rect 726 -4272 730 -4264
rect 735 -4272 739 -4264
rect 853 -4272 857 -4264
rect 862 -4272 866 -4264
rect 871 -4272 875 -4264
rect 879 -4272 883 -4264
rect 888 -4272 892 -4264
rect 897 -4272 901 -4264
rect 905 -4272 909 -4264
rect 923 -4272 927 -4264
rect 945 -4272 949 -4264
rect 957 -4272 961 -4264
rect 966 -4272 970 -4264
rect 975 -4272 979 -4264
rect 983 -4272 987 -4264
rect 1001 -4272 1005 -4264
rect 1023 -4272 1027 -4264
rect 1035 -4272 1039 -4264
rect 1047 -4272 1051 -4264
rect 1059 -4272 1063 -4264
rect 1067 -4272 1071 -4264
rect 1084 -4272 1088 -4264
rect 1093 -4272 1097 -4264
rect 1211 -4272 1215 -4264
rect 1220 -4272 1224 -4264
rect 1229 -4272 1233 -4264
rect 1237 -4272 1241 -4264
rect 1246 -4272 1250 -4264
rect 1255 -4272 1259 -4264
rect 1263 -4272 1267 -4264
rect 1281 -4272 1285 -4264
rect 1303 -4272 1307 -4264
rect 1315 -4272 1319 -4264
rect 1324 -4272 1328 -4264
rect 1333 -4272 1337 -4264
rect 1341 -4272 1345 -4264
rect 1359 -4272 1363 -4264
rect 1381 -4272 1385 -4264
rect 1393 -4272 1397 -4264
rect 1405 -4272 1409 -4264
rect 1417 -4272 1421 -4264
rect 1425 -4272 1429 -4264
rect 1442 -4272 1446 -4264
rect 1451 -4272 1455 -4264
rect -1814 -4395 -1810 -4387
rect -1805 -4395 -1801 -4387
rect -1796 -4395 -1792 -4387
rect -1788 -4395 -1784 -4387
rect -1780 -4395 -1776 -4387
rect -1768 -4395 -1764 -4387
rect -1756 -4395 -1752 -4387
rect -1747 -4395 -1743 -4387
rect -1738 -4395 -1734 -4387
rect -1726 -4395 -1722 -4387
rect -1714 -4395 -1710 -4387
rect -1705 -4395 -1701 -4387
rect -1696 -4395 -1692 -4387
rect -1684 -4395 -1680 -4387
rect -1672 -4395 -1668 -4387
rect -1663 -4395 -1659 -4387
rect -1654 -4395 -1650 -4387
rect -1642 -4395 -1638 -4387
rect -1630 -4395 -1626 -4387
rect -1622 -4395 -1618 -4387
rect -1551 -4395 -1547 -4387
rect -1542 -4395 -1538 -4387
rect -1533 -4395 -1529 -4387
rect -1525 -4395 -1521 -4387
rect -1517 -4395 -1513 -4387
rect -1505 -4395 -1501 -4387
rect -1493 -4395 -1489 -4387
rect -1484 -4395 -1480 -4387
rect -1475 -4395 -1471 -4387
rect -1463 -4395 -1459 -4387
rect -1451 -4395 -1447 -4387
rect -1442 -4395 -1438 -4387
rect -1433 -4395 -1429 -4387
rect -1421 -4395 -1417 -4387
rect -1409 -4395 -1405 -4387
rect -1400 -4395 -1396 -4387
rect -1391 -4395 -1387 -4387
rect -1379 -4395 -1375 -4387
rect -1367 -4395 -1363 -4387
rect -1359 -4395 -1355 -4387
rect -1234 -4395 -1230 -4387
rect -1225 -4395 -1221 -4387
rect -1216 -4395 -1212 -4387
rect -1208 -4395 -1204 -4387
rect -1200 -4395 -1196 -4387
rect -1188 -4395 -1184 -4387
rect -1176 -4395 -1172 -4387
rect -1167 -4395 -1163 -4387
rect -1158 -4395 -1154 -4387
rect -1146 -4395 -1142 -4387
rect -1134 -4395 -1130 -4387
rect -1125 -4395 -1121 -4387
rect -1116 -4395 -1112 -4387
rect -1104 -4395 -1100 -4387
rect -1092 -4395 -1088 -4387
rect -1083 -4395 -1079 -4387
rect -1074 -4395 -1070 -4387
rect -1062 -4395 -1058 -4387
rect -1050 -4395 -1046 -4387
rect -1042 -4395 -1038 -4387
rect -935 -4395 -931 -4387
rect -926 -4395 -922 -4387
rect -917 -4395 -913 -4387
rect -909 -4395 -905 -4387
rect -901 -4395 -897 -4387
rect -889 -4395 -885 -4387
rect -877 -4395 -873 -4387
rect -868 -4395 -864 -4387
rect -859 -4395 -855 -4387
rect -847 -4395 -843 -4387
rect -835 -4395 -831 -4387
rect -826 -4395 -822 -4387
rect -817 -4395 -813 -4387
rect -805 -4395 -801 -4387
rect -793 -4395 -789 -4387
rect -784 -4395 -780 -4387
rect -775 -4395 -771 -4387
rect -763 -4395 -759 -4387
rect -751 -4395 -747 -4387
rect -743 -4395 -739 -4387
rect -577 -4395 -573 -4387
rect -568 -4395 -564 -4387
rect -559 -4395 -555 -4387
rect -551 -4395 -547 -4387
rect -543 -4395 -539 -4387
rect -531 -4395 -527 -4387
rect -519 -4395 -515 -4387
rect -510 -4395 -506 -4387
rect -501 -4395 -497 -4387
rect -489 -4395 -485 -4387
rect -477 -4395 -473 -4387
rect -468 -4395 -464 -4387
rect -459 -4395 -455 -4387
rect -447 -4395 -443 -4387
rect -435 -4395 -431 -4387
rect -426 -4395 -422 -4387
rect -417 -4395 -413 -4387
rect -405 -4395 -401 -4387
rect -393 -4395 -389 -4387
rect -385 -4395 -381 -4387
rect -1814 -4566 -1810 -4558
rect -1805 -4566 -1801 -4558
rect -1796 -4566 -1792 -4558
rect -1788 -4566 -1784 -4558
rect -1780 -4566 -1776 -4558
rect -1768 -4566 -1764 -4558
rect -1756 -4566 -1752 -4558
rect -1747 -4566 -1743 -4558
rect -1738 -4566 -1734 -4558
rect -1726 -4566 -1722 -4558
rect -1714 -4566 -1710 -4558
rect -1705 -4566 -1701 -4558
rect -1696 -4566 -1692 -4558
rect -1684 -4566 -1680 -4558
rect -1672 -4566 -1668 -4558
rect -1663 -4566 -1659 -4558
rect -1654 -4566 -1650 -4558
rect -1642 -4566 -1638 -4558
rect -1630 -4566 -1626 -4558
rect -1622 -4566 -1618 -4558
rect -1551 -4566 -1547 -4558
rect -1542 -4566 -1538 -4558
rect -1533 -4566 -1529 -4558
rect -1525 -4566 -1521 -4558
rect -1517 -4566 -1513 -4558
rect -1505 -4566 -1501 -4558
rect -1493 -4566 -1489 -4558
rect -1484 -4566 -1480 -4558
rect -1475 -4566 -1471 -4558
rect -1463 -4566 -1459 -4558
rect -1451 -4566 -1447 -4558
rect -1442 -4566 -1438 -4558
rect -1433 -4566 -1429 -4558
rect -1421 -4566 -1417 -4558
rect -1409 -4566 -1405 -4558
rect -1400 -4566 -1396 -4558
rect -1391 -4566 -1387 -4558
rect -1379 -4566 -1375 -4558
rect -1367 -4566 -1363 -4558
rect -1359 -4566 -1355 -4558
rect -1234 -4566 -1230 -4558
rect -1225 -4566 -1221 -4558
rect -1216 -4566 -1212 -4558
rect -1208 -4566 -1204 -4558
rect -1200 -4566 -1196 -4558
rect -1188 -4566 -1184 -4558
rect -1176 -4566 -1172 -4558
rect -1167 -4566 -1163 -4558
rect -1158 -4566 -1154 -4558
rect -1146 -4566 -1142 -4558
rect -1134 -4566 -1130 -4558
rect -1125 -4566 -1121 -4558
rect -1116 -4566 -1112 -4558
rect -1104 -4566 -1100 -4558
rect -1092 -4566 -1088 -4558
rect -1083 -4566 -1079 -4558
rect -1074 -4566 -1070 -4558
rect -1062 -4566 -1058 -4558
rect -1050 -4566 -1046 -4558
rect -1042 -4566 -1038 -4558
rect -935 -4566 -931 -4558
rect -926 -4566 -922 -4558
rect -917 -4566 -913 -4558
rect -909 -4566 -905 -4558
rect -901 -4566 -897 -4558
rect -889 -4566 -885 -4558
rect -877 -4566 -873 -4558
rect -868 -4566 -864 -4558
rect -859 -4566 -855 -4558
rect -847 -4566 -843 -4558
rect -835 -4566 -831 -4558
rect -826 -4566 -822 -4558
rect -817 -4566 -813 -4558
rect -805 -4566 -801 -4558
rect -793 -4566 -789 -4558
rect -784 -4566 -780 -4558
rect -775 -4566 -771 -4558
rect -763 -4566 -759 -4558
rect -751 -4566 -747 -4558
rect -743 -4566 -739 -4558
rect -577 -4566 -573 -4558
rect -568 -4566 -564 -4558
rect -559 -4566 -555 -4558
rect -551 -4566 -547 -4558
rect -543 -4566 -539 -4558
rect -531 -4566 -527 -4558
rect -519 -4566 -515 -4558
rect -510 -4566 -506 -4558
rect -501 -4566 -497 -4558
rect -489 -4566 -485 -4558
rect -477 -4566 -473 -4558
rect -468 -4566 -464 -4558
rect -459 -4566 -455 -4558
rect -447 -4566 -443 -4558
rect -435 -4566 -431 -4558
rect -426 -4566 -422 -4558
rect -417 -4566 -413 -4558
rect -405 -4566 -401 -4558
rect -393 -4566 -389 -4558
rect -385 -4566 -381 -4558
rect -219 -4566 -215 -4558
rect -210 -4566 -206 -4558
rect -201 -4566 -197 -4558
rect -193 -4566 -189 -4558
rect -185 -4566 -181 -4558
rect -173 -4566 -169 -4558
rect -161 -4566 -157 -4558
rect -152 -4566 -148 -4558
rect -143 -4566 -139 -4558
rect -131 -4566 -127 -4558
rect -119 -4566 -115 -4558
rect -110 -4566 -106 -4558
rect -101 -4566 -97 -4558
rect -89 -4566 -85 -4558
rect -77 -4566 -73 -4558
rect -68 -4566 -64 -4558
rect -59 -4566 -55 -4558
rect -47 -4566 -43 -4558
rect -35 -4566 -31 -4558
rect -27 -4566 -23 -4558
rect 139 -4566 143 -4558
rect 148 -4566 152 -4558
rect 157 -4566 161 -4558
rect 165 -4566 169 -4558
rect 173 -4566 177 -4558
rect 185 -4566 189 -4558
rect 197 -4566 201 -4558
rect 206 -4566 210 -4558
rect 215 -4566 219 -4558
rect 227 -4566 231 -4558
rect 239 -4566 243 -4558
rect 248 -4566 252 -4558
rect 257 -4566 261 -4558
rect 269 -4566 273 -4558
rect 281 -4566 285 -4558
rect 290 -4566 294 -4558
rect 299 -4566 303 -4558
rect 311 -4566 315 -4558
rect 323 -4566 327 -4558
rect 331 -4566 335 -4558
rect 495 -4566 499 -4558
rect 504 -4566 508 -4558
rect 513 -4566 517 -4558
rect 521 -4566 525 -4558
rect 529 -4566 533 -4558
rect 541 -4566 545 -4558
rect 553 -4566 557 -4558
rect 562 -4566 566 -4558
rect 571 -4566 575 -4558
rect 583 -4566 587 -4558
rect 595 -4566 599 -4558
rect 604 -4566 608 -4558
rect 613 -4566 617 -4558
rect 625 -4566 629 -4558
rect 637 -4566 641 -4558
rect 646 -4566 650 -4558
rect 655 -4566 659 -4558
rect 667 -4566 671 -4558
rect 679 -4566 683 -4558
rect 687 -4566 691 -4558
rect 853 -4566 857 -4558
rect 862 -4566 866 -4558
rect 871 -4566 875 -4558
rect 879 -4566 883 -4558
rect 887 -4566 891 -4558
rect 899 -4566 903 -4558
rect 911 -4566 915 -4558
rect 920 -4566 924 -4558
rect 929 -4566 933 -4558
rect 941 -4566 945 -4558
rect 953 -4566 957 -4558
rect 962 -4566 966 -4558
rect 971 -4566 975 -4558
rect 983 -4566 987 -4558
rect 995 -4566 999 -4558
rect 1004 -4566 1008 -4558
rect 1013 -4566 1017 -4558
rect 1025 -4566 1029 -4558
rect 1037 -4566 1041 -4558
rect 1045 -4566 1049 -4558
rect 1211 -4566 1215 -4558
rect 1220 -4566 1224 -4558
rect 1229 -4566 1233 -4558
rect 1237 -4566 1241 -4558
rect 1245 -4566 1249 -4558
rect 1257 -4566 1261 -4558
rect 1269 -4566 1273 -4558
rect 1278 -4566 1282 -4558
rect 1287 -4566 1291 -4558
rect 1299 -4566 1303 -4558
rect 1311 -4566 1315 -4558
rect 1320 -4566 1324 -4558
rect 1329 -4566 1333 -4558
rect 1341 -4566 1345 -4558
rect 1353 -4566 1357 -4558
rect 1362 -4566 1366 -4558
rect 1371 -4566 1375 -4558
rect 1383 -4566 1387 -4558
rect 1395 -4566 1399 -4558
rect 1403 -4566 1407 -4558
rect -1551 -4737 -1547 -4729
rect -1542 -4737 -1538 -4729
rect -1533 -4737 -1529 -4729
rect -1525 -4737 -1521 -4729
rect -1517 -4737 -1513 -4729
rect -1505 -4737 -1501 -4729
rect -1493 -4737 -1489 -4729
rect -1484 -4737 -1480 -4729
rect -1475 -4737 -1471 -4729
rect -1463 -4737 -1459 -4729
rect -1451 -4737 -1447 -4729
rect -1442 -4737 -1438 -4729
rect -1433 -4737 -1429 -4729
rect -1421 -4737 -1417 -4729
rect -1409 -4737 -1405 -4729
rect -1400 -4737 -1396 -4729
rect -1391 -4737 -1387 -4729
rect -1379 -4737 -1375 -4729
rect -1367 -4737 -1363 -4729
rect -1359 -4737 -1355 -4729
rect -1234 -4737 -1230 -4729
rect -1225 -4737 -1221 -4729
rect -1216 -4737 -1212 -4729
rect -1208 -4737 -1204 -4729
rect -1200 -4737 -1196 -4729
rect -1188 -4737 -1184 -4729
rect -1176 -4737 -1172 -4729
rect -1167 -4737 -1163 -4729
rect -1158 -4737 -1154 -4729
rect -1146 -4737 -1142 -4729
rect -1134 -4737 -1130 -4729
rect -1125 -4737 -1121 -4729
rect -1116 -4737 -1112 -4729
rect -1104 -4737 -1100 -4729
rect -1092 -4737 -1088 -4729
rect -1083 -4737 -1079 -4729
rect -1074 -4737 -1070 -4729
rect -1062 -4737 -1058 -4729
rect -1050 -4737 -1046 -4729
rect -1042 -4737 -1038 -4729
rect -935 -4737 -931 -4729
rect -926 -4737 -922 -4729
rect -917 -4737 -913 -4729
rect -909 -4737 -905 -4729
rect -901 -4737 -897 -4729
rect -889 -4737 -885 -4729
rect -877 -4737 -873 -4729
rect -868 -4737 -864 -4729
rect -859 -4737 -855 -4729
rect -847 -4737 -843 -4729
rect -835 -4737 -831 -4729
rect -826 -4737 -822 -4729
rect -817 -4737 -813 -4729
rect -805 -4737 -801 -4729
rect -793 -4737 -789 -4729
rect -784 -4737 -780 -4729
rect -775 -4737 -771 -4729
rect -763 -4737 -759 -4729
rect -751 -4737 -747 -4729
rect -743 -4737 -739 -4729
rect -577 -4737 -573 -4729
rect -568 -4737 -564 -4729
rect -559 -4737 -555 -4729
rect -551 -4737 -547 -4729
rect -543 -4737 -539 -4729
rect -531 -4737 -527 -4729
rect -519 -4737 -515 -4729
rect -510 -4737 -506 -4729
rect -501 -4737 -497 -4729
rect -489 -4737 -485 -4729
rect -477 -4737 -473 -4729
rect -468 -4737 -464 -4729
rect -459 -4737 -455 -4729
rect -447 -4737 -443 -4729
rect -435 -4737 -431 -4729
rect -426 -4737 -422 -4729
rect -417 -4737 -413 -4729
rect -405 -4737 -401 -4729
rect -393 -4737 -389 -4729
rect -385 -4737 -381 -4729
rect -219 -4737 -215 -4729
rect -210 -4737 -206 -4729
rect -201 -4737 -197 -4729
rect -193 -4737 -189 -4729
rect -185 -4737 -181 -4729
rect -173 -4737 -169 -4729
rect -161 -4737 -157 -4729
rect -152 -4737 -148 -4729
rect -143 -4737 -139 -4729
rect -131 -4737 -127 -4729
rect -119 -4737 -115 -4729
rect -110 -4737 -106 -4729
rect -101 -4737 -97 -4729
rect -89 -4737 -85 -4729
rect -77 -4737 -73 -4729
rect -68 -4737 -64 -4729
rect -59 -4737 -55 -4729
rect -47 -4737 -43 -4729
rect -35 -4737 -31 -4729
rect -27 -4737 -23 -4729
rect 139 -4737 143 -4729
rect 148 -4737 152 -4729
rect 157 -4737 161 -4729
rect 165 -4737 169 -4729
rect 173 -4737 177 -4729
rect 185 -4737 189 -4729
rect 197 -4737 201 -4729
rect 206 -4737 210 -4729
rect 215 -4737 219 -4729
rect 227 -4737 231 -4729
rect 239 -4737 243 -4729
rect 248 -4737 252 -4729
rect 257 -4737 261 -4729
rect 269 -4737 273 -4729
rect 281 -4737 285 -4729
rect 290 -4737 294 -4729
rect 299 -4737 303 -4729
rect 311 -4737 315 -4729
rect 323 -4737 327 -4729
rect 331 -4737 335 -4729
rect 495 -4737 499 -4729
rect 504 -4737 508 -4729
rect 513 -4737 517 -4729
rect 521 -4737 525 -4729
rect 529 -4737 533 -4729
rect 541 -4737 545 -4729
rect 553 -4737 557 -4729
rect 562 -4737 566 -4729
rect 571 -4737 575 -4729
rect 583 -4737 587 -4729
rect 595 -4737 599 -4729
rect 604 -4737 608 -4729
rect 613 -4737 617 -4729
rect 625 -4737 629 -4729
rect 637 -4737 641 -4729
rect 646 -4737 650 -4729
rect 655 -4737 659 -4729
rect 667 -4737 671 -4729
rect 679 -4737 683 -4729
rect 687 -4737 691 -4729
rect 853 -4737 857 -4729
rect 862 -4737 866 -4729
rect 871 -4737 875 -4729
rect 879 -4737 883 -4729
rect 887 -4737 891 -4729
rect 899 -4737 903 -4729
rect 911 -4737 915 -4729
rect 920 -4737 924 -4729
rect 929 -4737 933 -4729
rect 941 -4737 945 -4729
rect 953 -4737 957 -4729
rect 962 -4737 966 -4729
rect 971 -4737 975 -4729
rect 983 -4737 987 -4729
rect 995 -4737 999 -4729
rect 1004 -4737 1008 -4729
rect 1013 -4737 1017 -4729
rect 1025 -4737 1029 -4729
rect 1037 -4737 1041 -4729
rect 1045 -4737 1049 -4729
rect 1211 -4737 1215 -4729
rect 1220 -4737 1224 -4729
rect 1229 -4737 1233 -4729
rect 1237 -4737 1241 -4729
rect 1245 -4737 1249 -4729
rect 1257 -4737 1261 -4729
rect 1269 -4737 1273 -4729
rect 1278 -4737 1282 -4729
rect 1287 -4737 1291 -4729
rect 1299 -4737 1303 -4729
rect 1311 -4737 1315 -4729
rect 1320 -4737 1324 -4729
rect 1329 -4737 1333 -4729
rect 1341 -4737 1345 -4729
rect 1353 -4737 1357 -4729
rect 1362 -4737 1366 -4729
rect 1371 -4737 1375 -4729
rect 1383 -4737 1387 -4729
rect 1395 -4737 1399 -4729
rect 1403 -4737 1407 -4729
rect -1309 -4852 -1305 -4844
rect -1301 -4852 -1297 -4844
rect -1292 -4852 -1288 -4844
rect -1283 -4852 -1279 -4844
rect -935 -4852 -931 -4844
rect -927 -4852 -923 -4844
rect -918 -4852 -914 -4844
rect -909 -4852 -905 -4844
rect -577 -4852 -573 -4844
rect -569 -4852 -565 -4844
rect -560 -4852 -556 -4844
rect -551 -4852 -547 -4844
rect -219 -4852 -215 -4844
rect -211 -4852 -207 -4844
rect -202 -4852 -198 -4844
rect -193 -4852 -189 -4844
rect 139 -4852 143 -4844
rect 147 -4852 151 -4844
rect 156 -4852 160 -4844
rect 165 -4852 169 -4844
rect 495 -4852 499 -4844
rect 503 -4852 507 -4844
rect 512 -4852 516 -4844
rect 521 -4852 525 -4844
rect 853 -4852 857 -4844
rect 861 -4852 865 -4844
rect 870 -4852 874 -4844
rect 879 -4852 883 -4844
rect 1211 -4852 1215 -4844
rect 1219 -4852 1223 -4844
rect 1228 -4852 1232 -4844
rect 1237 -4852 1241 -4844
rect -1234 -5011 -1230 -5003
rect -1225 -5011 -1221 -5003
rect -1216 -5011 -1212 -5003
rect -1208 -5011 -1204 -5003
rect -1190 -5011 -1186 -5003
rect -1168 -5011 -1164 -5003
rect -1156 -5011 -1152 -5003
rect -1147 -5011 -1143 -5003
rect -1138 -5011 -1134 -5003
rect -935 -5011 -931 -5003
rect -926 -5011 -922 -5003
rect -917 -5011 -913 -5003
rect -909 -5011 -905 -5003
rect -900 -5011 -896 -5003
rect -891 -5011 -887 -5003
rect -883 -5011 -879 -5003
rect -865 -5011 -861 -5003
rect -843 -5011 -839 -5003
rect -831 -5011 -827 -5003
rect -822 -5011 -818 -5003
rect -813 -5011 -809 -5003
rect -805 -5011 -801 -5003
rect -787 -5011 -783 -5003
rect -765 -5011 -761 -5003
rect -753 -5011 -749 -5003
rect -741 -5011 -737 -5003
rect -729 -5011 -725 -5003
rect -721 -5011 -717 -5003
rect -704 -5011 -700 -5003
rect -695 -5011 -691 -5003
rect -577 -5011 -573 -5003
rect -568 -5011 -564 -5003
rect -559 -5011 -555 -5003
rect -551 -5011 -547 -5003
rect -542 -5011 -538 -5003
rect -533 -5011 -529 -5003
rect -525 -5011 -521 -5003
rect -507 -5011 -503 -5003
rect -485 -5011 -481 -5003
rect -473 -5011 -469 -5003
rect -464 -5011 -460 -5003
rect -455 -5011 -451 -5003
rect -447 -5011 -443 -5003
rect -429 -5011 -425 -5003
rect -407 -5011 -403 -5003
rect -395 -5011 -391 -5003
rect -383 -5011 -379 -5003
rect -371 -5011 -367 -5003
rect -363 -5011 -359 -5003
rect -346 -5011 -342 -5003
rect -337 -5011 -333 -5003
rect -219 -5011 -215 -5003
rect -210 -5011 -206 -5003
rect -201 -5011 -197 -5003
rect -193 -5011 -189 -5003
rect -184 -5011 -180 -5003
rect -175 -5011 -171 -5003
rect -167 -5011 -163 -5003
rect -149 -5011 -145 -5003
rect -127 -5011 -123 -5003
rect -115 -5011 -111 -5003
rect -106 -5011 -102 -5003
rect -97 -5011 -93 -5003
rect -89 -5011 -85 -5003
rect -71 -5011 -67 -5003
rect -49 -5011 -45 -5003
rect -37 -5011 -33 -5003
rect -25 -5011 -21 -5003
rect -13 -5011 -9 -5003
rect -5 -5011 -1 -5003
rect 12 -5011 16 -5003
rect 21 -5011 25 -5003
rect 139 -5011 143 -5003
rect 148 -5011 152 -5003
rect 157 -5011 161 -5003
rect 165 -5011 169 -5003
rect 174 -5011 178 -5003
rect 183 -5011 187 -5003
rect 191 -5011 195 -5003
rect 209 -5011 213 -5003
rect 231 -5011 235 -5003
rect 243 -5011 247 -5003
rect 252 -5011 256 -5003
rect 261 -5011 265 -5003
rect 269 -5011 273 -5003
rect 287 -5011 291 -5003
rect 309 -5011 313 -5003
rect 321 -5011 325 -5003
rect 333 -5011 337 -5003
rect 345 -5011 349 -5003
rect 353 -5011 357 -5003
rect 370 -5011 374 -5003
rect 379 -5011 383 -5003
rect 495 -5011 499 -5003
rect 504 -5011 508 -5003
rect 513 -5011 517 -5003
rect 521 -5011 525 -5003
rect 530 -5011 534 -5003
rect 539 -5011 543 -5003
rect 547 -5011 551 -5003
rect 565 -5011 569 -5003
rect 587 -5011 591 -5003
rect 599 -5011 603 -5003
rect 608 -5011 612 -5003
rect 617 -5011 621 -5003
rect 625 -5011 629 -5003
rect 643 -5011 647 -5003
rect 665 -5011 669 -5003
rect 677 -5011 681 -5003
rect 689 -5011 693 -5003
rect 701 -5011 705 -5003
rect 709 -5011 713 -5003
rect 726 -5011 730 -5003
rect 735 -5011 739 -5003
rect 853 -5011 857 -5003
rect 862 -5011 866 -5003
rect 871 -5011 875 -5003
rect 879 -5011 883 -5003
rect 888 -5011 892 -5003
rect 897 -5011 901 -5003
rect 905 -5011 909 -5003
rect 923 -5011 927 -5003
rect 945 -5011 949 -5003
rect 957 -5011 961 -5003
rect 966 -5011 970 -5003
rect 975 -5011 979 -5003
rect 983 -5011 987 -5003
rect 1001 -5011 1005 -5003
rect 1023 -5011 1027 -5003
rect 1035 -5011 1039 -5003
rect 1047 -5011 1051 -5003
rect 1059 -5011 1063 -5003
rect 1067 -5011 1071 -5003
rect 1084 -5011 1088 -5003
rect 1093 -5011 1097 -5003
rect 1211 -5011 1215 -5003
rect 1220 -5011 1224 -5003
rect 1229 -5011 1233 -5003
rect 1237 -5011 1241 -5003
rect 1246 -5011 1250 -5003
rect 1255 -5011 1259 -5003
rect 1263 -5011 1267 -5003
rect 1281 -5011 1285 -5003
rect 1303 -5011 1307 -5003
rect 1315 -5011 1319 -5003
rect 1324 -5011 1328 -5003
rect 1333 -5011 1337 -5003
rect 1341 -5011 1345 -5003
rect 1359 -5011 1363 -5003
rect 1381 -5011 1385 -5003
rect 1393 -5011 1397 -5003
rect 1405 -5011 1409 -5003
rect 1417 -5011 1421 -5003
rect 1425 -5011 1429 -5003
rect 1442 -5011 1446 -5003
rect 1451 -5011 1455 -5003
rect -1810 -5130 -1806 -5122
rect -1801 -5130 -1797 -5122
rect -1792 -5130 -1788 -5122
rect -1784 -5130 -1780 -5122
rect -1776 -5130 -1772 -5122
rect -1764 -5130 -1760 -5122
rect -1752 -5130 -1748 -5122
rect -1743 -5130 -1739 -5122
rect -1734 -5130 -1730 -5122
rect -1722 -5130 -1718 -5122
rect -1710 -5130 -1706 -5122
rect -1701 -5130 -1697 -5122
rect -1692 -5130 -1688 -5122
rect -1680 -5130 -1676 -5122
rect -1668 -5130 -1664 -5122
rect -1659 -5130 -1655 -5122
rect -1650 -5130 -1646 -5122
rect -1638 -5130 -1634 -5122
rect -1626 -5130 -1622 -5122
rect -1618 -5130 -1614 -5122
rect -1547 -5130 -1543 -5122
rect -1538 -5130 -1534 -5122
rect -1529 -5130 -1525 -5122
rect -1521 -5130 -1517 -5122
rect -1513 -5130 -1509 -5122
rect -1501 -5130 -1497 -5122
rect -1489 -5130 -1485 -5122
rect -1480 -5130 -1476 -5122
rect -1471 -5130 -1467 -5122
rect -1459 -5130 -1455 -5122
rect -1447 -5130 -1443 -5122
rect -1438 -5130 -1434 -5122
rect -1429 -5130 -1425 -5122
rect -1417 -5130 -1413 -5122
rect -1405 -5130 -1401 -5122
rect -1396 -5130 -1392 -5122
rect -1387 -5130 -1383 -5122
rect -1375 -5130 -1371 -5122
rect -1363 -5130 -1359 -5122
rect -1355 -5130 -1351 -5122
rect -1234 -5130 -1230 -5122
rect -1225 -5130 -1221 -5122
rect -1216 -5130 -1212 -5122
rect -1208 -5130 -1204 -5122
rect -1200 -5130 -1196 -5122
rect -1188 -5130 -1184 -5122
rect -1176 -5130 -1172 -5122
rect -1167 -5130 -1163 -5122
rect -1158 -5130 -1154 -5122
rect -1146 -5130 -1142 -5122
rect -1134 -5130 -1130 -5122
rect -1125 -5130 -1121 -5122
rect -1116 -5130 -1112 -5122
rect -1104 -5130 -1100 -5122
rect -1092 -5130 -1088 -5122
rect -1083 -5130 -1079 -5122
rect -1074 -5130 -1070 -5122
rect -1062 -5130 -1058 -5122
rect -1050 -5130 -1046 -5122
rect -1042 -5130 -1038 -5122
rect -935 -5130 -931 -5122
rect -926 -5130 -922 -5122
rect -917 -5130 -913 -5122
rect -909 -5130 -905 -5122
rect -901 -5130 -897 -5122
rect -889 -5130 -885 -5122
rect -877 -5130 -873 -5122
rect -868 -5130 -864 -5122
rect -859 -5130 -855 -5122
rect -847 -5130 -843 -5122
rect -835 -5130 -831 -5122
rect -826 -5130 -822 -5122
rect -817 -5130 -813 -5122
rect -805 -5130 -801 -5122
rect -793 -5130 -789 -5122
rect -784 -5130 -780 -5122
rect -775 -5130 -771 -5122
rect -763 -5130 -759 -5122
rect -751 -5130 -747 -5122
rect -743 -5130 -739 -5122
rect -1810 -5301 -1806 -5293
rect -1801 -5301 -1797 -5293
rect -1792 -5301 -1788 -5293
rect -1784 -5301 -1780 -5293
rect -1776 -5301 -1772 -5293
rect -1764 -5301 -1760 -5293
rect -1752 -5301 -1748 -5293
rect -1743 -5301 -1739 -5293
rect -1734 -5301 -1730 -5293
rect -1722 -5301 -1718 -5293
rect -1710 -5301 -1706 -5293
rect -1701 -5301 -1697 -5293
rect -1692 -5301 -1688 -5293
rect -1680 -5301 -1676 -5293
rect -1668 -5301 -1664 -5293
rect -1659 -5301 -1655 -5293
rect -1650 -5301 -1646 -5293
rect -1638 -5301 -1634 -5293
rect -1626 -5301 -1622 -5293
rect -1618 -5301 -1614 -5293
rect -1547 -5301 -1543 -5293
rect -1538 -5301 -1534 -5293
rect -1529 -5301 -1525 -5293
rect -1521 -5301 -1517 -5293
rect -1513 -5301 -1509 -5293
rect -1501 -5301 -1497 -5293
rect -1489 -5301 -1485 -5293
rect -1480 -5301 -1476 -5293
rect -1471 -5301 -1467 -5293
rect -1459 -5301 -1455 -5293
rect -1447 -5301 -1443 -5293
rect -1438 -5301 -1434 -5293
rect -1429 -5301 -1425 -5293
rect -1417 -5301 -1413 -5293
rect -1405 -5301 -1401 -5293
rect -1396 -5301 -1392 -5293
rect -1387 -5301 -1383 -5293
rect -1375 -5301 -1371 -5293
rect -1363 -5301 -1359 -5293
rect -1355 -5301 -1351 -5293
rect -1234 -5301 -1230 -5293
rect -1225 -5301 -1221 -5293
rect -1216 -5301 -1212 -5293
rect -1208 -5301 -1204 -5293
rect -1200 -5301 -1196 -5293
rect -1188 -5301 -1184 -5293
rect -1176 -5301 -1172 -5293
rect -1167 -5301 -1163 -5293
rect -1158 -5301 -1154 -5293
rect -1146 -5301 -1142 -5293
rect -1134 -5301 -1130 -5293
rect -1125 -5301 -1121 -5293
rect -1116 -5301 -1112 -5293
rect -1104 -5301 -1100 -5293
rect -1092 -5301 -1088 -5293
rect -1083 -5301 -1079 -5293
rect -1074 -5301 -1070 -5293
rect -1062 -5301 -1058 -5293
rect -1050 -5301 -1046 -5293
rect -1042 -5301 -1038 -5293
rect -935 -5301 -931 -5293
rect -926 -5301 -922 -5293
rect -917 -5301 -913 -5293
rect -909 -5301 -905 -5293
rect -901 -5301 -897 -5293
rect -889 -5301 -885 -5293
rect -877 -5301 -873 -5293
rect -868 -5301 -864 -5293
rect -859 -5301 -855 -5293
rect -847 -5301 -843 -5293
rect -835 -5301 -831 -5293
rect -826 -5301 -822 -5293
rect -817 -5301 -813 -5293
rect -805 -5301 -801 -5293
rect -793 -5301 -789 -5293
rect -784 -5301 -780 -5293
rect -775 -5301 -771 -5293
rect -763 -5301 -759 -5293
rect -751 -5301 -747 -5293
rect -743 -5301 -739 -5293
rect -577 -5301 -573 -5293
rect -568 -5301 -564 -5293
rect -559 -5301 -555 -5293
rect -551 -5301 -547 -5293
rect -543 -5301 -539 -5293
rect -531 -5301 -527 -5293
rect -519 -5301 -515 -5293
rect -510 -5301 -506 -5293
rect -501 -5301 -497 -5293
rect -489 -5301 -485 -5293
rect -477 -5301 -473 -5293
rect -468 -5301 -464 -5293
rect -459 -5301 -455 -5293
rect -447 -5301 -443 -5293
rect -435 -5301 -431 -5293
rect -426 -5301 -422 -5293
rect -417 -5301 -413 -5293
rect -405 -5301 -401 -5293
rect -393 -5301 -389 -5293
rect -385 -5301 -381 -5293
rect -219 -5301 -215 -5293
rect -210 -5301 -206 -5293
rect -201 -5301 -197 -5293
rect -193 -5301 -189 -5293
rect -185 -5301 -181 -5293
rect -173 -5301 -169 -5293
rect -161 -5301 -157 -5293
rect -152 -5301 -148 -5293
rect -143 -5301 -139 -5293
rect -131 -5301 -127 -5293
rect -119 -5301 -115 -5293
rect -110 -5301 -106 -5293
rect -101 -5301 -97 -5293
rect -89 -5301 -85 -5293
rect -77 -5301 -73 -5293
rect -68 -5301 -64 -5293
rect -59 -5301 -55 -5293
rect -47 -5301 -43 -5293
rect -35 -5301 -31 -5293
rect -27 -5301 -23 -5293
rect 139 -5301 143 -5293
rect 148 -5301 152 -5293
rect 157 -5301 161 -5293
rect 165 -5301 169 -5293
rect 173 -5301 177 -5293
rect 185 -5301 189 -5293
rect 197 -5301 201 -5293
rect 206 -5301 210 -5293
rect 215 -5301 219 -5293
rect 227 -5301 231 -5293
rect 239 -5301 243 -5293
rect 248 -5301 252 -5293
rect 257 -5301 261 -5293
rect 269 -5301 273 -5293
rect 281 -5301 285 -5293
rect 290 -5301 294 -5293
rect 299 -5301 303 -5293
rect 311 -5301 315 -5293
rect 323 -5301 327 -5293
rect 331 -5301 335 -5293
rect 495 -5301 499 -5293
rect 504 -5301 508 -5293
rect 513 -5301 517 -5293
rect 521 -5301 525 -5293
rect 529 -5301 533 -5293
rect 541 -5301 545 -5293
rect 553 -5301 557 -5293
rect 562 -5301 566 -5293
rect 571 -5301 575 -5293
rect 583 -5301 587 -5293
rect 595 -5301 599 -5293
rect 604 -5301 608 -5293
rect 613 -5301 617 -5293
rect 625 -5301 629 -5293
rect 637 -5301 641 -5293
rect 646 -5301 650 -5293
rect 655 -5301 659 -5293
rect 667 -5301 671 -5293
rect 679 -5301 683 -5293
rect 687 -5301 691 -5293
rect 853 -5301 857 -5293
rect 862 -5301 866 -5293
rect 871 -5301 875 -5293
rect 879 -5301 883 -5293
rect 887 -5301 891 -5293
rect 899 -5301 903 -5293
rect 911 -5301 915 -5293
rect 920 -5301 924 -5293
rect 929 -5301 933 -5293
rect 941 -5301 945 -5293
rect 953 -5301 957 -5293
rect 962 -5301 966 -5293
rect 971 -5301 975 -5293
rect 983 -5301 987 -5293
rect 995 -5301 999 -5293
rect 1004 -5301 1008 -5293
rect 1013 -5301 1017 -5293
rect 1025 -5301 1029 -5293
rect 1037 -5301 1041 -5293
rect 1045 -5301 1049 -5293
rect 1211 -5301 1215 -5293
rect 1220 -5301 1224 -5293
rect 1229 -5301 1233 -5293
rect 1237 -5301 1241 -5293
rect 1245 -5301 1249 -5293
rect 1257 -5301 1261 -5293
rect 1269 -5301 1273 -5293
rect 1278 -5301 1282 -5293
rect 1287 -5301 1291 -5293
rect 1299 -5301 1303 -5293
rect 1311 -5301 1315 -5293
rect 1320 -5301 1324 -5293
rect 1329 -5301 1333 -5293
rect 1341 -5301 1345 -5293
rect 1353 -5301 1357 -5293
rect 1362 -5301 1366 -5293
rect 1371 -5301 1375 -5293
rect 1383 -5301 1387 -5293
rect 1395 -5301 1399 -5293
rect 1403 -5301 1407 -5293
rect -1810 -5461 -1806 -5453
rect -1801 -5461 -1797 -5453
rect -1792 -5461 -1788 -5453
rect -1784 -5461 -1780 -5453
rect -1776 -5461 -1772 -5453
rect -1764 -5461 -1760 -5453
rect -1752 -5461 -1748 -5453
rect -1743 -5461 -1739 -5453
rect -1734 -5461 -1730 -5453
rect -1722 -5461 -1718 -5453
rect -1710 -5461 -1706 -5453
rect -1701 -5461 -1697 -5453
rect -1692 -5461 -1688 -5453
rect -1680 -5461 -1676 -5453
rect -1668 -5461 -1664 -5453
rect -1659 -5461 -1655 -5453
rect -1650 -5461 -1646 -5453
rect -1638 -5461 -1634 -5453
rect -1626 -5461 -1622 -5453
rect -1618 -5461 -1614 -5453
rect -1547 -5461 -1543 -5453
rect -1538 -5461 -1534 -5453
rect -1529 -5461 -1525 -5453
rect -1521 -5461 -1517 -5453
rect -1513 -5461 -1509 -5453
rect -1501 -5461 -1497 -5453
rect -1489 -5461 -1485 -5453
rect -1480 -5461 -1476 -5453
rect -1471 -5461 -1467 -5453
rect -1459 -5461 -1455 -5453
rect -1447 -5461 -1443 -5453
rect -1438 -5461 -1434 -5453
rect -1429 -5461 -1425 -5453
rect -1417 -5461 -1413 -5453
rect -1405 -5461 -1401 -5453
rect -1396 -5461 -1392 -5453
rect -1387 -5461 -1383 -5453
rect -1375 -5461 -1371 -5453
rect -1363 -5461 -1359 -5453
rect -1355 -5461 -1351 -5453
rect -1234 -5461 -1230 -5453
rect -1225 -5461 -1221 -5453
rect -1216 -5461 -1212 -5453
rect -1208 -5461 -1204 -5453
rect -1200 -5461 -1196 -5453
rect -1188 -5461 -1184 -5453
rect -1176 -5461 -1172 -5453
rect -1167 -5461 -1163 -5453
rect -1158 -5461 -1154 -5453
rect -1146 -5461 -1142 -5453
rect -1134 -5461 -1130 -5453
rect -1125 -5461 -1121 -5453
rect -1116 -5461 -1112 -5453
rect -1104 -5461 -1100 -5453
rect -1092 -5461 -1088 -5453
rect -1083 -5461 -1079 -5453
rect -1074 -5461 -1070 -5453
rect -1062 -5461 -1058 -5453
rect -1050 -5461 -1046 -5453
rect -1042 -5461 -1038 -5453
rect -935 -5461 -931 -5453
rect -926 -5461 -922 -5453
rect -917 -5461 -913 -5453
rect -909 -5461 -905 -5453
rect -901 -5461 -897 -5453
rect -889 -5461 -885 -5453
rect -877 -5461 -873 -5453
rect -868 -5461 -864 -5453
rect -859 -5461 -855 -5453
rect -847 -5461 -843 -5453
rect -835 -5461 -831 -5453
rect -826 -5461 -822 -5453
rect -817 -5461 -813 -5453
rect -805 -5461 -801 -5453
rect -793 -5461 -789 -5453
rect -784 -5461 -780 -5453
rect -775 -5461 -771 -5453
rect -763 -5461 -759 -5453
rect -751 -5461 -747 -5453
rect -743 -5461 -739 -5453
rect -577 -5461 -573 -5453
rect -568 -5461 -564 -5453
rect -559 -5461 -555 -5453
rect -551 -5461 -547 -5453
rect -543 -5461 -539 -5453
rect -531 -5461 -527 -5453
rect -519 -5461 -515 -5453
rect -510 -5461 -506 -5453
rect -501 -5461 -497 -5453
rect -489 -5461 -485 -5453
rect -477 -5461 -473 -5453
rect -468 -5461 -464 -5453
rect -459 -5461 -455 -5453
rect -447 -5461 -443 -5453
rect -435 -5461 -431 -5453
rect -426 -5461 -422 -5453
rect -417 -5461 -413 -5453
rect -405 -5461 -401 -5453
rect -393 -5461 -389 -5453
rect -385 -5461 -381 -5453
rect -219 -5461 -215 -5453
rect -210 -5461 -206 -5453
rect -201 -5461 -197 -5453
rect -193 -5461 -189 -5453
rect -185 -5461 -181 -5453
rect -173 -5461 -169 -5453
rect -161 -5461 -157 -5453
rect -152 -5461 -148 -5453
rect -143 -5461 -139 -5453
rect -131 -5461 -127 -5453
rect -119 -5461 -115 -5453
rect -110 -5461 -106 -5453
rect -101 -5461 -97 -5453
rect -89 -5461 -85 -5453
rect -77 -5461 -73 -5453
rect -68 -5461 -64 -5453
rect -59 -5461 -55 -5453
rect -47 -5461 -43 -5453
rect -35 -5461 -31 -5453
rect -27 -5461 -23 -5453
rect 139 -5461 143 -5453
rect 148 -5461 152 -5453
rect 157 -5461 161 -5453
rect 165 -5461 169 -5453
rect 173 -5461 177 -5453
rect 185 -5461 189 -5453
rect 197 -5461 201 -5453
rect 206 -5461 210 -5453
rect 215 -5461 219 -5453
rect 227 -5461 231 -5453
rect 239 -5461 243 -5453
rect 248 -5461 252 -5453
rect 257 -5461 261 -5453
rect 269 -5461 273 -5453
rect 281 -5461 285 -5453
rect 290 -5461 294 -5453
rect 299 -5461 303 -5453
rect 311 -5461 315 -5453
rect 323 -5461 327 -5453
rect 331 -5461 335 -5453
rect 495 -5461 499 -5453
rect 504 -5461 508 -5453
rect 513 -5461 517 -5453
rect 521 -5461 525 -5453
rect 529 -5461 533 -5453
rect 541 -5461 545 -5453
rect 553 -5461 557 -5453
rect 562 -5461 566 -5453
rect 571 -5461 575 -5453
rect 583 -5461 587 -5453
rect 595 -5461 599 -5453
rect 604 -5461 608 -5453
rect 613 -5461 617 -5453
rect 625 -5461 629 -5453
rect 637 -5461 641 -5453
rect 646 -5461 650 -5453
rect 655 -5461 659 -5453
rect 667 -5461 671 -5453
rect 679 -5461 683 -5453
rect 687 -5461 691 -5453
rect 853 -5461 857 -5453
rect 862 -5461 866 -5453
rect 871 -5461 875 -5453
rect 879 -5461 883 -5453
rect 887 -5461 891 -5453
rect 899 -5461 903 -5453
rect 911 -5461 915 -5453
rect 920 -5461 924 -5453
rect 929 -5461 933 -5453
rect 941 -5461 945 -5453
rect 953 -5461 957 -5453
rect 962 -5461 966 -5453
rect 971 -5461 975 -5453
rect 983 -5461 987 -5453
rect 995 -5461 999 -5453
rect 1004 -5461 1008 -5453
rect 1013 -5461 1017 -5453
rect 1025 -5461 1029 -5453
rect 1037 -5461 1041 -5453
rect 1045 -5461 1049 -5453
rect 1211 -5461 1215 -5453
rect 1220 -5461 1224 -5453
rect 1229 -5461 1233 -5453
rect 1237 -5461 1241 -5453
rect 1245 -5461 1249 -5453
rect 1257 -5461 1261 -5453
rect 1269 -5461 1273 -5453
rect 1278 -5461 1282 -5453
rect 1287 -5461 1291 -5453
rect 1299 -5461 1303 -5453
rect 1311 -5461 1315 -5453
rect 1320 -5461 1324 -5453
rect 1329 -5461 1333 -5453
rect 1341 -5461 1345 -5453
rect 1353 -5461 1357 -5453
rect 1362 -5461 1366 -5453
rect 1371 -5461 1375 -5453
rect 1383 -5461 1387 -5453
rect 1395 -5461 1399 -5453
rect 1403 -5461 1407 -5453
rect -1309 -5575 -1305 -5567
rect -1301 -5575 -1297 -5567
rect -1292 -5575 -1288 -5567
rect -1283 -5575 -1279 -5567
rect -935 -5575 -931 -5567
rect -927 -5575 -923 -5567
rect -918 -5575 -914 -5567
rect -909 -5575 -905 -5567
rect -577 -5575 -573 -5567
rect -569 -5575 -565 -5567
rect -560 -5575 -556 -5567
rect -551 -5575 -547 -5567
rect -219 -5575 -215 -5567
rect -211 -5575 -207 -5567
rect -202 -5575 -198 -5567
rect -193 -5575 -189 -5567
rect 139 -5575 143 -5567
rect 147 -5575 151 -5567
rect 156 -5575 160 -5567
rect 165 -5575 169 -5567
rect 495 -5575 499 -5567
rect 503 -5575 507 -5567
rect 512 -5575 516 -5567
rect 521 -5575 525 -5567
rect 853 -5575 857 -5567
rect 861 -5575 865 -5567
rect 870 -5575 874 -5567
rect 879 -5575 883 -5567
rect 1211 -5575 1215 -5567
rect 1219 -5575 1223 -5567
rect 1228 -5575 1232 -5567
rect 1237 -5575 1241 -5567
rect -1234 -5734 -1230 -5726
rect -1225 -5734 -1221 -5726
rect -1216 -5734 -1212 -5726
rect -1208 -5734 -1204 -5726
rect -1190 -5734 -1186 -5726
rect -1168 -5734 -1164 -5726
rect -1156 -5734 -1152 -5726
rect -1147 -5734 -1143 -5726
rect -1138 -5734 -1134 -5726
rect -935 -5734 -931 -5726
rect -926 -5734 -922 -5726
rect -917 -5734 -913 -5726
rect -909 -5734 -905 -5726
rect -900 -5734 -896 -5726
rect -891 -5734 -887 -5726
rect -883 -5734 -879 -5726
rect -865 -5734 -861 -5726
rect -843 -5734 -839 -5726
rect -831 -5734 -827 -5726
rect -822 -5734 -818 -5726
rect -813 -5734 -809 -5726
rect -805 -5734 -801 -5726
rect -787 -5734 -783 -5726
rect -765 -5734 -761 -5726
rect -753 -5734 -749 -5726
rect -741 -5734 -737 -5726
rect -729 -5734 -725 -5726
rect -721 -5734 -717 -5726
rect -704 -5734 -700 -5726
rect -695 -5734 -691 -5726
rect -577 -5734 -573 -5726
rect -568 -5734 -564 -5726
rect -559 -5734 -555 -5726
rect -551 -5734 -547 -5726
rect -542 -5734 -538 -5726
rect -533 -5734 -529 -5726
rect -525 -5734 -521 -5726
rect -507 -5734 -503 -5726
rect -485 -5734 -481 -5726
rect -473 -5734 -469 -5726
rect -464 -5734 -460 -5726
rect -455 -5734 -451 -5726
rect -447 -5734 -443 -5726
rect -429 -5734 -425 -5726
rect -407 -5734 -403 -5726
rect -395 -5734 -391 -5726
rect -383 -5734 -379 -5726
rect -371 -5734 -367 -5726
rect -363 -5734 -359 -5726
rect -346 -5734 -342 -5726
rect -337 -5734 -333 -5726
rect -219 -5734 -215 -5726
rect -210 -5734 -206 -5726
rect -201 -5734 -197 -5726
rect -193 -5734 -189 -5726
rect -184 -5734 -180 -5726
rect -175 -5734 -171 -5726
rect -167 -5734 -163 -5726
rect -149 -5734 -145 -5726
rect -127 -5734 -123 -5726
rect -115 -5734 -111 -5726
rect -106 -5734 -102 -5726
rect -97 -5734 -93 -5726
rect -89 -5734 -85 -5726
rect -71 -5734 -67 -5726
rect -49 -5734 -45 -5726
rect -37 -5734 -33 -5726
rect -25 -5734 -21 -5726
rect -13 -5734 -9 -5726
rect -5 -5734 -1 -5726
rect 12 -5734 16 -5726
rect 21 -5734 25 -5726
rect 139 -5734 143 -5726
rect 148 -5734 152 -5726
rect 157 -5734 161 -5726
rect 165 -5734 169 -5726
rect 174 -5734 178 -5726
rect 183 -5734 187 -5726
rect 191 -5734 195 -5726
rect 209 -5734 213 -5726
rect 231 -5734 235 -5726
rect 243 -5734 247 -5726
rect 252 -5734 256 -5726
rect 261 -5734 265 -5726
rect 269 -5734 273 -5726
rect 287 -5734 291 -5726
rect 309 -5734 313 -5726
rect 321 -5734 325 -5726
rect 333 -5734 337 -5726
rect 345 -5734 349 -5726
rect 353 -5734 357 -5726
rect 370 -5734 374 -5726
rect 379 -5734 383 -5726
rect 495 -5734 499 -5726
rect 504 -5734 508 -5726
rect 513 -5734 517 -5726
rect 521 -5734 525 -5726
rect 530 -5734 534 -5726
rect 539 -5734 543 -5726
rect 547 -5734 551 -5726
rect 565 -5734 569 -5726
rect 587 -5734 591 -5726
rect 599 -5734 603 -5726
rect 608 -5734 612 -5726
rect 617 -5734 621 -5726
rect 625 -5734 629 -5726
rect 643 -5734 647 -5726
rect 665 -5734 669 -5726
rect 677 -5734 681 -5726
rect 689 -5734 693 -5726
rect 701 -5734 705 -5726
rect 709 -5734 713 -5726
rect 726 -5734 730 -5726
rect 735 -5734 739 -5726
rect 853 -5734 857 -5726
rect 862 -5734 866 -5726
rect 871 -5734 875 -5726
rect 879 -5734 883 -5726
rect 888 -5734 892 -5726
rect 897 -5734 901 -5726
rect 905 -5734 909 -5726
rect 923 -5734 927 -5726
rect 945 -5734 949 -5726
rect 957 -5734 961 -5726
rect 966 -5734 970 -5726
rect 975 -5734 979 -5726
rect 983 -5734 987 -5726
rect 1001 -5734 1005 -5726
rect 1023 -5734 1027 -5726
rect 1035 -5734 1039 -5726
rect 1047 -5734 1051 -5726
rect 1059 -5734 1063 -5726
rect 1067 -5734 1071 -5726
rect 1084 -5734 1088 -5726
rect 1093 -5734 1097 -5726
rect 1211 -5734 1215 -5726
rect 1220 -5734 1224 -5726
rect 1229 -5734 1233 -5726
rect 1237 -5734 1241 -5726
rect 1246 -5734 1250 -5726
rect 1255 -5734 1259 -5726
rect 1263 -5734 1267 -5726
rect 1281 -5734 1285 -5726
rect 1303 -5734 1307 -5726
rect 1315 -5734 1319 -5726
rect 1324 -5734 1328 -5726
rect 1333 -5734 1337 -5726
rect 1341 -5734 1345 -5726
rect 1359 -5734 1363 -5726
rect 1381 -5734 1385 -5726
rect 1393 -5734 1397 -5726
rect 1405 -5734 1409 -5726
rect 1417 -5734 1421 -5726
rect 1425 -5734 1429 -5726
rect 1442 -5734 1446 -5726
rect 1451 -5734 1455 -5726
rect -1234 -5857 -1230 -5849
rect -1225 -5857 -1221 -5849
rect -1216 -5857 -1212 -5849
rect -1208 -5857 -1204 -5849
rect -1200 -5857 -1196 -5849
rect -1188 -5857 -1184 -5849
rect -1176 -5857 -1172 -5849
rect -1167 -5857 -1163 -5849
rect -1158 -5857 -1154 -5849
rect -1146 -5857 -1142 -5849
rect -1134 -5857 -1130 -5849
rect -1125 -5857 -1121 -5849
rect -1116 -5857 -1112 -5849
rect -1104 -5857 -1100 -5849
rect -1092 -5857 -1088 -5849
rect -1083 -5857 -1079 -5849
rect -1074 -5857 -1070 -5849
rect -1062 -5857 -1058 -5849
rect -1050 -5857 -1046 -5849
rect -1042 -5857 -1038 -5849
rect -935 -5857 -931 -5849
rect -926 -5857 -922 -5849
rect -917 -5857 -913 -5849
rect -909 -5857 -905 -5849
rect -901 -5857 -897 -5849
rect -889 -5857 -885 -5849
rect -877 -5857 -873 -5849
rect -868 -5857 -864 -5849
rect -859 -5857 -855 -5849
rect -847 -5857 -843 -5849
rect -835 -5857 -831 -5849
rect -826 -5857 -822 -5849
rect -817 -5857 -813 -5849
rect -805 -5857 -801 -5849
rect -793 -5857 -789 -5849
rect -784 -5857 -780 -5849
rect -775 -5857 -771 -5849
rect -763 -5857 -759 -5849
rect -751 -5857 -747 -5849
rect -743 -5857 -739 -5849
rect -577 -5857 -573 -5849
rect -568 -5857 -564 -5849
rect -559 -5857 -555 -5849
rect -551 -5857 -547 -5849
rect -543 -5857 -539 -5849
rect -531 -5857 -527 -5849
rect -519 -5857 -515 -5849
rect -510 -5857 -506 -5849
rect -501 -5857 -497 -5849
rect -489 -5857 -485 -5849
rect -477 -5857 -473 -5849
rect -468 -5857 -464 -5849
rect -459 -5857 -455 -5849
rect -447 -5857 -443 -5849
rect -435 -5857 -431 -5849
rect -426 -5857 -422 -5849
rect -417 -5857 -413 -5849
rect -405 -5857 -401 -5849
rect -393 -5857 -389 -5849
rect -385 -5857 -381 -5849
rect -219 -5857 -215 -5849
rect -210 -5857 -206 -5849
rect -201 -5857 -197 -5849
rect -193 -5857 -189 -5849
rect -185 -5857 -181 -5849
rect -173 -5857 -169 -5849
rect -161 -5857 -157 -5849
rect -152 -5857 -148 -5849
rect -143 -5857 -139 -5849
rect -131 -5857 -127 -5849
rect -119 -5857 -115 -5849
rect -110 -5857 -106 -5849
rect -101 -5857 -97 -5849
rect -89 -5857 -85 -5849
rect -77 -5857 -73 -5849
rect -68 -5857 -64 -5849
rect -59 -5857 -55 -5849
rect -47 -5857 -43 -5849
rect -35 -5857 -31 -5849
rect -27 -5857 -23 -5849
rect 139 -5857 143 -5849
rect 148 -5857 152 -5849
rect 157 -5857 161 -5849
rect 165 -5857 169 -5849
rect 173 -5857 177 -5849
rect 185 -5857 189 -5849
rect 197 -5857 201 -5849
rect 206 -5857 210 -5849
rect 215 -5857 219 -5849
rect 227 -5857 231 -5849
rect 239 -5857 243 -5849
rect 248 -5857 252 -5849
rect 257 -5857 261 -5849
rect 269 -5857 273 -5849
rect 281 -5857 285 -5849
rect 290 -5857 294 -5849
rect 299 -5857 303 -5849
rect 311 -5857 315 -5849
rect 323 -5857 327 -5849
rect 331 -5857 335 -5849
rect 495 -5857 499 -5849
rect 504 -5857 508 -5849
rect 513 -5857 517 -5849
rect 521 -5857 525 -5849
rect 529 -5857 533 -5849
rect 541 -5857 545 -5849
rect 553 -5857 557 -5849
rect 562 -5857 566 -5849
rect 571 -5857 575 -5849
rect 583 -5857 587 -5849
rect 595 -5857 599 -5849
rect 604 -5857 608 -5849
rect 613 -5857 617 -5849
rect 625 -5857 629 -5849
rect 637 -5857 641 -5849
rect 646 -5857 650 -5849
rect 655 -5857 659 -5849
rect 667 -5857 671 -5849
rect 679 -5857 683 -5849
rect 687 -5857 691 -5849
rect 853 -5857 857 -5849
rect 862 -5857 866 -5849
rect 871 -5857 875 -5849
rect 879 -5857 883 -5849
rect 887 -5857 891 -5849
rect 899 -5857 903 -5849
rect 911 -5857 915 -5849
rect 920 -5857 924 -5849
rect 929 -5857 933 -5849
rect 941 -5857 945 -5849
rect 953 -5857 957 -5849
rect 962 -5857 966 -5849
rect 971 -5857 975 -5849
rect 983 -5857 987 -5849
rect 995 -5857 999 -5849
rect 1004 -5857 1008 -5849
rect 1013 -5857 1017 -5849
rect 1025 -5857 1029 -5849
rect 1037 -5857 1041 -5849
rect 1045 -5857 1049 -5849
rect 1211 -5857 1215 -5849
rect 1220 -5857 1224 -5849
rect 1229 -5857 1233 -5849
rect 1237 -5857 1241 -5849
rect 1245 -5857 1249 -5849
rect 1257 -5857 1261 -5849
rect 1269 -5857 1273 -5849
rect 1278 -5857 1282 -5849
rect 1287 -5857 1291 -5849
rect 1299 -5857 1303 -5849
rect 1311 -5857 1315 -5849
rect 1320 -5857 1324 -5849
rect 1329 -5857 1333 -5849
rect 1341 -5857 1345 -5849
rect 1353 -5857 1357 -5849
rect 1362 -5857 1366 -5849
rect 1371 -5857 1375 -5849
rect 1383 -5857 1387 -5849
rect 1395 -5857 1399 -5849
rect 1403 -5857 1407 -5849
rect 1555 -5857 1559 -5849
rect 1564 -5857 1568 -5849
rect 1573 -5857 1577 -5849
rect 1581 -5857 1585 -5849
rect 1589 -5857 1593 -5849
rect 1601 -5857 1605 -5849
rect 1613 -5857 1617 -5849
rect 1622 -5857 1626 -5849
rect 1631 -5857 1635 -5849
rect 1643 -5857 1647 -5849
rect 1655 -5857 1659 -5849
rect 1664 -5857 1668 -5849
rect 1673 -5857 1677 -5849
rect 1685 -5857 1689 -5849
rect 1697 -5857 1701 -5849
rect 1706 -5857 1710 -5849
rect 1715 -5857 1719 -5849
rect 1727 -5857 1731 -5849
rect 1739 -5857 1743 -5849
rect 1747 -5857 1751 -5849
<< m2contact >>
rect -1307 -784 -1303 -780
rect -1290 -784 -1286 -780
rect -936 -784 -932 -780
rect -919 -784 -915 -780
rect -964 -832 -960 -828
rect -1290 -876 -1286 -872
rect -1281 -1074 -1277 -1070
rect -1251 -840 -1247 -836
rect -1309 -1134 -1305 -1130
rect -1292 -1134 -1288 -1130
rect -1550 -1763 -1546 -1759
rect -1533 -1763 -1529 -1759
rect -1513 -1763 -1509 -1759
rect -1492 -1763 -1488 -1759
rect -1471 -1763 -1467 -1759
rect -1450 -1763 -1446 -1759
rect -1429 -1763 -1425 -1759
rect -1408 -1763 -1404 -1759
rect -1387 -1763 -1383 -1759
rect -1367 -1763 -1363 -1759
rect -1559 -1826 -1555 -1822
rect -1501 -1819 -1497 -1815
rect -1459 -1826 -1455 -1822
rect -1441 -1819 -1437 -1815
rect -1399 -1803 -1395 -1799
rect -1399 -1819 -1395 -1815
rect -1417 -1833 -1413 -1829
rect -1517 -1840 -1513 -1836
rect -1475 -1840 -1471 -1836
rect -1351 -1803 -1347 -1799
rect -1375 -1826 -1371 -1822
rect -1550 -1855 -1546 -1851
rect -1533 -1855 -1529 -1851
rect -1492 -1855 -1488 -1851
rect -1450 -1855 -1446 -1851
rect -1408 -1855 -1404 -1851
rect -1367 -1855 -1363 -1851
rect -1292 -1226 -1288 -1222
rect -1221 -1018 -1217 -1014
rect -1204 -1018 -1200 -1014
rect -1184 -1018 -1180 -1014
rect -1163 -1018 -1159 -1014
rect -1142 -1018 -1138 -1014
rect -1121 -1018 -1117 -1014
rect -1100 -1018 -1096 -1014
rect -1079 -1018 -1075 -1014
rect -1058 -1018 -1054 -1014
rect -1038 -1018 -1034 -1014
rect -1230 -1081 -1226 -1077
rect -1172 -1074 -1168 -1070
rect -1130 -1081 -1126 -1077
rect -1112 -1074 -1108 -1070
rect -1070 -1066 -1066 -1062
rect -1070 -1074 -1066 -1070
rect -1088 -1088 -1084 -1084
rect -1188 -1095 -1184 -1091
rect -1146 -1095 -1142 -1091
rect -1046 -1081 -1042 -1077
rect -1221 -1110 -1217 -1106
rect -1204 -1110 -1200 -1106
rect -1163 -1110 -1159 -1106
rect -1121 -1110 -1117 -1106
rect -1079 -1110 -1075 -1106
rect -1038 -1110 -1034 -1106
rect -976 -1187 -972 -1183
rect -1221 -1298 -1217 -1294
rect -1204 -1298 -1200 -1294
rect -1164 -1298 -1160 -1294
rect -1143 -1298 -1139 -1294
rect -1251 -1354 -1247 -1350
rect -1230 -1347 -1226 -1343
rect -1283 -1361 -1279 -1357
rect -1186 -1368 -1182 -1364
rect -1134 -1346 -1130 -1342
rect -1204 -1375 -1200 -1371
rect -1168 -1375 -1164 -1371
rect -964 -1338 -960 -1334
rect -577 -784 -573 -780
rect -560 -784 -556 -780
rect -910 -840 -906 -836
rect -605 -840 -601 -836
rect -919 -876 -915 -872
rect -926 -1018 -922 -1014
rect -909 -1018 -905 -1014
rect -889 -1018 -885 -1014
rect -868 -1018 -864 -1014
rect -847 -1018 -843 -1014
rect -826 -1018 -822 -1014
rect -805 -1018 -801 -1014
rect -784 -1018 -780 -1014
rect -763 -1018 -759 -1014
rect -743 -1018 -739 -1014
rect -935 -1081 -931 -1077
rect -877 -1074 -873 -1070
rect -835 -1081 -831 -1077
rect -817 -1074 -813 -1070
rect -775 -1066 -771 -1062
rect -775 -1074 -771 -1070
rect -793 -1088 -789 -1084
rect -893 -1095 -889 -1091
rect -851 -1095 -847 -1091
rect -751 -1081 -747 -1077
rect -926 -1110 -922 -1106
rect -909 -1110 -905 -1106
rect -868 -1110 -864 -1106
rect -826 -1110 -822 -1106
rect -784 -1110 -780 -1106
rect -743 -1110 -739 -1106
rect -935 -1134 -931 -1130
rect -918 -1134 -914 -1130
rect -976 -1353 -972 -1349
rect -1124 -1368 -1120 -1364
rect -1221 -1390 -1217 -1386
rect -1177 -1390 -1173 -1386
rect -1143 -1390 -1139 -1386
rect -1257 -1397 -1253 -1393
rect -1244 -1404 -1240 -1400
rect -1124 -1404 -1120 -1400
rect -976 -1404 -972 -1400
rect -1221 -1421 -1217 -1417
rect -1204 -1421 -1200 -1417
rect -1184 -1421 -1180 -1417
rect -1163 -1421 -1159 -1417
rect -1142 -1421 -1138 -1417
rect -1121 -1421 -1117 -1417
rect -1100 -1421 -1096 -1417
rect -1079 -1421 -1075 -1417
rect -1058 -1421 -1054 -1417
rect -1038 -1421 -1034 -1417
rect -1244 -1477 -1240 -1473
rect -1230 -1484 -1226 -1480
rect -1172 -1477 -1168 -1473
rect -1130 -1484 -1126 -1480
rect -1112 -1477 -1108 -1473
rect -1070 -1469 -1066 -1465
rect -1070 -1477 -1066 -1473
rect -1088 -1491 -1084 -1487
rect -1188 -1498 -1184 -1494
rect -1146 -1498 -1142 -1494
rect -1046 -1484 -1042 -1480
rect -1221 -1513 -1217 -1509
rect -1204 -1513 -1200 -1509
rect -1163 -1513 -1159 -1509
rect -1121 -1513 -1117 -1509
rect -1079 -1513 -1075 -1509
rect -1038 -1513 -1034 -1509
rect -1221 -1592 -1217 -1588
rect -1204 -1592 -1200 -1588
rect -1184 -1592 -1180 -1588
rect -1163 -1592 -1159 -1588
rect -1142 -1592 -1138 -1588
rect -1121 -1592 -1117 -1588
rect -1100 -1592 -1096 -1588
rect -1079 -1592 -1075 -1588
rect -1058 -1592 -1054 -1588
rect -1038 -1592 -1034 -1588
rect -1257 -1648 -1253 -1644
rect -1230 -1655 -1226 -1651
rect -1172 -1648 -1168 -1644
rect -1130 -1655 -1126 -1651
rect -1112 -1648 -1108 -1644
rect -1070 -1640 -1066 -1636
rect -1070 -1648 -1066 -1644
rect -1088 -1662 -1084 -1658
rect -1188 -1669 -1184 -1665
rect -1146 -1669 -1142 -1665
rect -1023 -1640 -1019 -1636
rect -1046 -1655 -1042 -1651
rect -1221 -1684 -1217 -1680
rect -1204 -1684 -1200 -1680
rect -1163 -1684 -1159 -1680
rect -1121 -1684 -1117 -1680
rect -1079 -1684 -1075 -1680
rect -1038 -1684 -1034 -1680
rect -976 -1648 -972 -1644
rect -1319 -1819 -1315 -1815
rect -1257 -1691 -1253 -1687
rect -1023 -1691 -1019 -1687
rect -1309 -1870 -1305 -1866
rect -1292 -1870 -1288 -1866
rect -1351 -1910 -1347 -1906
rect -1550 -2344 -1546 -2340
rect -1533 -2344 -1529 -2340
rect -1513 -2344 -1509 -2340
rect -1492 -2344 -1488 -2340
rect -1471 -2344 -1467 -2340
rect -1450 -2344 -1446 -2340
rect -1429 -2344 -1425 -2340
rect -1408 -2344 -1404 -2340
rect -1387 -2344 -1383 -2340
rect -1367 -2344 -1363 -2340
rect -1559 -2407 -1555 -2403
rect -1501 -2400 -1497 -2396
rect -1459 -2407 -1455 -2403
rect -1441 -2400 -1437 -2396
rect -1399 -2392 -1395 -2388
rect -1399 -2400 -1395 -2396
rect -1417 -2414 -1413 -2410
rect -1517 -2421 -1513 -2417
rect -1475 -2421 -1471 -2417
rect -1350 -2392 -1346 -2388
rect -1375 -2407 -1371 -2403
rect -1550 -2436 -1546 -2432
rect -1533 -2436 -1529 -2432
rect -1492 -2436 -1488 -2432
rect -1450 -2436 -1446 -2432
rect -1408 -2436 -1404 -2432
rect -1367 -2436 -1363 -2432
rect -1581 -2444 -1577 -2440
rect -1350 -2444 -1346 -2440
rect -1550 -2515 -1546 -2511
rect -1533 -2515 -1529 -2511
rect -1513 -2515 -1509 -2511
rect -1492 -2515 -1488 -2511
rect -1471 -2515 -1467 -2511
rect -1450 -2515 -1446 -2511
rect -1429 -2515 -1425 -2511
rect -1408 -2515 -1404 -2511
rect -1387 -2515 -1383 -2511
rect -1367 -2515 -1363 -2511
rect -1581 -2571 -1577 -2567
rect -1559 -2578 -1555 -2574
rect -1501 -2571 -1497 -2567
rect -1459 -2578 -1455 -2574
rect -1441 -2571 -1437 -2567
rect -1399 -2563 -1395 -2559
rect -1399 -2571 -1395 -2567
rect -1417 -2585 -1413 -2581
rect -1517 -2592 -1513 -2588
rect -1475 -2592 -1471 -2588
rect -1355 -2563 -1351 -2559
rect -1375 -2578 -1371 -2574
rect -1550 -2607 -1546 -2603
rect -1533 -2607 -1529 -2603
rect -1492 -2607 -1488 -2603
rect -1450 -2607 -1446 -2603
rect -1408 -2607 -1404 -2603
rect -1367 -2607 -1363 -2603
rect -1292 -1962 -1288 -1958
rect -976 -1692 -972 -1688
rect -1221 -1763 -1217 -1759
rect -1204 -1763 -1200 -1759
rect -1184 -1763 -1180 -1759
rect -1163 -1763 -1159 -1759
rect -1142 -1763 -1138 -1759
rect -1121 -1763 -1117 -1759
rect -1100 -1763 -1096 -1759
rect -1079 -1763 -1075 -1759
rect -1058 -1763 -1054 -1759
rect -1038 -1763 -1034 -1759
rect -1230 -1826 -1226 -1822
rect -1172 -1819 -1168 -1815
rect -1130 -1826 -1126 -1822
rect -1112 -1819 -1108 -1815
rect -1070 -1811 -1066 -1807
rect -1070 -1819 -1066 -1815
rect -1088 -1833 -1084 -1829
rect -1188 -1840 -1184 -1836
rect -1146 -1840 -1142 -1836
rect -1016 -1811 -1012 -1807
rect -1046 -1826 -1042 -1822
rect -1221 -1855 -1217 -1851
rect -1204 -1855 -1200 -1851
rect -1163 -1855 -1159 -1851
rect -1121 -1855 -1117 -1851
rect -1079 -1855 -1075 -1851
rect -1038 -1855 -1034 -1851
rect -1016 -1902 -1012 -1898
rect -1225 -2029 -1221 -2025
rect -1208 -2029 -1204 -2025
rect -1168 -2029 -1164 -2025
rect -1147 -2029 -1143 -2025
rect -1257 -2085 -1253 -2081
rect -1234 -2078 -1230 -2074
rect -1283 -2092 -1279 -2088
rect -1190 -2099 -1186 -2095
rect -909 -1187 -905 -1183
rect -618 -1187 -614 -1183
rect -918 -1226 -914 -1222
rect -926 -1298 -922 -1294
rect -900 -1298 -896 -1294
rect -883 -1298 -879 -1294
rect -843 -1298 -839 -1294
rect -822 -1298 -818 -1294
rect -805 -1298 -801 -1294
rect -765 -1298 -761 -1294
rect -741 -1298 -737 -1294
rect -704 -1298 -700 -1294
rect -935 -1331 -931 -1327
rect -917 -1324 -913 -1320
rect -891 -1346 -887 -1342
rect -909 -1353 -905 -1349
rect -865 -1338 -861 -1334
rect -813 -1331 -809 -1327
rect -883 -1375 -879 -1371
rect -847 -1375 -843 -1371
rect -787 -1346 -783 -1342
rect -805 -1375 -801 -1371
rect -769 -1375 -765 -1371
rect -695 -1338 -691 -1334
rect -688 -1346 -684 -1342
rect -926 -1390 -922 -1386
rect -900 -1390 -896 -1386
rect -857 -1390 -853 -1386
rect -822 -1390 -818 -1386
rect -778 -1390 -774 -1386
rect -761 -1390 -757 -1386
rect -725 -1390 -721 -1386
rect -704 -1390 -700 -1386
rect -605 -1338 -601 -1334
rect -219 -784 -215 -780
rect -202 -784 -198 -780
rect -551 -832 -547 -828
rect -244 -832 -240 -828
rect -560 -876 -556 -872
rect -568 -1018 -564 -1014
rect -551 -1018 -547 -1014
rect -531 -1018 -527 -1014
rect -510 -1018 -506 -1014
rect -489 -1018 -485 -1014
rect -468 -1018 -464 -1014
rect -447 -1018 -443 -1014
rect -426 -1018 -422 -1014
rect -405 -1018 -401 -1014
rect -385 -1018 -381 -1014
rect -577 -1081 -573 -1077
rect -519 -1074 -515 -1070
rect -477 -1081 -473 -1077
rect -459 -1074 -455 -1070
rect -417 -1066 -413 -1062
rect -417 -1074 -413 -1070
rect -435 -1088 -431 -1084
rect -535 -1095 -531 -1091
rect -493 -1095 -489 -1091
rect -393 -1081 -389 -1077
rect -568 -1110 -564 -1106
rect -551 -1110 -547 -1106
rect -510 -1110 -506 -1106
rect -468 -1110 -464 -1106
rect -426 -1110 -422 -1106
rect -385 -1110 -381 -1106
rect -577 -1134 -573 -1130
rect -560 -1134 -556 -1130
rect -618 -1353 -614 -1349
rect -688 -1397 -684 -1393
rect -605 -1411 -601 -1407
rect -926 -1421 -922 -1417
rect -909 -1421 -905 -1417
rect -889 -1421 -885 -1417
rect -868 -1421 -864 -1417
rect -847 -1421 -843 -1417
rect -826 -1421 -822 -1417
rect -805 -1421 -801 -1417
rect -784 -1421 -780 -1417
rect -763 -1421 -759 -1417
rect -743 -1421 -739 -1417
rect -935 -1484 -931 -1480
rect -877 -1477 -873 -1473
rect -835 -1484 -831 -1480
rect -817 -1477 -813 -1473
rect -775 -1469 -771 -1465
rect -775 -1477 -771 -1473
rect -793 -1491 -789 -1487
rect -893 -1498 -889 -1494
rect -851 -1498 -847 -1494
rect -751 -1484 -747 -1480
rect -926 -1513 -922 -1509
rect -909 -1513 -905 -1509
rect -868 -1513 -864 -1509
rect -826 -1513 -822 -1509
rect -784 -1513 -780 -1509
rect -743 -1513 -739 -1509
rect -926 -1592 -922 -1588
rect -909 -1592 -905 -1588
rect -889 -1592 -885 -1588
rect -868 -1592 -864 -1588
rect -847 -1592 -843 -1588
rect -826 -1592 -822 -1588
rect -805 -1592 -801 -1588
rect -784 -1592 -780 -1588
rect -763 -1592 -759 -1588
rect -743 -1592 -739 -1588
rect -935 -1655 -931 -1651
rect -877 -1648 -873 -1644
rect -835 -1655 -831 -1651
rect -817 -1648 -813 -1644
rect -775 -1640 -771 -1636
rect -775 -1648 -771 -1644
rect -793 -1662 -789 -1658
rect -893 -1669 -889 -1665
rect -851 -1669 -847 -1665
rect -730 -1640 -726 -1636
rect -751 -1655 -747 -1651
rect -926 -1684 -922 -1680
rect -909 -1684 -905 -1680
rect -868 -1684 -864 -1680
rect -826 -1684 -822 -1680
rect -784 -1684 -780 -1680
rect -743 -1684 -739 -1680
rect -605 -1648 -601 -1644
rect -730 -1692 -726 -1688
rect -605 -1692 -601 -1688
rect -926 -1763 -922 -1759
rect -909 -1763 -905 -1759
rect -889 -1763 -885 -1759
rect -868 -1763 -864 -1759
rect -847 -1763 -843 -1759
rect -826 -1763 -822 -1759
rect -805 -1763 -801 -1759
rect -784 -1763 -780 -1759
rect -763 -1763 -759 -1759
rect -743 -1763 -739 -1759
rect -949 -1819 -945 -1815
rect -935 -1826 -931 -1822
rect -877 -1819 -873 -1815
rect -835 -1826 -831 -1822
rect -817 -1819 -813 -1815
rect -775 -1811 -771 -1807
rect -775 -1819 -771 -1815
rect -793 -1833 -789 -1829
rect -893 -1840 -889 -1836
rect -851 -1840 -847 -1836
rect -723 -1811 -719 -1807
rect -751 -1826 -747 -1822
rect -926 -1855 -922 -1851
rect -909 -1855 -905 -1851
rect -868 -1855 -864 -1851
rect -826 -1855 -822 -1851
rect -784 -1855 -780 -1851
rect -743 -1855 -739 -1851
rect -935 -1870 -931 -1866
rect -918 -1870 -914 -1866
rect -976 -2069 -972 -2065
rect -968 -1923 -964 -1919
rect -1138 -2077 -1134 -2073
rect -1208 -2106 -1204 -2102
rect -1172 -2106 -1168 -2102
rect -968 -2084 -964 -2080
rect -1115 -2099 -1111 -2095
rect -1225 -2121 -1221 -2117
rect -1181 -2121 -1177 -2117
rect -1147 -2121 -1143 -2117
rect -1257 -2128 -1253 -2124
rect -1245 -2135 -1241 -2131
rect -1115 -2135 -1111 -2131
rect -963 -2135 -959 -2131
rect -1225 -2173 -1221 -2169
rect -1208 -2173 -1204 -2169
rect -1188 -2173 -1184 -2169
rect -1167 -2173 -1163 -2169
rect -1146 -2173 -1142 -2169
rect -1125 -2173 -1121 -2169
rect -1104 -2173 -1100 -2169
rect -1083 -2173 -1079 -2169
rect -1062 -2173 -1058 -2169
rect -1042 -2173 -1038 -2169
rect -1245 -2229 -1241 -2225
rect -1234 -2236 -1230 -2232
rect -1176 -2229 -1172 -2225
rect -1134 -2236 -1130 -2232
rect -1116 -2229 -1112 -2225
rect -1074 -2221 -1070 -2217
rect -1074 -2229 -1070 -2225
rect -1092 -2243 -1088 -2239
rect -1192 -2250 -1188 -2246
rect -1150 -2250 -1146 -2246
rect -1050 -2236 -1046 -2232
rect -1225 -2265 -1221 -2261
rect -1208 -2265 -1204 -2261
rect -1167 -2265 -1163 -2261
rect -1125 -2265 -1121 -2261
rect -1083 -2265 -1079 -2261
rect -1042 -2265 -1038 -2261
rect -1225 -2344 -1221 -2340
rect -1208 -2344 -1204 -2340
rect -1188 -2344 -1184 -2340
rect -1167 -2344 -1163 -2340
rect -1146 -2344 -1142 -2340
rect -1125 -2344 -1121 -2340
rect -1104 -2344 -1100 -2340
rect -1083 -2344 -1079 -2340
rect -1062 -2344 -1058 -2340
rect -1042 -2344 -1038 -2340
rect -1257 -2400 -1253 -2396
rect -1234 -2407 -1230 -2403
rect -1176 -2400 -1172 -2396
rect -1134 -2407 -1130 -2403
rect -1116 -2400 -1112 -2396
rect -1074 -2392 -1070 -2388
rect -1074 -2400 -1070 -2396
rect -1092 -2414 -1088 -2410
rect -1192 -2421 -1188 -2417
rect -1150 -2421 -1146 -2417
rect -1024 -2392 -1020 -2388
rect -1050 -2407 -1046 -2403
rect -1225 -2436 -1221 -2432
rect -1208 -2436 -1204 -2432
rect -1167 -2436 -1163 -2432
rect -1125 -2436 -1121 -2432
rect -1083 -2436 -1079 -2432
rect -1042 -2436 -1038 -2432
rect -963 -2400 -959 -2396
rect -1319 -2571 -1315 -2567
rect -1257 -2444 -1253 -2440
rect -1024 -2444 -1020 -2440
rect -963 -2443 -959 -2439
rect -1309 -2620 -1305 -2616
rect -1292 -2620 -1288 -2616
rect -1355 -2660 -1351 -2656
rect -1550 -2898 -1546 -2894
rect -1533 -2898 -1529 -2894
rect -1513 -2898 -1509 -2894
rect -1492 -2898 -1488 -2894
rect -1471 -2898 -1467 -2894
rect -1450 -2898 -1446 -2894
rect -1429 -2898 -1425 -2894
rect -1408 -2898 -1404 -2894
rect -1387 -2898 -1383 -2894
rect -1367 -2898 -1363 -2894
rect -1559 -2961 -1555 -2957
rect -1501 -2954 -1497 -2950
rect -1459 -2961 -1455 -2957
rect -1441 -2954 -1437 -2950
rect -1399 -2946 -1395 -2942
rect -1399 -2954 -1395 -2950
rect -1417 -2968 -1413 -2964
rect -1517 -2975 -1513 -2971
rect -1475 -2975 -1471 -2971
rect -1352 -2946 -1348 -2942
rect -1375 -2961 -1371 -2957
rect -1550 -2990 -1546 -2986
rect -1533 -2990 -1529 -2986
rect -1492 -2990 -1488 -2986
rect -1450 -2990 -1446 -2986
rect -1408 -2990 -1404 -2986
rect -1367 -2990 -1363 -2986
rect -1581 -2997 -1577 -2993
rect -1352 -2997 -1348 -2993
rect -1550 -3069 -1546 -3065
rect -1533 -3069 -1529 -3065
rect -1513 -3069 -1509 -3065
rect -1492 -3069 -1488 -3065
rect -1471 -3069 -1467 -3065
rect -1450 -3069 -1446 -3065
rect -1429 -3069 -1425 -3065
rect -1408 -3069 -1404 -3065
rect -1387 -3069 -1383 -3065
rect -1367 -3069 -1363 -3065
rect -1581 -3125 -1577 -3121
rect -1559 -3132 -1555 -3128
rect -1501 -3125 -1497 -3121
rect -1459 -3132 -1455 -3128
rect -1441 -3125 -1437 -3121
rect -1399 -3117 -1395 -3113
rect -1399 -3125 -1395 -3121
rect -1417 -3139 -1413 -3135
rect -1517 -3146 -1513 -3142
rect -1475 -3146 -1471 -3142
rect -1355 -3117 -1351 -3113
rect -1375 -3132 -1371 -3128
rect -1550 -3161 -1546 -3157
rect -1533 -3161 -1529 -3157
rect -1492 -3161 -1488 -3157
rect -1450 -3161 -1446 -3157
rect -1408 -3161 -1404 -3157
rect -1367 -3161 -1363 -3157
rect -1582 -3168 -1578 -3164
rect -1355 -3168 -1351 -3164
rect -1550 -3240 -1546 -3236
rect -1533 -3240 -1529 -3236
rect -1513 -3240 -1509 -3236
rect -1492 -3240 -1488 -3236
rect -1471 -3240 -1467 -3236
rect -1450 -3240 -1446 -3236
rect -1429 -3240 -1425 -3236
rect -1408 -3240 -1404 -3236
rect -1387 -3240 -1383 -3236
rect -1367 -3240 -1363 -3236
rect -1582 -3296 -1578 -3292
rect -1559 -3303 -1555 -3299
rect -1501 -3296 -1497 -3292
rect -1459 -3303 -1455 -3299
rect -1441 -3296 -1437 -3292
rect -1399 -3288 -1395 -3284
rect -1399 -3296 -1395 -3292
rect -1417 -3310 -1413 -3306
rect -1517 -3317 -1513 -3313
rect -1475 -3317 -1471 -3313
rect -1355 -3288 -1351 -3284
rect -1375 -3303 -1371 -3299
rect -1550 -3332 -1546 -3328
rect -1533 -3332 -1529 -3328
rect -1492 -3332 -1488 -3328
rect -1450 -3332 -1446 -3328
rect -1408 -3332 -1404 -3328
rect -1367 -3332 -1363 -3328
rect -1292 -2712 -1288 -2708
rect -1225 -2515 -1221 -2511
rect -1208 -2515 -1204 -2511
rect -1188 -2515 -1184 -2511
rect -1167 -2515 -1163 -2511
rect -1146 -2515 -1142 -2511
rect -1125 -2515 -1121 -2511
rect -1104 -2515 -1100 -2511
rect -1083 -2515 -1079 -2511
rect -1062 -2515 -1058 -2511
rect -1042 -2515 -1038 -2511
rect -1234 -2578 -1230 -2574
rect -1176 -2571 -1172 -2567
rect -1134 -2578 -1130 -2574
rect -1116 -2571 -1112 -2567
rect -1074 -2563 -1070 -2559
rect -1074 -2571 -1070 -2567
rect -1092 -2585 -1088 -2581
rect -1192 -2592 -1188 -2588
rect -1150 -2592 -1146 -2588
rect -1026 -2563 -1022 -2559
rect -1050 -2578 -1046 -2574
rect -1225 -2607 -1221 -2603
rect -1208 -2607 -1204 -2603
rect -1167 -2607 -1163 -2603
rect -1125 -2607 -1121 -2603
rect -1083 -2607 -1079 -2603
rect -1042 -2607 -1038 -2603
rect -1026 -2652 -1022 -2648
rect -979 -2673 -975 -2669
rect -1225 -2779 -1221 -2775
rect -1208 -2779 -1204 -2775
rect -1168 -2779 -1164 -2775
rect -1147 -2779 -1143 -2775
rect -1257 -2835 -1253 -2831
rect -1234 -2828 -1230 -2824
rect -1283 -2842 -1279 -2838
rect -1190 -2849 -1186 -2845
rect -979 -2819 -975 -2815
rect -1138 -2827 -1134 -2823
rect -1208 -2856 -1204 -2852
rect -1172 -2856 -1168 -2852
rect -723 -1902 -719 -1898
rect -909 -1923 -905 -1919
rect -618 -1923 -614 -1919
rect -918 -1962 -914 -1958
rect -926 -2029 -922 -2025
rect -900 -2029 -896 -2025
rect -883 -2029 -879 -2025
rect -843 -2029 -839 -2025
rect -822 -2029 -818 -2025
rect -805 -2029 -801 -2025
rect -765 -2029 -761 -2025
rect -741 -2029 -737 -2025
rect -704 -2029 -700 -2025
rect -935 -2062 -931 -2058
rect -917 -2055 -913 -2051
rect -891 -2077 -887 -2073
rect -909 -2084 -905 -2080
rect -865 -2069 -861 -2065
rect -813 -2062 -809 -2058
rect -883 -2106 -879 -2102
rect -847 -2106 -843 -2102
rect -787 -2077 -783 -2073
rect -805 -2106 -801 -2102
rect -769 -2106 -765 -2102
rect -695 -2069 -691 -2065
rect -687 -2077 -683 -2073
rect -926 -2121 -922 -2117
rect -900 -2121 -896 -2117
rect -857 -2121 -853 -2117
rect -822 -2121 -818 -2117
rect -778 -2121 -774 -2117
rect -761 -2121 -757 -2117
rect -725 -2121 -721 -2117
rect -704 -2121 -700 -2117
rect -551 -1187 -547 -1183
rect -267 -1187 -263 -1183
rect -560 -1226 -556 -1222
rect -568 -1298 -564 -1294
rect -542 -1298 -538 -1294
rect -525 -1298 -521 -1294
rect -485 -1298 -481 -1294
rect -464 -1298 -460 -1294
rect -447 -1298 -443 -1294
rect -407 -1298 -403 -1294
rect -383 -1298 -379 -1294
rect -346 -1298 -342 -1294
rect -577 -1331 -573 -1327
rect -559 -1324 -555 -1320
rect -533 -1346 -529 -1342
rect -551 -1353 -547 -1349
rect -507 -1338 -503 -1334
rect -455 -1331 -451 -1327
rect -525 -1375 -521 -1371
rect -489 -1375 -485 -1371
rect -429 -1346 -425 -1342
rect -447 -1375 -443 -1371
rect -411 -1375 -407 -1371
rect -337 -1338 -333 -1334
rect -328 -1346 -324 -1342
rect -568 -1390 -564 -1386
rect -542 -1390 -538 -1386
rect -499 -1390 -495 -1386
rect -464 -1390 -460 -1386
rect -420 -1390 -416 -1386
rect -403 -1390 -399 -1386
rect -367 -1390 -363 -1386
rect -346 -1390 -342 -1386
rect -244 -1338 -240 -1334
rect 138 -784 142 -780
rect 155 -784 159 -780
rect -193 -840 -189 -836
rect 107 -840 111 -836
rect -202 -876 -198 -872
rect -210 -1018 -206 -1014
rect -193 -1018 -189 -1014
rect -173 -1018 -169 -1014
rect -152 -1018 -148 -1014
rect -131 -1018 -127 -1014
rect -110 -1018 -106 -1014
rect -89 -1018 -85 -1014
rect -68 -1018 -64 -1014
rect -47 -1018 -43 -1014
rect -27 -1018 -23 -1014
rect -219 -1081 -215 -1077
rect -161 -1074 -157 -1070
rect -119 -1081 -115 -1077
rect -101 -1074 -97 -1070
rect -59 -1066 -55 -1062
rect -59 -1074 -55 -1070
rect -77 -1088 -73 -1084
rect -177 -1095 -173 -1091
rect -135 -1095 -131 -1091
rect -35 -1081 -31 -1077
rect -210 -1110 -206 -1106
rect -193 -1110 -189 -1106
rect -152 -1110 -148 -1106
rect -110 -1110 -106 -1106
rect -68 -1110 -64 -1106
rect -27 -1110 -23 -1106
rect -219 -1134 -215 -1130
rect -202 -1134 -198 -1130
rect -267 -1353 -263 -1349
rect -328 -1404 -324 -1400
rect -244 -1404 -240 -1400
rect -568 -1421 -564 -1417
rect -551 -1421 -547 -1417
rect -531 -1421 -527 -1417
rect -510 -1421 -506 -1417
rect -489 -1421 -485 -1417
rect -468 -1421 -464 -1417
rect -447 -1421 -443 -1417
rect -426 -1421 -422 -1417
rect -405 -1421 -401 -1417
rect -385 -1421 -381 -1417
rect -577 -1484 -573 -1480
rect -519 -1477 -515 -1473
rect -477 -1484 -473 -1480
rect -459 -1477 -455 -1473
rect -417 -1469 -413 -1465
rect -417 -1477 -413 -1473
rect -435 -1491 -431 -1487
rect -535 -1498 -531 -1494
rect -493 -1498 -489 -1494
rect -393 -1484 -389 -1480
rect -568 -1513 -564 -1509
rect -551 -1513 -547 -1509
rect -510 -1513 -506 -1509
rect -468 -1513 -464 -1509
rect -426 -1513 -422 -1509
rect -385 -1513 -381 -1509
rect -568 -1592 -564 -1588
rect -551 -1592 -547 -1588
rect -531 -1592 -527 -1588
rect -510 -1592 -506 -1588
rect -489 -1592 -485 -1588
rect -468 -1592 -464 -1588
rect -447 -1592 -443 -1588
rect -426 -1592 -422 -1588
rect -405 -1592 -401 -1588
rect -385 -1592 -381 -1588
rect -577 -1655 -573 -1651
rect -519 -1648 -515 -1644
rect -477 -1655 -473 -1651
rect -459 -1648 -455 -1644
rect -417 -1640 -413 -1636
rect -417 -1648 -413 -1644
rect -435 -1662 -431 -1658
rect -535 -1669 -531 -1665
rect -493 -1669 -489 -1665
rect -368 -1640 -364 -1636
rect -393 -1655 -389 -1651
rect -568 -1684 -564 -1680
rect -551 -1684 -547 -1680
rect -510 -1684 -506 -1680
rect -468 -1684 -464 -1680
rect -426 -1684 -422 -1680
rect -385 -1684 -381 -1680
rect -244 -1648 -240 -1644
rect -368 -1692 -364 -1688
rect -244 -1691 -240 -1687
rect -568 -1763 -564 -1759
rect -551 -1763 -547 -1759
rect -531 -1763 -527 -1759
rect -510 -1763 -506 -1759
rect -489 -1763 -485 -1759
rect -468 -1763 -464 -1759
rect -447 -1763 -443 -1759
rect -426 -1763 -422 -1759
rect -405 -1763 -401 -1759
rect -385 -1763 -381 -1759
rect -591 -1819 -587 -1815
rect -577 -1826 -573 -1822
rect -519 -1819 -515 -1815
rect -477 -1826 -473 -1822
rect -459 -1819 -455 -1815
rect -417 -1811 -413 -1807
rect -417 -1819 -413 -1815
rect -435 -1833 -431 -1829
rect -535 -1840 -531 -1836
rect -493 -1840 -489 -1836
rect -366 -1811 -362 -1807
rect -393 -1826 -389 -1822
rect -568 -1855 -564 -1851
rect -551 -1855 -547 -1851
rect -510 -1855 -506 -1851
rect -468 -1855 -464 -1851
rect -426 -1855 -422 -1851
rect -385 -1855 -381 -1851
rect -577 -1870 -573 -1866
rect -560 -1870 -556 -1866
rect -605 -2069 -601 -2065
rect -618 -2084 -614 -2080
rect -687 -2128 -683 -2124
rect -603 -2128 -599 -2124
rect -926 -2173 -922 -2169
rect -909 -2173 -905 -2169
rect -889 -2173 -885 -2169
rect -868 -2173 -864 -2169
rect -847 -2173 -843 -2169
rect -826 -2173 -822 -2169
rect -805 -2173 -801 -2169
rect -784 -2173 -780 -2169
rect -763 -2173 -759 -2169
rect -743 -2173 -739 -2169
rect -935 -2236 -931 -2232
rect -877 -2229 -873 -2225
rect -835 -2236 -831 -2232
rect -817 -2229 -813 -2225
rect -775 -2221 -771 -2217
rect -775 -2229 -771 -2225
rect -793 -2243 -789 -2239
rect -893 -2250 -889 -2246
rect -851 -2250 -847 -2246
rect -751 -2236 -747 -2232
rect -926 -2265 -922 -2261
rect -909 -2265 -905 -2261
rect -868 -2265 -864 -2261
rect -826 -2265 -822 -2261
rect -784 -2265 -780 -2261
rect -743 -2265 -739 -2261
rect -926 -2344 -922 -2340
rect -909 -2344 -905 -2340
rect -889 -2344 -885 -2340
rect -868 -2344 -864 -2340
rect -847 -2344 -843 -2340
rect -826 -2344 -822 -2340
rect -805 -2344 -801 -2340
rect -784 -2344 -780 -2340
rect -763 -2344 -759 -2340
rect -743 -2344 -739 -2340
rect -935 -2407 -931 -2403
rect -877 -2400 -873 -2396
rect -835 -2407 -831 -2403
rect -817 -2400 -813 -2396
rect -775 -2392 -771 -2388
rect -775 -2400 -771 -2396
rect -793 -2414 -789 -2410
rect -893 -2421 -889 -2417
rect -851 -2421 -847 -2417
rect -723 -2392 -719 -2388
rect -751 -2407 -747 -2403
rect -926 -2436 -922 -2432
rect -909 -2436 -905 -2432
rect -868 -2436 -864 -2432
rect -826 -2436 -822 -2432
rect -784 -2436 -780 -2432
rect -743 -2436 -739 -2432
rect -603 -2400 -599 -2396
rect -723 -2443 -719 -2439
rect -603 -2444 -599 -2440
rect -926 -2515 -922 -2511
rect -909 -2515 -905 -2511
rect -889 -2515 -885 -2511
rect -868 -2515 -864 -2511
rect -847 -2515 -843 -2511
rect -826 -2515 -822 -2511
rect -805 -2515 -801 -2511
rect -784 -2515 -780 -2511
rect -763 -2515 -759 -2511
rect -743 -2515 -739 -2511
rect -949 -2571 -945 -2567
rect -935 -2578 -931 -2574
rect -877 -2571 -873 -2567
rect -835 -2578 -831 -2574
rect -817 -2571 -813 -2567
rect -775 -2563 -771 -2559
rect -775 -2571 -771 -2567
rect -793 -2585 -789 -2581
rect -893 -2592 -889 -2588
rect -851 -2592 -847 -2588
rect -720 -2563 -716 -2559
rect -751 -2578 -747 -2574
rect -926 -2607 -922 -2603
rect -909 -2607 -905 -2603
rect -868 -2607 -864 -2603
rect -826 -2607 -822 -2603
rect -784 -2607 -780 -2603
rect -743 -2607 -739 -2603
rect -935 -2620 -931 -2616
rect -918 -2620 -914 -2616
rect -963 -2834 -959 -2830
rect -1117 -2849 -1113 -2845
rect -1225 -2871 -1221 -2867
rect -1181 -2871 -1177 -2867
rect -1147 -2871 -1143 -2867
rect -1257 -2878 -1253 -2874
rect -1246 -2886 -1242 -2882
rect -1117 -2886 -1113 -2882
rect -963 -2885 -959 -2881
rect -1225 -2898 -1221 -2894
rect -1208 -2898 -1204 -2894
rect -1188 -2898 -1184 -2894
rect -1167 -2898 -1163 -2894
rect -1146 -2898 -1142 -2894
rect -1125 -2898 -1121 -2894
rect -1104 -2898 -1100 -2894
rect -1083 -2898 -1079 -2894
rect -1062 -2898 -1058 -2894
rect -1042 -2898 -1038 -2894
rect -1246 -2954 -1242 -2950
rect -1234 -2961 -1230 -2957
rect -1176 -2954 -1172 -2950
rect -1134 -2961 -1130 -2957
rect -1116 -2954 -1112 -2950
rect -1074 -2946 -1070 -2942
rect -1074 -2954 -1070 -2950
rect -1092 -2968 -1088 -2964
rect -1192 -2975 -1188 -2971
rect -1150 -2975 -1146 -2971
rect -1050 -2961 -1046 -2957
rect -1225 -2990 -1221 -2986
rect -1208 -2990 -1204 -2986
rect -1167 -2990 -1163 -2986
rect -1125 -2990 -1121 -2986
rect -1083 -2990 -1079 -2986
rect -1042 -2990 -1038 -2986
rect -1225 -3069 -1221 -3065
rect -1208 -3069 -1204 -3065
rect -1188 -3069 -1184 -3065
rect -1167 -3069 -1163 -3065
rect -1146 -3069 -1142 -3065
rect -1125 -3069 -1121 -3065
rect -1104 -3069 -1100 -3065
rect -1083 -3069 -1079 -3065
rect -1062 -3069 -1058 -3065
rect -1042 -3069 -1038 -3065
rect -1257 -3125 -1253 -3121
rect -1234 -3132 -1230 -3128
rect -1176 -3125 -1172 -3121
rect -1134 -3132 -1130 -3128
rect -1116 -3125 -1112 -3121
rect -1074 -3117 -1070 -3113
rect -1074 -3125 -1070 -3121
rect -1092 -3139 -1088 -3135
rect -1192 -3146 -1188 -3142
rect -1150 -3146 -1146 -3142
rect -1026 -3117 -1022 -3113
rect -1050 -3132 -1046 -3128
rect -1225 -3161 -1221 -3157
rect -1208 -3161 -1204 -3157
rect -1167 -3161 -1163 -3157
rect -1125 -3161 -1121 -3157
rect -1083 -3161 -1079 -3157
rect -1042 -3161 -1038 -3157
rect -963 -3125 -959 -3121
rect -1319 -3296 -1315 -3292
rect -1257 -3169 -1253 -3165
rect -1026 -3169 -1022 -3165
rect -963 -3169 -959 -3165
rect -1309 -3351 -1305 -3347
rect -1292 -3351 -1288 -3347
rect -1355 -3391 -1351 -3387
rect -1813 -3640 -1809 -3636
rect -1796 -3640 -1792 -3636
rect -1776 -3640 -1772 -3636
rect -1755 -3640 -1751 -3636
rect -1734 -3640 -1730 -3636
rect -1713 -3640 -1709 -3636
rect -1692 -3640 -1688 -3636
rect -1671 -3640 -1667 -3636
rect -1650 -3640 -1646 -3636
rect -1630 -3640 -1626 -3636
rect -1550 -3640 -1546 -3636
rect -1533 -3640 -1529 -3636
rect -1513 -3640 -1509 -3636
rect -1492 -3640 -1488 -3636
rect -1471 -3640 -1467 -3636
rect -1450 -3640 -1446 -3636
rect -1429 -3640 -1425 -3636
rect -1408 -3640 -1404 -3636
rect -1387 -3640 -1383 -3636
rect -1367 -3640 -1363 -3636
rect -1822 -3703 -1818 -3699
rect -1764 -3696 -1760 -3692
rect -1722 -3703 -1718 -3699
rect -1704 -3696 -1700 -3692
rect -1662 -3688 -1658 -3684
rect -1662 -3696 -1658 -3692
rect -1680 -3710 -1676 -3706
rect -1780 -3717 -1776 -3713
rect -1738 -3717 -1734 -3713
rect -1638 -3703 -1634 -3699
rect -1559 -3703 -1555 -3699
rect -1501 -3696 -1497 -3692
rect -1459 -3703 -1455 -3699
rect -1441 -3696 -1437 -3692
rect -1399 -3688 -1395 -3684
rect -1399 -3696 -1395 -3692
rect -1417 -3710 -1413 -3706
rect -1517 -3717 -1513 -3713
rect -1475 -3717 -1471 -3713
rect -1353 -3688 -1349 -3684
rect -1375 -3703 -1371 -3699
rect -1813 -3732 -1809 -3728
rect -1796 -3732 -1792 -3728
rect -1755 -3732 -1751 -3728
rect -1713 -3732 -1709 -3728
rect -1671 -3732 -1667 -3728
rect -1630 -3732 -1626 -3728
rect -1550 -3732 -1546 -3728
rect -1533 -3732 -1529 -3728
rect -1492 -3732 -1488 -3728
rect -1450 -3732 -1446 -3728
rect -1408 -3732 -1404 -3728
rect -1367 -3732 -1363 -3728
rect -1572 -3740 -1568 -3736
rect -1353 -3740 -1349 -3736
rect -1550 -3811 -1546 -3807
rect -1533 -3811 -1529 -3807
rect -1513 -3811 -1509 -3807
rect -1492 -3811 -1488 -3807
rect -1471 -3811 -1467 -3807
rect -1450 -3811 -1446 -3807
rect -1429 -3811 -1425 -3807
rect -1408 -3811 -1404 -3807
rect -1387 -3811 -1383 -3807
rect -1367 -3811 -1363 -3807
rect -1572 -3867 -1568 -3863
rect -1559 -3874 -1555 -3870
rect -1501 -3867 -1497 -3863
rect -1459 -3874 -1455 -3870
rect -1441 -3867 -1437 -3863
rect -1399 -3859 -1395 -3855
rect -1399 -3867 -1395 -3863
rect -1417 -3881 -1413 -3877
rect -1517 -3888 -1513 -3884
rect -1475 -3888 -1471 -3884
rect -1355 -3859 -1351 -3855
rect -1375 -3874 -1371 -3870
rect -1550 -3903 -1546 -3899
rect -1533 -3903 -1529 -3899
rect -1492 -3903 -1488 -3899
rect -1450 -3903 -1446 -3899
rect -1408 -3903 -1404 -3899
rect -1367 -3903 -1363 -3899
rect -1575 -3911 -1571 -3907
rect -1355 -3911 -1351 -3907
rect -1550 -3986 -1546 -3982
rect -1533 -3986 -1529 -3982
rect -1513 -3986 -1509 -3982
rect -1492 -3986 -1488 -3982
rect -1471 -3986 -1467 -3982
rect -1450 -3986 -1446 -3982
rect -1429 -3986 -1425 -3982
rect -1408 -3986 -1404 -3982
rect -1387 -3986 -1383 -3982
rect -1367 -3986 -1363 -3982
rect -1575 -4042 -1571 -4038
rect -1559 -4049 -1555 -4045
rect -1501 -4042 -1497 -4038
rect -1459 -4049 -1455 -4045
rect -1441 -4042 -1437 -4038
rect -1399 -4034 -1395 -4030
rect -1399 -4042 -1395 -4038
rect -1417 -4056 -1413 -4052
rect -1517 -4063 -1513 -4059
rect -1475 -4063 -1471 -4059
rect -1357 -4034 -1353 -4030
rect -1375 -4049 -1371 -4045
rect -1550 -4078 -1546 -4074
rect -1533 -4078 -1529 -4074
rect -1492 -4078 -1488 -4074
rect -1450 -4078 -1446 -4074
rect -1408 -4078 -1404 -4074
rect -1367 -4078 -1363 -4074
rect -1292 -3443 -1288 -3439
rect -1225 -3240 -1221 -3236
rect -1208 -3240 -1204 -3236
rect -1188 -3240 -1184 -3236
rect -1167 -3240 -1163 -3236
rect -1146 -3240 -1142 -3236
rect -1125 -3240 -1121 -3236
rect -1104 -3240 -1100 -3236
rect -1083 -3240 -1079 -3236
rect -1062 -3240 -1058 -3236
rect -1042 -3240 -1038 -3236
rect -1234 -3303 -1230 -3299
rect -1176 -3296 -1172 -3292
rect -1134 -3303 -1130 -3299
rect -1116 -3296 -1112 -3292
rect -1074 -3288 -1070 -3284
rect -1074 -3296 -1070 -3292
rect -1092 -3310 -1088 -3306
rect -1192 -3317 -1188 -3313
rect -1150 -3317 -1146 -3313
rect -1026 -3288 -1022 -3284
rect -1050 -3303 -1046 -3299
rect -1225 -3332 -1221 -3328
rect -1208 -3332 -1204 -3328
rect -1167 -3332 -1163 -3328
rect -1125 -3332 -1121 -3328
rect -1083 -3332 -1079 -3328
rect -1042 -3332 -1038 -3328
rect -1026 -3383 -1022 -3379
rect -979 -3404 -975 -3400
rect -1225 -3510 -1221 -3506
rect -1208 -3510 -1204 -3506
rect -1168 -3510 -1164 -3506
rect -1147 -3510 -1143 -3506
rect -1257 -3566 -1253 -3562
rect -1234 -3559 -1230 -3555
rect -1283 -3573 -1279 -3569
rect -1190 -3580 -1186 -3576
rect -979 -3550 -975 -3546
rect -1138 -3558 -1134 -3554
rect -1208 -3587 -1204 -3583
rect -1172 -3587 -1168 -3583
rect -720 -2652 -716 -2648
rect -909 -2673 -905 -2669
rect -616 -2673 -612 -2669
rect -918 -2712 -914 -2708
rect -926 -2779 -922 -2775
rect -900 -2779 -896 -2775
rect -883 -2779 -879 -2775
rect -843 -2779 -839 -2775
rect -822 -2779 -818 -2775
rect -805 -2779 -801 -2775
rect -765 -2779 -761 -2775
rect -741 -2779 -737 -2775
rect -704 -2779 -700 -2775
rect -935 -2812 -931 -2808
rect -917 -2805 -913 -2801
rect -891 -2827 -887 -2823
rect -909 -2834 -905 -2830
rect -865 -2819 -861 -2815
rect -813 -2812 -809 -2808
rect -883 -2856 -879 -2852
rect -847 -2856 -843 -2852
rect -787 -2827 -783 -2823
rect -805 -2856 -801 -2852
rect -769 -2856 -765 -2852
rect -695 -2819 -691 -2815
rect -688 -2827 -684 -2823
rect -926 -2871 -922 -2867
rect -900 -2871 -896 -2867
rect -857 -2871 -853 -2867
rect -822 -2871 -818 -2867
rect -778 -2871 -774 -2867
rect -761 -2871 -757 -2867
rect -725 -2871 -721 -2867
rect -704 -2871 -700 -2867
rect -366 -1902 -362 -1898
rect -551 -1923 -547 -1919
rect -262 -1923 -258 -1919
rect -560 -1962 -556 -1958
rect -568 -2029 -564 -2025
rect -542 -2029 -538 -2025
rect -525 -2029 -521 -2025
rect -485 -2029 -481 -2025
rect -464 -2029 -460 -2025
rect -447 -2029 -443 -2025
rect -407 -2029 -403 -2025
rect -383 -2029 -379 -2025
rect -346 -2029 -342 -2025
rect -577 -2062 -573 -2058
rect -559 -2055 -555 -2051
rect -533 -2077 -529 -2073
rect -551 -2084 -547 -2080
rect -507 -2069 -503 -2065
rect -455 -2062 -451 -2058
rect -525 -2106 -521 -2102
rect -489 -2106 -485 -2102
rect -429 -2077 -425 -2073
rect -447 -2106 -443 -2102
rect -411 -2106 -407 -2102
rect -337 -2066 -333 -2062
rect -328 -2077 -324 -2073
rect -568 -2121 -564 -2117
rect -542 -2121 -538 -2117
rect -499 -2121 -495 -2117
rect -464 -2121 -460 -2117
rect -420 -2121 -416 -2117
rect -403 -2121 -399 -2117
rect -367 -2121 -363 -2117
rect -346 -2121 -342 -2117
rect -193 -1187 -189 -1183
rect 91 -1187 95 -1183
rect -202 -1226 -198 -1222
rect -210 -1298 -206 -1294
rect -184 -1298 -180 -1294
rect -167 -1298 -163 -1294
rect -127 -1298 -123 -1294
rect -106 -1298 -102 -1294
rect -89 -1298 -85 -1294
rect -49 -1298 -45 -1294
rect -25 -1298 -21 -1294
rect 12 -1298 16 -1294
rect -219 -1331 -215 -1327
rect -201 -1324 -197 -1320
rect -175 -1346 -171 -1342
rect -193 -1353 -189 -1349
rect -149 -1338 -145 -1334
rect -97 -1331 -93 -1327
rect -167 -1375 -163 -1371
rect -131 -1375 -127 -1371
rect -71 -1346 -67 -1342
rect -89 -1375 -85 -1371
rect -53 -1375 -49 -1371
rect 21 -1338 25 -1334
rect 29 -1346 33 -1342
rect -210 -1390 -206 -1386
rect -184 -1390 -180 -1386
rect -141 -1390 -137 -1386
rect -106 -1390 -102 -1386
rect -62 -1390 -58 -1386
rect -45 -1390 -41 -1386
rect -9 -1390 -5 -1386
rect 12 -1390 16 -1386
rect 107 -1338 111 -1334
rect 495 -784 499 -780
rect 512 -784 516 -780
rect 164 -832 168 -828
rect 470 -832 474 -828
rect 155 -876 159 -872
rect 148 -1018 152 -1014
rect 165 -1018 169 -1014
rect 185 -1018 189 -1014
rect 206 -1018 210 -1014
rect 227 -1018 231 -1014
rect 248 -1018 252 -1014
rect 269 -1018 273 -1014
rect 290 -1018 294 -1014
rect 311 -1018 315 -1014
rect 331 -1018 335 -1014
rect 139 -1081 143 -1077
rect 197 -1074 201 -1070
rect 239 -1081 243 -1077
rect 257 -1074 261 -1070
rect 299 -1066 303 -1062
rect 299 -1074 303 -1070
rect 281 -1088 285 -1084
rect 181 -1095 185 -1091
rect 223 -1095 227 -1091
rect 323 -1081 327 -1077
rect 148 -1110 152 -1106
rect 165 -1110 169 -1106
rect 206 -1110 210 -1106
rect 248 -1110 252 -1106
rect 290 -1110 294 -1106
rect 331 -1110 335 -1106
rect 139 -1134 143 -1130
rect 156 -1134 160 -1130
rect 91 -1353 95 -1349
rect 29 -1411 33 -1407
rect 107 -1411 111 -1407
rect -210 -1421 -206 -1417
rect -193 -1421 -189 -1417
rect -173 -1421 -169 -1417
rect -152 -1421 -148 -1417
rect -131 -1421 -127 -1417
rect -110 -1421 -106 -1417
rect -89 -1421 -85 -1417
rect -68 -1421 -64 -1417
rect -47 -1421 -43 -1417
rect -27 -1421 -23 -1417
rect -219 -1484 -215 -1480
rect -161 -1477 -157 -1473
rect -119 -1484 -115 -1480
rect -101 -1477 -97 -1473
rect -59 -1469 -55 -1465
rect -59 -1477 -55 -1473
rect -77 -1491 -73 -1487
rect -177 -1498 -173 -1494
rect -135 -1498 -131 -1494
rect -35 -1484 -31 -1480
rect -210 -1513 -206 -1509
rect -193 -1513 -189 -1509
rect -152 -1513 -148 -1509
rect -110 -1513 -106 -1509
rect -68 -1513 -64 -1509
rect -27 -1513 -23 -1509
rect -210 -1592 -206 -1588
rect -193 -1592 -189 -1588
rect -173 -1592 -169 -1588
rect -152 -1592 -148 -1588
rect -131 -1592 -127 -1588
rect -110 -1592 -106 -1588
rect -89 -1592 -85 -1588
rect -68 -1592 -64 -1588
rect -47 -1592 -43 -1588
rect -27 -1592 -23 -1588
rect -219 -1655 -215 -1651
rect -161 -1648 -157 -1644
rect -119 -1655 -115 -1651
rect -101 -1648 -97 -1644
rect -59 -1640 -55 -1636
rect -59 -1648 -55 -1644
rect -77 -1662 -73 -1658
rect -177 -1669 -173 -1665
rect -135 -1669 -131 -1665
rect -12 -1640 -8 -1636
rect -35 -1655 -31 -1651
rect -210 -1684 -206 -1680
rect -193 -1684 -189 -1680
rect -152 -1684 -148 -1680
rect -110 -1684 -106 -1680
rect -68 -1684 -64 -1680
rect -27 -1684 -23 -1680
rect 107 -1648 111 -1644
rect -12 -1691 -8 -1687
rect 107 -1692 111 -1688
rect -210 -1763 -206 -1759
rect -193 -1763 -189 -1759
rect -173 -1763 -169 -1759
rect -152 -1763 -148 -1759
rect -131 -1763 -127 -1759
rect -110 -1763 -106 -1759
rect -89 -1763 -85 -1759
rect -68 -1763 -64 -1759
rect -47 -1763 -43 -1759
rect -27 -1763 -23 -1759
rect -233 -1819 -229 -1815
rect -219 -1826 -215 -1822
rect -161 -1819 -157 -1815
rect -119 -1826 -115 -1822
rect -101 -1819 -97 -1815
rect -59 -1811 -55 -1807
rect -59 -1819 -55 -1815
rect -77 -1833 -73 -1829
rect -177 -1840 -173 -1836
rect -135 -1840 -131 -1836
rect -9 -1811 -5 -1807
rect -35 -1826 -31 -1822
rect -210 -1855 -206 -1851
rect -193 -1855 -189 -1851
rect -152 -1855 -148 -1851
rect -110 -1855 -106 -1851
rect -68 -1855 -64 -1851
rect -27 -1855 -23 -1851
rect -219 -1870 -215 -1866
rect -202 -1870 -198 -1866
rect -244 -2069 -240 -2065
rect -262 -2084 -258 -2080
rect -328 -2135 -324 -2131
rect -249 -2135 -245 -2131
rect -568 -2173 -564 -2169
rect -551 -2173 -547 -2169
rect -531 -2173 -527 -2169
rect -510 -2173 -506 -2169
rect -489 -2173 -485 -2169
rect -468 -2173 -464 -2169
rect -447 -2173 -443 -2169
rect -426 -2173 -422 -2169
rect -405 -2173 -401 -2169
rect -385 -2173 -381 -2169
rect -577 -2236 -573 -2232
rect -519 -2229 -515 -2225
rect -477 -2236 -473 -2232
rect -459 -2229 -455 -2225
rect -417 -2221 -413 -2217
rect -417 -2229 -413 -2225
rect -435 -2243 -431 -2239
rect -535 -2250 -531 -2246
rect -493 -2250 -489 -2246
rect -393 -2236 -389 -2232
rect -568 -2265 -564 -2261
rect -551 -2265 -547 -2261
rect -510 -2265 -506 -2261
rect -468 -2265 -464 -2261
rect -426 -2265 -422 -2261
rect -385 -2265 -381 -2261
rect -568 -2344 -564 -2340
rect -551 -2344 -547 -2340
rect -531 -2344 -527 -2340
rect -510 -2344 -506 -2340
rect -489 -2344 -485 -2340
rect -468 -2344 -464 -2340
rect -447 -2344 -443 -2340
rect -426 -2344 -422 -2340
rect -405 -2344 -401 -2340
rect -385 -2344 -381 -2340
rect -577 -2407 -573 -2403
rect -519 -2400 -515 -2396
rect -477 -2407 -473 -2403
rect -459 -2400 -455 -2396
rect -417 -2392 -413 -2388
rect -417 -2400 -413 -2396
rect -435 -2414 -431 -2410
rect -535 -2421 -531 -2417
rect -493 -2421 -489 -2417
rect -366 -2392 -362 -2388
rect -393 -2407 -389 -2403
rect -568 -2436 -564 -2432
rect -551 -2436 -547 -2432
rect -510 -2436 -506 -2432
rect -468 -2436 -464 -2432
rect -426 -2436 -422 -2432
rect -385 -2436 -381 -2432
rect -249 -2400 -245 -2396
rect -366 -2444 -362 -2440
rect -249 -2444 -245 -2440
rect -568 -2515 -564 -2511
rect -551 -2515 -547 -2511
rect -531 -2515 -527 -2511
rect -510 -2515 -506 -2511
rect -489 -2515 -485 -2511
rect -468 -2515 -464 -2511
rect -447 -2515 -443 -2511
rect -426 -2515 -422 -2511
rect -405 -2515 -401 -2511
rect -385 -2515 -381 -2511
rect -591 -2571 -587 -2567
rect -577 -2578 -573 -2574
rect -519 -2571 -515 -2567
rect -477 -2578 -473 -2574
rect -459 -2571 -455 -2567
rect -417 -2563 -413 -2559
rect -417 -2571 -413 -2567
rect -435 -2585 -431 -2581
rect -535 -2592 -531 -2588
rect -493 -2592 -489 -2588
rect -373 -2563 -369 -2559
rect -393 -2578 -389 -2574
rect -568 -2607 -564 -2603
rect -551 -2607 -547 -2603
rect -510 -2607 -506 -2603
rect -468 -2607 -464 -2603
rect -426 -2607 -422 -2603
rect -385 -2607 -381 -2603
rect -577 -2620 -573 -2616
rect -560 -2620 -556 -2616
rect -603 -2819 -599 -2815
rect -616 -2834 -612 -2830
rect -688 -2878 -684 -2874
rect -603 -2878 -599 -2874
rect -926 -2898 -922 -2894
rect -909 -2898 -905 -2894
rect -889 -2898 -885 -2894
rect -868 -2898 -864 -2894
rect -847 -2898 -843 -2894
rect -826 -2898 -822 -2894
rect -805 -2898 -801 -2894
rect -784 -2898 -780 -2894
rect -763 -2898 -759 -2894
rect -743 -2898 -739 -2894
rect -935 -2961 -931 -2957
rect -877 -2954 -873 -2950
rect -835 -2961 -831 -2957
rect -817 -2954 -813 -2950
rect -775 -2946 -771 -2942
rect -775 -2954 -771 -2950
rect -793 -2968 -789 -2964
rect -893 -2975 -889 -2971
rect -851 -2975 -847 -2971
rect -751 -2961 -747 -2957
rect -926 -2990 -922 -2986
rect -909 -2990 -905 -2986
rect -868 -2990 -864 -2986
rect -826 -2990 -822 -2986
rect -784 -2990 -780 -2986
rect -743 -2990 -739 -2986
rect -926 -3069 -922 -3065
rect -909 -3069 -905 -3065
rect -889 -3069 -885 -3065
rect -868 -3069 -864 -3065
rect -847 -3069 -843 -3065
rect -826 -3069 -822 -3065
rect -805 -3069 -801 -3065
rect -784 -3069 -780 -3065
rect -763 -3069 -759 -3065
rect -743 -3069 -739 -3065
rect -935 -3132 -931 -3128
rect -877 -3125 -873 -3121
rect -835 -3132 -831 -3128
rect -817 -3125 -813 -3121
rect -775 -3117 -771 -3113
rect -775 -3125 -771 -3121
rect -793 -3139 -789 -3135
rect -893 -3146 -889 -3142
rect -851 -3146 -847 -3142
rect -725 -3117 -721 -3113
rect -751 -3132 -747 -3128
rect -926 -3161 -922 -3157
rect -909 -3161 -905 -3157
rect -868 -3161 -864 -3157
rect -826 -3161 -822 -3157
rect -784 -3161 -780 -3157
rect -743 -3161 -739 -3157
rect -603 -3125 -599 -3121
rect -725 -3169 -721 -3165
rect -603 -3168 -599 -3164
rect -926 -3240 -922 -3236
rect -909 -3240 -905 -3236
rect -889 -3240 -885 -3236
rect -868 -3240 -864 -3236
rect -847 -3240 -843 -3236
rect -826 -3240 -822 -3236
rect -805 -3240 -801 -3236
rect -784 -3240 -780 -3236
rect -763 -3240 -759 -3236
rect -743 -3240 -739 -3236
rect -949 -3296 -945 -3292
rect -935 -3303 -931 -3299
rect -877 -3296 -873 -3292
rect -835 -3303 -831 -3299
rect -817 -3296 -813 -3292
rect -775 -3288 -771 -3284
rect -775 -3296 -771 -3292
rect -793 -3310 -789 -3306
rect -893 -3317 -889 -3313
rect -851 -3317 -847 -3313
rect -722 -3288 -718 -3284
rect -751 -3303 -747 -3299
rect -926 -3332 -922 -3328
rect -909 -3332 -905 -3328
rect -868 -3332 -864 -3328
rect -826 -3332 -822 -3328
rect -784 -3332 -780 -3328
rect -743 -3332 -739 -3328
rect -935 -3351 -931 -3347
rect -918 -3351 -914 -3347
rect -963 -3565 -959 -3561
rect -1113 -3580 -1109 -3576
rect -1225 -3602 -1221 -3598
rect -1181 -3602 -1177 -3598
rect -1147 -3602 -1143 -3598
rect -1257 -3609 -1253 -3605
rect -1246 -3616 -1242 -3612
rect -1113 -3616 -1109 -3612
rect -963 -3616 -959 -3612
rect -1225 -3640 -1221 -3636
rect -1208 -3640 -1204 -3636
rect -1188 -3640 -1184 -3636
rect -1167 -3640 -1163 -3636
rect -1146 -3640 -1142 -3636
rect -1125 -3640 -1121 -3636
rect -1104 -3640 -1100 -3636
rect -1083 -3640 -1079 -3636
rect -1062 -3640 -1058 -3636
rect -1042 -3640 -1038 -3636
rect -1246 -3696 -1242 -3692
rect -1234 -3703 -1230 -3699
rect -1176 -3696 -1172 -3692
rect -1134 -3703 -1130 -3699
rect -1116 -3696 -1112 -3692
rect -1074 -3688 -1070 -3684
rect -1074 -3696 -1070 -3692
rect -1092 -3710 -1088 -3706
rect -1192 -3717 -1188 -3713
rect -1150 -3717 -1146 -3713
rect -1050 -3703 -1046 -3699
rect -1225 -3732 -1221 -3728
rect -1208 -3732 -1204 -3728
rect -1167 -3732 -1163 -3728
rect -1125 -3732 -1121 -3728
rect -1083 -3732 -1079 -3728
rect -1042 -3732 -1038 -3728
rect -1225 -3811 -1221 -3807
rect -1208 -3811 -1204 -3807
rect -1188 -3811 -1184 -3807
rect -1167 -3811 -1163 -3807
rect -1146 -3811 -1142 -3807
rect -1125 -3811 -1121 -3807
rect -1104 -3811 -1100 -3807
rect -1083 -3811 -1079 -3807
rect -1062 -3811 -1058 -3807
rect -1042 -3811 -1038 -3807
rect -1257 -3867 -1253 -3863
rect -1234 -3874 -1230 -3870
rect -1176 -3867 -1172 -3863
rect -1134 -3874 -1130 -3870
rect -1116 -3867 -1112 -3863
rect -1074 -3859 -1070 -3855
rect -1074 -3867 -1070 -3863
rect -1092 -3881 -1088 -3877
rect -1192 -3888 -1188 -3884
rect -1150 -3888 -1146 -3884
rect -1028 -3859 -1024 -3855
rect -1050 -3874 -1046 -3870
rect -1225 -3903 -1221 -3899
rect -1208 -3903 -1204 -3899
rect -1167 -3903 -1163 -3899
rect -1125 -3903 -1121 -3899
rect -1083 -3903 -1079 -3899
rect -1042 -3903 -1038 -3899
rect -963 -3867 -959 -3863
rect -1319 -4042 -1315 -4038
rect -1257 -3910 -1253 -3906
rect -1028 -3910 -1024 -3906
rect -1309 -4101 -1305 -4097
rect -1292 -4101 -1288 -4097
rect -1357 -4141 -1353 -4137
rect -1805 -4383 -1801 -4379
rect -1788 -4383 -1784 -4379
rect -1768 -4383 -1764 -4379
rect -1747 -4383 -1743 -4379
rect -1726 -4383 -1722 -4379
rect -1705 -4383 -1701 -4379
rect -1684 -4383 -1680 -4379
rect -1663 -4383 -1659 -4379
rect -1642 -4383 -1638 -4379
rect -1622 -4383 -1618 -4379
rect -1542 -4383 -1538 -4379
rect -1525 -4383 -1521 -4379
rect -1505 -4383 -1501 -4379
rect -1484 -4383 -1480 -4379
rect -1463 -4383 -1459 -4379
rect -1442 -4383 -1438 -4379
rect -1421 -4383 -1417 -4379
rect -1400 -4383 -1396 -4379
rect -1379 -4383 -1375 -4379
rect -1359 -4383 -1355 -4379
rect -1814 -4446 -1810 -4442
rect -1756 -4439 -1752 -4435
rect -1714 -4446 -1710 -4442
rect -1696 -4439 -1692 -4435
rect -1654 -4431 -1650 -4427
rect -1654 -4439 -1650 -4435
rect -1672 -4453 -1668 -4449
rect -1772 -4460 -1768 -4456
rect -1730 -4460 -1726 -4456
rect -1630 -4446 -1626 -4442
rect -1551 -4446 -1547 -4442
rect -1493 -4439 -1489 -4435
rect -1451 -4446 -1447 -4442
rect -1433 -4439 -1429 -4435
rect -1391 -4431 -1387 -4427
rect -1391 -4439 -1387 -4435
rect -1409 -4453 -1405 -4449
rect -1509 -4460 -1505 -4456
rect -1467 -4460 -1463 -4456
rect -1346 -4431 -1342 -4427
rect -1367 -4446 -1363 -4442
rect -1805 -4475 -1801 -4471
rect -1788 -4475 -1784 -4471
rect -1747 -4475 -1743 -4471
rect -1705 -4475 -1701 -4471
rect -1663 -4475 -1659 -4471
rect -1622 -4475 -1618 -4471
rect -1542 -4475 -1538 -4471
rect -1525 -4475 -1521 -4471
rect -1484 -4475 -1480 -4471
rect -1442 -4475 -1438 -4471
rect -1400 -4475 -1396 -4471
rect -1359 -4475 -1355 -4471
rect -1831 -4482 -1827 -4478
rect -1346 -4482 -1342 -4478
rect -1805 -4554 -1801 -4550
rect -1788 -4554 -1784 -4550
rect -1768 -4554 -1764 -4550
rect -1747 -4554 -1743 -4550
rect -1726 -4554 -1722 -4550
rect -1705 -4554 -1701 -4550
rect -1684 -4554 -1680 -4550
rect -1663 -4554 -1659 -4550
rect -1642 -4554 -1638 -4550
rect -1622 -4554 -1618 -4550
rect -1542 -4554 -1538 -4550
rect -1525 -4554 -1521 -4550
rect -1505 -4554 -1501 -4550
rect -1484 -4554 -1480 -4550
rect -1463 -4554 -1459 -4550
rect -1442 -4554 -1438 -4550
rect -1421 -4554 -1417 -4550
rect -1400 -4554 -1396 -4550
rect -1379 -4554 -1375 -4550
rect -1359 -4554 -1355 -4550
rect -1831 -4610 -1827 -4606
rect -1814 -4617 -1810 -4613
rect -1756 -4610 -1752 -4606
rect -1714 -4617 -1710 -4613
rect -1696 -4610 -1692 -4606
rect -1654 -4602 -1650 -4598
rect -1654 -4610 -1650 -4606
rect -1672 -4624 -1668 -4620
rect -1772 -4631 -1768 -4627
rect -1730 -4631 -1726 -4627
rect -1630 -4617 -1626 -4613
rect -1551 -4617 -1547 -4613
rect -1493 -4610 -1489 -4606
rect -1451 -4617 -1447 -4613
rect -1433 -4610 -1429 -4606
rect -1391 -4602 -1387 -4598
rect -1391 -4610 -1387 -4606
rect -1409 -4624 -1405 -4620
rect -1509 -4631 -1505 -4627
rect -1467 -4631 -1463 -4627
rect -1347 -4602 -1343 -4598
rect -1367 -4617 -1363 -4613
rect -1805 -4646 -1801 -4642
rect -1788 -4646 -1784 -4642
rect -1747 -4646 -1743 -4642
rect -1705 -4646 -1701 -4642
rect -1663 -4646 -1659 -4642
rect -1622 -4646 -1618 -4642
rect -1542 -4646 -1538 -4642
rect -1525 -4646 -1521 -4642
rect -1484 -4646 -1480 -4642
rect -1442 -4646 -1438 -4642
rect -1400 -4646 -1396 -4642
rect -1359 -4646 -1355 -4642
rect -1566 -4654 -1562 -4650
rect -1347 -4654 -1343 -4650
rect -1542 -4725 -1538 -4721
rect -1525 -4725 -1521 -4721
rect -1505 -4725 -1501 -4721
rect -1484 -4725 -1480 -4721
rect -1463 -4725 -1459 -4721
rect -1442 -4725 -1438 -4721
rect -1421 -4725 -1417 -4721
rect -1400 -4725 -1396 -4721
rect -1379 -4725 -1375 -4721
rect -1359 -4725 -1355 -4721
rect -1566 -4781 -1562 -4777
rect -1551 -4788 -1547 -4784
rect -1493 -4781 -1489 -4777
rect -1451 -4788 -1447 -4784
rect -1433 -4781 -1429 -4777
rect -1391 -4773 -1387 -4769
rect -1391 -4781 -1387 -4777
rect -1409 -4795 -1405 -4791
rect -1509 -4802 -1505 -4798
rect -1467 -4802 -1463 -4798
rect -1346 -4773 -1342 -4769
rect -1367 -4788 -1363 -4784
rect -1542 -4817 -1538 -4813
rect -1525 -4817 -1521 -4813
rect -1484 -4817 -1480 -4813
rect -1442 -4817 -1438 -4813
rect -1400 -4817 -1396 -4813
rect -1359 -4817 -1355 -4813
rect -1292 -4193 -1288 -4189
rect -963 -3911 -959 -3907
rect -1225 -3986 -1221 -3982
rect -1208 -3986 -1204 -3982
rect -1188 -3986 -1184 -3982
rect -1167 -3986 -1163 -3982
rect -1146 -3986 -1142 -3982
rect -1125 -3986 -1121 -3982
rect -1104 -3986 -1100 -3982
rect -1083 -3986 -1079 -3982
rect -1062 -3986 -1058 -3982
rect -1042 -3986 -1038 -3982
rect -1234 -4049 -1230 -4045
rect -1176 -4042 -1172 -4038
rect -1134 -4049 -1130 -4045
rect -1116 -4042 -1112 -4038
rect -1074 -4034 -1070 -4030
rect -1074 -4042 -1070 -4038
rect -1092 -4056 -1088 -4052
rect -1192 -4063 -1188 -4059
rect -1150 -4063 -1146 -4059
rect -1024 -4034 -1020 -4030
rect -1050 -4049 -1046 -4045
rect -1225 -4078 -1221 -4074
rect -1208 -4078 -1204 -4074
rect -1167 -4078 -1163 -4074
rect -1125 -4078 -1121 -4074
rect -1083 -4078 -1079 -4074
rect -1042 -4078 -1038 -4074
rect -1024 -4133 -1020 -4129
rect -979 -4154 -975 -4150
rect -1225 -4260 -1221 -4256
rect -1208 -4260 -1204 -4256
rect -1168 -4260 -1164 -4256
rect -1147 -4260 -1143 -4256
rect -1257 -4316 -1253 -4312
rect -1234 -4309 -1230 -4305
rect -1283 -4323 -1279 -4319
rect -1190 -4330 -1186 -4326
rect -979 -4300 -975 -4296
rect -1138 -4308 -1134 -4304
rect -1208 -4337 -1204 -4333
rect -1172 -4337 -1168 -4333
rect -722 -3383 -718 -3379
rect -909 -3404 -905 -3400
rect -616 -3404 -612 -3400
rect -918 -3443 -914 -3439
rect -926 -3510 -922 -3506
rect -900 -3510 -896 -3506
rect -883 -3510 -879 -3506
rect -843 -3510 -839 -3506
rect -822 -3510 -818 -3506
rect -805 -3510 -801 -3506
rect -765 -3510 -761 -3506
rect -741 -3510 -737 -3506
rect -704 -3510 -700 -3506
rect -935 -3543 -931 -3539
rect -917 -3536 -913 -3532
rect -891 -3558 -887 -3554
rect -909 -3565 -905 -3561
rect -865 -3550 -861 -3546
rect -813 -3543 -809 -3539
rect -883 -3587 -879 -3583
rect -847 -3587 -843 -3583
rect -787 -3558 -783 -3554
rect -805 -3587 -801 -3583
rect -769 -3587 -765 -3583
rect -695 -3550 -691 -3546
rect -687 -3558 -683 -3554
rect -926 -3602 -922 -3598
rect -900 -3602 -896 -3598
rect -857 -3602 -853 -3598
rect -822 -3602 -818 -3598
rect -778 -3602 -774 -3598
rect -761 -3602 -757 -3598
rect -725 -3602 -721 -3598
rect -704 -3602 -700 -3598
rect -373 -2652 -369 -2648
rect -551 -2673 -547 -2669
rect -263 -2673 -259 -2669
rect -560 -2712 -556 -2708
rect -568 -2779 -564 -2775
rect -542 -2779 -538 -2775
rect -525 -2779 -521 -2775
rect -485 -2779 -481 -2775
rect -464 -2779 -460 -2775
rect -447 -2779 -443 -2775
rect -407 -2779 -403 -2775
rect -383 -2779 -379 -2775
rect -346 -2779 -342 -2775
rect -577 -2812 -573 -2808
rect -559 -2805 -555 -2801
rect -533 -2827 -529 -2823
rect -551 -2834 -547 -2830
rect -507 -2819 -503 -2815
rect -455 -2812 -451 -2808
rect -525 -2856 -521 -2852
rect -489 -2856 -485 -2852
rect -429 -2827 -425 -2823
rect -447 -2856 -443 -2852
rect -411 -2856 -407 -2852
rect -337 -2818 -333 -2814
rect -329 -2827 -325 -2823
rect -568 -2871 -564 -2867
rect -542 -2871 -538 -2867
rect -499 -2871 -495 -2867
rect -464 -2871 -460 -2867
rect -420 -2871 -416 -2867
rect -403 -2871 -399 -2867
rect -367 -2871 -363 -2867
rect -346 -2871 -342 -2867
rect -9 -1902 -5 -1898
rect -193 -1923 -189 -1919
rect 93 -1923 97 -1919
rect -202 -1962 -198 -1958
rect -210 -2029 -206 -2025
rect -184 -2029 -180 -2025
rect -167 -2029 -163 -2025
rect -127 -2029 -123 -2025
rect -106 -2029 -102 -2025
rect -89 -2029 -85 -2025
rect -49 -2029 -45 -2025
rect -25 -2029 -21 -2025
rect 12 -2029 16 -2025
rect -219 -2062 -215 -2058
rect -201 -2055 -197 -2051
rect -175 -2077 -171 -2073
rect -193 -2084 -189 -2080
rect -149 -2069 -145 -2065
rect -97 -2062 -93 -2058
rect -167 -2106 -163 -2102
rect -131 -2106 -127 -2102
rect -71 -2077 -67 -2073
rect -89 -2106 -85 -2102
rect -53 -2106 -49 -2102
rect 21 -2069 25 -2065
rect 29 -2077 33 -2073
rect -210 -2121 -206 -2117
rect -184 -2121 -180 -2117
rect -141 -2121 -137 -2117
rect -106 -2121 -102 -2117
rect -62 -2121 -58 -2117
rect -45 -2121 -41 -2117
rect -9 -2121 -5 -2117
rect 12 -2121 16 -2117
rect 165 -1187 169 -1183
rect 447 -1187 451 -1183
rect 156 -1226 160 -1222
rect 148 -1298 152 -1294
rect 174 -1298 178 -1294
rect 191 -1298 195 -1294
rect 231 -1298 235 -1294
rect 252 -1298 256 -1294
rect 269 -1298 273 -1294
rect 309 -1298 313 -1294
rect 333 -1298 337 -1294
rect 370 -1298 374 -1294
rect 139 -1331 143 -1327
rect 157 -1324 161 -1320
rect 183 -1346 187 -1342
rect 165 -1353 169 -1349
rect 209 -1338 213 -1334
rect 261 -1331 265 -1327
rect 191 -1375 195 -1371
rect 227 -1375 231 -1371
rect 287 -1346 291 -1342
rect 269 -1375 273 -1371
rect 305 -1375 309 -1371
rect 379 -1338 383 -1334
rect 386 -1346 390 -1342
rect 148 -1390 152 -1386
rect 174 -1390 178 -1386
rect 217 -1390 221 -1386
rect 252 -1390 256 -1386
rect 296 -1390 300 -1386
rect 313 -1390 317 -1386
rect 349 -1390 353 -1386
rect 370 -1390 374 -1386
rect 470 -1338 474 -1334
rect 853 -784 857 -780
rect 870 -784 874 -780
rect 521 -840 525 -836
rect 821 -840 825 -836
rect 512 -876 516 -872
rect 504 -1018 508 -1014
rect 521 -1018 525 -1014
rect 541 -1018 545 -1014
rect 562 -1018 566 -1014
rect 583 -1018 587 -1014
rect 604 -1018 608 -1014
rect 625 -1018 629 -1014
rect 646 -1018 650 -1014
rect 667 -1018 671 -1014
rect 687 -1018 691 -1014
rect 495 -1081 499 -1077
rect 553 -1074 557 -1070
rect 595 -1081 599 -1077
rect 613 -1074 617 -1070
rect 655 -1066 659 -1062
rect 655 -1074 659 -1070
rect 637 -1088 641 -1084
rect 537 -1095 541 -1091
rect 579 -1095 583 -1091
rect 679 -1081 683 -1077
rect 504 -1110 508 -1106
rect 521 -1110 525 -1106
rect 562 -1110 566 -1106
rect 604 -1110 608 -1106
rect 646 -1110 650 -1106
rect 687 -1110 691 -1106
rect 495 -1134 499 -1130
rect 512 -1134 516 -1130
rect 447 -1353 451 -1349
rect 386 -1404 390 -1400
rect 470 -1404 474 -1400
rect 148 -1421 152 -1417
rect 165 -1421 169 -1417
rect 185 -1421 189 -1417
rect 206 -1421 210 -1417
rect 227 -1421 231 -1417
rect 248 -1421 252 -1417
rect 269 -1421 273 -1417
rect 290 -1421 294 -1417
rect 311 -1421 315 -1417
rect 331 -1421 335 -1417
rect 139 -1484 143 -1480
rect 197 -1477 201 -1473
rect 239 -1484 243 -1480
rect 257 -1477 261 -1473
rect 299 -1469 303 -1465
rect 299 -1477 303 -1473
rect 281 -1491 285 -1487
rect 181 -1498 185 -1494
rect 223 -1498 227 -1494
rect 323 -1484 327 -1480
rect 148 -1513 152 -1509
rect 165 -1513 169 -1509
rect 206 -1513 210 -1509
rect 248 -1513 252 -1509
rect 290 -1513 294 -1509
rect 331 -1513 335 -1509
rect 148 -1592 152 -1588
rect 165 -1592 169 -1588
rect 185 -1592 189 -1588
rect 206 -1592 210 -1588
rect 227 -1592 231 -1588
rect 248 -1592 252 -1588
rect 269 -1592 273 -1588
rect 290 -1592 294 -1588
rect 311 -1592 315 -1588
rect 331 -1592 335 -1588
rect 139 -1655 143 -1651
rect 197 -1648 201 -1644
rect 239 -1655 243 -1651
rect 257 -1648 261 -1644
rect 299 -1640 303 -1636
rect 299 -1648 303 -1644
rect 281 -1662 285 -1658
rect 181 -1669 185 -1665
rect 223 -1669 227 -1665
rect 346 -1640 350 -1636
rect 323 -1655 327 -1651
rect 148 -1684 152 -1680
rect 165 -1684 169 -1680
rect 206 -1684 210 -1680
rect 248 -1684 252 -1680
rect 290 -1684 294 -1680
rect 331 -1684 335 -1680
rect 470 -1648 474 -1644
rect 346 -1692 350 -1688
rect 470 -1691 474 -1687
rect 148 -1763 152 -1759
rect 165 -1763 169 -1759
rect 185 -1763 189 -1759
rect 206 -1763 210 -1759
rect 227 -1763 231 -1759
rect 248 -1763 252 -1759
rect 269 -1763 273 -1759
rect 290 -1763 294 -1759
rect 311 -1763 315 -1759
rect 331 -1763 335 -1759
rect 125 -1819 129 -1815
rect 139 -1826 143 -1822
rect 197 -1819 201 -1815
rect 239 -1826 243 -1822
rect 257 -1819 261 -1815
rect 299 -1811 303 -1807
rect 299 -1819 303 -1815
rect 281 -1833 285 -1829
rect 181 -1840 185 -1836
rect 223 -1840 227 -1836
rect 350 -1811 354 -1807
rect 323 -1826 327 -1822
rect 148 -1855 152 -1851
rect 165 -1855 169 -1851
rect 206 -1855 210 -1851
rect 248 -1855 252 -1851
rect 290 -1855 294 -1851
rect 331 -1855 335 -1851
rect 139 -1870 143 -1866
rect 156 -1870 160 -1866
rect 107 -2069 111 -2065
rect 93 -2084 97 -2080
rect 29 -2128 33 -2124
rect 111 -2128 115 -2124
rect -210 -2173 -206 -2169
rect -193 -2173 -189 -2169
rect -173 -2173 -169 -2169
rect -152 -2173 -148 -2169
rect -131 -2173 -127 -2169
rect -110 -2173 -106 -2169
rect -89 -2173 -85 -2169
rect -68 -2173 -64 -2169
rect -47 -2173 -43 -2169
rect -27 -2173 -23 -2169
rect -219 -2236 -215 -2232
rect -161 -2229 -157 -2225
rect -119 -2236 -115 -2232
rect -101 -2229 -97 -2225
rect -59 -2221 -55 -2217
rect -59 -2229 -55 -2225
rect -77 -2243 -73 -2239
rect -177 -2250 -173 -2246
rect -135 -2250 -131 -2246
rect -35 -2236 -31 -2232
rect -210 -2265 -206 -2261
rect -193 -2265 -189 -2261
rect -152 -2265 -148 -2261
rect -110 -2265 -106 -2261
rect -68 -2265 -64 -2261
rect -27 -2265 -23 -2261
rect -210 -2344 -206 -2340
rect -193 -2344 -189 -2340
rect -173 -2344 -169 -2340
rect -152 -2344 -148 -2340
rect -131 -2344 -127 -2340
rect -110 -2344 -106 -2340
rect -89 -2344 -85 -2340
rect -68 -2344 -64 -2340
rect -47 -2344 -43 -2340
rect -27 -2344 -23 -2340
rect -219 -2407 -215 -2403
rect -161 -2400 -157 -2396
rect -119 -2407 -115 -2403
rect -101 -2400 -97 -2396
rect -59 -2392 -55 -2388
rect -59 -2400 -55 -2396
rect -77 -2414 -73 -2410
rect -177 -2421 -173 -2417
rect -135 -2421 -131 -2417
rect -8 -2392 -4 -2388
rect -35 -2407 -31 -2403
rect -210 -2436 -206 -2432
rect -193 -2436 -189 -2432
rect -152 -2436 -148 -2432
rect -110 -2436 -106 -2432
rect -68 -2436 -64 -2432
rect -27 -2436 -23 -2432
rect 111 -2400 115 -2396
rect -8 -2444 -4 -2440
rect 111 -2443 115 -2439
rect -211 -2515 -207 -2511
rect -194 -2515 -190 -2511
rect -174 -2515 -170 -2511
rect -153 -2515 -149 -2511
rect -132 -2515 -128 -2511
rect -111 -2515 -107 -2511
rect -90 -2515 -86 -2511
rect -69 -2515 -65 -2511
rect -48 -2515 -44 -2511
rect -28 -2515 -24 -2511
rect -233 -2571 -229 -2567
rect -220 -2578 -216 -2574
rect -162 -2571 -158 -2567
rect -120 -2578 -116 -2574
rect -102 -2571 -98 -2567
rect -60 -2563 -56 -2559
rect -60 -2571 -56 -2567
rect -78 -2585 -74 -2581
rect -178 -2592 -174 -2588
rect -136 -2592 -132 -2588
rect -12 -2563 -8 -2559
rect -36 -2578 -32 -2574
rect -211 -2607 -207 -2603
rect -194 -2607 -190 -2603
rect -153 -2607 -149 -2603
rect -111 -2607 -107 -2603
rect -69 -2607 -65 -2603
rect -28 -2607 -24 -2603
rect -219 -2620 -215 -2616
rect -202 -2620 -198 -2616
rect -249 -2819 -245 -2815
rect -263 -2834 -259 -2830
rect -329 -2885 -325 -2881
rect -249 -2885 -245 -2881
rect -568 -2898 -564 -2894
rect -551 -2898 -547 -2894
rect -531 -2898 -527 -2894
rect -510 -2898 -506 -2894
rect -489 -2898 -485 -2894
rect -468 -2898 -464 -2894
rect -447 -2898 -443 -2894
rect -426 -2898 -422 -2894
rect -405 -2898 -401 -2894
rect -385 -2898 -381 -2894
rect -577 -2961 -573 -2957
rect -519 -2954 -515 -2950
rect -477 -2961 -473 -2957
rect -459 -2954 -455 -2950
rect -417 -2946 -413 -2942
rect -417 -2954 -413 -2950
rect -435 -2968 -431 -2964
rect -535 -2975 -531 -2971
rect -493 -2975 -489 -2971
rect -393 -2961 -389 -2957
rect -568 -2990 -564 -2986
rect -551 -2990 -547 -2986
rect -510 -2990 -506 -2986
rect -468 -2990 -464 -2986
rect -426 -2990 -422 -2986
rect -385 -2990 -381 -2986
rect -568 -3069 -564 -3065
rect -551 -3069 -547 -3065
rect -531 -3069 -527 -3065
rect -510 -3069 -506 -3065
rect -489 -3069 -485 -3065
rect -468 -3069 -464 -3065
rect -447 -3069 -443 -3065
rect -426 -3069 -422 -3065
rect -405 -3069 -401 -3065
rect -385 -3069 -381 -3065
rect -577 -3132 -573 -3128
rect -519 -3125 -515 -3121
rect -477 -3132 -473 -3128
rect -459 -3125 -455 -3121
rect -417 -3117 -413 -3113
rect -417 -3125 -413 -3121
rect -435 -3139 -431 -3135
rect -535 -3146 -531 -3142
rect -493 -3146 -489 -3142
rect -367 -3117 -363 -3113
rect -393 -3132 -389 -3128
rect -568 -3161 -564 -3157
rect -551 -3161 -547 -3157
rect -510 -3161 -506 -3157
rect -468 -3161 -464 -3157
rect -426 -3161 -422 -3157
rect -385 -3161 -381 -3157
rect -249 -3125 -245 -3121
rect -367 -3168 -363 -3164
rect -249 -3169 -245 -3165
rect -568 -3240 -564 -3236
rect -551 -3240 -547 -3236
rect -531 -3240 -527 -3236
rect -510 -3240 -506 -3236
rect -489 -3240 -485 -3236
rect -468 -3240 -464 -3236
rect -447 -3240 -443 -3236
rect -426 -3240 -422 -3236
rect -405 -3240 -401 -3236
rect -385 -3240 -381 -3236
rect -591 -3296 -587 -3292
rect -577 -3303 -573 -3299
rect -519 -3296 -515 -3292
rect -477 -3303 -473 -3299
rect -459 -3296 -455 -3292
rect -417 -3288 -413 -3284
rect -417 -3296 -413 -3292
rect -435 -3310 -431 -3306
rect -535 -3317 -531 -3313
rect -493 -3317 -489 -3313
rect -369 -3288 -365 -3284
rect -393 -3303 -389 -3299
rect -568 -3332 -564 -3328
rect -551 -3332 -547 -3328
rect -510 -3332 -506 -3328
rect -468 -3332 -464 -3328
rect -426 -3332 -422 -3328
rect -385 -3332 -381 -3328
rect -577 -3351 -573 -3347
rect -560 -3351 -556 -3347
rect -603 -3550 -599 -3546
rect -616 -3565 -612 -3561
rect -687 -3609 -683 -3605
rect -603 -3609 -599 -3605
rect -925 -3640 -921 -3636
rect -908 -3640 -904 -3636
rect -888 -3640 -884 -3636
rect -867 -3640 -863 -3636
rect -846 -3640 -842 -3636
rect -825 -3640 -821 -3636
rect -804 -3640 -800 -3636
rect -783 -3640 -779 -3636
rect -762 -3640 -758 -3636
rect -742 -3640 -738 -3636
rect -934 -3703 -930 -3699
rect -876 -3696 -872 -3692
rect -834 -3703 -830 -3699
rect -816 -3696 -812 -3692
rect -774 -3688 -770 -3684
rect -774 -3696 -770 -3692
rect -792 -3710 -788 -3706
rect -892 -3717 -888 -3713
rect -850 -3717 -846 -3713
rect -750 -3703 -746 -3699
rect -925 -3732 -921 -3728
rect -908 -3732 -904 -3728
rect -867 -3732 -863 -3728
rect -825 -3732 -821 -3728
rect -783 -3732 -779 -3728
rect -742 -3732 -738 -3728
rect -925 -3811 -921 -3807
rect -908 -3811 -904 -3807
rect -888 -3811 -884 -3807
rect -867 -3811 -863 -3807
rect -846 -3811 -842 -3807
rect -825 -3811 -821 -3807
rect -804 -3811 -800 -3807
rect -783 -3811 -779 -3807
rect -762 -3811 -758 -3807
rect -742 -3811 -738 -3807
rect -934 -3874 -930 -3870
rect -876 -3867 -872 -3863
rect -834 -3874 -830 -3870
rect -816 -3867 -812 -3863
rect -774 -3859 -770 -3855
rect -774 -3867 -770 -3863
rect -792 -3881 -788 -3877
rect -892 -3888 -888 -3884
rect -850 -3888 -846 -3884
rect -723 -3859 -719 -3855
rect -750 -3874 -746 -3870
rect -925 -3903 -921 -3899
rect -908 -3903 -904 -3899
rect -867 -3903 -863 -3899
rect -825 -3903 -821 -3899
rect -783 -3903 -779 -3899
rect -742 -3903 -738 -3899
rect -603 -3867 -599 -3863
rect -723 -3911 -719 -3907
rect -603 -3910 -599 -3906
rect -926 -3986 -922 -3982
rect -909 -3986 -905 -3982
rect -889 -3986 -885 -3982
rect -868 -3986 -864 -3982
rect -847 -3986 -843 -3982
rect -826 -3986 -822 -3982
rect -805 -3986 -801 -3982
rect -784 -3986 -780 -3982
rect -763 -3986 -759 -3982
rect -743 -3986 -739 -3982
rect -949 -4042 -945 -4038
rect -935 -4049 -931 -4045
rect -877 -4042 -873 -4038
rect -835 -4049 -831 -4045
rect -817 -4042 -813 -4038
rect -775 -4034 -771 -4030
rect -775 -4042 -771 -4038
rect -793 -4056 -789 -4052
rect -893 -4063 -889 -4059
rect -851 -4063 -847 -4059
rect -719 -4034 -715 -4030
rect -751 -4049 -747 -4045
rect -926 -4078 -922 -4074
rect -909 -4078 -905 -4074
rect -868 -4078 -864 -4074
rect -826 -4078 -822 -4074
rect -784 -4078 -780 -4074
rect -743 -4078 -739 -4074
rect -935 -4101 -931 -4097
rect -918 -4101 -914 -4097
rect -963 -4315 -959 -4311
rect -1114 -4330 -1110 -4326
rect -1225 -4352 -1221 -4348
rect -1181 -4352 -1177 -4348
rect -1147 -4352 -1143 -4348
rect -1257 -4359 -1253 -4355
rect -1246 -4366 -1242 -4362
rect -1114 -4366 -1110 -4362
rect -963 -4366 -959 -4362
rect -1225 -4383 -1221 -4379
rect -1208 -4383 -1204 -4379
rect -1188 -4383 -1184 -4379
rect -1167 -4383 -1163 -4379
rect -1146 -4383 -1142 -4379
rect -1125 -4383 -1121 -4379
rect -1104 -4383 -1100 -4379
rect -1083 -4383 -1079 -4379
rect -1062 -4383 -1058 -4379
rect -1042 -4383 -1038 -4379
rect -1246 -4439 -1242 -4435
rect -1234 -4446 -1230 -4442
rect -1176 -4439 -1172 -4435
rect -1134 -4446 -1130 -4442
rect -1116 -4439 -1112 -4435
rect -1074 -4431 -1070 -4427
rect -1074 -4439 -1070 -4435
rect -1092 -4453 -1088 -4449
rect -1192 -4460 -1188 -4456
rect -1150 -4460 -1146 -4456
rect -1050 -4446 -1046 -4442
rect -1225 -4475 -1221 -4471
rect -1208 -4475 -1204 -4471
rect -1167 -4475 -1163 -4471
rect -1125 -4475 -1121 -4471
rect -1083 -4475 -1079 -4471
rect -1042 -4475 -1038 -4471
rect -1225 -4554 -1221 -4550
rect -1208 -4554 -1204 -4550
rect -1188 -4554 -1184 -4550
rect -1167 -4554 -1163 -4550
rect -1146 -4554 -1142 -4550
rect -1125 -4554 -1121 -4550
rect -1104 -4554 -1100 -4550
rect -1083 -4554 -1079 -4550
rect -1062 -4554 -1058 -4550
rect -1042 -4554 -1038 -4550
rect -1257 -4610 -1253 -4606
rect -1234 -4617 -1230 -4613
rect -1176 -4610 -1172 -4606
rect -1134 -4617 -1130 -4613
rect -1116 -4610 -1112 -4606
rect -1074 -4602 -1070 -4598
rect -1074 -4610 -1070 -4606
rect -1092 -4624 -1088 -4620
rect -1192 -4631 -1188 -4627
rect -1150 -4631 -1146 -4627
rect -1023 -4602 -1019 -4598
rect -1050 -4617 -1046 -4613
rect -1225 -4646 -1221 -4642
rect -1208 -4646 -1204 -4642
rect -1167 -4646 -1163 -4642
rect -1125 -4646 -1121 -4642
rect -1083 -4646 -1079 -4642
rect -1042 -4646 -1038 -4642
rect -963 -4610 -959 -4606
rect -1319 -4781 -1315 -4777
rect -1257 -4654 -1253 -4650
rect -1023 -4654 -1019 -4650
rect -963 -4653 -959 -4649
rect -1309 -4840 -1305 -4836
rect -1292 -4840 -1288 -4836
rect -1346 -4880 -1342 -4876
rect -1801 -5118 -1797 -5114
rect -1784 -5118 -1780 -5114
rect -1764 -5118 -1760 -5114
rect -1743 -5118 -1739 -5114
rect -1722 -5118 -1718 -5114
rect -1701 -5118 -1697 -5114
rect -1680 -5118 -1676 -5114
rect -1659 -5118 -1655 -5114
rect -1638 -5118 -1634 -5114
rect -1618 -5118 -1614 -5114
rect -1538 -5118 -1534 -5114
rect -1521 -5118 -1517 -5114
rect -1501 -5118 -1497 -5114
rect -1480 -5118 -1476 -5114
rect -1459 -5118 -1455 -5114
rect -1438 -5118 -1434 -5114
rect -1417 -5118 -1413 -5114
rect -1396 -5118 -1392 -5114
rect -1375 -5118 -1371 -5114
rect -1355 -5118 -1351 -5114
rect -1810 -5181 -1806 -5177
rect -1752 -5174 -1748 -5170
rect -1710 -5181 -1706 -5177
rect -1692 -5174 -1688 -5170
rect -1650 -5166 -1646 -5162
rect -1650 -5174 -1646 -5170
rect -1668 -5188 -1664 -5184
rect -1768 -5195 -1764 -5191
rect -1726 -5195 -1722 -5191
rect -1626 -5181 -1622 -5177
rect -1547 -5181 -1543 -5177
rect -1489 -5174 -1485 -5170
rect -1447 -5181 -1443 -5177
rect -1429 -5174 -1425 -5170
rect -1387 -5166 -1383 -5162
rect -1387 -5174 -1383 -5170
rect -1405 -5188 -1401 -5184
rect -1505 -5195 -1501 -5191
rect -1463 -5195 -1459 -5191
rect -1340 -5166 -1336 -5162
rect -1363 -5181 -1359 -5177
rect -1801 -5210 -1797 -5206
rect -1784 -5210 -1780 -5206
rect -1743 -5210 -1739 -5206
rect -1701 -5210 -1697 -5206
rect -1659 -5210 -1655 -5206
rect -1618 -5210 -1614 -5206
rect -1538 -5210 -1534 -5206
rect -1521 -5210 -1517 -5206
rect -1480 -5210 -1476 -5206
rect -1438 -5210 -1434 -5206
rect -1396 -5210 -1392 -5206
rect -1355 -5210 -1351 -5206
rect -1825 -5218 -1821 -5214
rect -1340 -5218 -1336 -5214
rect -1801 -5289 -1797 -5285
rect -1784 -5289 -1780 -5285
rect -1764 -5289 -1760 -5285
rect -1743 -5289 -1739 -5285
rect -1722 -5289 -1718 -5285
rect -1701 -5289 -1697 -5285
rect -1680 -5289 -1676 -5285
rect -1659 -5289 -1655 -5285
rect -1638 -5289 -1634 -5285
rect -1618 -5289 -1614 -5285
rect -1538 -5289 -1534 -5285
rect -1521 -5289 -1517 -5285
rect -1501 -5289 -1497 -5285
rect -1480 -5289 -1476 -5285
rect -1459 -5289 -1455 -5285
rect -1438 -5289 -1434 -5285
rect -1417 -5289 -1413 -5285
rect -1396 -5289 -1392 -5285
rect -1375 -5289 -1371 -5285
rect -1355 -5289 -1351 -5285
rect -1825 -5345 -1821 -5341
rect -1810 -5352 -1806 -5348
rect -1752 -5345 -1748 -5341
rect -1710 -5352 -1706 -5348
rect -1692 -5345 -1688 -5341
rect -1650 -5337 -1646 -5333
rect -1650 -5345 -1646 -5341
rect -1668 -5359 -1664 -5355
rect -1768 -5366 -1764 -5362
rect -1726 -5366 -1722 -5362
rect -1626 -5352 -1622 -5348
rect -1547 -5352 -1543 -5348
rect -1489 -5345 -1485 -5341
rect -1447 -5352 -1443 -5348
rect -1429 -5345 -1425 -5341
rect -1387 -5337 -1383 -5333
rect -1387 -5345 -1383 -5341
rect -1405 -5359 -1401 -5355
rect -1505 -5366 -1501 -5362
rect -1463 -5366 -1459 -5362
rect -1340 -5337 -1336 -5333
rect -1363 -5352 -1359 -5348
rect -1801 -5381 -1797 -5377
rect -1784 -5381 -1780 -5377
rect -1743 -5381 -1739 -5377
rect -1701 -5381 -1697 -5377
rect -1659 -5381 -1655 -5377
rect -1618 -5381 -1614 -5377
rect -1538 -5381 -1534 -5377
rect -1521 -5381 -1517 -5377
rect -1480 -5381 -1476 -5377
rect -1438 -5381 -1434 -5377
rect -1396 -5381 -1392 -5377
rect -1355 -5381 -1351 -5377
rect -1826 -5389 -1822 -5385
rect -1340 -5389 -1336 -5385
rect -1801 -5449 -1797 -5445
rect -1784 -5449 -1780 -5445
rect -1764 -5449 -1760 -5445
rect -1743 -5449 -1739 -5445
rect -1722 -5449 -1718 -5445
rect -1701 -5449 -1697 -5445
rect -1680 -5449 -1676 -5445
rect -1659 -5449 -1655 -5445
rect -1638 -5449 -1634 -5445
rect -1618 -5449 -1614 -5445
rect -1538 -5449 -1534 -5445
rect -1521 -5449 -1517 -5445
rect -1501 -5449 -1497 -5445
rect -1480 -5449 -1476 -5445
rect -1459 -5449 -1455 -5445
rect -1438 -5449 -1434 -5445
rect -1417 -5449 -1413 -5445
rect -1396 -5449 -1392 -5445
rect -1375 -5449 -1371 -5445
rect -1355 -5449 -1351 -5445
rect -1826 -5505 -1822 -5501
rect -1810 -5512 -1806 -5508
rect -1752 -5505 -1748 -5501
rect -1710 -5512 -1706 -5508
rect -1692 -5505 -1688 -5501
rect -1650 -5497 -1646 -5493
rect -1650 -5505 -1646 -5501
rect -1668 -5519 -1664 -5515
rect -1768 -5526 -1764 -5522
rect -1726 -5526 -1722 -5522
rect -1626 -5512 -1622 -5508
rect -1547 -5512 -1543 -5508
rect -1489 -5505 -1485 -5501
rect -1447 -5512 -1443 -5508
rect -1429 -5505 -1425 -5501
rect -1387 -5497 -1383 -5493
rect -1387 -5505 -1383 -5501
rect -1405 -5519 -1401 -5515
rect -1505 -5526 -1501 -5522
rect -1463 -5526 -1459 -5522
rect -1342 -5497 -1338 -5493
rect -1363 -5512 -1359 -5508
rect -1801 -5541 -1797 -5537
rect -1784 -5541 -1780 -5537
rect -1743 -5541 -1739 -5537
rect -1701 -5541 -1697 -5537
rect -1659 -5541 -1655 -5537
rect -1618 -5541 -1614 -5537
rect -1538 -5541 -1534 -5537
rect -1521 -5541 -1517 -5537
rect -1480 -5541 -1476 -5537
rect -1438 -5541 -1434 -5537
rect -1396 -5541 -1392 -5537
rect -1355 -5541 -1351 -5537
rect -1292 -4932 -1288 -4928
rect -1225 -4725 -1221 -4721
rect -1208 -4725 -1204 -4721
rect -1188 -4725 -1184 -4721
rect -1167 -4725 -1163 -4721
rect -1146 -4725 -1142 -4721
rect -1125 -4725 -1121 -4721
rect -1104 -4725 -1100 -4721
rect -1083 -4725 -1079 -4721
rect -1062 -4725 -1058 -4721
rect -1042 -4725 -1038 -4721
rect -1234 -4788 -1230 -4784
rect -1176 -4781 -1172 -4777
rect -1134 -4788 -1130 -4784
rect -1116 -4781 -1112 -4777
rect -1074 -4773 -1070 -4769
rect -1074 -4781 -1070 -4777
rect -1092 -4795 -1088 -4791
rect -1192 -4802 -1188 -4798
rect -1150 -4802 -1146 -4798
rect -1022 -4773 -1018 -4769
rect -1050 -4788 -1046 -4784
rect -1225 -4817 -1221 -4813
rect -1208 -4817 -1204 -4813
rect -1167 -4817 -1163 -4813
rect -1125 -4817 -1121 -4813
rect -1083 -4817 -1079 -4813
rect -1042 -4817 -1038 -4813
rect -1022 -4872 -1018 -4868
rect -979 -4893 -975 -4889
rect -1225 -4999 -1221 -4995
rect -1208 -4999 -1204 -4995
rect -1168 -4999 -1164 -4995
rect -1147 -4999 -1143 -4995
rect -1257 -5055 -1253 -5051
rect -1234 -5048 -1230 -5044
rect -1283 -5062 -1279 -5058
rect -1190 -5069 -1186 -5065
rect -979 -5039 -975 -5035
rect -1138 -5047 -1134 -5043
rect -1208 -5076 -1204 -5072
rect -1172 -5076 -1168 -5072
rect -719 -4133 -715 -4129
rect -909 -4154 -905 -4150
rect -616 -4154 -612 -4150
rect -918 -4193 -914 -4189
rect -926 -4260 -922 -4256
rect -900 -4260 -896 -4256
rect -883 -4260 -879 -4256
rect -843 -4260 -839 -4256
rect -822 -4260 -818 -4256
rect -805 -4260 -801 -4256
rect -765 -4260 -761 -4256
rect -741 -4260 -737 -4256
rect -704 -4260 -700 -4256
rect -935 -4293 -931 -4289
rect -917 -4286 -913 -4282
rect -891 -4308 -887 -4304
rect -909 -4315 -905 -4311
rect -865 -4300 -861 -4296
rect -813 -4293 -809 -4289
rect -883 -4337 -879 -4333
rect -847 -4337 -843 -4333
rect -787 -4308 -783 -4304
rect -805 -4337 -801 -4333
rect -769 -4337 -765 -4333
rect -695 -4300 -691 -4296
rect -687 -4308 -683 -4304
rect -926 -4352 -922 -4348
rect -900 -4352 -896 -4348
rect -857 -4352 -853 -4348
rect -822 -4352 -818 -4348
rect -778 -4352 -774 -4348
rect -761 -4352 -757 -4348
rect -725 -4352 -721 -4348
rect -704 -4352 -700 -4348
rect -369 -3383 -365 -3379
rect -551 -3404 -547 -3400
rect -263 -3404 -259 -3400
rect -560 -3443 -556 -3439
rect -568 -3510 -564 -3506
rect -542 -3510 -538 -3506
rect -525 -3510 -521 -3506
rect -485 -3510 -481 -3506
rect -464 -3510 -460 -3506
rect -447 -3510 -443 -3506
rect -407 -3510 -403 -3506
rect -383 -3510 -379 -3506
rect -346 -3510 -342 -3506
rect -577 -3543 -573 -3539
rect -559 -3536 -555 -3532
rect -533 -3558 -529 -3554
rect -551 -3565 -547 -3561
rect -507 -3550 -503 -3546
rect -455 -3543 -451 -3539
rect -525 -3587 -521 -3583
rect -489 -3587 -485 -3583
rect -429 -3558 -425 -3554
rect -447 -3587 -443 -3583
rect -411 -3587 -407 -3583
rect -337 -3549 -333 -3545
rect -328 -3558 -324 -3554
rect -568 -3602 -564 -3598
rect -542 -3602 -538 -3598
rect -499 -3602 -495 -3598
rect -464 -3602 -460 -3598
rect -420 -3602 -416 -3598
rect -403 -3602 -399 -3598
rect -367 -3602 -363 -3598
rect -346 -3602 -342 -3598
rect -12 -2652 -8 -2648
rect -193 -2673 -189 -2669
rect 97 -2673 101 -2669
rect -202 -2712 -198 -2708
rect -210 -2779 -206 -2775
rect -184 -2779 -180 -2775
rect -167 -2779 -163 -2775
rect -127 -2779 -123 -2775
rect -106 -2779 -102 -2775
rect -89 -2779 -85 -2775
rect -49 -2779 -45 -2775
rect -25 -2779 -21 -2775
rect 12 -2779 16 -2775
rect -219 -2812 -215 -2808
rect -201 -2805 -197 -2801
rect -175 -2827 -171 -2823
rect -193 -2834 -189 -2830
rect -149 -2819 -145 -2815
rect -97 -2812 -93 -2808
rect -167 -2856 -163 -2852
rect -131 -2856 -127 -2852
rect -71 -2827 -67 -2823
rect -89 -2856 -85 -2852
rect -53 -2856 -49 -2852
rect 21 -2819 25 -2815
rect 28 -2827 32 -2823
rect -210 -2871 -206 -2867
rect -184 -2871 -180 -2867
rect -141 -2871 -137 -2867
rect -106 -2871 -102 -2867
rect -62 -2871 -58 -2867
rect -45 -2871 -41 -2867
rect -9 -2871 -5 -2867
rect 12 -2871 16 -2867
rect 350 -1902 354 -1898
rect 165 -1923 169 -1919
rect 451 -1923 455 -1919
rect 156 -1962 160 -1958
rect 148 -2029 152 -2025
rect 174 -2029 178 -2025
rect 191 -2029 195 -2025
rect 231 -2029 235 -2025
rect 252 -2029 256 -2025
rect 269 -2029 273 -2025
rect 309 -2029 313 -2025
rect 333 -2029 337 -2025
rect 370 -2029 374 -2025
rect 139 -2062 143 -2058
rect 157 -2055 161 -2051
rect 183 -2077 187 -2073
rect 165 -2084 169 -2080
rect 209 -2069 213 -2065
rect 261 -2062 265 -2058
rect 191 -2106 195 -2102
rect 227 -2106 231 -2102
rect 287 -2077 291 -2073
rect 269 -2106 273 -2102
rect 305 -2106 309 -2102
rect 379 -2069 383 -2065
rect 388 -2077 392 -2073
rect 148 -2121 152 -2117
rect 174 -2121 178 -2117
rect 217 -2121 221 -2117
rect 252 -2121 256 -2117
rect 296 -2121 300 -2117
rect 313 -2121 317 -2117
rect 349 -2121 353 -2117
rect 370 -2121 374 -2117
rect 521 -1187 525 -1183
rect 805 -1187 809 -1183
rect 512 -1226 516 -1222
rect 504 -1298 508 -1294
rect 530 -1298 534 -1294
rect 547 -1298 551 -1294
rect 587 -1298 591 -1294
rect 608 -1298 612 -1294
rect 625 -1298 629 -1294
rect 665 -1298 669 -1294
rect 689 -1298 693 -1294
rect 726 -1298 730 -1294
rect 495 -1331 499 -1327
rect 513 -1324 517 -1320
rect 539 -1346 543 -1342
rect 521 -1353 525 -1349
rect 565 -1338 569 -1334
rect 617 -1331 621 -1327
rect 547 -1375 551 -1371
rect 583 -1375 587 -1371
rect 643 -1346 647 -1342
rect 625 -1375 629 -1371
rect 661 -1375 665 -1371
rect 735 -1338 739 -1334
rect 742 -1346 746 -1342
rect 504 -1390 508 -1386
rect 530 -1390 534 -1386
rect 573 -1390 577 -1386
rect 608 -1390 612 -1386
rect 652 -1390 656 -1386
rect 669 -1390 673 -1386
rect 705 -1390 709 -1386
rect 726 -1390 730 -1386
rect 821 -1338 825 -1334
rect 879 -832 883 -828
rect 1211 -784 1215 -780
rect 1228 -784 1232 -780
rect 870 -876 874 -872
rect 862 -1018 866 -1014
rect 879 -1018 883 -1014
rect 899 -1018 903 -1014
rect 920 -1018 924 -1014
rect 941 -1018 945 -1014
rect 962 -1018 966 -1014
rect 983 -1018 987 -1014
rect 1004 -1018 1008 -1014
rect 1025 -1018 1029 -1014
rect 1045 -1018 1049 -1014
rect 853 -1081 857 -1077
rect 911 -1074 915 -1070
rect 953 -1081 957 -1077
rect 971 -1074 975 -1070
rect 1013 -1066 1017 -1062
rect 1013 -1074 1017 -1070
rect 995 -1088 999 -1084
rect 895 -1095 899 -1091
rect 937 -1095 941 -1091
rect 1037 -1081 1041 -1077
rect 862 -1110 866 -1106
rect 879 -1110 883 -1106
rect 920 -1110 924 -1106
rect 962 -1110 966 -1106
rect 1004 -1110 1008 -1106
rect 1045 -1110 1049 -1106
rect 853 -1134 857 -1130
rect 870 -1134 874 -1130
rect 805 -1353 809 -1349
rect 742 -1411 746 -1407
rect 823 -1411 827 -1407
rect 504 -1421 508 -1417
rect 521 -1421 525 -1417
rect 541 -1421 545 -1417
rect 562 -1421 566 -1417
rect 583 -1421 587 -1417
rect 604 -1421 608 -1417
rect 625 -1421 629 -1417
rect 646 -1421 650 -1417
rect 667 -1421 671 -1417
rect 687 -1421 691 -1417
rect 495 -1484 499 -1480
rect 553 -1477 557 -1473
rect 595 -1484 599 -1480
rect 613 -1477 617 -1473
rect 655 -1469 659 -1465
rect 655 -1477 659 -1473
rect 637 -1491 641 -1487
rect 537 -1498 541 -1494
rect 579 -1498 583 -1494
rect 679 -1484 683 -1480
rect 504 -1513 508 -1509
rect 521 -1513 525 -1509
rect 562 -1513 566 -1509
rect 604 -1513 608 -1509
rect 646 -1513 650 -1509
rect 687 -1513 691 -1509
rect 504 -1592 508 -1588
rect 521 -1592 525 -1588
rect 541 -1592 545 -1588
rect 562 -1592 566 -1588
rect 583 -1592 587 -1588
rect 604 -1592 608 -1588
rect 625 -1592 629 -1588
rect 646 -1592 650 -1588
rect 667 -1592 671 -1588
rect 687 -1592 691 -1588
rect 495 -1655 499 -1651
rect 553 -1648 557 -1644
rect 595 -1655 599 -1651
rect 613 -1648 617 -1644
rect 655 -1640 659 -1636
rect 655 -1648 659 -1644
rect 637 -1662 641 -1658
rect 537 -1669 541 -1665
rect 579 -1669 583 -1665
rect 704 -1640 708 -1636
rect 679 -1655 683 -1651
rect 504 -1684 508 -1680
rect 521 -1684 525 -1680
rect 562 -1684 566 -1680
rect 604 -1684 608 -1680
rect 646 -1684 650 -1680
rect 687 -1684 691 -1680
rect 823 -1648 827 -1644
rect 704 -1691 708 -1687
rect 823 -1691 827 -1687
rect 504 -1763 508 -1759
rect 521 -1763 525 -1759
rect 541 -1763 545 -1759
rect 562 -1763 566 -1759
rect 583 -1763 587 -1759
rect 604 -1763 608 -1759
rect 625 -1763 629 -1759
rect 646 -1763 650 -1759
rect 667 -1763 671 -1759
rect 687 -1763 691 -1759
rect 481 -1819 485 -1815
rect 495 -1826 499 -1822
rect 553 -1819 557 -1815
rect 595 -1826 599 -1822
rect 613 -1819 617 -1815
rect 655 -1811 659 -1807
rect 655 -1819 659 -1815
rect 637 -1833 641 -1829
rect 537 -1840 541 -1836
rect 579 -1840 583 -1836
rect 703 -1811 707 -1807
rect 679 -1826 683 -1822
rect 504 -1855 508 -1851
rect 521 -1855 525 -1851
rect 562 -1855 566 -1851
rect 604 -1855 608 -1851
rect 646 -1855 650 -1851
rect 687 -1855 691 -1851
rect 495 -1870 499 -1866
rect 512 -1870 516 -1866
rect 470 -2069 474 -2065
rect 451 -2084 455 -2080
rect 388 -2135 392 -2131
rect 465 -2135 469 -2131
rect 148 -2173 152 -2169
rect 165 -2173 169 -2169
rect 185 -2173 189 -2169
rect 206 -2173 210 -2169
rect 227 -2173 231 -2169
rect 248 -2173 252 -2169
rect 269 -2173 273 -2169
rect 290 -2173 294 -2169
rect 311 -2173 315 -2169
rect 331 -2173 335 -2169
rect 139 -2236 143 -2232
rect 197 -2229 201 -2225
rect 239 -2236 243 -2232
rect 257 -2229 261 -2225
rect 299 -2221 303 -2217
rect 299 -2229 303 -2225
rect 281 -2243 285 -2239
rect 181 -2250 185 -2246
rect 223 -2250 227 -2246
rect 323 -2236 327 -2232
rect 148 -2265 152 -2261
rect 165 -2265 169 -2261
rect 206 -2265 210 -2261
rect 248 -2265 252 -2261
rect 290 -2265 294 -2261
rect 331 -2265 335 -2261
rect 148 -2344 152 -2340
rect 165 -2344 169 -2340
rect 185 -2344 189 -2340
rect 206 -2344 210 -2340
rect 227 -2344 231 -2340
rect 248 -2344 252 -2340
rect 269 -2344 273 -2340
rect 290 -2344 294 -2340
rect 311 -2344 315 -2340
rect 331 -2344 335 -2340
rect 139 -2407 143 -2403
rect 197 -2400 201 -2396
rect 239 -2407 243 -2403
rect 257 -2400 261 -2396
rect 299 -2392 303 -2388
rect 299 -2400 303 -2396
rect 281 -2414 285 -2410
rect 181 -2421 185 -2417
rect 223 -2421 227 -2417
rect 346 -2392 350 -2388
rect 323 -2407 327 -2403
rect 148 -2436 152 -2432
rect 165 -2436 169 -2432
rect 206 -2436 210 -2432
rect 248 -2436 252 -2432
rect 290 -2436 294 -2432
rect 331 -2436 335 -2432
rect 465 -2400 469 -2396
rect 346 -2443 350 -2439
rect 465 -2443 469 -2439
rect 148 -2515 152 -2511
rect 165 -2515 169 -2511
rect 185 -2515 189 -2511
rect 206 -2515 210 -2511
rect 227 -2515 231 -2511
rect 248 -2515 252 -2511
rect 269 -2515 273 -2511
rect 290 -2515 294 -2511
rect 311 -2515 315 -2511
rect 331 -2515 335 -2511
rect 125 -2571 129 -2567
rect 139 -2578 143 -2574
rect 197 -2571 201 -2567
rect 239 -2578 243 -2574
rect 257 -2571 261 -2567
rect 299 -2563 303 -2559
rect 299 -2571 303 -2567
rect 281 -2585 285 -2581
rect 181 -2592 185 -2588
rect 223 -2592 227 -2588
rect 347 -2563 351 -2559
rect 323 -2578 327 -2574
rect 148 -2607 152 -2603
rect 165 -2607 169 -2603
rect 206 -2607 210 -2603
rect 248 -2607 252 -2603
rect 290 -2607 294 -2603
rect 331 -2607 335 -2603
rect 139 -2620 143 -2616
rect 156 -2620 160 -2616
rect 111 -2819 115 -2815
rect 97 -2834 101 -2830
rect 28 -2878 32 -2874
rect 111 -2878 115 -2874
rect -210 -2898 -206 -2894
rect -193 -2898 -189 -2894
rect -173 -2898 -169 -2894
rect -152 -2898 -148 -2894
rect -131 -2898 -127 -2894
rect -110 -2898 -106 -2894
rect -89 -2898 -85 -2894
rect -68 -2898 -64 -2894
rect -47 -2898 -43 -2894
rect -27 -2898 -23 -2894
rect -219 -2961 -215 -2957
rect -161 -2954 -157 -2950
rect -119 -2961 -115 -2957
rect -101 -2954 -97 -2950
rect -59 -2946 -55 -2942
rect -59 -2954 -55 -2950
rect -77 -2968 -73 -2964
rect -177 -2975 -173 -2971
rect -135 -2975 -131 -2971
rect -35 -2961 -31 -2957
rect -210 -2990 -206 -2986
rect -193 -2990 -189 -2986
rect -152 -2990 -148 -2986
rect -110 -2990 -106 -2986
rect -68 -2990 -64 -2986
rect -27 -2990 -23 -2986
rect -210 -3069 -206 -3065
rect -193 -3069 -189 -3065
rect -173 -3069 -169 -3065
rect -152 -3069 -148 -3065
rect -131 -3069 -127 -3065
rect -110 -3069 -106 -3065
rect -89 -3069 -85 -3065
rect -68 -3069 -64 -3065
rect -47 -3069 -43 -3065
rect -27 -3069 -23 -3065
rect -219 -3132 -215 -3128
rect -161 -3125 -157 -3121
rect -119 -3132 -115 -3128
rect -101 -3125 -97 -3121
rect -59 -3117 -55 -3113
rect -59 -3125 -55 -3121
rect -77 -3139 -73 -3135
rect -177 -3146 -173 -3142
rect -135 -3146 -131 -3142
rect -13 -3117 -9 -3113
rect -35 -3132 -31 -3128
rect -210 -3161 -206 -3157
rect -193 -3161 -189 -3157
rect -152 -3161 -148 -3157
rect -110 -3161 -106 -3157
rect -68 -3161 -64 -3157
rect -27 -3161 -23 -3157
rect 111 -3125 115 -3121
rect -13 -3169 -9 -3165
rect 111 -3168 115 -3164
rect -210 -3240 -206 -3236
rect -193 -3240 -189 -3236
rect -173 -3240 -169 -3236
rect -152 -3240 -148 -3236
rect -131 -3240 -127 -3236
rect -110 -3240 -106 -3236
rect -89 -3240 -85 -3236
rect -68 -3240 -64 -3236
rect -47 -3240 -43 -3236
rect -27 -3240 -23 -3236
rect -233 -3296 -229 -3292
rect -219 -3303 -215 -3299
rect -161 -3296 -157 -3292
rect -119 -3303 -115 -3299
rect -101 -3296 -97 -3292
rect -59 -3288 -55 -3284
rect -59 -3296 -55 -3292
rect -77 -3310 -73 -3306
rect -177 -3317 -173 -3313
rect -135 -3317 -131 -3313
rect -13 -3288 -9 -3284
rect -35 -3303 -31 -3299
rect -210 -3332 -206 -3328
rect -193 -3332 -189 -3328
rect -152 -3332 -148 -3328
rect -110 -3332 -106 -3328
rect -68 -3332 -64 -3328
rect -27 -3332 -23 -3328
rect -219 -3351 -215 -3347
rect -202 -3351 -198 -3347
rect -249 -3550 -245 -3546
rect -263 -3565 -259 -3561
rect -328 -3616 -324 -3612
rect -249 -3616 -245 -3612
rect -568 -3640 -564 -3636
rect -551 -3640 -547 -3636
rect -531 -3640 -527 -3636
rect -510 -3640 -506 -3636
rect -489 -3640 -485 -3636
rect -468 -3640 -464 -3636
rect -447 -3640 -443 -3636
rect -426 -3640 -422 -3636
rect -405 -3640 -401 -3636
rect -385 -3640 -381 -3636
rect -577 -3703 -573 -3699
rect -519 -3696 -515 -3692
rect -477 -3703 -473 -3699
rect -459 -3696 -455 -3692
rect -417 -3688 -413 -3684
rect -417 -3696 -413 -3692
rect -435 -3710 -431 -3706
rect -535 -3717 -531 -3713
rect -493 -3717 -489 -3713
rect -393 -3703 -389 -3699
rect -568 -3732 -564 -3728
rect -551 -3732 -547 -3728
rect -510 -3732 -506 -3728
rect -468 -3732 -464 -3728
rect -426 -3732 -422 -3728
rect -385 -3732 -381 -3728
rect -568 -3811 -564 -3807
rect -551 -3811 -547 -3807
rect -531 -3811 -527 -3807
rect -510 -3811 -506 -3807
rect -489 -3811 -485 -3807
rect -468 -3811 -464 -3807
rect -447 -3811 -443 -3807
rect -426 -3811 -422 -3807
rect -405 -3811 -401 -3807
rect -385 -3811 -381 -3807
rect -577 -3874 -573 -3870
rect -519 -3867 -515 -3863
rect -477 -3874 -473 -3870
rect -459 -3867 -455 -3863
rect -417 -3859 -413 -3855
rect -417 -3867 -413 -3863
rect -435 -3881 -431 -3877
rect -535 -3888 -531 -3884
rect -493 -3888 -489 -3884
rect -369 -3859 -365 -3855
rect -393 -3874 -389 -3870
rect -568 -3903 -564 -3899
rect -551 -3903 -547 -3899
rect -510 -3903 -506 -3899
rect -468 -3903 -464 -3899
rect -426 -3903 -422 -3899
rect -385 -3903 -381 -3899
rect -249 -3867 -245 -3863
rect -369 -3910 -365 -3906
rect -249 -3910 -245 -3906
rect -568 -3986 -564 -3982
rect -551 -3986 -547 -3982
rect -531 -3986 -527 -3982
rect -510 -3986 -506 -3982
rect -489 -3986 -485 -3982
rect -468 -3986 -464 -3982
rect -447 -3986 -443 -3982
rect -426 -3986 -422 -3982
rect -405 -3986 -401 -3982
rect -385 -3986 -381 -3982
rect -591 -4042 -587 -4038
rect -577 -4049 -573 -4045
rect -519 -4042 -515 -4038
rect -477 -4049 -473 -4045
rect -459 -4042 -455 -4038
rect -417 -4034 -413 -4030
rect -417 -4042 -413 -4038
rect -435 -4056 -431 -4052
rect -535 -4063 -531 -4059
rect -493 -4063 -489 -4059
rect -369 -4034 -365 -4030
rect -393 -4049 -389 -4045
rect -568 -4078 -564 -4074
rect -551 -4078 -547 -4074
rect -510 -4078 -506 -4074
rect -468 -4078 -464 -4074
rect -426 -4078 -422 -4074
rect -385 -4078 -381 -4074
rect -577 -4101 -573 -4097
rect -560 -4101 -556 -4097
rect -603 -4300 -599 -4296
rect -616 -4315 -612 -4311
rect -687 -4359 -683 -4355
rect -603 -4359 -599 -4355
rect -926 -4383 -922 -4379
rect -909 -4383 -905 -4379
rect -889 -4383 -885 -4379
rect -868 -4383 -864 -4379
rect -847 -4383 -843 -4379
rect -826 -4383 -822 -4379
rect -805 -4383 -801 -4379
rect -784 -4383 -780 -4379
rect -763 -4383 -759 -4379
rect -743 -4383 -739 -4379
rect -935 -4446 -931 -4442
rect -877 -4439 -873 -4435
rect -835 -4446 -831 -4442
rect -817 -4439 -813 -4435
rect -775 -4431 -771 -4427
rect -775 -4439 -771 -4435
rect -793 -4453 -789 -4449
rect -893 -4460 -889 -4456
rect -851 -4460 -847 -4456
rect -751 -4446 -747 -4442
rect -926 -4475 -922 -4471
rect -909 -4475 -905 -4471
rect -868 -4475 -864 -4471
rect -826 -4475 -822 -4471
rect -784 -4475 -780 -4471
rect -743 -4475 -739 -4471
rect -926 -4554 -922 -4550
rect -909 -4554 -905 -4550
rect -889 -4554 -885 -4550
rect -868 -4554 -864 -4550
rect -847 -4554 -843 -4550
rect -826 -4554 -822 -4550
rect -805 -4554 -801 -4550
rect -784 -4554 -780 -4550
rect -763 -4554 -759 -4550
rect -743 -4554 -739 -4550
rect -935 -4617 -931 -4613
rect -877 -4610 -873 -4606
rect -835 -4617 -831 -4613
rect -817 -4610 -813 -4606
rect -775 -4602 -771 -4598
rect -775 -4610 -771 -4606
rect -793 -4624 -789 -4620
rect -893 -4631 -889 -4627
rect -851 -4631 -847 -4627
rect -729 -4602 -725 -4598
rect -751 -4617 -747 -4613
rect -926 -4646 -922 -4642
rect -909 -4646 -905 -4642
rect -868 -4646 -864 -4642
rect -826 -4646 -822 -4642
rect -784 -4646 -780 -4642
rect -743 -4646 -739 -4642
rect -603 -4610 -599 -4606
rect -729 -4653 -725 -4649
rect -603 -4653 -599 -4649
rect -926 -4725 -922 -4721
rect -909 -4725 -905 -4721
rect -889 -4725 -885 -4721
rect -868 -4725 -864 -4721
rect -847 -4725 -843 -4721
rect -826 -4725 -822 -4721
rect -805 -4725 -801 -4721
rect -784 -4725 -780 -4721
rect -763 -4725 -759 -4721
rect -743 -4725 -739 -4721
rect -949 -4781 -945 -4777
rect -935 -4788 -931 -4784
rect -877 -4781 -873 -4777
rect -835 -4788 -831 -4784
rect -817 -4781 -813 -4777
rect -775 -4773 -771 -4769
rect -775 -4781 -771 -4777
rect -793 -4795 -789 -4791
rect -893 -4802 -889 -4798
rect -851 -4802 -847 -4798
rect -722 -4773 -718 -4769
rect -751 -4788 -747 -4784
rect -926 -4817 -922 -4813
rect -909 -4817 -905 -4813
rect -868 -4817 -864 -4813
rect -826 -4817 -822 -4813
rect -784 -4817 -780 -4813
rect -743 -4817 -739 -4813
rect -935 -4840 -931 -4836
rect -918 -4840 -914 -4836
rect -963 -5054 -959 -5050
rect -1102 -5069 -1098 -5065
rect -1225 -5091 -1221 -5087
rect -1181 -5091 -1177 -5087
rect -1147 -5091 -1143 -5087
rect -1257 -5098 -1253 -5094
rect -1246 -5106 -1242 -5102
rect -1102 -5106 -1098 -5102
rect -963 -5105 -959 -5101
rect -1225 -5118 -1221 -5114
rect -1208 -5118 -1204 -5114
rect -1188 -5118 -1184 -5114
rect -1167 -5118 -1163 -5114
rect -1146 -5118 -1142 -5114
rect -1125 -5118 -1121 -5114
rect -1104 -5118 -1100 -5114
rect -1083 -5118 -1079 -5114
rect -1062 -5118 -1058 -5114
rect -1042 -5118 -1038 -5114
rect -1246 -5174 -1242 -5170
rect -1234 -5181 -1230 -5177
rect -1176 -5174 -1172 -5170
rect -1134 -5181 -1130 -5177
rect -1116 -5174 -1112 -5170
rect -1074 -5166 -1070 -5162
rect -1074 -5174 -1070 -5170
rect -1092 -5188 -1088 -5184
rect -1192 -5195 -1188 -5191
rect -1150 -5195 -1146 -5191
rect -1050 -5181 -1046 -5177
rect -1225 -5210 -1221 -5206
rect -1208 -5210 -1204 -5206
rect -1167 -5210 -1163 -5206
rect -1125 -5210 -1121 -5206
rect -1083 -5210 -1079 -5206
rect -1042 -5210 -1038 -5206
rect -1225 -5289 -1221 -5285
rect -1208 -5289 -1204 -5285
rect -1188 -5289 -1184 -5285
rect -1167 -5289 -1163 -5285
rect -1146 -5289 -1142 -5285
rect -1125 -5289 -1121 -5285
rect -1104 -5289 -1100 -5285
rect -1083 -5289 -1079 -5285
rect -1062 -5289 -1058 -5285
rect -1042 -5289 -1038 -5285
rect -1257 -5345 -1253 -5341
rect -1234 -5352 -1230 -5348
rect -1176 -5345 -1172 -5341
rect -1134 -5352 -1130 -5348
rect -1116 -5345 -1112 -5341
rect -1074 -5337 -1070 -5333
rect -1074 -5345 -1070 -5341
rect -1092 -5359 -1088 -5355
rect -1192 -5366 -1188 -5362
rect -1150 -5366 -1146 -5362
rect -1024 -5337 -1020 -5333
rect -1050 -5352 -1046 -5348
rect -1225 -5381 -1221 -5377
rect -1208 -5381 -1204 -5377
rect -1167 -5381 -1163 -5377
rect -1125 -5381 -1121 -5377
rect -1083 -5381 -1079 -5377
rect -1042 -5381 -1038 -5377
rect -963 -5345 -959 -5341
rect -1319 -5505 -1315 -5501
rect -1257 -5388 -1253 -5384
rect -1024 -5388 -1020 -5384
rect -963 -5388 -959 -5384
rect -1309 -5563 -1305 -5559
rect -1292 -5563 -1288 -5559
rect -1342 -5603 -1338 -5599
rect -1292 -5655 -1288 -5651
rect -1225 -5449 -1221 -5445
rect -1208 -5449 -1204 -5445
rect -1188 -5449 -1184 -5445
rect -1167 -5449 -1163 -5445
rect -1146 -5449 -1142 -5445
rect -1125 -5449 -1121 -5445
rect -1104 -5449 -1100 -5445
rect -1083 -5449 -1079 -5445
rect -1062 -5449 -1058 -5445
rect -1042 -5449 -1038 -5445
rect -1234 -5512 -1230 -5508
rect -1176 -5505 -1172 -5501
rect -1134 -5512 -1130 -5508
rect -1116 -5505 -1112 -5501
rect -1074 -5497 -1070 -5493
rect -1074 -5505 -1070 -5501
rect -1092 -5519 -1088 -5515
rect -1192 -5526 -1188 -5522
rect -1150 -5526 -1146 -5522
rect -1020 -5497 -1016 -5493
rect -1050 -5512 -1046 -5508
rect -1225 -5541 -1221 -5537
rect -1208 -5541 -1204 -5537
rect -1167 -5541 -1163 -5537
rect -1125 -5541 -1121 -5537
rect -1083 -5541 -1079 -5537
rect -1042 -5541 -1038 -5537
rect -1020 -5595 -1016 -5591
rect -979 -5616 -975 -5612
rect -1225 -5722 -1221 -5718
rect -1208 -5722 -1204 -5718
rect -1168 -5722 -1164 -5718
rect -1147 -5722 -1143 -5718
rect -1257 -5778 -1253 -5774
rect -1234 -5771 -1230 -5767
rect -1283 -5785 -1279 -5781
rect -1190 -5792 -1186 -5788
rect -979 -5762 -975 -5758
rect -1138 -5770 -1134 -5766
rect -1208 -5799 -1204 -5795
rect -1172 -5799 -1168 -5795
rect -722 -4872 -718 -4868
rect -909 -4893 -905 -4889
rect -616 -4893 -612 -4889
rect -918 -4932 -914 -4928
rect -926 -4999 -922 -4995
rect -900 -4999 -896 -4995
rect -883 -4999 -879 -4995
rect -843 -4999 -839 -4995
rect -822 -4999 -818 -4995
rect -805 -4999 -801 -4995
rect -765 -4999 -761 -4995
rect -741 -4999 -737 -4995
rect -704 -4999 -700 -4995
rect -935 -5032 -931 -5028
rect -917 -5025 -913 -5021
rect -891 -5047 -887 -5043
rect -909 -5054 -905 -5050
rect -865 -5039 -861 -5035
rect -813 -5032 -809 -5028
rect -883 -5076 -879 -5072
rect -847 -5076 -843 -5072
rect -787 -5047 -783 -5043
rect -805 -5076 -801 -5072
rect -769 -5076 -765 -5072
rect -695 -5039 -691 -5035
rect -687 -5047 -683 -5043
rect -926 -5091 -922 -5087
rect -900 -5091 -896 -5087
rect -857 -5091 -853 -5087
rect -822 -5091 -818 -5087
rect -778 -5091 -774 -5087
rect -761 -5091 -757 -5087
rect -725 -5091 -721 -5087
rect -704 -5091 -700 -5087
rect -369 -4133 -365 -4129
rect -551 -4154 -547 -4150
rect -263 -4154 -259 -4150
rect -560 -4193 -556 -4189
rect -568 -4260 -564 -4256
rect -542 -4260 -538 -4256
rect -525 -4260 -521 -4256
rect -485 -4260 -481 -4256
rect -464 -4260 -460 -4256
rect -447 -4260 -443 -4256
rect -407 -4260 -403 -4256
rect -383 -4260 -379 -4256
rect -346 -4260 -342 -4256
rect -577 -4293 -573 -4289
rect -559 -4286 -555 -4282
rect -533 -4308 -529 -4304
rect -551 -4315 -547 -4311
rect -507 -4300 -503 -4296
rect -455 -4293 -451 -4289
rect -525 -4337 -521 -4333
rect -489 -4337 -485 -4333
rect -429 -4308 -425 -4304
rect -447 -4337 -443 -4333
rect -411 -4337 -407 -4333
rect -337 -4299 -333 -4295
rect -328 -4308 -324 -4304
rect -568 -4352 -564 -4348
rect -542 -4352 -538 -4348
rect -499 -4352 -495 -4348
rect -464 -4352 -460 -4348
rect -420 -4352 -416 -4348
rect -403 -4352 -399 -4348
rect -367 -4352 -363 -4348
rect -346 -4352 -342 -4348
rect -13 -3383 -9 -3379
rect -193 -3404 -189 -3400
rect 97 -3404 101 -3400
rect -202 -3443 -198 -3439
rect -210 -3510 -206 -3506
rect -184 -3510 -180 -3506
rect -167 -3510 -163 -3506
rect -127 -3510 -123 -3506
rect -106 -3510 -102 -3506
rect -89 -3510 -85 -3506
rect -49 -3510 -45 -3506
rect -25 -3510 -21 -3506
rect 12 -3510 16 -3506
rect -219 -3543 -215 -3539
rect -201 -3536 -197 -3532
rect -175 -3558 -171 -3554
rect -193 -3565 -189 -3561
rect -149 -3550 -145 -3546
rect -97 -3543 -93 -3539
rect -167 -3587 -163 -3583
rect -131 -3587 -127 -3583
rect -71 -3558 -67 -3554
rect -89 -3587 -85 -3583
rect -53 -3587 -49 -3583
rect 21 -3550 25 -3546
rect 29 -3558 33 -3554
rect -210 -3602 -206 -3598
rect -184 -3602 -180 -3598
rect -141 -3602 -137 -3598
rect -106 -3602 -102 -3598
rect -62 -3602 -58 -3598
rect -45 -3602 -41 -3598
rect -9 -3602 -5 -3598
rect 12 -3602 16 -3598
rect 347 -2652 351 -2648
rect 165 -2673 169 -2669
rect 451 -2673 455 -2669
rect 156 -2712 160 -2708
rect 148 -2779 152 -2775
rect 174 -2779 178 -2775
rect 191 -2779 195 -2775
rect 231 -2779 235 -2775
rect 252 -2779 256 -2775
rect 269 -2779 273 -2775
rect 309 -2779 313 -2775
rect 333 -2779 337 -2775
rect 370 -2779 374 -2775
rect 139 -2812 143 -2808
rect 157 -2805 161 -2801
rect 183 -2827 187 -2823
rect 165 -2834 169 -2830
rect 209 -2819 213 -2815
rect 261 -2812 265 -2808
rect 191 -2856 195 -2852
rect 227 -2856 231 -2852
rect 287 -2827 291 -2823
rect 269 -2856 273 -2852
rect 305 -2856 309 -2852
rect 379 -2819 383 -2815
rect 389 -2827 393 -2823
rect 148 -2871 152 -2867
rect 174 -2871 178 -2867
rect 217 -2871 221 -2867
rect 252 -2871 256 -2867
rect 296 -2871 300 -2867
rect 313 -2871 317 -2867
rect 349 -2871 353 -2867
rect 370 -2871 374 -2867
rect 703 -1902 707 -1898
rect 521 -1923 525 -1919
rect 809 -1923 813 -1919
rect 512 -1962 516 -1958
rect 504 -2029 508 -2025
rect 530 -2029 534 -2025
rect 547 -2029 551 -2025
rect 587 -2029 591 -2025
rect 608 -2029 612 -2025
rect 625 -2029 629 -2025
rect 665 -2029 669 -2025
rect 689 -2029 693 -2025
rect 726 -2029 730 -2025
rect 495 -2062 499 -2058
rect 513 -2055 517 -2051
rect 539 -2077 543 -2073
rect 521 -2084 525 -2080
rect 565 -2069 569 -2065
rect 617 -2062 621 -2058
rect 547 -2106 551 -2102
rect 583 -2106 587 -2102
rect 643 -2077 647 -2073
rect 625 -2106 629 -2102
rect 661 -2106 665 -2102
rect 735 -2069 739 -2065
rect 743 -2077 747 -2073
rect 504 -2121 508 -2117
rect 530 -2121 534 -2117
rect 573 -2121 577 -2117
rect 608 -2121 612 -2117
rect 652 -2121 656 -2117
rect 669 -2121 673 -2117
rect 705 -2121 709 -2117
rect 726 -2121 730 -2117
rect 1237 -840 1241 -836
rect 1228 -876 1232 -872
rect 1211 -1134 1215 -1130
rect 1228 -1134 1232 -1130
rect 879 -1187 883 -1183
rect 1163 -1187 1167 -1183
rect 870 -1226 874 -1222
rect 862 -1298 866 -1294
rect 888 -1298 892 -1294
rect 905 -1298 909 -1294
rect 945 -1298 949 -1294
rect 966 -1298 970 -1294
rect 983 -1298 987 -1294
rect 1023 -1298 1027 -1294
rect 1047 -1298 1051 -1294
rect 1084 -1298 1088 -1294
rect 853 -1331 857 -1327
rect 871 -1324 875 -1320
rect 897 -1346 901 -1342
rect 879 -1353 883 -1349
rect 923 -1338 927 -1334
rect 975 -1331 979 -1327
rect 905 -1375 909 -1371
rect 941 -1375 945 -1371
rect 1001 -1346 1005 -1342
rect 983 -1375 987 -1371
rect 1019 -1375 1023 -1371
rect 1093 -1354 1097 -1350
rect 1100 -1346 1104 -1342
rect 862 -1390 866 -1386
rect 888 -1390 892 -1386
rect 931 -1390 935 -1386
rect 966 -1390 970 -1386
rect 1010 -1390 1014 -1386
rect 1027 -1390 1031 -1386
rect 1063 -1390 1067 -1386
rect 1084 -1390 1088 -1386
rect 1163 -1361 1167 -1357
rect 1100 -1404 1104 -1400
rect 1184 -1404 1188 -1400
rect 862 -1421 866 -1417
rect 879 -1421 883 -1417
rect 899 -1421 903 -1417
rect 920 -1421 924 -1417
rect 941 -1421 945 -1417
rect 962 -1421 966 -1417
rect 983 -1421 987 -1417
rect 1004 -1421 1008 -1417
rect 1025 -1421 1029 -1417
rect 1045 -1421 1049 -1417
rect 853 -1484 857 -1480
rect 911 -1477 915 -1473
rect 953 -1484 957 -1480
rect 971 -1477 975 -1473
rect 1013 -1469 1017 -1465
rect 1013 -1477 1017 -1473
rect 995 -1491 999 -1487
rect 895 -1498 899 -1494
rect 937 -1498 941 -1494
rect 1037 -1484 1041 -1480
rect 862 -1513 866 -1509
rect 879 -1513 883 -1509
rect 920 -1513 924 -1509
rect 962 -1513 966 -1509
rect 1004 -1513 1008 -1509
rect 1045 -1513 1049 -1509
rect 862 -1592 866 -1588
rect 879 -1592 883 -1588
rect 899 -1592 903 -1588
rect 920 -1592 924 -1588
rect 941 -1592 945 -1588
rect 962 -1592 966 -1588
rect 983 -1592 987 -1588
rect 1004 -1592 1008 -1588
rect 1025 -1592 1029 -1588
rect 1045 -1592 1049 -1588
rect 853 -1655 857 -1651
rect 911 -1648 915 -1644
rect 953 -1655 957 -1651
rect 971 -1648 975 -1644
rect 1013 -1640 1017 -1636
rect 1013 -1648 1017 -1644
rect 995 -1662 999 -1658
rect 895 -1669 899 -1665
rect 937 -1669 941 -1665
rect 1063 -1640 1067 -1636
rect 1037 -1655 1041 -1651
rect 862 -1684 866 -1680
rect 879 -1684 883 -1680
rect 920 -1684 924 -1680
rect 962 -1684 966 -1680
rect 1004 -1684 1008 -1680
rect 1045 -1684 1049 -1680
rect 1184 -1648 1188 -1644
rect 1063 -1691 1067 -1687
rect 1184 -1692 1188 -1688
rect 862 -1763 866 -1759
rect 879 -1763 883 -1759
rect 899 -1763 903 -1759
rect 920 -1763 924 -1759
rect 941 -1763 945 -1759
rect 962 -1763 966 -1759
rect 983 -1763 987 -1759
rect 1004 -1763 1008 -1759
rect 1025 -1763 1029 -1759
rect 1045 -1763 1049 -1759
rect 839 -1819 843 -1815
rect 853 -1826 857 -1822
rect 911 -1819 915 -1815
rect 953 -1826 957 -1822
rect 971 -1819 975 -1815
rect 1013 -1811 1017 -1807
rect 1013 -1819 1017 -1815
rect 995 -1833 999 -1829
rect 895 -1840 899 -1836
rect 937 -1840 941 -1836
rect 1060 -1811 1064 -1807
rect 1037 -1826 1041 -1822
rect 862 -1855 866 -1851
rect 879 -1855 883 -1851
rect 920 -1855 924 -1851
rect 962 -1855 966 -1851
rect 1004 -1855 1008 -1851
rect 1045 -1855 1049 -1851
rect 853 -1870 857 -1866
rect 870 -1870 874 -1866
rect 823 -2069 827 -2065
rect 809 -2084 813 -2080
rect 743 -2128 747 -2124
rect 824 -2128 828 -2124
rect 504 -2173 508 -2169
rect 521 -2173 525 -2169
rect 541 -2173 545 -2169
rect 562 -2173 566 -2169
rect 583 -2173 587 -2169
rect 604 -2173 608 -2169
rect 625 -2173 629 -2169
rect 646 -2173 650 -2169
rect 667 -2173 671 -2169
rect 687 -2173 691 -2169
rect 495 -2236 499 -2232
rect 553 -2229 557 -2225
rect 595 -2236 599 -2232
rect 613 -2229 617 -2225
rect 655 -2221 659 -2217
rect 655 -2229 659 -2225
rect 637 -2243 641 -2239
rect 537 -2250 541 -2246
rect 579 -2250 583 -2246
rect 679 -2236 683 -2232
rect 504 -2265 508 -2261
rect 521 -2265 525 -2261
rect 562 -2265 566 -2261
rect 604 -2265 608 -2261
rect 646 -2265 650 -2261
rect 687 -2265 691 -2261
rect 504 -2344 508 -2340
rect 521 -2344 525 -2340
rect 541 -2344 545 -2340
rect 562 -2344 566 -2340
rect 583 -2344 587 -2340
rect 604 -2344 608 -2340
rect 625 -2344 629 -2340
rect 646 -2344 650 -2340
rect 667 -2344 671 -2340
rect 687 -2344 691 -2340
rect 495 -2407 499 -2403
rect 553 -2400 557 -2396
rect 595 -2407 599 -2403
rect 613 -2400 617 -2396
rect 655 -2392 659 -2388
rect 655 -2400 659 -2396
rect 637 -2414 641 -2410
rect 537 -2421 541 -2417
rect 579 -2421 583 -2417
rect 705 -2392 709 -2388
rect 679 -2407 683 -2403
rect 504 -2436 508 -2432
rect 521 -2436 525 -2432
rect 562 -2436 566 -2432
rect 604 -2436 608 -2432
rect 646 -2436 650 -2432
rect 687 -2436 691 -2432
rect 824 -2400 828 -2396
rect 705 -2443 709 -2439
rect 824 -2444 828 -2440
rect 504 -2515 508 -2511
rect 521 -2515 525 -2511
rect 541 -2515 545 -2511
rect 562 -2515 566 -2511
rect 583 -2515 587 -2511
rect 604 -2515 608 -2511
rect 625 -2515 629 -2511
rect 646 -2515 650 -2511
rect 667 -2515 671 -2511
rect 687 -2515 691 -2511
rect 481 -2571 485 -2567
rect 495 -2578 499 -2574
rect 553 -2571 557 -2567
rect 595 -2578 599 -2574
rect 613 -2571 617 -2567
rect 655 -2563 659 -2559
rect 655 -2571 659 -2567
rect 637 -2585 641 -2581
rect 537 -2592 541 -2588
rect 579 -2592 583 -2588
rect 703 -2563 707 -2559
rect 679 -2578 683 -2574
rect 504 -2607 508 -2603
rect 521 -2607 525 -2603
rect 562 -2607 566 -2603
rect 604 -2607 608 -2603
rect 646 -2607 650 -2603
rect 687 -2607 691 -2603
rect 495 -2620 499 -2616
rect 512 -2620 516 -2616
rect 465 -2819 469 -2815
rect 451 -2834 455 -2830
rect 389 -2885 393 -2881
rect 465 -2885 469 -2881
rect 148 -2898 152 -2894
rect 165 -2898 169 -2894
rect 185 -2898 189 -2894
rect 206 -2898 210 -2894
rect 227 -2898 231 -2894
rect 248 -2898 252 -2894
rect 269 -2898 273 -2894
rect 290 -2898 294 -2894
rect 311 -2898 315 -2894
rect 331 -2898 335 -2894
rect 139 -2961 143 -2957
rect 197 -2954 201 -2950
rect 239 -2961 243 -2957
rect 257 -2954 261 -2950
rect 299 -2946 303 -2942
rect 299 -2954 303 -2950
rect 281 -2968 285 -2964
rect 181 -2975 185 -2971
rect 223 -2975 227 -2971
rect 323 -2961 327 -2957
rect 148 -2990 152 -2986
rect 165 -2990 169 -2986
rect 206 -2990 210 -2986
rect 248 -2990 252 -2986
rect 290 -2990 294 -2986
rect 331 -2990 335 -2986
rect 148 -3069 152 -3065
rect 165 -3069 169 -3065
rect 185 -3069 189 -3065
rect 206 -3069 210 -3065
rect 227 -3069 231 -3065
rect 248 -3069 252 -3065
rect 269 -3069 273 -3065
rect 290 -3069 294 -3065
rect 311 -3069 315 -3065
rect 331 -3069 335 -3065
rect 139 -3132 143 -3128
rect 197 -3125 201 -3121
rect 239 -3132 243 -3128
rect 257 -3125 261 -3121
rect 299 -3117 303 -3113
rect 299 -3125 303 -3121
rect 281 -3139 285 -3135
rect 181 -3146 185 -3142
rect 223 -3146 227 -3142
rect 345 -3117 349 -3113
rect 323 -3132 327 -3128
rect 148 -3161 152 -3157
rect 165 -3161 169 -3157
rect 206 -3161 210 -3157
rect 248 -3161 252 -3157
rect 290 -3161 294 -3157
rect 331 -3161 335 -3157
rect 465 -3125 469 -3121
rect 345 -3168 349 -3164
rect 465 -3168 469 -3164
rect 148 -3240 152 -3236
rect 165 -3240 169 -3236
rect 185 -3240 189 -3236
rect 206 -3240 210 -3236
rect 227 -3240 231 -3236
rect 248 -3240 252 -3236
rect 269 -3240 273 -3236
rect 290 -3240 294 -3236
rect 311 -3240 315 -3236
rect 331 -3240 335 -3236
rect 125 -3296 129 -3292
rect 139 -3303 143 -3299
rect 197 -3296 201 -3292
rect 239 -3303 243 -3299
rect 257 -3296 261 -3292
rect 299 -3288 303 -3284
rect 299 -3296 303 -3292
rect 281 -3310 285 -3306
rect 181 -3317 185 -3313
rect 223 -3317 227 -3313
rect 347 -3288 351 -3284
rect 323 -3303 327 -3299
rect 148 -3332 152 -3328
rect 165 -3332 169 -3328
rect 206 -3332 210 -3328
rect 248 -3332 252 -3328
rect 290 -3332 294 -3328
rect 331 -3332 335 -3328
rect 139 -3351 143 -3347
rect 156 -3351 160 -3347
rect 111 -3550 115 -3546
rect 97 -3565 101 -3561
rect 29 -3609 33 -3605
rect 111 -3609 115 -3605
rect -210 -3640 -206 -3636
rect -193 -3640 -189 -3636
rect -173 -3640 -169 -3636
rect -152 -3640 -148 -3636
rect -131 -3640 -127 -3636
rect -110 -3640 -106 -3636
rect -89 -3640 -85 -3636
rect -68 -3640 -64 -3636
rect -47 -3640 -43 -3636
rect -27 -3640 -23 -3636
rect -219 -3703 -215 -3699
rect -161 -3696 -157 -3692
rect -119 -3703 -115 -3699
rect -101 -3696 -97 -3692
rect -59 -3688 -55 -3684
rect -59 -3696 -55 -3692
rect -77 -3710 -73 -3706
rect -177 -3717 -173 -3713
rect -135 -3717 -131 -3713
rect -35 -3703 -31 -3699
rect -210 -3732 -206 -3728
rect -193 -3732 -189 -3728
rect -152 -3732 -148 -3728
rect -110 -3732 -106 -3728
rect -68 -3732 -64 -3728
rect -27 -3732 -23 -3728
rect -210 -3811 -206 -3807
rect -193 -3811 -189 -3807
rect -173 -3811 -169 -3807
rect -152 -3811 -148 -3807
rect -131 -3811 -127 -3807
rect -110 -3811 -106 -3807
rect -89 -3811 -85 -3807
rect -68 -3811 -64 -3807
rect -47 -3811 -43 -3807
rect -27 -3811 -23 -3807
rect -219 -3874 -215 -3870
rect -161 -3867 -157 -3863
rect -119 -3874 -115 -3870
rect -101 -3867 -97 -3863
rect -59 -3859 -55 -3855
rect -59 -3867 -55 -3863
rect -77 -3881 -73 -3877
rect -177 -3888 -173 -3884
rect -135 -3888 -131 -3884
rect -9 -3859 -5 -3855
rect -35 -3874 -31 -3870
rect -210 -3903 -206 -3899
rect -193 -3903 -189 -3899
rect -152 -3903 -148 -3899
rect -110 -3903 -106 -3899
rect -68 -3903 -64 -3899
rect -27 -3903 -23 -3899
rect 111 -3867 115 -3863
rect -9 -3910 -5 -3906
rect 111 -3910 115 -3906
rect -210 -3986 -206 -3982
rect -193 -3986 -189 -3982
rect -173 -3986 -169 -3982
rect -152 -3986 -148 -3982
rect -131 -3986 -127 -3982
rect -110 -3986 -106 -3982
rect -89 -3986 -85 -3982
rect -68 -3986 -64 -3982
rect -47 -3986 -43 -3982
rect -27 -3986 -23 -3982
rect -233 -4042 -229 -4038
rect -219 -4049 -215 -4045
rect -161 -4042 -157 -4038
rect -119 -4049 -115 -4045
rect -101 -4042 -97 -4038
rect -59 -4034 -55 -4030
rect -59 -4042 -55 -4038
rect -77 -4056 -73 -4052
rect -177 -4063 -173 -4059
rect -135 -4063 -131 -4059
rect -9 -4034 -5 -4030
rect -35 -4049 -31 -4045
rect -210 -4078 -206 -4074
rect -193 -4078 -189 -4074
rect -152 -4078 -148 -4074
rect -110 -4078 -106 -4074
rect -68 -4078 -64 -4074
rect -27 -4078 -23 -4074
rect -219 -4101 -215 -4097
rect -202 -4101 -198 -4097
rect -249 -4300 -245 -4296
rect -263 -4315 -259 -4311
rect -328 -4366 -324 -4362
rect -249 -4366 -245 -4362
rect -568 -4383 -564 -4379
rect -551 -4383 -547 -4379
rect -531 -4383 -527 -4379
rect -510 -4383 -506 -4379
rect -489 -4383 -485 -4379
rect -468 -4383 -464 -4379
rect -447 -4383 -443 -4379
rect -426 -4383 -422 -4379
rect -405 -4383 -401 -4379
rect -385 -4383 -381 -4379
rect -577 -4446 -573 -4442
rect -519 -4439 -515 -4435
rect -477 -4446 -473 -4442
rect -459 -4439 -455 -4435
rect -417 -4431 -413 -4427
rect -417 -4439 -413 -4435
rect -435 -4453 -431 -4449
rect -535 -4460 -531 -4456
rect -493 -4460 -489 -4456
rect -393 -4446 -389 -4442
rect -568 -4475 -564 -4471
rect -551 -4475 -547 -4471
rect -510 -4475 -506 -4471
rect -468 -4475 -464 -4471
rect -426 -4475 -422 -4471
rect -385 -4475 -381 -4471
rect -568 -4554 -564 -4550
rect -551 -4554 -547 -4550
rect -531 -4554 -527 -4550
rect -510 -4554 -506 -4550
rect -489 -4554 -485 -4550
rect -468 -4554 -464 -4550
rect -447 -4554 -443 -4550
rect -426 -4554 -422 -4550
rect -405 -4554 -401 -4550
rect -385 -4554 -381 -4550
rect -577 -4617 -573 -4613
rect -519 -4610 -515 -4606
rect -477 -4617 -473 -4613
rect -459 -4610 -455 -4606
rect -417 -4602 -413 -4598
rect -417 -4610 -413 -4606
rect -435 -4624 -431 -4620
rect -535 -4631 -531 -4627
rect -493 -4631 -489 -4627
rect -370 -4602 -366 -4598
rect -393 -4617 -389 -4613
rect -568 -4646 -564 -4642
rect -551 -4646 -547 -4642
rect -510 -4646 -506 -4642
rect -468 -4646 -464 -4642
rect -426 -4646 -422 -4642
rect -385 -4646 -381 -4642
rect -249 -4610 -245 -4606
rect -370 -4653 -366 -4649
rect -249 -4653 -245 -4649
rect -568 -4725 -564 -4721
rect -551 -4725 -547 -4721
rect -531 -4725 -527 -4721
rect -510 -4725 -506 -4721
rect -489 -4725 -485 -4721
rect -468 -4725 -464 -4721
rect -447 -4725 -443 -4721
rect -426 -4725 -422 -4721
rect -405 -4725 -401 -4721
rect -385 -4725 -381 -4721
rect -591 -4781 -587 -4777
rect -577 -4788 -573 -4784
rect -519 -4781 -515 -4777
rect -477 -4788 -473 -4784
rect -459 -4781 -455 -4777
rect -417 -4773 -413 -4769
rect -417 -4781 -413 -4777
rect -435 -4795 -431 -4791
rect -535 -4802 -531 -4798
rect -493 -4802 -489 -4798
rect -369 -4773 -365 -4769
rect -393 -4788 -389 -4784
rect -568 -4817 -564 -4813
rect -551 -4817 -547 -4813
rect -510 -4817 -506 -4813
rect -468 -4817 -464 -4813
rect -426 -4817 -422 -4813
rect -385 -4817 -381 -4813
rect -577 -4840 -573 -4836
rect -560 -4840 -556 -4836
rect -603 -5039 -599 -5035
rect -616 -5054 -612 -5050
rect -687 -5098 -683 -5094
rect -603 -5098 -599 -5094
rect -926 -5118 -922 -5114
rect -909 -5118 -905 -5114
rect -889 -5118 -885 -5114
rect -868 -5118 -864 -5114
rect -847 -5118 -843 -5114
rect -826 -5118 -822 -5114
rect -805 -5118 -801 -5114
rect -784 -5118 -780 -5114
rect -763 -5118 -759 -5114
rect -743 -5118 -739 -5114
rect -935 -5181 -931 -5177
rect -877 -5174 -873 -5170
rect -835 -5181 -831 -5177
rect -817 -5174 -813 -5170
rect -775 -5166 -771 -5162
rect -775 -5174 -771 -5170
rect -793 -5188 -789 -5184
rect -893 -5195 -889 -5191
rect -851 -5195 -847 -5191
rect -751 -5181 -747 -5177
rect -926 -5210 -922 -5206
rect -909 -5210 -905 -5206
rect -868 -5210 -864 -5206
rect -826 -5210 -822 -5206
rect -784 -5210 -780 -5206
rect -743 -5210 -739 -5206
rect -926 -5289 -922 -5285
rect -909 -5289 -905 -5285
rect -889 -5289 -885 -5285
rect -868 -5289 -864 -5285
rect -847 -5289 -843 -5285
rect -826 -5289 -822 -5285
rect -805 -5289 -801 -5285
rect -784 -5289 -780 -5285
rect -763 -5289 -759 -5285
rect -743 -5289 -739 -5285
rect -935 -5352 -931 -5348
rect -877 -5345 -873 -5341
rect -835 -5352 -831 -5348
rect -817 -5345 -813 -5341
rect -775 -5337 -771 -5333
rect -775 -5345 -771 -5341
rect -793 -5359 -789 -5355
rect -893 -5366 -889 -5362
rect -851 -5366 -847 -5362
rect -725 -5337 -721 -5333
rect -751 -5352 -747 -5348
rect -926 -5381 -922 -5377
rect -909 -5381 -905 -5377
rect -868 -5381 -864 -5377
rect -826 -5381 -822 -5377
rect -784 -5381 -780 -5377
rect -743 -5381 -739 -5377
rect -603 -5345 -599 -5341
rect -725 -5388 -721 -5384
rect -603 -5389 -599 -5385
rect -926 -5449 -922 -5445
rect -909 -5449 -905 -5445
rect -889 -5449 -885 -5445
rect -868 -5449 -864 -5445
rect -847 -5449 -843 -5445
rect -826 -5449 -822 -5445
rect -805 -5449 -801 -5445
rect -784 -5449 -780 -5445
rect -763 -5449 -759 -5445
rect -743 -5449 -739 -5445
rect -949 -5505 -945 -5501
rect -935 -5512 -931 -5508
rect -877 -5505 -873 -5501
rect -835 -5512 -831 -5508
rect -817 -5505 -813 -5501
rect -775 -5497 -771 -5493
rect -775 -5505 -771 -5501
rect -793 -5519 -789 -5515
rect -893 -5526 -889 -5522
rect -851 -5526 -847 -5522
rect -725 -5497 -721 -5493
rect -751 -5512 -747 -5508
rect -926 -5541 -922 -5537
rect -909 -5541 -905 -5537
rect -868 -5541 -864 -5537
rect -826 -5541 -822 -5537
rect -784 -5541 -780 -5537
rect -743 -5541 -739 -5537
rect -935 -5563 -931 -5559
rect -918 -5563 -914 -5559
rect -725 -5595 -721 -5591
rect -909 -5616 -905 -5612
rect -616 -5616 -612 -5612
rect -918 -5655 -914 -5651
rect -926 -5722 -922 -5718
rect -900 -5722 -896 -5718
rect -883 -5722 -879 -5718
rect -843 -5722 -839 -5718
rect -822 -5722 -818 -5718
rect -805 -5722 -801 -5718
rect -765 -5722 -761 -5718
rect -741 -5722 -737 -5718
rect -704 -5722 -700 -5718
rect -963 -5777 -959 -5773
rect -935 -5755 -931 -5751
rect -1103 -5792 -1099 -5788
rect -1225 -5814 -1221 -5810
rect -1181 -5814 -1177 -5810
rect -1147 -5814 -1143 -5810
rect -917 -5748 -913 -5744
rect -891 -5770 -887 -5766
rect -909 -5777 -905 -5773
rect -865 -5762 -861 -5758
rect -813 -5755 -809 -5751
rect -883 -5799 -879 -5795
rect -847 -5799 -843 -5795
rect -787 -5770 -783 -5766
rect -805 -5799 -801 -5795
rect -769 -5799 -765 -5795
rect -695 -5762 -691 -5758
rect -683 -5770 -679 -5766
rect -926 -5814 -922 -5810
rect -900 -5814 -896 -5810
rect -857 -5814 -853 -5810
rect -822 -5814 -818 -5810
rect -778 -5814 -774 -5810
rect -761 -5814 -757 -5810
rect -725 -5814 -721 -5810
rect -704 -5814 -700 -5810
rect -369 -4872 -365 -4868
rect -551 -4893 -547 -4889
rect -263 -4893 -259 -4889
rect -560 -4932 -556 -4928
rect -568 -4999 -564 -4995
rect -542 -4999 -538 -4995
rect -525 -4999 -521 -4995
rect -485 -4999 -481 -4995
rect -464 -4999 -460 -4995
rect -447 -4999 -443 -4995
rect -407 -4999 -403 -4995
rect -383 -4999 -379 -4995
rect -346 -4999 -342 -4995
rect -577 -5032 -573 -5028
rect -559 -5025 -555 -5021
rect -533 -5047 -529 -5043
rect -551 -5054 -547 -5050
rect -507 -5039 -503 -5035
rect -455 -5032 -451 -5028
rect -525 -5076 -521 -5072
rect -489 -5076 -485 -5072
rect -429 -5047 -425 -5043
rect -447 -5076 -443 -5072
rect -411 -5076 -407 -5072
rect -337 -5038 -333 -5034
rect -328 -5047 -324 -5043
rect -568 -5091 -564 -5087
rect -542 -5091 -538 -5087
rect -499 -5091 -495 -5087
rect -464 -5091 -460 -5087
rect -420 -5091 -416 -5087
rect -403 -5091 -399 -5087
rect -367 -5091 -363 -5087
rect -346 -5091 -342 -5087
rect -9 -4133 -5 -4129
rect -193 -4154 -189 -4150
rect 97 -4154 101 -4150
rect -202 -4193 -198 -4189
rect -210 -4260 -206 -4256
rect -184 -4260 -180 -4256
rect -167 -4260 -163 -4256
rect -127 -4260 -123 -4256
rect -106 -4260 -102 -4256
rect -89 -4260 -85 -4256
rect -49 -4260 -45 -4256
rect -25 -4260 -21 -4256
rect 12 -4260 16 -4256
rect -219 -4293 -215 -4289
rect -201 -4286 -197 -4282
rect -175 -4308 -171 -4304
rect -193 -4315 -189 -4311
rect -149 -4300 -145 -4296
rect -97 -4293 -93 -4289
rect -167 -4337 -163 -4333
rect -131 -4337 -127 -4333
rect -71 -4308 -67 -4304
rect -89 -4337 -85 -4333
rect -53 -4337 -49 -4333
rect 21 -4300 25 -4296
rect 29 -4308 33 -4304
rect -210 -4352 -206 -4348
rect -184 -4352 -180 -4348
rect -141 -4352 -137 -4348
rect -106 -4352 -102 -4348
rect -62 -4352 -58 -4348
rect -45 -4352 -41 -4348
rect -9 -4352 -5 -4348
rect 12 -4352 16 -4348
rect 347 -3383 351 -3379
rect 165 -3404 169 -3400
rect 451 -3404 455 -3400
rect 156 -3443 160 -3439
rect 148 -3510 152 -3506
rect 174 -3510 178 -3506
rect 191 -3510 195 -3506
rect 231 -3510 235 -3506
rect 252 -3510 256 -3506
rect 269 -3510 273 -3506
rect 309 -3510 313 -3506
rect 333 -3510 337 -3506
rect 370 -3510 374 -3506
rect 139 -3543 143 -3539
rect 157 -3536 161 -3532
rect 183 -3558 187 -3554
rect 165 -3565 169 -3561
rect 209 -3550 213 -3546
rect 261 -3543 265 -3539
rect 191 -3587 195 -3583
rect 227 -3587 231 -3583
rect 287 -3558 291 -3554
rect 269 -3587 273 -3583
rect 305 -3587 309 -3583
rect 379 -3550 383 -3546
rect 388 -3558 392 -3554
rect 148 -3602 152 -3598
rect 174 -3602 178 -3598
rect 217 -3602 221 -3598
rect 252 -3602 256 -3598
rect 296 -3602 300 -3598
rect 313 -3602 317 -3598
rect 349 -3602 353 -3598
rect 370 -3602 374 -3598
rect 703 -2652 707 -2648
rect 521 -2673 525 -2669
rect 810 -2673 814 -2669
rect 512 -2712 516 -2708
rect 504 -2779 508 -2775
rect 530 -2779 534 -2775
rect 547 -2779 551 -2775
rect 587 -2779 591 -2775
rect 608 -2779 612 -2775
rect 625 -2779 629 -2775
rect 665 -2779 669 -2775
rect 689 -2779 693 -2775
rect 726 -2779 730 -2775
rect 495 -2812 499 -2808
rect 513 -2805 517 -2801
rect 539 -2827 543 -2823
rect 521 -2834 525 -2830
rect 565 -2819 569 -2815
rect 617 -2812 621 -2808
rect 547 -2856 551 -2852
rect 583 -2856 587 -2852
rect 643 -2827 647 -2823
rect 625 -2856 629 -2852
rect 661 -2856 665 -2852
rect 735 -2819 739 -2815
rect 742 -2827 746 -2823
rect 504 -2871 508 -2867
rect 530 -2871 534 -2867
rect 573 -2871 577 -2867
rect 608 -2871 612 -2867
rect 652 -2871 656 -2867
rect 669 -2871 673 -2867
rect 705 -2871 709 -2867
rect 726 -2871 730 -2867
rect 1060 -1902 1064 -1898
rect 879 -1923 883 -1919
rect 1167 -1923 1171 -1919
rect 870 -1962 874 -1958
rect 862 -2029 866 -2025
rect 888 -2029 892 -2025
rect 905 -2029 909 -2025
rect 945 -2029 949 -2025
rect 966 -2029 970 -2025
rect 983 -2029 987 -2025
rect 1023 -2029 1027 -2025
rect 1047 -2029 1051 -2025
rect 1084 -2029 1088 -2025
rect 853 -2062 857 -2058
rect 871 -2055 875 -2051
rect 897 -2077 901 -2073
rect 879 -2084 883 -2080
rect 923 -2069 927 -2065
rect 975 -2062 979 -2058
rect 905 -2106 909 -2102
rect 941 -2106 945 -2102
rect 1001 -2077 1005 -2073
rect 983 -2106 987 -2102
rect 1019 -2106 1023 -2102
rect 1093 -2067 1097 -2063
rect 1167 -2069 1171 -2065
rect 1093 -2085 1097 -2081
rect 1101 -2077 1105 -2073
rect 862 -2121 866 -2117
rect 888 -2121 892 -2117
rect 931 -2121 935 -2117
rect 966 -2121 970 -2117
rect 1010 -2121 1014 -2117
rect 1027 -2121 1031 -2117
rect 1063 -2121 1067 -2117
rect 1084 -2121 1088 -2117
rect 1237 -1187 1241 -1183
rect 1228 -1226 1232 -1222
rect 1220 -1298 1224 -1294
rect 1237 -1298 1241 -1294
rect 1277 -1298 1281 -1294
rect 1298 -1298 1302 -1294
rect 1211 -1347 1215 -1343
rect 1255 -1368 1259 -1364
rect 1307 -1346 1311 -1342
rect 1237 -1375 1241 -1371
rect 1273 -1375 1277 -1371
rect 1322 -1368 1326 -1364
rect 1220 -1390 1224 -1386
rect 1264 -1390 1268 -1386
rect 1298 -1390 1302 -1386
rect 1329 -1404 1333 -1400
rect 1322 -1411 1326 -1407
rect 1220 -1592 1224 -1588
rect 1237 -1592 1241 -1588
rect 1257 -1592 1261 -1588
rect 1278 -1592 1282 -1588
rect 1299 -1592 1303 -1588
rect 1320 -1592 1324 -1588
rect 1341 -1592 1345 -1588
rect 1362 -1592 1366 -1588
rect 1383 -1592 1387 -1588
rect 1403 -1592 1407 -1588
rect 1211 -1655 1215 -1651
rect 1269 -1648 1273 -1644
rect 1311 -1655 1315 -1651
rect 1329 -1648 1333 -1644
rect 1371 -1640 1375 -1636
rect 1371 -1648 1375 -1644
rect 1353 -1662 1357 -1658
rect 1253 -1669 1257 -1665
rect 1295 -1669 1299 -1665
rect 1424 -1640 1428 -1636
rect 1395 -1655 1399 -1651
rect 1220 -1684 1224 -1680
rect 1237 -1684 1241 -1680
rect 1278 -1684 1282 -1680
rect 1320 -1684 1324 -1680
rect 1362 -1684 1366 -1680
rect 1403 -1684 1407 -1680
rect 1424 -1692 1428 -1688
rect 1220 -1763 1224 -1759
rect 1237 -1763 1241 -1759
rect 1257 -1763 1261 -1759
rect 1278 -1763 1282 -1759
rect 1299 -1763 1303 -1759
rect 1320 -1763 1324 -1759
rect 1341 -1763 1345 -1759
rect 1362 -1763 1366 -1759
rect 1383 -1763 1387 -1759
rect 1403 -1763 1407 -1759
rect 1197 -1819 1201 -1815
rect 1211 -1826 1215 -1822
rect 1269 -1819 1273 -1815
rect 1311 -1826 1315 -1822
rect 1329 -1819 1333 -1815
rect 1371 -1811 1375 -1807
rect 1371 -1819 1375 -1815
rect 1353 -1833 1357 -1829
rect 1253 -1840 1257 -1836
rect 1295 -1840 1299 -1836
rect 1419 -1811 1423 -1807
rect 1395 -1826 1399 -1822
rect 1220 -1855 1224 -1851
rect 1237 -1855 1241 -1851
rect 1278 -1855 1282 -1851
rect 1320 -1855 1324 -1851
rect 1362 -1855 1366 -1851
rect 1403 -1855 1407 -1851
rect 1211 -1870 1215 -1866
rect 1228 -1870 1232 -1866
rect 1184 -2084 1188 -2080
rect 1101 -2135 1105 -2131
rect 1184 -2135 1188 -2131
rect 862 -2344 866 -2340
rect 879 -2344 883 -2340
rect 899 -2344 903 -2340
rect 920 -2344 924 -2340
rect 941 -2344 945 -2340
rect 962 -2344 966 -2340
rect 983 -2344 987 -2340
rect 1004 -2344 1008 -2340
rect 1025 -2344 1029 -2340
rect 1045 -2344 1049 -2340
rect 853 -2407 857 -2403
rect 911 -2400 915 -2396
rect 953 -2407 957 -2403
rect 971 -2400 975 -2396
rect 1013 -2392 1017 -2388
rect 1013 -2400 1017 -2396
rect 995 -2414 999 -2410
rect 895 -2421 899 -2417
rect 937 -2421 941 -2417
rect 1062 -2392 1066 -2388
rect 1037 -2407 1041 -2403
rect 862 -2436 866 -2432
rect 879 -2436 883 -2432
rect 920 -2436 924 -2432
rect 962 -2436 966 -2432
rect 1004 -2436 1008 -2432
rect 1045 -2436 1049 -2432
rect 1184 -2400 1188 -2396
rect 1062 -2444 1066 -2440
rect 1184 -2444 1188 -2440
rect 862 -2515 866 -2511
rect 879 -2515 883 -2511
rect 899 -2515 903 -2511
rect 920 -2515 924 -2511
rect 941 -2515 945 -2511
rect 962 -2515 966 -2511
rect 983 -2515 987 -2511
rect 1004 -2515 1008 -2511
rect 1025 -2515 1029 -2511
rect 1045 -2515 1049 -2511
rect 839 -2571 843 -2567
rect 853 -2578 857 -2574
rect 911 -2571 915 -2567
rect 953 -2578 957 -2574
rect 971 -2571 975 -2567
rect 1013 -2563 1017 -2559
rect 1013 -2571 1017 -2567
rect 995 -2585 999 -2581
rect 895 -2592 899 -2588
rect 937 -2592 941 -2588
rect 1062 -2563 1066 -2559
rect 1037 -2578 1041 -2574
rect 862 -2607 866 -2603
rect 879 -2607 883 -2603
rect 920 -2607 924 -2603
rect 962 -2607 966 -2603
rect 1004 -2607 1008 -2603
rect 1045 -2607 1049 -2603
rect 853 -2620 857 -2616
rect 870 -2620 874 -2616
rect 824 -2819 828 -2815
rect 810 -2834 814 -2830
rect 742 -2878 746 -2874
rect 823 -2878 827 -2874
rect 504 -3069 508 -3065
rect 521 -3069 525 -3065
rect 541 -3069 545 -3065
rect 562 -3069 566 -3065
rect 583 -3069 587 -3065
rect 604 -3069 608 -3065
rect 625 -3069 629 -3065
rect 646 -3069 650 -3065
rect 667 -3069 671 -3065
rect 687 -3069 691 -3065
rect 495 -3132 499 -3128
rect 553 -3125 557 -3121
rect 595 -3132 599 -3128
rect 613 -3125 617 -3121
rect 655 -3117 659 -3113
rect 655 -3125 659 -3121
rect 637 -3139 641 -3135
rect 537 -3146 541 -3142
rect 579 -3146 583 -3142
rect 701 -3117 705 -3113
rect 679 -3132 683 -3128
rect 504 -3161 508 -3157
rect 521 -3161 525 -3157
rect 562 -3161 566 -3157
rect 604 -3161 608 -3157
rect 646 -3161 650 -3157
rect 687 -3161 691 -3157
rect 823 -3125 827 -3121
rect 701 -3168 705 -3164
rect 823 -3168 827 -3164
rect 504 -3240 508 -3236
rect 521 -3240 525 -3236
rect 541 -3240 545 -3236
rect 562 -3240 566 -3236
rect 583 -3240 587 -3236
rect 604 -3240 608 -3236
rect 625 -3240 629 -3236
rect 646 -3240 650 -3236
rect 667 -3240 671 -3236
rect 687 -3240 691 -3236
rect 481 -3296 485 -3292
rect 495 -3303 499 -3299
rect 553 -3296 557 -3292
rect 595 -3303 599 -3299
rect 613 -3296 617 -3292
rect 655 -3288 659 -3284
rect 655 -3296 659 -3292
rect 637 -3310 641 -3306
rect 537 -3317 541 -3313
rect 579 -3317 583 -3313
rect 705 -3288 709 -3284
rect 679 -3303 683 -3299
rect 504 -3332 508 -3328
rect 521 -3332 525 -3328
rect 562 -3332 566 -3328
rect 604 -3332 608 -3328
rect 646 -3332 650 -3328
rect 687 -3332 691 -3328
rect 495 -3351 499 -3347
rect 512 -3351 516 -3347
rect 465 -3550 469 -3546
rect 451 -3565 455 -3561
rect 388 -3616 392 -3612
rect 465 -3616 469 -3612
rect 148 -3811 152 -3807
rect 165 -3811 169 -3807
rect 185 -3811 189 -3807
rect 206 -3811 210 -3807
rect 227 -3811 231 -3807
rect 248 -3811 252 -3807
rect 269 -3811 273 -3807
rect 290 -3811 294 -3807
rect 311 -3811 315 -3807
rect 331 -3811 335 -3807
rect 139 -3874 143 -3870
rect 197 -3867 201 -3863
rect 239 -3874 243 -3870
rect 257 -3867 261 -3863
rect 299 -3859 303 -3855
rect 299 -3867 303 -3863
rect 281 -3881 285 -3877
rect 181 -3888 185 -3884
rect 223 -3888 227 -3884
rect 349 -3859 353 -3855
rect 323 -3874 327 -3870
rect 148 -3903 152 -3899
rect 165 -3903 169 -3899
rect 206 -3903 210 -3899
rect 248 -3903 252 -3899
rect 290 -3903 294 -3899
rect 331 -3903 335 -3899
rect 465 -3867 469 -3863
rect 349 -3910 353 -3906
rect 465 -3911 469 -3907
rect 148 -3986 152 -3982
rect 165 -3986 169 -3982
rect 185 -3986 189 -3982
rect 206 -3986 210 -3982
rect 227 -3986 231 -3982
rect 248 -3986 252 -3982
rect 269 -3986 273 -3982
rect 290 -3986 294 -3982
rect 311 -3986 315 -3982
rect 331 -3986 335 -3982
rect 125 -4042 129 -4038
rect 139 -4049 143 -4045
rect 197 -4042 201 -4038
rect 239 -4049 243 -4045
rect 257 -4042 261 -4038
rect 299 -4034 303 -4030
rect 299 -4042 303 -4038
rect 281 -4056 285 -4052
rect 181 -4063 185 -4059
rect 223 -4063 227 -4059
rect 348 -4034 352 -4030
rect 323 -4049 327 -4045
rect 148 -4078 152 -4074
rect 165 -4078 169 -4074
rect 206 -4078 210 -4074
rect 248 -4078 252 -4074
rect 290 -4078 294 -4074
rect 331 -4078 335 -4074
rect 139 -4101 143 -4097
rect 156 -4101 160 -4097
rect 111 -4300 115 -4296
rect 97 -4315 101 -4311
rect 29 -4359 33 -4355
rect 111 -4359 115 -4355
rect -210 -4554 -206 -4550
rect -193 -4554 -189 -4550
rect -173 -4554 -169 -4550
rect -152 -4554 -148 -4550
rect -131 -4554 -127 -4550
rect -110 -4554 -106 -4550
rect -89 -4554 -85 -4550
rect -68 -4554 -64 -4550
rect -47 -4554 -43 -4550
rect -27 -4554 -23 -4550
rect -219 -4617 -215 -4613
rect -161 -4610 -157 -4606
rect -119 -4617 -115 -4613
rect -101 -4610 -97 -4606
rect -59 -4602 -55 -4598
rect -59 -4610 -55 -4606
rect -77 -4624 -73 -4620
rect -177 -4631 -173 -4627
rect -135 -4631 -131 -4627
rect -9 -4602 -5 -4598
rect -35 -4617 -31 -4613
rect -210 -4646 -206 -4642
rect -193 -4646 -189 -4642
rect -152 -4646 -148 -4642
rect -110 -4646 -106 -4642
rect -68 -4646 -64 -4642
rect -27 -4646 -23 -4642
rect 111 -4610 115 -4606
rect -9 -4653 -5 -4649
rect 111 -4655 115 -4651
rect -210 -4725 -206 -4721
rect -193 -4725 -189 -4721
rect -173 -4725 -169 -4721
rect -152 -4725 -148 -4721
rect -131 -4725 -127 -4721
rect -110 -4725 -106 -4721
rect -89 -4725 -85 -4721
rect -68 -4725 -64 -4721
rect -47 -4725 -43 -4721
rect -27 -4725 -23 -4721
rect -233 -4781 -229 -4777
rect -219 -4788 -215 -4784
rect -161 -4781 -157 -4777
rect -119 -4788 -115 -4784
rect -101 -4781 -97 -4777
rect -59 -4773 -55 -4769
rect -59 -4781 -55 -4777
rect -77 -4795 -73 -4791
rect -177 -4802 -173 -4798
rect -135 -4802 -131 -4798
rect -11 -4773 -7 -4769
rect -35 -4788 -31 -4784
rect -210 -4817 -206 -4813
rect -193 -4817 -189 -4813
rect -152 -4817 -148 -4813
rect -110 -4817 -106 -4813
rect -68 -4817 -64 -4813
rect -27 -4817 -23 -4813
rect -219 -4840 -215 -4836
rect -202 -4840 -198 -4836
rect -249 -5039 -245 -5035
rect -263 -5054 -259 -5050
rect -328 -5105 -324 -5101
rect -249 -5105 -245 -5101
rect -568 -5289 -564 -5285
rect -551 -5289 -547 -5285
rect -531 -5289 -527 -5285
rect -510 -5289 -506 -5285
rect -489 -5289 -485 -5285
rect -468 -5289 -464 -5285
rect -447 -5289 -443 -5285
rect -426 -5289 -422 -5285
rect -405 -5289 -401 -5285
rect -385 -5289 -381 -5285
rect -577 -5352 -573 -5348
rect -519 -5345 -515 -5341
rect -477 -5352 -473 -5348
rect -459 -5345 -455 -5341
rect -417 -5337 -413 -5333
rect -417 -5345 -413 -5341
rect -435 -5359 -431 -5355
rect -535 -5366 -531 -5362
rect -493 -5366 -489 -5362
rect -369 -5337 -365 -5333
rect -393 -5352 -389 -5348
rect -568 -5381 -564 -5377
rect -551 -5381 -547 -5377
rect -510 -5381 -506 -5377
rect -468 -5381 -464 -5377
rect -426 -5381 -422 -5377
rect -385 -5381 -381 -5377
rect -249 -5345 -245 -5341
rect -369 -5389 -365 -5385
rect -249 -5388 -245 -5384
rect -568 -5449 -564 -5445
rect -551 -5449 -547 -5445
rect -531 -5449 -527 -5445
rect -510 -5449 -506 -5445
rect -489 -5449 -485 -5445
rect -468 -5449 -464 -5445
rect -447 -5449 -443 -5445
rect -426 -5449 -422 -5445
rect -405 -5449 -401 -5445
rect -385 -5449 -381 -5445
rect -591 -5505 -587 -5501
rect -577 -5512 -573 -5508
rect -519 -5505 -515 -5501
rect -477 -5512 -473 -5508
rect -459 -5505 -455 -5501
rect -417 -5497 -413 -5493
rect -417 -5505 -413 -5501
rect -435 -5519 -431 -5515
rect -535 -5526 -531 -5522
rect -493 -5526 -489 -5522
rect -368 -5497 -364 -5493
rect -393 -5512 -389 -5508
rect -568 -5541 -564 -5537
rect -551 -5541 -547 -5537
rect -510 -5541 -506 -5537
rect -468 -5541 -464 -5537
rect -426 -5541 -422 -5537
rect -385 -5541 -381 -5537
rect -577 -5563 -573 -5559
rect -560 -5563 -556 -5559
rect -368 -5595 -364 -5591
rect -551 -5616 -547 -5612
rect -263 -5616 -259 -5612
rect -560 -5655 -556 -5651
rect -568 -5722 -564 -5718
rect -542 -5722 -538 -5718
rect -525 -5722 -521 -5718
rect -485 -5722 -481 -5718
rect -464 -5722 -460 -5718
rect -447 -5722 -443 -5718
rect -407 -5722 -403 -5718
rect -383 -5722 -379 -5718
rect -346 -5722 -342 -5718
rect -603 -5762 -599 -5758
rect -577 -5755 -573 -5751
rect -616 -5777 -612 -5773
rect -559 -5748 -555 -5744
rect -533 -5770 -529 -5766
rect -551 -5777 -547 -5773
rect -507 -5762 -503 -5758
rect -455 -5755 -451 -5751
rect -525 -5799 -521 -5795
rect -489 -5799 -485 -5795
rect -429 -5770 -425 -5766
rect -447 -5799 -443 -5795
rect -411 -5799 -407 -5795
rect -337 -5761 -333 -5757
rect -326 -5770 -322 -5766
rect -568 -5814 -564 -5810
rect -542 -5814 -538 -5810
rect -499 -5814 -495 -5810
rect -464 -5814 -460 -5810
rect -420 -5814 -416 -5810
rect -403 -5814 -399 -5810
rect -367 -5814 -363 -5810
rect -346 -5814 -342 -5810
rect -11 -4872 -7 -4868
rect -193 -4893 -189 -4889
rect 97 -4893 101 -4889
rect -202 -4932 -198 -4928
rect -210 -4999 -206 -4995
rect -184 -4999 -180 -4995
rect -167 -4999 -163 -4995
rect -127 -4999 -123 -4995
rect -106 -4999 -102 -4995
rect -89 -4999 -85 -4995
rect -49 -4999 -45 -4995
rect -25 -4999 -21 -4995
rect 12 -4999 16 -4995
rect -219 -5032 -215 -5028
rect -201 -5025 -197 -5021
rect -175 -5047 -171 -5043
rect -193 -5054 -189 -5050
rect -149 -5039 -145 -5035
rect -97 -5032 -93 -5028
rect -167 -5076 -163 -5072
rect -131 -5076 -127 -5072
rect -71 -5047 -67 -5043
rect -89 -5076 -85 -5072
rect -53 -5076 -49 -5072
rect 21 -5039 25 -5035
rect 29 -5047 33 -5043
rect -210 -5091 -206 -5087
rect -184 -5091 -180 -5087
rect -141 -5091 -137 -5087
rect -106 -5091 -102 -5087
rect -62 -5091 -58 -5087
rect -45 -5091 -41 -5087
rect -9 -5091 -5 -5087
rect 12 -5091 16 -5087
rect 348 -4133 352 -4129
rect 165 -4154 169 -4150
rect 451 -4154 455 -4150
rect 156 -4193 160 -4189
rect 148 -4260 152 -4256
rect 174 -4260 178 -4256
rect 191 -4260 195 -4256
rect 231 -4260 235 -4256
rect 252 -4260 256 -4256
rect 269 -4260 273 -4256
rect 309 -4260 313 -4256
rect 333 -4260 337 -4256
rect 370 -4260 374 -4256
rect 139 -4293 143 -4289
rect 157 -4286 161 -4282
rect 183 -4308 187 -4304
rect 165 -4315 169 -4311
rect 209 -4300 213 -4296
rect 261 -4293 265 -4289
rect 191 -4337 195 -4333
rect 227 -4337 231 -4333
rect 287 -4308 291 -4304
rect 269 -4337 273 -4333
rect 305 -4337 309 -4333
rect 379 -4300 383 -4296
rect 388 -4308 392 -4304
rect 148 -4352 152 -4348
rect 174 -4352 178 -4348
rect 217 -4352 221 -4348
rect 252 -4352 256 -4348
rect 296 -4352 300 -4348
rect 313 -4352 317 -4348
rect 349 -4352 353 -4348
rect 370 -4352 374 -4348
rect 705 -3383 709 -3379
rect 521 -3404 525 -3400
rect 809 -3404 813 -3400
rect 512 -3443 516 -3439
rect 1062 -2652 1066 -2648
rect 879 -2673 883 -2669
rect 1167 -2673 1171 -2669
rect 870 -2712 874 -2708
rect 862 -2779 866 -2775
rect 888 -2779 892 -2775
rect 905 -2779 909 -2775
rect 945 -2779 949 -2775
rect 966 -2779 970 -2775
rect 983 -2779 987 -2775
rect 1023 -2779 1027 -2775
rect 1047 -2779 1051 -2775
rect 1084 -2779 1088 -2775
rect 853 -2812 857 -2808
rect 871 -2805 875 -2801
rect 897 -2827 901 -2823
rect 879 -2834 883 -2830
rect 923 -2819 927 -2815
rect 975 -2812 979 -2808
rect 905 -2856 909 -2852
rect 941 -2856 945 -2852
rect 1001 -2827 1005 -2823
rect 983 -2856 987 -2852
rect 1019 -2856 1023 -2852
rect 1093 -2817 1097 -2813
rect 1167 -2819 1171 -2815
rect 1093 -2835 1097 -2831
rect 1103 -2827 1107 -2823
rect 862 -2871 866 -2867
rect 888 -2871 892 -2867
rect 931 -2871 935 -2867
rect 966 -2871 970 -2867
rect 1010 -2871 1014 -2867
rect 1027 -2871 1031 -2867
rect 1063 -2871 1067 -2867
rect 1084 -2871 1088 -2867
rect 1419 -1902 1423 -1898
rect 1237 -1923 1241 -1919
rect 1228 -1962 1232 -1958
rect 1220 -2029 1224 -2025
rect 1246 -2029 1250 -2025
rect 1263 -2029 1267 -2025
rect 1303 -2029 1307 -2025
rect 1324 -2029 1328 -2025
rect 1341 -2029 1345 -2025
rect 1381 -2029 1385 -2025
rect 1405 -2029 1409 -2025
rect 1442 -2029 1446 -2025
rect 1211 -2062 1215 -2058
rect 1229 -2055 1233 -2051
rect 1255 -2077 1259 -2073
rect 1237 -2084 1241 -2080
rect 1281 -2069 1285 -2065
rect 1333 -2062 1337 -2058
rect 1263 -2106 1267 -2102
rect 1299 -2106 1303 -2102
rect 1359 -2077 1363 -2073
rect 1341 -2106 1345 -2102
rect 1377 -2106 1381 -2102
rect 1220 -2121 1224 -2117
rect 1246 -2121 1250 -2117
rect 1289 -2121 1293 -2117
rect 1324 -2121 1328 -2117
rect 1368 -2121 1372 -2117
rect 1385 -2121 1389 -2117
rect 1421 -2121 1425 -2117
rect 1442 -2121 1446 -2117
rect 1466 -2077 1470 -2073
rect 1466 -2128 1470 -2124
rect 1451 -2135 1455 -2131
rect 1220 -2344 1224 -2340
rect 1237 -2344 1241 -2340
rect 1257 -2344 1261 -2340
rect 1278 -2344 1282 -2340
rect 1299 -2344 1303 -2340
rect 1320 -2344 1324 -2340
rect 1341 -2344 1345 -2340
rect 1362 -2344 1366 -2340
rect 1383 -2344 1387 -2340
rect 1403 -2344 1407 -2340
rect 1211 -2407 1215 -2403
rect 1269 -2400 1273 -2396
rect 1311 -2407 1315 -2403
rect 1329 -2400 1333 -2396
rect 1371 -2392 1375 -2388
rect 1371 -2400 1375 -2396
rect 1353 -2414 1357 -2410
rect 1253 -2421 1257 -2417
rect 1295 -2421 1299 -2417
rect 1421 -2392 1425 -2388
rect 1395 -2407 1399 -2403
rect 1220 -2436 1224 -2432
rect 1237 -2436 1241 -2432
rect 1278 -2436 1282 -2432
rect 1320 -2436 1324 -2432
rect 1362 -2436 1366 -2432
rect 1403 -2436 1407 -2432
rect 1421 -2444 1425 -2440
rect 1220 -2515 1224 -2511
rect 1237 -2515 1241 -2511
rect 1257 -2515 1261 -2511
rect 1278 -2515 1282 -2511
rect 1299 -2515 1303 -2511
rect 1320 -2515 1324 -2511
rect 1341 -2515 1345 -2511
rect 1362 -2515 1366 -2511
rect 1383 -2515 1387 -2511
rect 1403 -2515 1407 -2511
rect 1197 -2571 1201 -2567
rect 1211 -2578 1215 -2574
rect 1269 -2571 1273 -2567
rect 1311 -2578 1315 -2574
rect 1329 -2571 1333 -2567
rect 1371 -2563 1375 -2559
rect 1371 -2571 1375 -2567
rect 1353 -2585 1357 -2581
rect 1253 -2592 1257 -2588
rect 1295 -2592 1299 -2588
rect 1419 -2563 1423 -2559
rect 1395 -2578 1399 -2574
rect 1220 -2607 1224 -2603
rect 1237 -2607 1241 -2603
rect 1278 -2607 1282 -2603
rect 1320 -2607 1324 -2603
rect 1362 -2607 1366 -2603
rect 1403 -2607 1407 -2603
rect 1211 -2620 1215 -2616
rect 1228 -2620 1232 -2616
rect 1184 -2834 1188 -2830
rect 1103 -2885 1107 -2881
rect 1184 -2885 1188 -2881
rect 862 -3069 866 -3065
rect 879 -3069 883 -3065
rect 899 -3069 903 -3065
rect 920 -3069 924 -3065
rect 941 -3069 945 -3065
rect 962 -3069 966 -3065
rect 983 -3069 987 -3065
rect 1004 -3069 1008 -3065
rect 1025 -3069 1029 -3065
rect 1045 -3069 1049 -3065
rect 853 -3132 857 -3128
rect 911 -3125 915 -3121
rect 953 -3132 957 -3128
rect 971 -3125 975 -3121
rect 1013 -3117 1017 -3113
rect 1013 -3125 1017 -3121
rect 995 -3139 999 -3135
rect 895 -3146 899 -3142
rect 937 -3146 941 -3142
rect 1060 -3117 1064 -3113
rect 1037 -3132 1041 -3128
rect 862 -3161 866 -3157
rect 879 -3161 883 -3157
rect 920 -3161 924 -3157
rect 962 -3161 966 -3157
rect 1004 -3161 1008 -3157
rect 1045 -3161 1049 -3157
rect 1184 -3125 1188 -3121
rect 1060 -3168 1064 -3164
rect 1184 -3169 1188 -3165
rect 862 -3240 866 -3236
rect 879 -3240 883 -3236
rect 899 -3240 903 -3236
rect 920 -3240 924 -3236
rect 941 -3240 945 -3236
rect 962 -3240 966 -3236
rect 983 -3240 987 -3236
rect 1004 -3240 1008 -3236
rect 1025 -3240 1029 -3236
rect 1045 -3240 1049 -3236
rect 839 -3296 843 -3292
rect 853 -3303 857 -3299
rect 911 -3296 915 -3292
rect 953 -3303 957 -3299
rect 971 -3296 975 -3292
rect 1013 -3288 1017 -3284
rect 1013 -3296 1017 -3292
rect 995 -3310 999 -3306
rect 895 -3317 899 -3313
rect 937 -3317 941 -3313
rect 1066 -3288 1070 -3284
rect 1037 -3303 1041 -3299
rect 862 -3332 866 -3328
rect 879 -3332 883 -3328
rect 920 -3332 924 -3328
rect 962 -3332 966 -3328
rect 1004 -3332 1008 -3328
rect 1045 -3332 1049 -3328
rect 853 -3351 857 -3347
rect 870 -3351 874 -3347
rect 504 -3510 508 -3506
rect 530 -3510 534 -3506
rect 547 -3510 551 -3506
rect 587 -3510 591 -3506
rect 608 -3510 612 -3506
rect 625 -3510 629 -3506
rect 665 -3510 669 -3506
rect 689 -3510 693 -3506
rect 726 -3510 730 -3506
rect 495 -3543 499 -3539
rect 513 -3536 517 -3532
rect 539 -3558 543 -3554
rect 521 -3565 525 -3561
rect 565 -3550 569 -3546
rect 617 -3543 621 -3539
rect 547 -3587 551 -3583
rect 583 -3587 587 -3583
rect 643 -3558 647 -3554
rect 625 -3587 629 -3583
rect 661 -3587 665 -3583
rect 735 -3550 739 -3546
rect 743 -3558 747 -3554
rect 504 -3602 508 -3598
rect 530 -3602 534 -3598
rect 573 -3602 577 -3598
rect 608 -3602 612 -3598
rect 652 -3602 656 -3598
rect 669 -3602 673 -3598
rect 705 -3602 709 -3598
rect 726 -3602 730 -3598
rect 824 -3550 828 -3546
rect 810 -3565 814 -3561
rect 743 -3609 747 -3605
rect 824 -3609 828 -3605
rect 504 -3811 508 -3807
rect 521 -3811 525 -3807
rect 541 -3811 545 -3807
rect 562 -3811 566 -3807
rect 583 -3811 587 -3807
rect 604 -3811 608 -3807
rect 625 -3811 629 -3807
rect 646 -3811 650 -3807
rect 667 -3811 671 -3807
rect 687 -3811 691 -3807
rect 495 -3874 499 -3870
rect 553 -3867 557 -3863
rect 595 -3874 599 -3870
rect 613 -3867 617 -3863
rect 655 -3859 659 -3855
rect 655 -3867 659 -3863
rect 637 -3881 641 -3877
rect 537 -3888 541 -3884
rect 579 -3888 583 -3884
rect 702 -3859 706 -3855
rect 679 -3874 683 -3870
rect 504 -3903 508 -3899
rect 521 -3903 525 -3899
rect 562 -3903 566 -3899
rect 604 -3903 608 -3899
rect 646 -3903 650 -3899
rect 687 -3903 691 -3899
rect 824 -3867 828 -3863
rect 702 -3911 706 -3907
rect 824 -3910 828 -3906
rect 504 -3986 508 -3982
rect 521 -3986 525 -3982
rect 541 -3986 545 -3982
rect 562 -3986 566 -3982
rect 583 -3986 587 -3982
rect 604 -3986 608 -3982
rect 625 -3986 629 -3982
rect 646 -3986 650 -3982
rect 667 -3986 671 -3982
rect 687 -3986 691 -3982
rect 481 -4042 485 -4038
rect 495 -4049 499 -4045
rect 553 -4042 557 -4038
rect 595 -4049 599 -4045
rect 613 -4042 617 -4038
rect 655 -4034 659 -4030
rect 655 -4042 659 -4038
rect 637 -4056 641 -4052
rect 537 -4063 541 -4059
rect 579 -4063 583 -4059
rect 705 -4034 709 -4030
rect 679 -4049 683 -4045
rect 504 -4078 508 -4074
rect 521 -4078 525 -4074
rect 562 -4078 566 -4074
rect 604 -4078 608 -4074
rect 646 -4078 650 -4074
rect 687 -4078 691 -4074
rect 495 -4101 499 -4097
rect 512 -4101 516 -4097
rect 465 -4300 469 -4296
rect 451 -4315 455 -4311
rect 388 -4366 392 -4362
rect 465 -4366 469 -4362
rect 148 -4554 152 -4550
rect 165 -4554 169 -4550
rect 185 -4554 189 -4550
rect 206 -4554 210 -4550
rect 227 -4554 231 -4550
rect 248 -4554 252 -4550
rect 269 -4554 273 -4550
rect 290 -4554 294 -4550
rect 311 -4554 315 -4550
rect 331 -4554 335 -4550
rect 139 -4617 143 -4613
rect 197 -4610 201 -4606
rect 239 -4617 243 -4613
rect 257 -4610 261 -4606
rect 299 -4602 303 -4598
rect 299 -4610 303 -4606
rect 281 -4624 285 -4620
rect 181 -4631 185 -4627
rect 223 -4631 227 -4627
rect 348 -4602 352 -4598
rect 323 -4617 327 -4613
rect 148 -4646 152 -4642
rect 165 -4646 169 -4642
rect 206 -4646 210 -4642
rect 248 -4646 252 -4642
rect 290 -4646 294 -4642
rect 331 -4646 335 -4642
rect 465 -4610 469 -4606
rect 348 -4655 352 -4651
rect 465 -4654 469 -4650
rect 148 -4725 152 -4721
rect 165 -4725 169 -4721
rect 185 -4725 189 -4721
rect 206 -4725 210 -4721
rect 227 -4725 231 -4721
rect 248 -4725 252 -4721
rect 269 -4725 273 -4721
rect 290 -4725 294 -4721
rect 311 -4725 315 -4721
rect 331 -4725 335 -4721
rect 125 -4781 129 -4777
rect 139 -4788 143 -4784
rect 197 -4781 201 -4777
rect 239 -4788 243 -4784
rect 257 -4781 261 -4777
rect 299 -4773 303 -4769
rect 299 -4781 303 -4777
rect 281 -4795 285 -4791
rect 181 -4802 185 -4798
rect 223 -4802 227 -4798
rect 347 -4773 351 -4769
rect 323 -4788 327 -4784
rect 148 -4817 152 -4813
rect 165 -4817 169 -4813
rect 206 -4817 210 -4813
rect 248 -4817 252 -4813
rect 290 -4817 294 -4813
rect 331 -4817 335 -4813
rect 139 -4840 143 -4836
rect 156 -4840 160 -4836
rect 111 -5039 115 -5035
rect 97 -5054 101 -5050
rect 29 -5098 33 -5094
rect 108 -5098 112 -5094
rect -210 -5289 -206 -5285
rect -193 -5289 -189 -5285
rect -173 -5289 -169 -5285
rect -152 -5289 -148 -5285
rect -131 -5289 -127 -5285
rect -110 -5289 -106 -5285
rect -89 -5289 -85 -5285
rect -68 -5289 -64 -5285
rect -47 -5289 -43 -5285
rect -27 -5289 -23 -5285
rect -219 -5352 -215 -5348
rect -161 -5345 -157 -5341
rect -119 -5352 -115 -5348
rect -101 -5345 -97 -5341
rect -59 -5337 -55 -5333
rect -59 -5345 -55 -5341
rect -77 -5359 -73 -5355
rect -177 -5366 -173 -5362
rect -135 -5366 -131 -5362
rect -7 -5337 -3 -5333
rect -35 -5352 -31 -5348
rect -210 -5381 -206 -5377
rect -193 -5381 -189 -5377
rect -152 -5381 -148 -5377
rect -110 -5381 -106 -5377
rect -68 -5381 -64 -5377
rect -27 -5381 -23 -5377
rect 108 -5345 112 -5341
rect -7 -5388 -3 -5384
rect 108 -5388 112 -5384
rect -210 -5449 -206 -5445
rect -193 -5449 -189 -5445
rect -173 -5449 -169 -5445
rect -152 -5449 -148 -5445
rect -131 -5449 -127 -5445
rect -110 -5449 -106 -5445
rect -89 -5449 -85 -5445
rect -68 -5449 -64 -5445
rect -47 -5449 -43 -5445
rect -27 -5449 -23 -5445
rect -233 -5505 -229 -5501
rect -219 -5512 -215 -5508
rect -161 -5505 -157 -5501
rect -119 -5512 -115 -5508
rect -101 -5505 -97 -5501
rect -59 -5497 -55 -5493
rect -59 -5505 -55 -5501
rect -77 -5519 -73 -5515
rect -177 -5526 -173 -5522
rect -135 -5526 -131 -5522
rect -12 -5497 -8 -5493
rect -35 -5512 -31 -5508
rect -210 -5541 -206 -5537
rect -193 -5541 -189 -5537
rect -152 -5541 -148 -5537
rect -110 -5541 -106 -5537
rect -68 -5541 -64 -5537
rect -27 -5541 -23 -5537
rect -219 -5563 -215 -5559
rect -202 -5563 -198 -5559
rect -12 -5595 -8 -5591
rect -193 -5616 -189 -5612
rect 97 -5616 101 -5612
rect -202 -5655 -198 -5651
rect -210 -5722 -206 -5718
rect -184 -5722 -180 -5718
rect -167 -5722 -163 -5718
rect -127 -5722 -123 -5718
rect -106 -5722 -102 -5718
rect -89 -5722 -85 -5718
rect -49 -5722 -45 -5718
rect -25 -5722 -21 -5718
rect 12 -5722 16 -5718
rect -249 -5762 -245 -5758
rect -219 -5755 -215 -5751
rect -263 -5777 -259 -5773
rect -201 -5748 -197 -5744
rect -175 -5770 -171 -5766
rect -193 -5777 -189 -5773
rect -149 -5762 -145 -5758
rect -97 -5755 -93 -5751
rect -167 -5799 -163 -5795
rect -131 -5799 -127 -5795
rect -71 -5770 -67 -5766
rect -89 -5799 -85 -5795
rect -53 -5799 -49 -5795
rect 21 -5762 25 -5758
rect 33 -5770 37 -5766
rect -210 -5814 -206 -5810
rect -184 -5814 -180 -5810
rect -141 -5814 -137 -5810
rect -106 -5814 -102 -5810
rect -62 -5814 -58 -5810
rect -45 -5814 -41 -5810
rect -9 -5814 -5 -5810
rect 12 -5814 16 -5810
rect 347 -4872 351 -4868
rect 165 -4893 169 -4889
rect 451 -4893 455 -4889
rect 156 -4932 160 -4928
rect 148 -4999 152 -4995
rect 174 -4999 178 -4995
rect 191 -4999 195 -4995
rect 231 -4999 235 -4995
rect 252 -4999 256 -4995
rect 269 -4999 273 -4995
rect 309 -4999 313 -4995
rect 333 -4999 337 -4995
rect 370 -4999 374 -4995
rect 139 -5032 143 -5028
rect 157 -5025 161 -5021
rect 183 -5047 187 -5043
rect 165 -5054 169 -5050
rect 209 -5039 213 -5035
rect 261 -5032 265 -5028
rect 191 -5076 195 -5072
rect 227 -5076 231 -5072
rect 287 -5047 291 -5043
rect 269 -5076 273 -5072
rect 305 -5076 309 -5072
rect 379 -5039 383 -5035
rect 388 -5047 392 -5043
rect 148 -5091 152 -5087
rect 174 -5091 178 -5087
rect 217 -5091 221 -5087
rect 252 -5091 256 -5087
rect 296 -5091 300 -5087
rect 313 -5091 317 -5087
rect 349 -5091 353 -5087
rect 370 -5091 374 -5087
rect 705 -4133 709 -4129
rect 521 -4154 525 -4150
rect 810 -4154 814 -4150
rect 512 -4193 516 -4189
rect 504 -4260 508 -4256
rect 530 -4260 534 -4256
rect 547 -4260 551 -4256
rect 587 -4260 591 -4256
rect 608 -4260 612 -4256
rect 625 -4260 629 -4256
rect 665 -4260 669 -4256
rect 689 -4260 693 -4256
rect 726 -4260 730 -4256
rect 495 -4293 499 -4289
rect 513 -4286 517 -4282
rect 539 -4308 543 -4304
rect 521 -4315 525 -4311
rect 565 -4300 569 -4296
rect 617 -4293 621 -4289
rect 547 -4337 551 -4333
rect 583 -4337 587 -4333
rect 643 -4308 647 -4304
rect 625 -4337 629 -4333
rect 661 -4337 665 -4333
rect 735 -4300 739 -4296
rect 743 -4308 747 -4304
rect 504 -4352 508 -4348
rect 530 -4352 534 -4348
rect 573 -4352 577 -4348
rect 608 -4352 612 -4348
rect 652 -4352 656 -4348
rect 669 -4352 673 -4348
rect 705 -4352 709 -4348
rect 726 -4352 730 -4348
rect 1066 -3383 1070 -3379
rect 879 -3404 883 -3400
rect 1167 -3404 1171 -3400
rect 870 -3443 874 -3439
rect 862 -3510 866 -3506
rect 888 -3510 892 -3506
rect 905 -3510 909 -3506
rect 945 -3510 949 -3506
rect 966 -3510 970 -3506
rect 983 -3510 987 -3506
rect 1023 -3510 1027 -3506
rect 1047 -3510 1051 -3506
rect 1084 -3510 1088 -3506
rect 853 -3543 857 -3539
rect 871 -3536 875 -3532
rect 897 -3558 901 -3554
rect 879 -3565 883 -3561
rect 923 -3550 927 -3546
rect 975 -3543 979 -3539
rect 905 -3587 909 -3583
rect 941 -3587 945 -3583
rect 1001 -3558 1005 -3554
rect 983 -3587 987 -3583
rect 1019 -3587 1023 -3583
rect 1093 -3548 1097 -3544
rect 1167 -3550 1171 -3546
rect 1101 -3558 1105 -3554
rect 862 -3602 866 -3598
rect 888 -3602 892 -3598
rect 931 -3602 935 -3598
rect 966 -3602 970 -3598
rect 1010 -3602 1014 -3598
rect 1027 -3602 1031 -3598
rect 1063 -3602 1067 -3598
rect 1084 -3602 1088 -3598
rect 1419 -2652 1423 -2648
rect 1237 -2673 1241 -2669
rect 1228 -2712 1232 -2708
rect 1220 -2779 1224 -2775
rect 1246 -2779 1250 -2775
rect 1263 -2779 1267 -2775
rect 1303 -2779 1307 -2775
rect 1324 -2779 1328 -2775
rect 1341 -2779 1345 -2775
rect 1381 -2779 1385 -2775
rect 1405 -2779 1409 -2775
rect 1442 -2779 1446 -2775
rect 1211 -2812 1215 -2808
rect 1229 -2805 1233 -2801
rect 1255 -2827 1259 -2823
rect 1237 -2834 1241 -2830
rect 1281 -2819 1285 -2815
rect 1333 -2812 1337 -2808
rect 1263 -2856 1267 -2852
rect 1299 -2856 1303 -2852
rect 1359 -2827 1363 -2823
rect 1341 -2856 1345 -2852
rect 1377 -2856 1381 -2852
rect 1220 -2871 1224 -2867
rect 1246 -2871 1250 -2867
rect 1289 -2871 1293 -2867
rect 1324 -2871 1328 -2867
rect 1368 -2871 1372 -2867
rect 1385 -2871 1389 -2867
rect 1421 -2871 1425 -2867
rect 1442 -2871 1446 -2867
rect 1467 -2827 1471 -2823
rect 1467 -2878 1471 -2874
rect 1451 -2885 1455 -2881
rect 1220 -3069 1224 -3065
rect 1237 -3069 1241 -3065
rect 1257 -3069 1261 -3065
rect 1278 -3069 1282 -3065
rect 1299 -3069 1303 -3065
rect 1320 -3069 1324 -3065
rect 1341 -3069 1345 -3065
rect 1362 -3069 1366 -3065
rect 1383 -3069 1387 -3065
rect 1403 -3069 1407 -3065
rect 1211 -3132 1215 -3128
rect 1269 -3125 1273 -3121
rect 1311 -3132 1315 -3128
rect 1329 -3125 1333 -3121
rect 1371 -3117 1375 -3113
rect 1371 -3125 1375 -3121
rect 1353 -3139 1357 -3135
rect 1253 -3146 1257 -3142
rect 1295 -3146 1299 -3142
rect 1419 -3117 1423 -3113
rect 1395 -3132 1399 -3128
rect 1220 -3161 1224 -3157
rect 1237 -3161 1241 -3157
rect 1278 -3161 1282 -3157
rect 1320 -3161 1324 -3157
rect 1362 -3161 1366 -3157
rect 1403 -3161 1407 -3157
rect 1419 -3169 1423 -3165
rect 1220 -3240 1224 -3236
rect 1237 -3240 1241 -3236
rect 1257 -3240 1261 -3236
rect 1278 -3240 1282 -3236
rect 1299 -3240 1303 -3236
rect 1320 -3240 1324 -3236
rect 1341 -3240 1345 -3236
rect 1362 -3240 1366 -3236
rect 1383 -3240 1387 -3236
rect 1403 -3240 1407 -3236
rect 1197 -3296 1201 -3292
rect 1211 -3303 1215 -3299
rect 1269 -3296 1273 -3292
rect 1311 -3303 1315 -3299
rect 1329 -3296 1333 -3292
rect 1371 -3288 1375 -3284
rect 1371 -3296 1375 -3292
rect 1353 -3310 1357 -3306
rect 1253 -3317 1257 -3313
rect 1295 -3317 1299 -3313
rect 1422 -3288 1426 -3284
rect 1395 -3303 1399 -3299
rect 1220 -3332 1224 -3328
rect 1237 -3332 1241 -3328
rect 1278 -3332 1282 -3328
rect 1320 -3332 1324 -3328
rect 1362 -3332 1366 -3328
rect 1403 -3332 1407 -3328
rect 1211 -3351 1215 -3347
rect 1228 -3351 1232 -3347
rect 1184 -3565 1188 -3561
rect 1101 -3616 1105 -3612
rect 1184 -3616 1188 -3612
rect 862 -3811 866 -3807
rect 879 -3811 883 -3807
rect 899 -3811 903 -3807
rect 920 -3811 924 -3807
rect 941 -3811 945 -3807
rect 962 -3811 966 -3807
rect 983 -3811 987 -3807
rect 1004 -3811 1008 -3807
rect 1025 -3811 1029 -3807
rect 1045 -3811 1049 -3807
rect 853 -3874 857 -3870
rect 911 -3867 915 -3863
rect 953 -3874 957 -3870
rect 971 -3867 975 -3863
rect 1013 -3859 1017 -3855
rect 1013 -3867 1017 -3863
rect 995 -3881 999 -3877
rect 895 -3888 899 -3884
rect 937 -3888 941 -3884
rect 1060 -3859 1064 -3855
rect 1037 -3874 1041 -3870
rect 862 -3903 866 -3899
rect 879 -3903 883 -3899
rect 920 -3903 924 -3899
rect 962 -3903 966 -3899
rect 1004 -3903 1008 -3899
rect 1045 -3903 1049 -3899
rect 1184 -3867 1188 -3863
rect 1060 -3910 1064 -3906
rect 1184 -3910 1188 -3906
rect 862 -3986 866 -3982
rect 879 -3986 883 -3982
rect 899 -3986 903 -3982
rect 920 -3986 924 -3982
rect 941 -3986 945 -3982
rect 962 -3986 966 -3982
rect 983 -3986 987 -3982
rect 1004 -3986 1008 -3982
rect 1025 -3986 1029 -3982
rect 1045 -3986 1049 -3982
rect 839 -4042 843 -4038
rect 853 -4049 857 -4045
rect 911 -4042 915 -4038
rect 953 -4049 957 -4045
rect 971 -4042 975 -4038
rect 1013 -4034 1017 -4030
rect 1013 -4042 1017 -4038
rect 995 -4056 999 -4052
rect 895 -4063 899 -4059
rect 937 -4063 941 -4059
rect 1063 -4034 1067 -4030
rect 1037 -4049 1041 -4045
rect 862 -4078 866 -4074
rect 879 -4078 883 -4074
rect 920 -4078 924 -4074
rect 962 -4078 966 -4074
rect 1004 -4078 1008 -4074
rect 1045 -4078 1049 -4074
rect 853 -4101 857 -4097
rect 870 -4101 874 -4097
rect 824 -4300 828 -4296
rect 810 -4315 814 -4311
rect 743 -4359 747 -4355
rect 824 -4359 828 -4355
rect 504 -4554 508 -4550
rect 521 -4554 525 -4550
rect 541 -4554 545 -4550
rect 562 -4554 566 -4550
rect 583 -4554 587 -4550
rect 604 -4554 608 -4550
rect 625 -4554 629 -4550
rect 646 -4554 650 -4550
rect 667 -4554 671 -4550
rect 687 -4554 691 -4550
rect 495 -4617 499 -4613
rect 553 -4610 557 -4606
rect 595 -4617 599 -4613
rect 613 -4610 617 -4606
rect 655 -4602 659 -4598
rect 655 -4610 659 -4606
rect 637 -4624 641 -4620
rect 537 -4631 541 -4627
rect 579 -4631 583 -4627
rect 700 -4602 704 -4598
rect 679 -4617 683 -4613
rect 504 -4646 508 -4642
rect 521 -4646 525 -4642
rect 562 -4646 566 -4642
rect 604 -4646 608 -4642
rect 646 -4646 650 -4642
rect 687 -4646 691 -4642
rect 824 -4610 828 -4606
rect 700 -4654 704 -4650
rect 824 -4653 828 -4649
rect 504 -4725 508 -4721
rect 521 -4725 525 -4721
rect 541 -4725 545 -4721
rect 562 -4725 566 -4721
rect 583 -4725 587 -4721
rect 604 -4725 608 -4721
rect 625 -4725 629 -4721
rect 646 -4725 650 -4721
rect 667 -4725 671 -4721
rect 687 -4725 691 -4721
rect 481 -4781 485 -4777
rect 495 -4788 499 -4784
rect 553 -4781 557 -4777
rect 595 -4788 599 -4784
rect 613 -4781 617 -4777
rect 655 -4773 659 -4769
rect 655 -4781 659 -4777
rect 637 -4795 641 -4791
rect 537 -4802 541 -4798
rect 579 -4802 583 -4798
rect 706 -4773 710 -4769
rect 679 -4788 683 -4784
rect 504 -4817 508 -4813
rect 521 -4817 525 -4813
rect 562 -4817 566 -4813
rect 604 -4817 608 -4813
rect 646 -4817 650 -4813
rect 687 -4817 691 -4813
rect 495 -4840 499 -4836
rect 512 -4840 516 -4836
rect 465 -5039 469 -5035
rect 451 -5054 455 -5050
rect 388 -5105 392 -5101
rect 464 -5105 468 -5101
rect 148 -5289 152 -5285
rect 165 -5289 169 -5285
rect 185 -5289 189 -5285
rect 206 -5289 210 -5285
rect 227 -5289 231 -5285
rect 248 -5289 252 -5285
rect 269 -5289 273 -5285
rect 290 -5289 294 -5285
rect 311 -5289 315 -5285
rect 331 -5289 335 -5285
rect 139 -5352 143 -5348
rect 197 -5345 201 -5341
rect 239 -5352 243 -5348
rect 257 -5345 261 -5341
rect 299 -5337 303 -5333
rect 299 -5345 303 -5341
rect 281 -5359 285 -5355
rect 181 -5366 185 -5362
rect 223 -5366 227 -5362
rect 349 -5337 353 -5333
rect 323 -5352 327 -5348
rect 148 -5381 152 -5377
rect 165 -5381 169 -5377
rect 206 -5381 210 -5377
rect 248 -5381 252 -5377
rect 290 -5381 294 -5377
rect 331 -5381 335 -5377
rect 464 -5345 468 -5341
rect 349 -5388 353 -5384
rect 464 -5390 468 -5386
rect 148 -5449 152 -5445
rect 165 -5449 169 -5445
rect 185 -5449 189 -5445
rect 206 -5449 210 -5445
rect 227 -5449 231 -5445
rect 248 -5449 252 -5445
rect 269 -5449 273 -5445
rect 290 -5449 294 -5445
rect 311 -5449 315 -5445
rect 331 -5449 335 -5445
rect 125 -5505 129 -5501
rect 139 -5512 143 -5508
rect 197 -5505 201 -5501
rect 239 -5512 243 -5508
rect 257 -5505 261 -5501
rect 299 -5497 303 -5493
rect 299 -5505 303 -5501
rect 281 -5519 285 -5515
rect 181 -5526 185 -5522
rect 223 -5526 227 -5522
rect 348 -5497 352 -5493
rect 323 -5512 327 -5508
rect 148 -5541 152 -5537
rect 165 -5541 169 -5537
rect 206 -5541 210 -5537
rect 248 -5541 252 -5537
rect 290 -5541 294 -5537
rect 331 -5541 335 -5537
rect 139 -5563 143 -5559
rect 156 -5563 160 -5559
rect 348 -5595 352 -5591
rect 165 -5616 169 -5612
rect 451 -5616 455 -5612
rect 156 -5655 160 -5651
rect 148 -5722 152 -5718
rect 174 -5722 178 -5718
rect 191 -5722 195 -5718
rect 231 -5722 235 -5718
rect 252 -5722 256 -5718
rect 269 -5722 273 -5718
rect 309 -5722 313 -5718
rect 333 -5722 337 -5718
rect 370 -5722 374 -5718
rect 108 -5762 112 -5758
rect 139 -5755 143 -5751
rect 97 -5777 101 -5773
rect 157 -5748 161 -5744
rect 183 -5770 187 -5766
rect 165 -5777 169 -5773
rect 209 -5762 213 -5758
rect 261 -5755 265 -5751
rect 191 -5799 195 -5795
rect 227 -5799 231 -5795
rect 287 -5770 291 -5766
rect 269 -5799 273 -5795
rect 305 -5799 309 -5795
rect 379 -5762 383 -5758
rect 392 -5770 396 -5766
rect 148 -5814 152 -5810
rect 174 -5814 178 -5810
rect 217 -5814 221 -5810
rect 252 -5814 256 -5810
rect 296 -5814 300 -5810
rect 313 -5814 317 -5810
rect 349 -5814 353 -5810
rect 370 -5814 374 -5810
rect -1246 -5824 -1242 -5820
rect -1103 -5824 -1099 -5820
rect -949 -5821 -945 -5817
rect -683 -5821 -679 -5817
rect -586 -5821 -582 -5817
rect -326 -5821 -322 -5817
rect -233 -5821 -229 -5817
rect 33 -5821 37 -5817
rect 706 -4872 710 -4868
rect 521 -4893 525 -4889
rect 810 -4893 814 -4889
rect 512 -4932 516 -4928
rect 504 -4999 508 -4995
rect 530 -4999 534 -4995
rect 547 -4999 551 -4995
rect 587 -4999 591 -4995
rect 608 -4999 612 -4995
rect 625 -4999 629 -4995
rect 665 -4999 669 -4995
rect 689 -4999 693 -4995
rect 726 -4999 730 -4995
rect 495 -5032 499 -5028
rect 513 -5025 517 -5021
rect 539 -5047 543 -5043
rect 521 -5054 525 -5050
rect 565 -5039 569 -5035
rect 617 -5032 621 -5028
rect 547 -5076 551 -5072
rect 583 -5076 587 -5072
rect 643 -5047 647 -5043
rect 625 -5076 629 -5072
rect 661 -5076 665 -5072
rect 735 -5039 739 -5035
rect 743 -5047 747 -5043
rect 504 -5091 508 -5087
rect 530 -5091 534 -5087
rect 573 -5091 577 -5087
rect 608 -5091 612 -5087
rect 652 -5091 656 -5087
rect 669 -5091 673 -5087
rect 705 -5091 709 -5087
rect 726 -5091 730 -5087
rect 1063 -4133 1067 -4129
rect 879 -4154 883 -4150
rect 1167 -4154 1171 -4150
rect 870 -4193 874 -4189
rect 862 -4260 866 -4256
rect 888 -4260 892 -4256
rect 905 -4260 909 -4256
rect 945 -4260 949 -4256
rect 966 -4260 970 -4256
rect 983 -4260 987 -4256
rect 1023 -4260 1027 -4256
rect 1047 -4260 1051 -4256
rect 1084 -4260 1088 -4256
rect 853 -4293 857 -4289
rect 871 -4286 875 -4282
rect 897 -4308 901 -4304
rect 879 -4315 883 -4311
rect 923 -4300 927 -4296
rect 975 -4293 979 -4289
rect 905 -4337 909 -4333
rect 941 -4337 945 -4333
rect 1001 -4308 1005 -4304
rect 983 -4337 987 -4333
rect 1019 -4337 1023 -4333
rect 1093 -4298 1097 -4294
rect 1167 -4300 1171 -4296
rect 1101 -4308 1105 -4304
rect 862 -4352 866 -4348
rect 888 -4352 892 -4348
rect 931 -4352 935 -4348
rect 966 -4352 970 -4348
rect 1010 -4352 1014 -4348
rect 1027 -4352 1031 -4348
rect 1063 -4352 1067 -4348
rect 1084 -4352 1088 -4348
rect 1422 -3383 1426 -3379
rect 1237 -3404 1241 -3400
rect 1228 -3443 1232 -3439
rect 1220 -3510 1224 -3506
rect 1246 -3510 1250 -3506
rect 1263 -3510 1267 -3506
rect 1303 -3510 1307 -3506
rect 1324 -3510 1328 -3506
rect 1341 -3510 1345 -3506
rect 1381 -3510 1385 -3506
rect 1405 -3510 1409 -3506
rect 1442 -3510 1446 -3506
rect 1211 -3543 1215 -3539
rect 1229 -3536 1233 -3532
rect 1255 -3558 1259 -3554
rect 1237 -3565 1241 -3561
rect 1281 -3550 1285 -3546
rect 1333 -3543 1337 -3539
rect 1263 -3587 1267 -3583
rect 1299 -3587 1303 -3583
rect 1359 -3558 1363 -3554
rect 1341 -3587 1345 -3583
rect 1377 -3587 1381 -3583
rect 1220 -3602 1224 -3598
rect 1246 -3602 1250 -3598
rect 1289 -3602 1293 -3598
rect 1324 -3602 1328 -3598
rect 1368 -3602 1372 -3598
rect 1385 -3602 1389 -3598
rect 1421 -3602 1425 -3598
rect 1442 -3602 1446 -3598
rect 1464 -3558 1468 -3554
rect 1464 -3609 1468 -3605
rect 1451 -3616 1455 -3612
rect 1220 -3811 1224 -3807
rect 1237 -3811 1241 -3807
rect 1257 -3811 1261 -3807
rect 1278 -3811 1282 -3807
rect 1299 -3811 1303 -3807
rect 1320 -3811 1324 -3807
rect 1341 -3811 1345 -3807
rect 1362 -3811 1366 -3807
rect 1383 -3811 1387 -3807
rect 1403 -3811 1407 -3807
rect 1211 -3874 1215 -3870
rect 1269 -3867 1273 -3863
rect 1311 -3874 1315 -3870
rect 1329 -3867 1333 -3863
rect 1371 -3859 1375 -3855
rect 1371 -3867 1375 -3863
rect 1353 -3881 1357 -3877
rect 1253 -3888 1257 -3884
rect 1295 -3888 1299 -3884
rect 1424 -3859 1428 -3855
rect 1395 -3874 1399 -3870
rect 1220 -3903 1224 -3899
rect 1237 -3903 1241 -3899
rect 1278 -3903 1282 -3899
rect 1320 -3903 1324 -3899
rect 1362 -3903 1366 -3899
rect 1403 -3903 1407 -3899
rect 1424 -3910 1428 -3906
rect 1220 -3986 1224 -3982
rect 1237 -3986 1241 -3982
rect 1257 -3986 1261 -3982
rect 1278 -3986 1282 -3982
rect 1299 -3986 1303 -3982
rect 1320 -3986 1324 -3982
rect 1341 -3986 1345 -3982
rect 1362 -3986 1366 -3982
rect 1383 -3986 1387 -3982
rect 1403 -3986 1407 -3982
rect 1197 -4042 1201 -4038
rect 1211 -4049 1215 -4045
rect 1269 -4042 1273 -4038
rect 1311 -4049 1315 -4045
rect 1329 -4042 1333 -4038
rect 1371 -4034 1375 -4030
rect 1371 -4042 1375 -4038
rect 1353 -4056 1357 -4052
rect 1253 -4063 1257 -4059
rect 1295 -4063 1299 -4059
rect 1418 -4034 1422 -4030
rect 1395 -4049 1399 -4045
rect 1220 -4078 1224 -4074
rect 1237 -4078 1241 -4074
rect 1278 -4078 1282 -4074
rect 1320 -4078 1324 -4074
rect 1362 -4078 1366 -4074
rect 1403 -4078 1407 -4074
rect 1211 -4101 1215 -4097
rect 1228 -4101 1232 -4097
rect 1184 -4315 1188 -4311
rect 1101 -4366 1105 -4362
rect 1184 -4366 1188 -4362
rect 862 -4554 866 -4550
rect 879 -4554 883 -4550
rect 899 -4554 903 -4550
rect 920 -4554 924 -4550
rect 941 -4554 945 -4550
rect 962 -4554 966 -4550
rect 983 -4554 987 -4550
rect 1004 -4554 1008 -4550
rect 1025 -4554 1029 -4550
rect 1045 -4554 1049 -4550
rect 853 -4617 857 -4613
rect 911 -4610 915 -4606
rect 953 -4617 957 -4613
rect 971 -4610 975 -4606
rect 1013 -4602 1017 -4598
rect 1013 -4610 1017 -4606
rect 995 -4624 999 -4620
rect 895 -4631 899 -4627
rect 937 -4631 941 -4627
rect 1059 -4602 1063 -4598
rect 1037 -4617 1041 -4613
rect 862 -4646 866 -4642
rect 879 -4646 883 -4642
rect 920 -4646 924 -4642
rect 962 -4646 966 -4642
rect 1004 -4646 1008 -4642
rect 1045 -4646 1049 -4642
rect 1184 -4610 1188 -4606
rect 1059 -4653 1063 -4649
rect 1184 -4653 1188 -4649
rect 862 -4725 866 -4721
rect 879 -4725 883 -4721
rect 899 -4725 903 -4721
rect 920 -4725 924 -4721
rect 941 -4725 945 -4721
rect 962 -4725 966 -4721
rect 983 -4725 987 -4721
rect 1004 -4725 1008 -4721
rect 1025 -4725 1029 -4721
rect 1045 -4725 1049 -4721
rect 839 -4781 843 -4777
rect 853 -4788 857 -4784
rect 911 -4781 915 -4777
rect 953 -4788 957 -4784
rect 971 -4781 975 -4777
rect 1013 -4773 1017 -4769
rect 1013 -4781 1017 -4777
rect 995 -4795 999 -4791
rect 895 -4802 899 -4798
rect 937 -4802 941 -4798
rect 1062 -4773 1066 -4769
rect 1037 -4788 1041 -4784
rect 862 -4817 866 -4813
rect 879 -4817 883 -4813
rect 920 -4817 924 -4813
rect 962 -4817 966 -4813
rect 1004 -4817 1008 -4813
rect 1045 -4817 1049 -4813
rect 853 -4840 857 -4836
rect 870 -4840 874 -4836
rect 824 -5039 828 -5035
rect 810 -5054 814 -5050
rect 743 -5098 747 -5094
rect 822 -5098 826 -5094
rect 504 -5289 508 -5285
rect 521 -5289 525 -5285
rect 541 -5289 545 -5285
rect 562 -5289 566 -5285
rect 583 -5289 587 -5285
rect 604 -5289 608 -5285
rect 625 -5289 629 -5285
rect 646 -5289 650 -5285
rect 667 -5289 671 -5285
rect 687 -5289 691 -5285
rect 495 -5352 499 -5348
rect 553 -5345 557 -5341
rect 595 -5352 599 -5348
rect 613 -5345 617 -5341
rect 655 -5337 659 -5333
rect 655 -5345 659 -5341
rect 637 -5359 641 -5355
rect 537 -5366 541 -5362
rect 579 -5366 583 -5362
rect 705 -5337 709 -5333
rect 679 -5352 683 -5348
rect 504 -5381 508 -5377
rect 521 -5381 525 -5377
rect 562 -5381 566 -5377
rect 604 -5381 608 -5377
rect 646 -5381 650 -5377
rect 687 -5381 691 -5377
rect 822 -5345 826 -5341
rect 705 -5390 709 -5386
rect 822 -5389 826 -5385
rect 504 -5449 508 -5445
rect 521 -5449 525 -5445
rect 541 -5449 545 -5445
rect 562 -5449 566 -5445
rect 583 -5449 587 -5445
rect 604 -5449 608 -5445
rect 625 -5449 629 -5445
rect 646 -5449 650 -5445
rect 667 -5449 671 -5445
rect 687 -5449 691 -5445
rect 481 -5505 485 -5501
rect 495 -5512 499 -5508
rect 553 -5505 557 -5501
rect 595 -5512 599 -5508
rect 613 -5505 617 -5501
rect 655 -5497 659 -5493
rect 655 -5505 659 -5501
rect 637 -5519 641 -5515
rect 537 -5526 541 -5522
rect 579 -5526 583 -5522
rect 705 -5497 709 -5493
rect 679 -5512 683 -5508
rect 504 -5541 508 -5537
rect 521 -5541 525 -5537
rect 562 -5541 566 -5537
rect 604 -5541 608 -5537
rect 646 -5541 650 -5537
rect 687 -5541 691 -5537
rect 495 -5563 499 -5559
rect 512 -5563 516 -5559
rect 705 -5595 709 -5591
rect 521 -5616 525 -5612
rect 810 -5616 814 -5612
rect 512 -5655 516 -5651
rect 504 -5722 508 -5718
rect 530 -5722 534 -5718
rect 547 -5722 551 -5718
rect 587 -5722 591 -5718
rect 608 -5722 612 -5718
rect 625 -5722 629 -5718
rect 665 -5722 669 -5718
rect 689 -5722 693 -5718
rect 726 -5722 730 -5718
rect 464 -5762 468 -5758
rect 495 -5755 499 -5751
rect 451 -5777 455 -5773
rect 513 -5748 517 -5744
rect 539 -5770 543 -5766
rect 521 -5777 525 -5773
rect 565 -5762 569 -5758
rect 617 -5755 621 -5751
rect 547 -5799 551 -5795
rect 583 -5799 587 -5795
rect 643 -5770 647 -5766
rect 625 -5799 629 -5795
rect 661 -5799 665 -5795
rect 735 -5762 739 -5758
rect 748 -5770 752 -5766
rect 504 -5814 508 -5810
rect 530 -5814 534 -5810
rect 573 -5814 577 -5810
rect 608 -5814 612 -5810
rect 652 -5814 656 -5810
rect 669 -5814 673 -5810
rect 705 -5814 709 -5810
rect 726 -5814 730 -5810
rect 1062 -4872 1066 -4868
rect 879 -4893 883 -4889
rect 1167 -4893 1171 -4889
rect 870 -4932 874 -4928
rect 862 -4999 866 -4995
rect 888 -4999 892 -4995
rect 905 -4999 909 -4995
rect 945 -4999 949 -4995
rect 966 -4999 970 -4995
rect 983 -4999 987 -4995
rect 1023 -4999 1027 -4995
rect 1047 -4999 1051 -4995
rect 1084 -4999 1088 -4995
rect 853 -5032 857 -5028
rect 871 -5025 875 -5021
rect 897 -5047 901 -5043
rect 879 -5054 883 -5050
rect 923 -5039 927 -5035
rect 975 -5032 979 -5028
rect 905 -5076 909 -5072
rect 941 -5076 945 -5072
rect 1001 -5047 1005 -5043
rect 983 -5076 987 -5072
rect 1019 -5076 1023 -5072
rect 1093 -5037 1097 -5033
rect 1167 -5039 1171 -5035
rect 1101 -5047 1105 -5043
rect 862 -5091 866 -5087
rect 888 -5091 892 -5087
rect 931 -5091 935 -5087
rect 966 -5091 970 -5087
rect 1010 -5091 1014 -5087
rect 1027 -5091 1031 -5087
rect 1063 -5091 1067 -5087
rect 1084 -5091 1088 -5087
rect 1418 -4133 1422 -4129
rect 1237 -4154 1241 -4150
rect 1228 -4193 1232 -4189
rect 1220 -4260 1224 -4256
rect 1246 -4260 1250 -4256
rect 1263 -4260 1267 -4256
rect 1303 -4260 1307 -4256
rect 1324 -4260 1328 -4256
rect 1341 -4260 1345 -4256
rect 1381 -4260 1385 -4256
rect 1405 -4260 1409 -4256
rect 1442 -4260 1446 -4256
rect 1211 -4293 1215 -4289
rect 1229 -4286 1233 -4282
rect 1255 -4308 1259 -4304
rect 1237 -4315 1241 -4311
rect 1281 -4300 1285 -4296
rect 1333 -4293 1337 -4289
rect 1263 -4337 1267 -4333
rect 1299 -4337 1303 -4333
rect 1359 -4308 1363 -4304
rect 1341 -4337 1345 -4333
rect 1377 -4337 1381 -4333
rect 1220 -4352 1224 -4348
rect 1246 -4352 1250 -4348
rect 1289 -4352 1293 -4348
rect 1324 -4352 1328 -4348
rect 1368 -4352 1372 -4348
rect 1385 -4352 1389 -4348
rect 1421 -4352 1425 -4348
rect 1442 -4352 1446 -4348
rect 1464 -4308 1468 -4304
rect 1464 -4359 1468 -4355
rect 1451 -4366 1455 -4362
rect 1220 -4554 1224 -4550
rect 1237 -4554 1241 -4550
rect 1257 -4554 1261 -4550
rect 1278 -4554 1282 -4550
rect 1299 -4554 1303 -4550
rect 1320 -4554 1324 -4550
rect 1341 -4554 1345 -4550
rect 1362 -4554 1366 -4550
rect 1383 -4554 1387 -4550
rect 1403 -4554 1407 -4550
rect 1211 -4617 1215 -4613
rect 1269 -4610 1273 -4606
rect 1311 -4617 1315 -4613
rect 1329 -4610 1333 -4606
rect 1371 -4602 1375 -4598
rect 1371 -4610 1375 -4606
rect 1353 -4624 1357 -4620
rect 1253 -4631 1257 -4627
rect 1295 -4631 1299 -4627
rect 1419 -4602 1423 -4598
rect 1395 -4617 1399 -4613
rect 1220 -4646 1224 -4642
rect 1237 -4646 1241 -4642
rect 1278 -4646 1282 -4642
rect 1320 -4646 1324 -4642
rect 1362 -4646 1366 -4642
rect 1403 -4646 1407 -4642
rect 1419 -4653 1423 -4649
rect 1220 -4725 1224 -4721
rect 1237 -4725 1241 -4721
rect 1257 -4725 1261 -4721
rect 1278 -4725 1282 -4721
rect 1299 -4725 1303 -4721
rect 1320 -4725 1324 -4721
rect 1341 -4725 1345 -4721
rect 1362 -4725 1366 -4721
rect 1383 -4725 1387 -4721
rect 1403 -4725 1407 -4721
rect 1197 -4781 1201 -4777
rect 1211 -4788 1215 -4784
rect 1269 -4781 1273 -4777
rect 1311 -4788 1315 -4784
rect 1329 -4781 1333 -4777
rect 1371 -4773 1375 -4769
rect 1371 -4781 1375 -4777
rect 1353 -4795 1357 -4791
rect 1253 -4802 1257 -4798
rect 1295 -4802 1299 -4798
rect 1420 -4773 1424 -4769
rect 1395 -4788 1399 -4784
rect 1220 -4817 1224 -4813
rect 1237 -4817 1241 -4813
rect 1278 -4817 1282 -4813
rect 1320 -4817 1324 -4813
rect 1362 -4817 1366 -4813
rect 1403 -4817 1407 -4813
rect 1211 -4840 1215 -4836
rect 1228 -4840 1232 -4836
rect 1184 -5054 1188 -5050
rect 1101 -5105 1105 -5101
rect 1177 -5105 1181 -5101
rect 862 -5289 866 -5285
rect 879 -5289 883 -5285
rect 899 -5289 903 -5285
rect 920 -5289 924 -5285
rect 941 -5289 945 -5285
rect 962 -5289 966 -5285
rect 983 -5289 987 -5285
rect 1004 -5289 1008 -5285
rect 1025 -5289 1029 -5285
rect 1045 -5289 1049 -5285
rect 853 -5352 857 -5348
rect 911 -5345 915 -5341
rect 953 -5352 957 -5348
rect 971 -5345 975 -5341
rect 1013 -5337 1017 -5333
rect 1013 -5345 1017 -5341
rect 995 -5359 999 -5355
rect 895 -5366 899 -5362
rect 937 -5366 941 -5362
rect 1061 -5337 1065 -5333
rect 1037 -5352 1041 -5348
rect 862 -5381 866 -5377
rect 879 -5381 883 -5377
rect 920 -5381 924 -5377
rect 962 -5381 966 -5377
rect 1004 -5381 1008 -5377
rect 1045 -5381 1049 -5377
rect 1177 -5345 1181 -5341
rect 1061 -5389 1065 -5385
rect 1177 -5388 1181 -5384
rect 862 -5449 866 -5445
rect 879 -5449 883 -5445
rect 899 -5449 903 -5445
rect 920 -5449 924 -5445
rect 941 -5449 945 -5445
rect 962 -5449 966 -5445
rect 983 -5449 987 -5445
rect 1004 -5449 1008 -5445
rect 1025 -5449 1029 -5445
rect 1045 -5449 1049 -5445
rect 839 -5505 843 -5501
rect 853 -5512 857 -5508
rect 911 -5505 915 -5501
rect 953 -5512 957 -5508
rect 971 -5505 975 -5501
rect 1013 -5497 1017 -5493
rect 1013 -5505 1017 -5501
rect 995 -5519 999 -5515
rect 895 -5526 899 -5522
rect 937 -5526 941 -5522
rect 1062 -5497 1066 -5493
rect 1037 -5512 1041 -5508
rect 862 -5541 866 -5537
rect 879 -5541 883 -5537
rect 920 -5541 924 -5537
rect 962 -5541 966 -5537
rect 1004 -5541 1008 -5537
rect 1045 -5541 1049 -5537
rect 853 -5563 857 -5559
rect 870 -5563 874 -5559
rect 1062 -5595 1066 -5591
rect 879 -5616 883 -5612
rect 1167 -5616 1171 -5612
rect 870 -5655 874 -5651
rect 862 -5722 866 -5718
rect 888 -5722 892 -5718
rect 905 -5722 909 -5718
rect 945 -5722 949 -5718
rect 966 -5722 970 -5718
rect 983 -5722 987 -5718
rect 1023 -5722 1027 -5718
rect 1047 -5722 1051 -5718
rect 1084 -5722 1088 -5718
rect 822 -5762 826 -5758
rect 853 -5755 857 -5751
rect 810 -5777 814 -5773
rect 871 -5748 875 -5744
rect 897 -5770 901 -5766
rect 879 -5777 883 -5773
rect 923 -5762 927 -5758
rect 975 -5755 979 -5751
rect 905 -5799 909 -5795
rect 941 -5799 945 -5795
rect 1001 -5770 1005 -5766
rect 983 -5799 987 -5795
rect 1019 -5799 1023 -5795
rect 1093 -5760 1097 -5756
rect 1167 -5762 1171 -5758
rect 1106 -5770 1110 -5766
rect 862 -5814 866 -5810
rect 888 -5814 892 -5810
rect 931 -5814 935 -5810
rect 966 -5814 970 -5810
rect 1010 -5814 1014 -5810
rect 1027 -5814 1031 -5810
rect 1063 -5814 1067 -5810
rect 1084 -5814 1088 -5810
rect 1420 -4872 1424 -4868
rect 1237 -4893 1241 -4889
rect 1228 -4932 1232 -4928
rect 1220 -4999 1224 -4995
rect 1246 -4999 1250 -4995
rect 1263 -4999 1267 -4995
rect 1303 -4999 1307 -4995
rect 1324 -4999 1328 -4995
rect 1341 -4999 1345 -4995
rect 1381 -4999 1385 -4995
rect 1405 -4999 1409 -4995
rect 1442 -4999 1446 -4995
rect 1211 -5032 1215 -5028
rect 1229 -5025 1233 -5021
rect 1255 -5047 1259 -5043
rect 1237 -5054 1241 -5050
rect 1281 -5039 1285 -5035
rect 1333 -5032 1337 -5028
rect 1263 -5076 1267 -5072
rect 1299 -5076 1303 -5072
rect 1359 -5047 1363 -5043
rect 1341 -5076 1345 -5072
rect 1377 -5076 1381 -5072
rect 1220 -5091 1224 -5087
rect 1246 -5091 1250 -5087
rect 1289 -5091 1293 -5087
rect 1324 -5091 1328 -5087
rect 1368 -5091 1372 -5087
rect 1385 -5091 1389 -5087
rect 1421 -5091 1425 -5087
rect 1442 -5091 1446 -5087
rect 1464 -5047 1468 -5043
rect 1464 -5098 1468 -5094
rect 1451 -5105 1455 -5101
rect 1220 -5289 1224 -5285
rect 1237 -5289 1241 -5285
rect 1257 -5289 1261 -5285
rect 1278 -5289 1282 -5285
rect 1299 -5289 1303 -5285
rect 1320 -5289 1324 -5285
rect 1341 -5289 1345 -5285
rect 1362 -5289 1366 -5285
rect 1383 -5289 1387 -5285
rect 1403 -5289 1407 -5285
rect 1211 -5352 1215 -5348
rect 1269 -5345 1273 -5341
rect 1311 -5352 1315 -5348
rect 1329 -5345 1333 -5341
rect 1371 -5337 1375 -5333
rect 1371 -5345 1375 -5341
rect 1353 -5359 1357 -5355
rect 1253 -5366 1257 -5362
rect 1295 -5366 1299 -5362
rect 1423 -5337 1427 -5333
rect 1395 -5352 1399 -5348
rect 1220 -5381 1224 -5377
rect 1237 -5381 1241 -5377
rect 1278 -5381 1282 -5377
rect 1320 -5381 1324 -5377
rect 1362 -5381 1366 -5377
rect 1403 -5381 1407 -5377
rect 1423 -5388 1427 -5384
rect 1220 -5449 1224 -5445
rect 1237 -5449 1241 -5445
rect 1257 -5449 1261 -5445
rect 1278 -5449 1282 -5445
rect 1299 -5449 1303 -5445
rect 1320 -5449 1324 -5445
rect 1341 -5449 1345 -5445
rect 1362 -5449 1366 -5445
rect 1383 -5449 1387 -5445
rect 1403 -5449 1407 -5445
rect 1197 -5505 1201 -5501
rect 1211 -5512 1215 -5508
rect 1269 -5505 1273 -5501
rect 1311 -5512 1315 -5508
rect 1329 -5505 1333 -5501
rect 1371 -5497 1375 -5493
rect 1371 -5505 1375 -5501
rect 1353 -5519 1357 -5515
rect 1253 -5526 1257 -5522
rect 1295 -5526 1299 -5522
rect 1423 -5497 1427 -5493
rect 1395 -5512 1399 -5508
rect 1220 -5541 1224 -5537
rect 1237 -5541 1241 -5537
rect 1278 -5541 1282 -5537
rect 1320 -5541 1324 -5537
rect 1362 -5541 1366 -5537
rect 1403 -5541 1407 -5537
rect 1211 -5563 1215 -5559
rect 1228 -5563 1232 -5559
rect 1423 -5595 1427 -5591
rect 1237 -5616 1241 -5612
rect 1228 -5655 1232 -5651
rect 1220 -5722 1224 -5718
rect 1246 -5722 1250 -5718
rect 1263 -5722 1267 -5718
rect 1303 -5722 1307 -5718
rect 1324 -5722 1328 -5718
rect 1341 -5722 1345 -5718
rect 1381 -5722 1385 -5718
rect 1405 -5722 1409 -5718
rect 1442 -5722 1446 -5718
rect 1177 -5777 1181 -5773
rect 1211 -5755 1215 -5751
rect 1229 -5748 1233 -5744
rect 1255 -5770 1259 -5766
rect 1237 -5777 1241 -5773
rect 1281 -5762 1285 -5758
rect 1333 -5755 1337 -5751
rect 1263 -5799 1267 -5795
rect 1299 -5799 1303 -5795
rect 1359 -5770 1363 -5766
rect 1341 -5799 1345 -5795
rect 1377 -5799 1381 -5795
rect 1220 -5814 1224 -5810
rect 1246 -5814 1250 -5810
rect 1289 -5814 1293 -5810
rect 1324 -5814 1328 -5810
rect 1368 -5814 1372 -5810
rect 1385 -5814 1389 -5810
rect 1421 -5814 1425 -5810
rect 1442 -5814 1446 -5810
rect -1225 -5845 -1221 -5841
rect -1208 -5845 -1204 -5841
rect -1188 -5845 -1184 -5841
rect -1167 -5845 -1163 -5841
rect -1146 -5845 -1142 -5841
rect -1125 -5845 -1121 -5841
rect -1104 -5845 -1100 -5841
rect -1083 -5845 -1079 -5841
rect -1062 -5845 -1058 -5841
rect -1042 -5845 -1038 -5841
rect -1246 -5901 -1242 -5897
rect -1234 -5908 -1230 -5904
rect -1176 -5901 -1172 -5897
rect -1134 -5908 -1130 -5904
rect -1116 -5901 -1112 -5897
rect -1074 -5893 -1070 -5889
rect -1074 -5901 -1070 -5897
rect -1092 -5915 -1088 -5911
rect -1192 -5922 -1188 -5918
rect -1150 -5922 -1146 -5918
rect -926 -5845 -922 -5841
rect -909 -5845 -905 -5841
rect -889 -5845 -885 -5841
rect -868 -5845 -864 -5841
rect -847 -5845 -843 -5841
rect -826 -5845 -822 -5841
rect -805 -5845 -801 -5841
rect -784 -5845 -780 -5841
rect -763 -5845 -759 -5841
rect -743 -5845 -739 -5841
rect -949 -5901 -945 -5897
rect -1050 -5908 -1046 -5904
rect -935 -5908 -931 -5904
rect -877 -5901 -873 -5897
rect -835 -5908 -831 -5904
rect -817 -5901 -813 -5897
rect -775 -5893 -771 -5889
rect -775 -5901 -771 -5897
rect -793 -5915 -789 -5911
rect -893 -5922 -889 -5918
rect -851 -5922 -847 -5918
rect -568 -5845 -564 -5841
rect -551 -5845 -547 -5841
rect -531 -5845 -527 -5841
rect -510 -5845 -506 -5841
rect -489 -5845 -485 -5841
rect -468 -5845 -464 -5841
rect -447 -5845 -443 -5841
rect -426 -5845 -422 -5841
rect -405 -5845 -401 -5841
rect -385 -5845 -381 -5841
rect -586 -5901 -582 -5897
rect -751 -5908 -747 -5904
rect -577 -5908 -573 -5904
rect -519 -5901 -515 -5897
rect -477 -5908 -473 -5904
rect -459 -5901 -455 -5897
rect -417 -5893 -413 -5889
rect -417 -5901 -413 -5897
rect -435 -5915 -431 -5911
rect -535 -5922 -531 -5918
rect -493 -5922 -489 -5918
rect 129 -5822 133 -5818
rect 392 -5822 396 -5818
rect 484 -5821 488 -5817
rect 748 -5821 752 -5817
rect 842 -5821 846 -5817
rect 1106 -5821 1110 -5817
rect 1199 -5821 1203 -5817
rect -210 -5845 -206 -5841
rect -193 -5845 -189 -5841
rect -173 -5845 -169 -5841
rect -152 -5845 -148 -5841
rect -131 -5845 -127 -5841
rect -110 -5845 -106 -5841
rect -89 -5845 -85 -5841
rect -68 -5845 -64 -5841
rect -47 -5845 -43 -5841
rect -27 -5845 -23 -5841
rect -233 -5901 -229 -5897
rect -393 -5908 -389 -5904
rect -219 -5908 -215 -5904
rect -161 -5901 -157 -5897
rect -119 -5908 -115 -5904
rect -101 -5901 -97 -5897
rect -59 -5893 -55 -5889
rect -59 -5901 -55 -5897
rect -77 -5915 -73 -5911
rect -177 -5922 -173 -5918
rect -135 -5922 -131 -5918
rect 148 -5845 152 -5841
rect 165 -5845 169 -5841
rect 185 -5845 189 -5841
rect 206 -5845 210 -5841
rect 227 -5845 231 -5841
rect 248 -5845 252 -5841
rect 269 -5845 273 -5841
rect 290 -5845 294 -5841
rect 311 -5845 315 -5841
rect 331 -5845 335 -5841
rect 129 -5901 133 -5897
rect -35 -5908 -31 -5904
rect 139 -5908 143 -5904
rect 197 -5901 201 -5897
rect 239 -5908 243 -5904
rect 257 -5901 261 -5897
rect 299 -5893 303 -5889
rect 299 -5901 303 -5897
rect 281 -5915 285 -5911
rect 181 -5922 185 -5918
rect 223 -5922 227 -5918
rect 504 -5845 508 -5841
rect 521 -5845 525 -5841
rect 541 -5845 545 -5841
rect 562 -5845 566 -5841
rect 583 -5845 587 -5841
rect 604 -5845 608 -5841
rect 625 -5845 629 -5841
rect 646 -5845 650 -5841
rect 667 -5845 671 -5841
rect 687 -5845 691 -5841
rect 484 -5901 488 -5897
rect 323 -5908 327 -5904
rect 495 -5908 499 -5904
rect 553 -5901 557 -5897
rect 595 -5908 599 -5904
rect 613 -5901 617 -5897
rect 655 -5893 659 -5889
rect 655 -5901 659 -5897
rect 637 -5915 641 -5911
rect 537 -5922 541 -5918
rect 579 -5922 583 -5918
rect 862 -5845 866 -5841
rect 879 -5845 883 -5841
rect 899 -5845 903 -5841
rect 920 -5845 924 -5841
rect 941 -5845 945 -5841
rect 962 -5845 966 -5841
rect 983 -5845 987 -5841
rect 1004 -5845 1008 -5841
rect 1025 -5845 1029 -5841
rect 1045 -5845 1049 -5841
rect 842 -5901 846 -5897
rect 679 -5908 683 -5904
rect 853 -5908 857 -5904
rect 911 -5901 915 -5897
rect 953 -5908 957 -5904
rect 971 -5901 975 -5897
rect 1013 -5893 1017 -5889
rect 1013 -5901 1017 -5897
rect 995 -5915 999 -5911
rect 895 -5922 899 -5918
rect 937 -5922 941 -5918
rect 1220 -5845 1224 -5841
rect 1237 -5845 1241 -5841
rect 1257 -5845 1261 -5841
rect 1278 -5845 1282 -5841
rect 1299 -5845 1303 -5841
rect 1320 -5845 1324 -5841
rect 1341 -5845 1345 -5841
rect 1362 -5845 1366 -5841
rect 1383 -5845 1387 -5841
rect 1403 -5845 1407 -5841
rect 1199 -5901 1203 -5897
rect 1037 -5908 1041 -5904
rect 1211 -5908 1215 -5904
rect 1269 -5901 1273 -5897
rect 1311 -5908 1315 -5904
rect 1329 -5901 1333 -5897
rect 1371 -5893 1375 -5889
rect 1371 -5901 1375 -5897
rect 1353 -5915 1357 -5911
rect 1253 -5922 1257 -5918
rect 1295 -5922 1299 -5918
rect 1466 -5770 1470 -5766
rect 1466 -5821 1470 -5817
rect 1564 -5845 1568 -5841
rect 1581 -5845 1585 -5841
rect 1601 -5845 1605 -5841
rect 1622 -5845 1626 -5841
rect 1643 -5845 1647 -5841
rect 1664 -5845 1668 -5841
rect 1685 -5845 1689 -5841
rect 1706 -5845 1710 -5841
rect 1727 -5845 1731 -5841
rect 1747 -5845 1751 -5841
rect 1451 -5901 1455 -5897
rect 1395 -5908 1399 -5904
rect 1555 -5908 1559 -5904
rect 1613 -5901 1617 -5897
rect 1655 -5908 1659 -5904
rect 1673 -5901 1677 -5897
rect 1715 -5893 1719 -5889
rect 1715 -5901 1719 -5897
rect 1697 -5915 1701 -5911
rect 1597 -5922 1601 -5918
rect 1639 -5922 1643 -5918
rect 1739 -5908 1743 -5904
rect -1225 -5937 -1221 -5933
rect -1208 -5937 -1204 -5933
rect -1167 -5937 -1163 -5933
rect -1125 -5937 -1121 -5933
rect -1083 -5937 -1079 -5933
rect -1042 -5937 -1038 -5933
rect -926 -5937 -922 -5933
rect -909 -5937 -905 -5933
rect -868 -5937 -864 -5933
rect -826 -5937 -822 -5933
rect -784 -5937 -780 -5933
rect -743 -5937 -739 -5933
rect -568 -5937 -564 -5933
rect -551 -5937 -547 -5933
rect -510 -5937 -506 -5933
rect -468 -5937 -464 -5933
rect -426 -5937 -422 -5933
rect -385 -5937 -381 -5933
rect -210 -5937 -206 -5933
rect -193 -5937 -189 -5933
rect -152 -5937 -148 -5933
rect -110 -5937 -106 -5933
rect -68 -5937 -64 -5933
rect -27 -5937 -23 -5933
rect 148 -5937 152 -5933
rect 165 -5937 169 -5933
rect 206 -5937 210 -5933
rect 248 -5937 252 -5933
rect 290 -5937 294 -5933
rect 331 -5937 335 -5933
rect 504 -5937 508 -5933
rect 521 -5937 525 -5933
rect 562 -5937 566 -5933
rect 604 -5937 608 -5933
rect 646 -5937 650 -5933
rect 687 -5937 691 -5933
rect 862 -5937 866 -5933
rect 879 -5937 883 -5933
rect 920 -5937 924 -5933
rect 962 -5937 966 -5933
rect 1004 -5937 1008 -5933
rect 1045 -5937 1049 -5933
rect 1220 -5937 1224 -5933
rect 1237 -5937 1241 -5933
rect 1278 -5937 1282 -5933
rect 1320 -5937 1324 -5933
rect 1362 -5937 1366 -5933
rect 1403 -5937 1407 -5933
rect 1564 -5937 1568 -5933
rect 1581 -5937 1585 -5933
rect 1622 -5937 1626 -5933
rect 1664 -5937 1668 -5933
rect 1706 -5937 1710 -5933
rect 1747 -5937 1751 -5933
<< pad >>
rect -1295 -824 -1291 -820
rect -924 -824 -920 -820
rect -565 -824 -561 -820
rect -207 -824 -203 -820
rect 150 -824 154 -820
rect 507 -824 511 -820
rect 865 -824 869 -820
rect 1223 -824 1227 -820
rect -1203 -1066 -1199 -1062
rect -1165 -1066 -1161 -1062
rect -1105 -1066 -1101 -1062
rect -1081 -1066 -1077 -1062
rect -908 -1066 -904 -1062
rect -870 -1066 -866 -1062
rect -810 -1066 -806 -1062
rect -786 -1066 -782 -1062
rect -550 -1066 -546 -1062
rect -512 -1066 -508 -1062
rect -452 -1066 -448 -1062
rect -428 -1066 -424 -1062
rect -192 -1066 -188 -1062
rect -154 -1066 -150 -1062
rect -94 -1066 -90 -1062
rect -70 -1066 -66 -1062
rect 166 -1066 170 -1062
rect 204 -1066 208 -1062
rect 264 -1066 268 -1062
rect 288 -1066 292 -1062
rect 522 -1066 526 -1062
rect 560 -1066 564 -1062
rect 620 -1066 624 -1062
rect 644 -1066 648 -1062
rect 880 -1066 884 -1062
rect 918 -1066 922 -1062
rect 978 -1066 982 -1062
rect 1002 -1066 1006 -1062
rect -1223 -1074 -1219 -1070
rect -1189 -1074 -1185 -1070
rect -1137 -1074 -1133 -1070
rect -1077 -1074 -1073 -1070
rect -1039 -1074 -1035 -1070
rect -928 -1074 -924 -1070
rect -894 -1074 -890 -1070
rect -842 -1074 -838 -1070
rect -782 -1074 -778 -1070
rect -744 -1074 -740 -1070
rect -570 -1074 -566 -1070
rect -536 -1074 -532 -1070
rect -484 -1074 -480 -1070
rect -424 -1074 -420 -1070
rect -386 -1074 -382 -1070
rect -212 -1074 -208 -1070
rect -178 -1074 -174 -1070
rect -126 -1074 -122 -1070
rect -66 -1074 -62 -1070
rect -28 -1074 -24 -1070
rect 146 -1074 150 -1070
rect 180 -1074 184 -1070
rect 232 -1074 236 -1070
rect 292 -1074 296 -1070
rect 330 -1074 334 -1070
rect 502 -1074 506 -1070
rect 536 -1074 540 -1070
rect 588 -1074 592 -1070
rect 648 -1074 652 -1070
rect 686 -1074 690 -1070
rect 860 -1074 864 -1070
rect 894 -1074 898 -1070
rect 946 -1074 950 -1070
rect 1006 -1074 1010 -1070
rect 1044 -1074 1048 -1070
rect -1179 -1081 -1175 -1077
rect -1147 -1081 -1143 -1077
rect -1095 -1081 -1091 -1077
rect -1063 -1081 -1059 -1077
rect -884 -1081 -880 -1077
rect -852 -1081 -848 -1077
rect -800 -1081 -796 -1077
rect -768 -1081 -764 -1077
rect -526 -1081 -522 -1077
rect -494 -1081 -490 -1077
rect -442 -1081 -438 -1077
rect -410 -1081 -406 -1077
rect -168 -1081 -164 -1077
rect -136 -1081 -132 -1077
rect -84 -1081 -80 -1077
rect -52 -1081 -48 -1077
rect 190 -1081 194 -1077
rect 222 -1081 226 -1077
rect 274 -1081 278 -1077
rect 306 -1081 310 -1077
rect 546 -1081 550 -1077
rect 578 -1081 582 -1077
rect 630 -1081 634 -1077
rect 662 -1081 666 -1077
rect 904 -1081 908 -1077
rect 936 -1081 940 -1077
rect 988 -1081 992 -1077
rect 1020 -1081 1024 -1077
rect -1219 -1088 -1215 -1084
rect -1105 -1088 -1101 -1084
rect -1053 -1088 -1049 -1084
rect -924 -1088 -920 -1084
rect -810 -1088 -806 -1084
rect -758 -1088 -754 -1084
rect -566 -1088 -562 -1084
rect -452 -1088 -448 -1084
rect -400 -1088 -396 -1084
rect -208 -1088 -204 -1084
rect -94 -1088 -90 -1084
rect -42 -1088 -38 -1084
rect 150 -1088 154 -1084
rect 264 -1088 268 -1084
rect 316 -1088 320 -1084
rect 506 -1088 510 -1084
rect 620 -1088 624 -1084
rect 672 -1088 676 -1084
rect 864 -1088 868 -1084
rect 978 -1088 982 -1084
rect 1030 -1088 1034 -1084
rect -1161 -1095 -1157 -1091
rect -1123 -1095 -1119 -1091
rect -866 -1095 -862 -1091
rect -828 -1095 -824 -1091
rect -508 -1095 -504 -1091
rect -470 -1095 -466 -1091
rect -150 -1095 -146 -1091
rect -112 -1095 -108 -1091
rect 208 -1095 212 -1091
rect 246 -1095 250 -1091
rect 564 -1095 568 -1091
rect 602 -1095 606 -1091
rect 922 -1095 926 -1091
rect 960 -1095 964 -1091
rect -1297 -1174 -1293 -1170
rect -923 -1174 -919 -1170
rect -565 -1174 -561 -1170
rect -207 -1174 -203 -1170
rect 151 -1174 155 -1170
rect 507 -1174 511 -1170
rect 865 -1174 869 -1170
rect 1223 -1174 1227 -1170
rect -924 -1317 -920 -1313
rect -858 -1317 -854 -1313
rect -824 -1317 -820 -1313
rect -780 -1317 -776 -1313
rect -746 -1317 -742 -1313
rect -566 -1317 -562 -1313
rect -500 -1317 -496 -1313
rect -466 -1317 -462 -1313
rect -422 -1317 -418 -1313
rect -388 -1317 -384 -1313
rect -208 -1317 -204 -1313
rect -142 -1317 -138 -1313
rect -108 -1317 -104 -1313
rect -64 -1317 -60 -1313
rect -30 -1317 -26 -1313
rect 150 -1317 154 -1313
rect 216 -1317 220 -1313
rect 250 -1317 254 -1313
rect 294 -1317 298 -1313
rect 328 -1317 332 -1313
rect 506 -1317 510 -1313
rect 572 -1317 576 -1313
rect 606 -1317 610 -1313
rect 650 -1317 654 -1313
rect 684 -1317 688 -1313
rect 864 -1317 868 -1313
rect 930 -1317 934 -1313
rect 964 -1317 968 -1313
rect 1008 -1317 1012 -1313
rect 1042 -1317 1046 -1313
rect -882 -1324 -878 -1320
rect -524 -1324 -520 -1320
rect -166 -1324 -162 -1320
rect 192 -1324 196 -1320
rect 548 -1324 552 -1320
rect 906 -1324 910 -1320
rect -848 -1331 -844 -1327
rect -706 -1331 -702 -1327
rect -490 -1331 -486 -1327
rect -348 -1331 -344 -1327
rect -132 -1331 -128 -1327
rect 10 -1331 14 -1327
rect 226 -1331 230 -1327
rect 368 -1331 372 -1327
rect 582 -1331 586 -1327
rect 724 -1331 728 -1327
rect 940 -1331 944 -1327
rect 1082 -1331 1086 -1327
rect -928 -1338 -924 -1334
rect -898 -1338 -894 -1334
rect -780 -1338 -776 -1334
rect -570 -1338 -566 -1334
rect -540 -1338 -536 -1334
rect -422 -1338 -418 -1334
rect -212 -1338 -208 -1334
rect -182 -1338 -178 -1334
rect -64 -1338 -60 -1334
rect 146 -1338 150 -1334
rect 176 -1338 180 -1334
rect 294 -1338 298 -1334
rect 502 -1338 506 -1334
rect 532 -1338 536 -1334
rect 650 -1338 654 -1334
rect 860 -1338 864 -1334
rect 890 -1338 894 -1334
rect 1008 -1338 1012 -1334
rect -1169 -1347 -1165 -1343
rect -902 -1346 -898 -1342
rect -804 -1346 -800 -1342
rect -544 -1346 -540 -1342
rect -446 -1346 -442 -1342
rect -186 -1346 -182 -1342
rect -88 -1346 -84 -1342
rect 172 -1346 176 -1342
rect 270 -1346 274 -1342
rect 528 -1346 532 -1342
rect 626 -1346 630 -1342
rect 886 -1346 890 -1342
rect 984 -1346 988 -1342
rect 1272 -1347 1276 -1343
rect -1219 -1354 -1215 -1350
rect -1179 -1354 -1175 -1350
rect -1159 -1354 -1155 -1350
rect -924 -1353 -920 -1349
rect -776 -1353 -772 -1349
rect -566 -1353 -562 -1349
rect -418 -1353 -414 -1349
rect -208 -1353 -204 -1349
rect -60 -1353 -56 -1349
rect 150 -1353 154 -1349
rect 298 -1353 302 -1349
rect 506 -1353 510 -1349
rect 654 -1353 658 -1349
rect 864 -1353 868 -1349
rect 1012 -1353 1016 -1349
rect 1222 -1354 1226 -1350
rect 1262 -1354 1266 -1350
rect 1282 -1354 1286 -1350
rect -1223 -1361 -1219 -1357
rect -1193 -1361 -1189 -1357
rect -1145 -1361 -1141 -1357
rect -902 -1360 -898 -1356
rect -794 -1360 -790 -1356
rect -760 -1360 -756 -1356
rect -544 -1360 -540 -1356
rect -436 -1360 -432 -1356
rect -402 -1360 -398 -1356
rect -186 -1360 -182 -1356
rect -78 -1360 -74 -1356
rect -44 -1360 -40 -1356
rect 172 -1360 176 -1356
rect 280 -1360 284 -1356
rect 314 -1360 318 -1356
rect 528 -1360 532 -1356
rect 636 -1360 640 -1356
rect 670 -1360 674 -1356
rect 886 -1360 890 -1356
rect 994 -1360 998 -1356
rect 1028 -1360 1032 -1356
rect 1218 -1361 1222 -1357
rect 1248 -1361 1252 -1357
rect 1296 -1361 1300 -1357
rect -928 -1367 -924 -1363
rect -872 -1367 -868 -1363
rect -838 -1367 -834 -1363
rect -570 -1367 -566 -1363
rect -514 -1367 -510 -1363
rect -480 -1367 -476 -1363
rect -212 -1367 -208 -1363
rect -156 -1367 -152 -1363
rect -122 -1367 -118 -1363
rect 146 -1367 150 -1363
rect 202 -1367 206 -1363
rect 236 -1367 240 -1363
rect 502 -1367 506 -1363
rect 558 -1367 562 -1363
rect 592 -1367 596 -1363
rect 860 -1367 864 -1363
rect 916 -1367 920 -1363
rect 950 -1367 954 -1363
rect -1203 -1469 -1199 -1465
rect -1165 -1469 -1161 -1465
rect -1105 -1469 -1101 -1465
rect -1081 -1469 -1077 -1465
rect -908 -1469 -904 -1465
rect -870 -1469 -866 -1465
rect -810 -1469 -806 -1465
rect -786 -1469 -782 -1465
rect -550 -1469 -546 -1465
rect -512 -1469 -508 -1465
rect -452 -1469 -448 -1465
rect -428 -1469 -424 -1465
rect -192 -1469 -188 -1465
rect -154 -1469 -150 -1465
rect -94 -1469 -90 -1465
rect -70 -1469 -66 -1465
rect 166 -1469 170 -1465
rect 204 -1469 208 -1465
rect 264 -1469 268 -1465
rect 288 -1469 292 -1465
rect 522 -1469 526 -1465
rect 560 -1469 564 -1465
rect 620 -1469 624 -1465
rect 644 -1469 648 -1465
rect 880 -1469 884 -1465
rect 918 -1469 922 -1465
rect 978 -1469 982 -1465
rect 1002 -1469 1006 -1465
rect -1223 -1477 -1219 -1473
rect -1189 -1477 -1185 -1473
rect -1137 -1477 -1133 -1473
rect -1077 -1477 -1073 -1473
rect -1039 -1477 -1035 -1473
rect -928 -1477 -924 -1473
rect -894 -1477 -890 -1473
rect -842 -1477 -838 -1473
rect -782 -1477 -778 -1473
rect -744 -1477 -740 -1473
rect -570 -1477 -566 -1473
rect -536 -1477 -532 -1473
rect -484 -1477 -480 -1473
rect -424 -1477 -420 -1473
rect -386 -1477 -382 -1473
rect -212 -1477 -208 -1473
rect -178 -1477 -174 -1473
rect -126 -1477 -122 -1473
rect -66 -1477 -62 -1473
rect -28 -1477 -24 -1473
rect 146 -1477 150 -1473
rect 180 -1477 184 -1473
rect 232 -1477 236 -1473
rect 292 -1477 296 -1473
rect 330 -1477 334 -1473
rect 502 -1477 506 -1473
rect 536 -1477 540 -1473
rect 588 -1477 592 -1473
rect 648 -1477 652 -1473
rect 686 -1477 690 -1473
rect 860 -1477 864 -1473
rect 894 -1477 898 -1473
rect 946 -1477 950 -1473
rect 1006 -1477 1010 -1473
rect 1044 -1477 1048 -1473
rect -1179 -1484 -1175 -1480
rect -1147 -1484 -1143 -1480
rect -1095 -1484 -1091 -1480
rect -1063 -1484 -1059 -1480
rect -884 -1484 -880 -1480
rect -852 -1484 -848 -1480
rect -800 -1484 -796 -1480
rect -768 -1484 -764 -1480
rect -526 -1484 -522 -1480
rect -494 -1484 -490 -1480
rect -442 -1484 -438 -1480
rect -410 -1484 -406 -1480
rect -168 -1484 -164 -1480
rect -136 -1484 -132 -1480
rect -84 -1484 -80 -1480
rect -52 -1484 -48 -1480
rect 190 -1484 194 -1480
rect 222 -1484 226 -1480
rect 274 -1484 278 -1480
rect 306 -1484 310 -1480
rect 546 -1484 550 -1480
rect 578 -1484 582 -1480
rect 630 -1484 634 -1480
rect 662 -1484 666 -1480
rect 904 -1484 908 -1480
rect 936 -1484 940 -1480
rect 988 -1484 992 -1480
rect 1020 -1484 1024 -1480
rect -1219 -1491 -1215 -1487
rect -1105 -1491 -1101 -1487
rect -1053 -1491 -1049 -1487
rect -924 -1491 -920 -1487
rect -810 -1491 -806 -1487
rect -758 -1491 -754 -1487
rect -566 -1491 -562 -1487
rect -452 -1491 -448 -1487
rect -400 -1491 -396 -1487
rect -208 -1491 -204 -1487
rect -94 -1491 -90 -1487
rect -42 -1491 -38 -1487
rect 150 -1491 154 -1487
rect 264 -1491 268 -1487
rect 316 -1491 320 -1487
rect 506 -1491 510 -1487
rect 620 -1491 624 -1487
rect 672 -1491 676 -1487
rect 864 -1491 868 -1487
rect 978 -1491 982 -1487
rect 1030 -1491 1034 -1487
rect -1161 -1498 -1157 -1494
rect -1123 -1498 -1119 -1494
rect -866 -1498 -862 -1494
rect -828 -1498 -824 -1494
rect -508 -1498 -504 -1494
rect -470 -1498 -466 -1494
rect -150 -1498 -146 -1494
rect -112 -1498 -108 -1494
rect 208 -1498 212 -1494
rect 246 -1498 250 -1494
rect 564 -1498 568 -1494
rect 602 -1498 606 -1494
rect 922 -1498 926 -1494
rect 960 -1498 964 -1494
rect -1203 -1640 -1199 -1636
rect -1165 -1640 -1161 -1636
rect -1105 -1640 -1101 -1636
rect -1081 -1640 -1077 -1636
rect -908 -1640 -904 -1636
rect -870 -1640 -866 -1636
rect -810 -1640 -806 -1636
rect -786 -1640 -782 -1636
rect -550 -1640 -546 -1636
rect -512 -1640 -508 -1636
rect -452 -1640 -448 -1636
rect -428 -1640 -424 -1636
rect -192 -1640 -188 -1636
rect -154 -1640 -150 -1636
rect -94 -1640 -90 -1636
rect -70 -1640 -66 -1636
rect 166 -1640 170 -1636
rect 204 -1640 208 -1636
rect 264 -1640 268 -1636
rect 288 -1640 292 -1636
rect 522 -1640 526 -1636
rect 560 -1640 564 -1636
rect 620 -1640 624 -1636
rect 644 -1640 648 -1636
rect 880 -1640 884 -1636
rect 918 -1640 922 -1636
rect 978 -1640 982 -1636
rect 1002 -1640 1006 -1636
rect 1238 -1640 1242 -1636
rect 1276 -1640 1280 -1636
rect 1336 -1640 1340 -1636
rect 1360 -1640 1364 -1636
rect -1223 -1648 -1219 -1644
rect -1189 -1648 -1185 -1644
rect -1137 -1648 -1133 -1644
rect -1077 -1648 -1073 -1644
rect -1039 -1648 -1035 -1644
rect -928 -1648 -924 -1644
rect -894 -1648 -890 -1644
rect -842 -1648 -838 -1644
rect -782 -1648 -778 -1644
rect -744 -1648 -740 -1644
rect -570 -1648 -566 -1644
rect -536 -1648 -532 -1644
rect -484 -1648 -480 -1644
rect -424 -1648 -420 -1644
rect -386 -1648 -382 -1644
rect -212 -1648 -208 -1644
rect -178 -1648 -174 -1644
rect -126 -1648 -122 -1644
rect -66 -1648 -62 -1644
rect -28 -1648 -24 -1644
rect 146 -1648 150 -1644
rect 180 -1648 184 -1644
rect 232 -1648 236 -1644
rect 292 -1648 296 -1644
rect 330 -1648 334 -1644
rect 502 -1648 506 -1644
rect 536 -1648 540 -1644
rect 588 -1648 592 -1644
rect 648 -1648 652 -1644
rect 686 -1648 690 -1644
rect 860 -1648 864 -1644
rect 894 -1648 898 -1644
rect 946 -1648 950 -1644
rect 1006 -1648 1010 -1644
rect 1044 -1648 1048 -1644
rect 1218 -1648 1222 -1644
rect 1252 -1648 1256 -1644
rect 1304 -1648 1308 -1644
rect 1364 -1648 1368 -1644
rect 1402 -1648 1406 -1644
rect -1179 -1655 -1175 -1651
rect -1147 -1655 -1143 -1651
rect -1095 -1655 -1091 -1651
rect -1063 -1655 -1059 -1651
rect -884 -1655 -880 -1651
rect -852 -1655 -848 -1651
rect -800 -1655 -796 -1651
rect -768 -1655 -764 -1651
rect -526 -1655 -522 -1651
rect -494 -1655 -490 -1651
rect -442 -1655 -438 -1651
rect -410 -1655 -406 -1651
rect -168 -1655 -164 -1651
rect -136 -1655 -132 -1651
rect -84 -1655 -80 -1651
rect -52 -1655 -48 -1651
rect 190 -1655 194 -1651
rect 222 -1655 226 -1651
rect 274 -1655 278 -1651
rect 306 -1655 310 -1651
rect 546 -1655 550 -1651
rect 578 -1655 582 -1651
rect 630 -1655 634 -1651
rect 662 -1655 666 -1651
rect 904 -1655 908 -1651
rect 936 -1655 940 -1651
rect 988 -1655 992 -1651
rect 1020 -1655 1024 -1651
rect 1262 -1655 1266 -1651
rect 1294 -1655 1298 -1651
rect 1346 -1655 1350 -1651
rect 1378 -1655 1382 -1651
rect -1219 -1662 -1215 -1658
rect -1105 -1662 -1101 -1658
rect -1053 -1662 -1049 -1658
rect -924 -1662 -920 -1658
rect -810 -1662 -806 -1658
rect -758 -1662 -754 -1658
rect -566 -1662 -562 -1658
rect -452 -1662 -448 -1658
rect -400 -1662 -396 -1658
rect -208 -1662 -204 -1658
rect -94 -1662 -90 -1658
rect -42 -1662 -38 -1658
rect 150 -1662 154 -1658
rect 264 -1662 268 -1658
rect 316 -1662 320 -1658
rect 506 -1662 510 -1658
rect 620 -1662 624 -1658
rect 672 -1662 676 -1658
rect 864 -1662 868 -1658
rect 978 -1662 982 -1658
rect 1030 -1662 1034 -1658
rect 1222 -1662 1226 -1658
rect 1336 -1662 1340 -1658
rect 1388 -1662 1392 -1658
rect -1161 -1669 -1157 -1665
rect -1123 -1669 -1119 -1665
rect -866 -1669 -862 -1665
rect -828 -1669 -824 -1665
rect -508 -1669 -504 -1665
rect -470 -1669 -466 -1665
rect -150 -1669 -146 -1665
rect -112 -1669 -108 -1665
rect 208 -1669 212 -1665
rect 246 -1669 250 -1665
rect 564 -1669 568 -1665
rect 602 -1669 606 -1665
rect 922 -1669 926 -1665
rect 960 -1669 964 -1665
rect 1280 -1669 1284 -1665
rect 1318 -1669 1322 -1665
rect -1532 -1811 -1528 -1807
rect -1494 -1811 -1490 -1807
rect -1434 -1811 -1430 -1807
rect -1410 -1811 -1406 -1807
rect -1203 -1811 -1199 -1807
rect -1165 -1811 -1161 -1807
rect -1105 -1811 -1101 -1807
rect -1081 -1811 -1077 -1807
rect -908 -1811 -904 -1807
rect -870 -1811 -866 -1807
rect -810 -1811 -806 -1807
rect -786 -1811 -782 -1807
rect -550 -1811 -546 -1807
rect -512 -1811 -508 -1807
rect -452 -1811 -448 -1807
rect -428 -1811 -424 -1807
rect -192 -1811 -188 -1807
rect -154 -1811 -150 -1807
rect -94 -1811 -90 -1807
rect -70 -1811 -66 -1807
rect 166 -1811 170 -1807
rect 204 -1811 208 -1807
rect 264 -1811 268 -1807
rect 288 -1811 292 -1807
rect 522 -1811 526 -1807
rect 560 -1811 564 -1807
rect 620 -1811 624 -1807
rect 644 -1811 648 -1807
rect 880 -1811 884 -1807
rect 918 -1811 922 -1807
rect 978 -1811 982 -1807
rect 1002 -1811 1006 -1807
rect 1238 -1811 1242 -1807
rect 1276 -1811 1280 -1807
rect 1336 -1811 1340 -1807
rect 1360 -1811 1364 -1807
rect -1552 -1819 -1548 -1815
rect -1518 -1819 -1514 -1815
rect -1466 -1819 -1462 -1815
rect -1406 -1819 -1402 -1815
rect -1368 -1819 -1364 -1815
rect -1223 -1819 -1219 -1815
rect -1189 -1819 -1185 -1815
rect -1137 -1819 -1133 -1815
rect -1077 -1819 -1073 -1815
rect -1039 -1819 -1035 -1815
rect -928 -1819 -924 -1815
rect -894 -1819 -890 -1815
rect -842 -1819 -838 -1815
rect -782 -1819 -778 -1815
rect -744 -1819 -740 -1815
rect -570 -1819 -566 -1815
rect -536 -1819 -532 -1815
rect -484 -1819 -480 -1815
rect -424 -1819 -420 -1815
rect -386 -1819 -382 -1815
rect -212 -1819 -208 -1815
rect -178 -1819 -174 -1815
rect -126 -1819 -122 -1815
rect -66 -1819 -62 -1815
rect -28 -1819 -24 -1815
rect 146 -1819 150 -1815
rect 180 -1819 184 -1815
rect 232 -1819 236 -1815
rect 292 -1819 296 -1815
rect 330 -1819 334 -1815
rect 502 -1819 506 -1815
rect 536 -1819 540 -1815
rect 588 -1819 592 -1815
rect 648 -1819 652 -1815
rect 686 -1819 690 -1815
rect 860 -1819 864 -1815
rect 894 -1819 898 -1815
rect 946 -1819 950 -1815
rect 1006 -1819 1010 -1815
rect 1044 -1819 1048 -1815
rect 1218 -1819 1222 -1815
rect 1252 -1819 1256 -1815
rect 1304 -1819 1308 -1815
rect 1364 -1819 1368 -1815
rect 1402 -1819 1406 -1815
rect -1508 -1826 -1504 -1822
rect -1476 -1826 -1472 -1822
rect -1424 -1826 -1420 -1822
rect -1392 -1826 -1388 -1822
rect -1179 -1826 -1175 -1822
rect -1147 -1826 -1143 -1822
rect -1095 -1826 -1091 -1822
rect -1063 -1826 -1059 -1822
rect -884 -1826 -880 -1822
rect -852 -1826 -848 -1822
rect -800 -1826 -796 -1822
rect -768 -1826 -764 -1822
rect -526 -1826 -522 -1822
rect -494 -1826 -490 -1822
rect -442 -1826 -438 -1822
rect -410 -1826 -406 -1822
rect -168 -1826 -164 -1822
rect -136 -1826 -132 -1822
rect -84 -1826 -80 -1822
rect -52 -1826 -48 -1822
rect 190 -1826 194 -1822
rect 222 -1826 226 -1822
rect 274 -1826 278 -1822
rect 306 -1826 310 -1822
rect 546 -1826 550 -1822
rect 578 -1826 582 -1822
rect 630 -1826 634 -1822
rect 662 -1826 666 -1822
rect 904 -1826 908 -1822
rect 936 -1826 940 -1822
rect 988 -1826 992 -1822
rect 1020 -1826 1024 -1822
rect 1262 -1826 1266 -1822
rect 1294 -1826 1298 -1822
rect 1346 -1826 1350 -1822
rect 1378 -1826 1382 -1822
rect -1548 -1833 -1544 -1829
rect -1434 -1833 -1430 -1829
rect -1382 -1833 -1378 -1829
rect -1219 -1833 -1215 -1829
rect -1105 -1833 -1101 -1829
rect -1053 -1833 -1049 -1829
rect -924 -1833 -920 -1829
rect -810 -1833 -806 -1829
rect -758 -1833 -754 -1829
rect -566 -1833 -562 -1829
rect -452 -1833 -448 -1829
rect -400 -1833 -396 -1829
rect -208 -1833 -204 -1829
rect -94 -1833 -90 -1829
rect -42 -1833 -38 -1829
rect 150 -1833 154 -1829
rect 264 -1833 268 -1829
rect 316 -1833 320 -1829
rect 506 -1833 510 -1829
rect 620 -1833 624 -1829
rect 672 -1833 676 -1829
rect 864 -1833 868 -1829
rect 978 -1833 982 -1829
rect 1030 -1833 1034 -1829
rect 1222 -1833 1226 -1829
rect 1336 -1833 1340 -1829
rect 1388 -1833 1392 -1829
rect -1490 -1840 -1486 -1836
rect -1452 -1840 -1448 -1836
rect -1161 -1840 -1157 -1836
rect -1123 -1840 -1119 -1836
rect -866 -1840 -862 -1836
rect -828 -1840 -824 -1836
rect -508 -1840 -504 -1836
rect -470 -1840 -466 -1836
rect -150 -1840 -146 -1836
rect -112 -1840 -108 -1836
rect 208 -1840 212 -1836
rect 246 -1840 250 -1836
rect 564 -1840 568 -1836
rect 602 -1840 606 -1836
rect 922 -1840 926 -1836
rect 960 -1840 964 -1836
rect 1280 -1840 1284 -1836
rect 1318 -1840 1322 -1836
rect -1308 -1902 -1304 -1898
rect -934 -1902 -930 -1898
rect -576 -1902 -572 -1898
rect -218 -1902 -214 -1898
rect 140 -1902 144 -1898
rect 496 -1902 500 -1898
rect 854 -1902 858 -1898
rect 1212 -1902 1216 -1898
rect -1297 -1910 -1293 -1906
rect -923 -1910 -919 -1906
rect -565 -1910 -561 -1906
rect -207 -1910 -203 -1906
rect 151 -1910 155 -1906
rect 507 -1910 511 -1906
rect 865 -1910 869 -1906
rect 1223 -1910 1227 -1906
rect -924 -2048 -920 -2044
rect -858 -2048 -854 -2044
rect -824 -2048 -820 -2044
rect -780 -2048 -776 -2044
rect -746 -2048 -742 -2044
rect -566 -2048 -562 -2044
rect -500 -2048 -496 -2044
rect -466 -2048 -462 -2044
rect -422 -2048 -418 -2044
rect -388 -2048 -384 -2044
rect -208 -2048 -204 -2044
rect -142 -2048 -138 -2044
rect -108 -2048 -104 -2044
rect -64 -2048 -60 -2044
rect -30 -2048 -26 -2044
rect 150 -2048 154 -2044
rect 216 -2048 220 -2044
rect 250 -2048 254 -2044
rect 294 -2048 298 -2044
rect 328 -2048 332 -2044
rect 506 -2048 510 -2044
rect 572 -2048 576 -2044
rect 606 -2048 610 -2044
rect 650 -2048 654 -2044
rect 684 -2048 688 -2044
rect 864 -2048 868 -2044
rect 930 -2048 934 -2044
rect 964 -2048 968 -2044
rect 1008 -2048 1012 -2044
rect 1042 -2048 1046 -2044
rect 1222 -2048 1226 -2044
rect 1288 -2048 1292 -2044
rect 1322 -2048 1326 -2044
rect 1366 -2048 1370 -2044
rect 1400 -2048 1404 -2044
rect -882 -2055 -878 -2051
rect -524 -2055 -520 -2051
rect -166 -2055 -162 -2051
rect 192 -2055 196 -2051
rect 548 -2055 552 -2051
rect 906 -2055 910 -2051
rect 1264 -2055 1268 -2051
rect -848 -2062 -844 -2058
rect -706 -2062 -702 -2058
rect -490 -2062 -486 -2058
rect -348 -2062 -344 -2058
rect -132 -2062 -128 -2058
rect 10 -2062 14 -2058
rect 226 -2062 230 -2058
rect 368 -2062 372 -2058
rect 582 -2062 586 -2058
rect 724 -2062 728 -2058
rect 940 -2062 944 -2058
rect 1082 -2062 1086 -2058
rect 1298 -2062 1302 -2058
rect 1440 -2062 1444 -2058
rect -928 -2069 -924 -2065
rect -898 -2069 -894 -2065
rect -780 -2069 -776 -2065
rect -570 -2069 -566 -2065
rect -540 -2069 -536 -2065
rect -422 -2069 -418 -2065
rect -212 -2069 -208 -2065
rect -182 -2069 -178 -2065
rect -64 -2069 -60 -2065
rect 146 -2069 150 -2065
rect 176 -2069 180 -2065
rect 294 -2069 298 -2065
rect 502 -2069 506 -2065
rect 532 -2069 536 -2065
rect 650 -2069 654 -2065
rect 860 -2069 864 -2065
rect 890 -2069 894 -2065
rect 1008 -2069 1012 -2065
rect 1218 -2069 1222 -2065
rect 1248 -2069 1252 -2065
rect 1366 -2069 1370 -2065
rect -1173 -2078 -1169 -2074
rect -902 -2077 -898 -2073
rect -804 -2077 -800 -2073
rect -544 -2077 -540 -2073
rect -446 -2077 -442 -2073
rect -186 -2077 -182 -2073
rect -88 -2077 -84 -2073
rect 172 -2077 176 -2073
rect 270 -2077 274 -2073
rect 528 -2077 532 -2073
rect 626 -2077 630 -2073
rect 886 -2077 890 -2073
rect 984 -2077 988 -2073
rect 1244 -2077 1248 -2073
rect 1342 -2077 1346 -2073
rect -1223 -2085 -1219 -2081
rect -1183 -2085 -1179 -2081
rect -1163 -2085 -1159 -2081
rect -924 -2084 -920 -2080
rect -776 -2084 -772 -2080
rect -566 -2084 -562 -2080
rect -418 -2084 -414 -2080
rect -208 -2084 -204 -2080
rect -60 -2084 -56 -2080
rect 150 -2084 154 -2080
rect 298 -2084 302 -2080
rect 506 -2084 510 -2080
rect 654 -2084 658 -2080
rect 864 -2084 868 -2080
rect 1012 -2084 1016 -2080
rect 1222 -2084 1226 -2080
rect 1370 -2084 1374 -2080
rect -1227 -2092 -1223 -2088
rect -1197 -2092 -1193 -2088
rect -1149 -2092 -1145 -2088
rect -902 -2091 -898 -2087
rect -794 -2091 -790 -2087
rect -760 -2091 -756 -2087
rect -544 -2091 -540 -2087
rect -436 -2091 -432 -2087
rect -402 -2091 -398 -2087
rect -186 -2091 -182 -2087
rect -78 -2091 -74 -2087
rect -44 -2091 -40 -2087
rect 172 -2091 176 -2087
rect 280 -2091 284 -2087
rect 314 -2091 318 -2087
rect 528 -2091 532 -2087
rect 636 -2091 640 -2087
rect 670 -2091 674 -2087
rect 886 -2091 890 -2087
rect 994 -2091 998 -2087
rect 1028 -2091 1032 -2087
rect 1244 -2091 1248 -2087
rect 1352 -2091 1356 -2087
rect 1386 -2091 1390 -2087
rect -928 -2098 -924 -2094
rect -872 -2098 -868 -2094
rect -838 -2098 -834 -2094
rect -570 -2098 -566 -2094
rect -514 -2098 -510 -2094
rect -480 -2098 -476 -2094
rect -212 -2098 -208 -2094
rect -156 -2098 -152 -2094
rect -122 -2098 -118 -2094
rect 146 -2098 150 -2094
rect 202 -2098 206 -2094
rect 236 -2098 240 -2094
rect 502 -2098 506 -2094
rect 558 -2098 562 -2094
rect 592 -2098 596 -2094
rect 860 -2098 864 -2094
rect 916 -2098 920 -2094
rect 950 -2098 954 -2094
rect 1218 -2098 1222 -2094
rect 1274 -2098 1278 -2094
rect 1308 -2098 1312 -2094
rect -1207 -2221 -1203 -2217
rect -1169 -2221 -1165 -2217
rect -1109 -2221 -1105 -2217
rect -1085 -2221 -1081 -2217
rect -908 -2221 -904 -2217
rect -870 -2221 -866 -2217
rect -810 -2221 -806 -2217
rect -786 -2221 -782 -2217
rect -550 -2221 -546 -2217
rect -512 -2221 -508 -2217
rect -452 -2221 -448 -2217
rect -428 -2221 -424 -2217
rect -192 -2221 -188 -2217
rect -154 -2221 -150 -2217
rect -94 -2221 -90 -2217
rect -70 -2221 -66 -2217
rect 166 -2221 170 -2217
rect 204 -2221 208 -2217
rect 264 -2221 268 -2217
rect 288 -2221 292 -2217
rect 522 -2221 526 -2217
rect 560 -2221 564 -2217
rect 620 -2221 624 -2217
rect 644 -2221 648 -2217
rect -1227 -2229 -1223 -2225
rect -1193 -2229 -1189 -2225
rect -1141 -2229 -1137 -2225
rect -1081 -2229 -1077 -2225
rect -1043 -2229 -1039 -2225
rect -928 -2229 -924 -2225
rect -894 -2229 -890 -2225
rect -842 -2229 -838 -2225
rect -782 -2229 -778 -2225
rect -744 -2229 -740 -2225
rect -570 -2229 -566 -2225
rect -536 -2229 -532 -2225
rect -484 -2229 -480 -2225
rect -424 -2229 -420 -2225
rect -386 -2229 -382 -2225
rect -212 -2229 -208 -2225
rect -178 -2229 -174 -2225
rect -126 -2229 -122 -2225
rect -66 -2229 -62 -2225
rect -28 -2229 -24 -2225
rect 146 -2229 150 -2225
rect 180 -2229 184 -2225
rect 232 -2229 236 -2225
rect 292 -2229 296 -2225
rect 330 -2229 334 -2225
rect 502 -2229 506 -2225
rect 536 -2229 540 -2225
rect 588 -2229 592 -2225
rect 648 -2229 652 -2225
rect 686 -2229 690 -2225
rect -1183 -2236 -1179 -2232
rect -1151 -2236 -1147 -2232
rect -1099 -2236 -1095 -2232
rect -1067 -2236 -1063 -2232
rect -884 -2236 -880 -2232
rect -852 -2236 -848 -2232
rect -800 -2236 -796 -2232
rect -768 -2236 -764 -2232
rect -526 -2236 -522 -2232
rect -494 -2236 -490 -2232
rect -442 -2236 -438 -2232
rect -410 -2236 -406 -2232
rect -168 -2236 -164 -2232
rect -136 -2236 -132 -2232
rect -84 -2236 -80 -2232
rect -52 -2236 -48 -2232
rect 190 -2236 194 -2232
rect 222 -2236 226 -2232
rect 274 -2236 278 -2232
rect 306 -2236 310 -2232
rect 546 -2236 550 -2232
rect 578 -2236 582 -2232
rect 630 -2236 634 -2232
rect 662 -2236 666 -2232
rect -1223 -2243 -1219 -2239
rect -1109 -2243 -1105 -2239
rect -1057 -2243 -1053 -2239
rect -924 -2243 -920 -2239
rect -810 -2243 -806 -2239
rect -758 -2243 -754 -2239
rect -566 -2243 -562 -2239
rect -452 -2243 -448 -2239
rect -400 -2243 -396 -2239
rect -208 -2243 -204 -2239
rect -94 -2243 -90 -2239
rect -42 -2243 -38 -2239
rect 150 -2243 154 -2239
rect 264 -2243 268 -2239
rect 316 -2243 320 -2239
rect 506 -2243 510 -2239
rect 620 -2243 624 -2239
rect 672 -2243 676 -2239
rect -1165 -2250 -1161 -2246
rect -1127 -2250 -1123 -2246
rect -866 -2250 -862 -2246
rect -828 -2250 -824 -2246
rect -508 -2250 -504 -2246
rect -470 -2250 -466 -2246
rect -150 -2250 -146 -2246
rect -112 -2250 -108 -2246
rect 208 -2250 212 -2246
rect 246 -2250 250 -2246
rect 564 -2250 568 -2246
rect 602 -2250 606 -2246
rect -1532 -2392 -1528 -2388
rect -1494 -2392 -1490 -2388
rect -1434 -2392 -1430 -2388
rect -1410 -2392 -1406 -2388
rect -1207 -2392 -1203 -2388
rect -1169 -2392 -1165 -2388
rect -1109 -2392 -1105 -2388
rect -1085 -2392 -1081 -2388
rect -908 -2392 -904 -2388
rect -870 -2392 -866 -2388
rect -810 -2392 -806 -2388
rect -786 -2392 -782 -2388
rect -550 -2392 -546 -2388
rect -512 -2392 -508 -2388
rect -452 -2392 -448 -2388
rect -428 -2392 -424 -2388
rect -192 -2392 -188 -2388
rect -154 -2392 -150 -2388
rect -94 -2392 -90 -2388
rect -70 -2392 -66 -2388
rect 166 -2392 170 -2388
rect 204 -2392 208 -2388
rect 264 -2392 268 -2388
rect 288 -2392 292 -2388
rect 522 -2392 526 -2388
rect 560 -2392 564 -2388
rect 620 -2392 624 -2388
rect 644 -2392 648 -2388
rect 880 -2392 884 -2388
rect 918 -2392 922 -2388
rect 978 -2392 982 -2388
rect 1002 -2392 1006 -2388
rect 1238 -2392 1242 -2388
rect 1276 -2392 1280 -2388
rect 1336 -2392 1340 -2388
rect 1360 -2392 1364 -2388
rect -1552 -2400 -1548 -2396
rect -1518 -2400 -1514 -2396
rect -1466 -2400 -1462 -2396
rect -1406 -2400 -1402 -2396
rect -1368 -2400 -1364 -2396
rect -1227 -2400 -1223 -2396
rect -1193 -2400 -1189 -2396
rect -1141 -2400 -1137 -2396
rect -1081 -2400 -1077 -2396
rect -1043 -2400 -1039 -2396
rect -928 -2400 -924 -2396
rect -894 -2400 -890 -2396
rect -842 -2400 -838 -2396
rect -782 -2400 -778 -2396
rect -744 -2400 -740 -2396
rect -570 -2400 -566 -2396
rect -536 -2400 -532 -2396
rect -484 -2400 -480 -2396
rect -424 -2400 -420 -2396
rect -386 -2400 -382 -2396
rect -212 -2400 -208 -2396
rect -178 -2400 -174 -2396
rect -126 -2400 -122 -2396
rect -66 -2400 -62 -2396
rect -28 -2400 -24 -2396
rect 146 -2400 150 -2396
rect 180 -2400 184 -2396
rect 232 -2400 236 -2396
rect 292 -2400 296 -2396
rect 330 -2400 334 -2396
rect 502 -2400 506 -2396
rect 536 -2400 540 -2396
rect 588 -2400 592 -2396
rect 648 -2400 652 -2396
rect 686 -2400 690 -2396
rect 860 -2400 864 -2396
rect 894 -2400 898 -2396
rect 946 -2400 950 -2396
rect 1006 -2400 1010 -2396
rect 1044 -2400 1048 -2396
rect 1218 -2400 1222 -2396
rect 1252 -2400 1256 -2396
rect 1304 -2400 1308 -2396
rect 1364 -2400 1368 -2396
rect 1402 -2400 1406 -2396
rect -1508 -2407 -1504 -2403
rect -1476 -2407 -1472 -2403
rect -1424 -2407 -1420 -2403
rect -1392 -2407 -1388 -2403
rect -1183 -2407 -1179 -2403
rect -1151 -2407 -1147 -2403
rect -1099 -2407 -1095 -2403
rect -1067 -2407 -1063 -2403
rect -884 -2407 -880 -2403
rect -852 -2407 -848 -2403
rect -800 -2407 -796 -2403
rect -768 -2407 -764 -2403
rect -526 -2407 -522 -2403
rect -494 -2407 -490 -2403
rect -442 -2407 -438 -2403
rect -410 -2407 -406 -2403
rect -168 -2407 -164 -2403
rect -136 -2407 -132 -2403
rect -84 -2407 -80 -2403
rect -52 -2407 -48 -2403
rect 190 -2407 194 -2403
rect 222 -2407 226 -2403
rect 274 -2407 278 -2403
rect 306 -2407 310 -2403
rect 546 -2407 550 -2403
rect 578 -2407 582 -2403
rect 630 -2407 634 -2403
rect 662 -2407 666 -2403
rect 904 -2407 908 -2403
rect 936 -2407 940 -2403
rect 988 -2407 992 -2403
rect 1020 -2407 1024 -2403
rect 1262 -2407 1266 -2403
rect 1294 -2407 1298 -2403
rect 1346 -2407 1350 -2403
rect 1378 -2407 1382 -2403
rect -1548 -2414 -1544 -2410
rect -1434 -2414 -1430 -2410
rect -1382 -2414 -1378 -2410
rect -1223 -2414 -1219 -2410
rect -1109 -2414 -1105 -2410
rect -1057 -2414 -1053 -2410
rect -924 -2414 -920 -2410
rect -810 -2414 -806 -2410
rect -758 -2414 -754 -2410
rect -566 -2414 -562 -2410
rect -452 -2414 -448 -2410
rect -400 -2414 -396 -2410
rect -208 -2414 -204 -2410
rect -94 -2414 -90 -2410
rect -42 -2414 -38 -2410
rect 150 -2414 154 -2410
rect 264 -2414 268 -2410
rect 316 -2414 320 -2410
rect 506 -2414 510 -2410
rect 620 -2414 624 -2410
rect 672 -2414 676 -2410
rect 864 -2414 868 -2410
rect 978 -2414 982 -2410
rect 1030 -2414 1034 -2410
rect 1222 -2414 1226 -2410
rect 1336 -2414 1340 -2410
rect 1388 -2414 1392 -2410
rect -1490 -2421 -1486 -2417
rect -1452 -2421 -1448 -2417
rect -1165 -2421 -1161 -2417
rect -1127 -2421 -1123 -2417
rect -866 -2421 -862 -2417
rect -828 -2421 -824 -2417
rect -508 -2421 -504 -2417
rect -470 -2421 -466 -2417
rect -150 -2421 -146 -2417
rect -112 -2421 -108 -2417
rect 208 -2421 212 -2417
rect 246 -2421 250 -2417
rect 564 -2421 568 -2417
rect 602 -2421 606 -2417
rect 922 -2421 926 -2417
rect 960 -2421 964 -2417
rect 1280 -2421 1284 -2417
rect 1318 -2421 1322 -2417
rect -1532 -2563 -1528 -2559
rect -1494 -2563 -1490 -2559
rect -1434 -2563 -1430 -2559
rect -1410 -2563 -1406 -2559
rect -1207 -2563 -1203 -2559
rect -1169 -2563 -1165 -2559
rect -1109 -2563 -1105 -2559
rect -1085 -2563 -1081 -2559
rect -908 -2563 -904 -2559
rect -870 -2563 -866 -2559
rect -810 -2563 -806 -2559
rect -786 -2563 -782 -2559
rect -550 -2563 -546 -2559
rect -512 -2563 -508 -2559
rect -452 -2563 -448 -2559
rect -428 -2563 -424 -2559
rect -193 -2563 -189 -2559
rect -155 -2563 -151 -2559
rect -95 -2563 -91 -2559
rect -71 -2563 -67 -2559
rect 166 -2563 170 -2559
rect 204 -2563 208 -2559
rect 264 -2563 268 -2559
rect 288 -2563 292 -2559
rect 522 -2563 526 -2559
rect 560 -2563 564 -2559
rect 620 -2563 624 -2559
rect 644 -2563 648 -2559
rect 880 -2563 884 -2559
rect 918 -2563 922 -2559
rect 978 -2563 982 -2559
rect 1002 -2563 1006 -2559
rect 1238 -2563 1242 -2559
rect 1276 -2563 1280 -2559
rect 1336 -2563 1340 -2559
rect 1360 -2563 1364 -2559
rect -1552 -2571 -1548 -2567
rect -1518 -2571 -1514 -2567
rect -1466 -2571 -1462 -2567
rect -1406 -2571 -1402 -2567
rect -1368 -2571 -1364 -2567
rect -1227 -2571 -1223 -2567
rect -1193 -2571 -1189 -2567
rect -1141 -2571 -1137 -2567
rect -1081 -2571 -1077 -2567
rect -1043 -2571 -1039 -2567
rect -928 -2571 -924 -2567
rect -894 -2571 -890 -2567
rect -842 -2571 -838 -2567
rect -782 -2571 -778 -2567
rect -744 -2571 -740 -2567
rect -570 -2571 -566 -2567
rect -536 -2571 -532 -2567
rect -484 -2571 -480 -2567
rect -424 -2571 -420 -2567
rect -386 -2571 -382 -2567
rect -213 -2571 -209 -2567
rect -179 -2571 -175 -2567
rect -127 -2571 -123 -2567
rect -67 -2571 -63 -2567
rect -29 -2571 -25 -2567
rect 146 -2571 150 -2567
rect 180 -2571 184 -2567
rect 232 -2571 236 -2567
rect 292 -2571 296 -2567
rect 330 -2571 334 -2567
rect 502 -2571 506 -2567
rect 536 -2571 540 -2567
rect 588 -2571 592 -2567
rect 648 -2571 652 -2567
rect 686 -2571 690 -2567
rect 860 -2571 864 -2567
rect 894 -2571 898 -2567
rect 946 -2571 950 -2567
rect 1006 -2571 1010 -2567
rect 1044 -2571 1048 -2567
rect 1218 -2571 1222 -2567
rect 1252 -2571 1256 -2567
rect 1304 -2571 1308 -2567
rect 1364 -2571 1368 -2567
rect 1402 -2571 1406 -2567
rect -1508 -2578 -1504 -2574
rect -1476 -2578 -1472 -2574
rect -1424 -2578 -1420 -2574
rect -1392 -2578 -1388 -2574
rect -1183 -2578 -1179 -2574
rect -1151 -2578 -1147 -2574
rect -1099 -2578 -1095 -2574
rect -1067 -2578 -1063 -2574
rect -884 -2578 -880 -2574
rect -852 -2578 -848 -2574
rect -800 -2578 -796 -2574
rect -768 -2578 -764 -2574
rect -526 -2578 -522 -2574
rect -494 -2578 -490 -2574
rect -442 -2578 -438 -2574
rect -410 -2578 -406 -2574
rect -169 -2578 -165 -2574
rect -137 -2578 -133 -2574
rect -85 -2578 -81 -2574
rect -53 -2578 -49 -2574
rect 190 -2578 194 -2574
rect 222 -2578 226 -2574
rect 274 -2578 278 -2574
rect 306 -2578 310 -2574
rect 546 -2578 550 -2574
rect 578 -2578 582 -2574
rect 630 -2578 634 -2574
rect 662 -2578 666 -2574
rect 904 -2578 908 -2574
rect 936 -2578 940 -2574
rect 988 -2578 992 -2574
rect 1020 -2578 1024 -2574
rect 1262 -2578 1266 -2574
rect 1294 -2578 1298 -2574
rect 1346 -2578 1350 -2574
rect 1378 -2578 1382 -2574
rect -1548 -2585 -1544 -2581
rect -1434 -2585 -1430 -2581
rect -1382 -2585 -1378 -2581
rect -1223 -2585 -1219 -2581
rect -1109 -2585 -1105 -2581
rect -1057 -2585 -1053 -2581
rect -924 -2585 -920 -2581
rect -810 -2585 -806 -2581
rect -758 -2585 -754 -2581
rect -566 -2585 -562 -2581
rect -452 -2585 -448 -2581
rect -400 -2585 -396 -2581
rect -209 -2585 -205 -2581
rect -95 -2585 -91 -2581
rect -43 -2585 -39 -2581
rect 150 -2585 154 -2581
rect 264 -2585 268 -2581
rect 316 -2585 320 -2581
rect 506 -2585 510 -2581
rect 620 -2585 624 -2581
rect 672 -2585 676 -2581
rect 864 -2585 868 -2581
rect 978 -2585 982 -2581
rect 1030 -2585 1034 -2581
rect 1222 -2585 1226 -2581
rect 1336 -2585 1340 -2581
rect 1388 -2585 1392 -2581
rect -1490 -2592 -1486 -2588
rect -1452 -2592 -1448 -2588
rect -1165 -2592 -1161 -2588
rect -1127 -2592 -1123 -2588
rect -866 -2592 -862 -2588
rect -828 -2592 -824 -2588
rect -508 -2592 -504 -2588
rect -470 -2592 -466 -2588
rect -151 -2592 -147 -2588
rect -113 -2592 -109 -2588
rect 208 -2592 212 -2588
rect 246 -2592 250 -2588
rect 564 -2592 568 -2588
rect 602 -2592 606 -2588
rect 922 -2592 926 -2588
rect 960 -2592 964 -2588
rect 1280 -2592 1284 -2588
rect 1318 -2592 1322 -2588
rect -1308 -2652 -1304 -2648
rect -934 -2652 -930 -2648
rect -576 -2652 -572 -2648
rect -218 -2652 -214 -2648
rect 140 -2652 144 -2648
rect 496 -2652 500 -2648
rect 854 -2652 858 -2648
rect 1212 -2652 1216 -2648
rect -1297 -2660 -1293 -2656
rect -923 -2660 -919 -2656
rect -565 -2660 -561 -2656
rect -207 -2660 -203 -2656
rect 151 -2660 155 -2656
rect 507 -2660 511 -2656
rect 865 -2660 869 -2656
rect 1223 -2660 1227 -2656
rect -924 -2798 -920 -2794
rect -858 -2798 -854 -2794
rect -824 -2798 -820 -2794
rect -780 -2798 -776 -2794
rect -746 -2798 -742 -2794
rect -566 -2798 -562 -2794
rect -500 -2798 -496 -2794
rect -466 -2798 -462 -2794
rect -422 -2798 -418 -2794
rect -388 -2798 -384 -2794
rect -208 -2798 -204 -2794
rect -142 -2798 -138 -2794
rect -108 -2798 -104 -2794
rect -64 -2798 -60 -2794
rect -30 -2798 -26 -2794
rect 150 -2798 154 -2794
rect 216 -2798 220 -2794
rect 250 -2798 254 -2794
rect 294 -2798 298 -2794
rect 328 -2798 332 -2794
rect 506 -2798 510 -2794
rect 572 -2798 576 -2794
rect 606 -2798 610 -2794
rect 650 -2798 654 -2794
rect 684 -2798 688 -2794
rect 864 -2798 868 -2794
rect 930 -2798 934 -2794
rect 964 -2798 968 -2794
rect 1008 -2798 1012 -2794
rect 1042 -2798 1046 -2794
rect 1222 -2798 1226 -2794
rect 1288 -2798 1292 -2794
rect 1322 -2798 1326 -2794
rect 1366 -2798 1370 -2794
rect 1400 -2798 1404 -2794
rect -882 -2805 -878 -2801
rect -524 -2805 -520 -2801
rect -166 -2805 -162 -2801
rect 192 -2805 196 -2801
rect 548 -2805 552 -2801
rect 906 -2805 910 -2801
rect 1264 -2805 1268 -2801
rect -848 -2812 -844 -2808
rect -706 -2812 -702 -2808
rect -490 -2812 -486 -2808
rect -348 -2812 -344 -2808
rect -132 -2812 -128 -2808
rect 10 -2812 14 -2808
rect 226 -2812 230 -2808
rect 368 -2812 372 -2808
rect 582 -2812 586 -2808
rect 724 -2812 728 -2808
rect 940 -2812 944 -2808
rect 1082 -2812 1086 -2808
rect 1298 -2812 1302 -2808
rect 1440 -2812 1444 -2808
rect -928 -2819 -924 -2815
rect -898 -2819 -894 -2815
rect -780 -2819 -776 -2815
rect -570 -2819 -566 -2815
rect -540 -2819 -536 -2815
rect -422 -2819 -418 -2815
rect -212 -2819 -208 -2815
rect -182 -2819 -178 -2815
rect -64 -2819 -60 -2815
rect 146 -2819 150 -2815
rect 176 -2819 180 -2815
rect 294 -2819 298 -2815
rect 502 -2819 506 -2815
rect 532 -2819 536 -2815
rect 650 -2819 654 -2815
rect 860 -2819 864 -2815
rect 890 -2819 894 -2815
rect 1008 -2819 1012 -2815
rect 1218 -2819 1222 -2815
rect 1248 -2819 1252 -2815
rect 1366 -2819 1370 -2815
rect -1173 -2828 -1169 -2824
rect -902 -2827 -898 -2823
rect -804 -2827 -800 -2823
rect -544 -2827 -540 -2823
rect -446 -2827 -442 -2823
rect -186 -2827 -182 -2823
rect -88 -2827 -84 -2823
rect 172 -2827 176 -2823
rect 270 -2827 274 -2823
rect 528 -2827 532 -2823
rect 626 -2827 630 -2823
rect 886 -2827 890 -2823
rect 984 -2827 988 -2823
rect 1244 -2827 1248 -2823
rect 1342 -2827 1346 -2823
rect -1223 -2835 -1219 -2831
rect -1183 -2835 -1179 -2831
rect -1163 -2835 -1159 -2831
rect -924 -2834 -920 -2830
rect -776 -2834 -772 -2830
rect -566 -2834 -562 -2830
rect -418 -2834 -414 -2830
rect -208 -2834 -204 -2830
rect -60 -2834 -56 -2830
rect 150 -2834 154 -2830
rect 298 -2834 302 -2830
rect 506 -2834 510 -2830
rect 654 -2834 658 -2830
rect 864 -2834 868 -2830
rect 1012 -2834 1016 -2830
rect 1222 -2834 1226 -2830
rect 1370 -2834 1374 -2830
rect -1227 -2842 -1223 -2838
rect -1197 -2842 -1193 -2838
rect -1149 -2842 -1145 -2838
rect -902 -2841 -898 -2837
rect -794 -2841 -790 -2837
rect -760 -2841 -756 -2837
rect -544 -2841 -540 -2837
rect -436 -2841 -432 -2837
rect -402 -2841 -398 -2837
rect -186 -2841 -182 -2837
rect -78 -2841 -74 -2837
rect -44 -2841 -40 -2837
rect 172 -2841 176 -2837
rect 280 -2841 284 -2837
rect 314 -2841 318 -2837
rect 528 -2841 532 -2837
rect 636 -2841 640 -2837
rect 670 -2841 674 -2837
rect 886 -2841 890 -2837
rect 994 -2841 998 -2837
rect 1028 -2841 1032 -2837
rect 1244 -2841 1248 -2837
rect 1352 -2841 1356 -2837
rect 1386 -2841 1390 -2837
rect -928 -2848 -924 -2844
rect -872 -2848 -868 -2844
rect -838 -2848 -834 -2844
rect -570 -2848 -566 -2844
rect -514 -2848 -510 -2844
rect -480 -2848 -476 -2844
rect -212 -2848 -208 -2844
rect -156 -2848 -152 -2844
rect -122 -2848 -118 -2844
rect 146 -2848 150 -2844
rect 202 -2848 206 -2844
rect 236 -2848 240 -2844
rect 502 -2848 506 -2844
rect 558 -2848 562 -2844
rect 592 -2848 596 -2844
rect 860 -2848 864 -2844
rect 916 -2848 920 -2844
rect 950 -2848 954 -2844
rect 1218 -2848 1222 -2844
rect 1274 -2848 1278 -2844
rect 1308 -2848 1312 -2844
rect -1532 -2946 -1528 -2942
rect -1494 -2946 -1490 -2942
rect -1434 -2946 -1430 -2942
rect -1410 -2946 -1406 -2942
rect -1207 -2946 -1203 -2942
rect -1169 -2946 -1165 -2942
rect -1109 -2946 -1105 -2942
rect -1085 -2946 -1081 -2942
rect -908 -2946 -904 -2942
rect -870 -2946 -866 -2942
rect -810 -2946 -806 -2942
rect -786 -2946 -782 -2942
rect -550 -2946 -546 -2942
rect -512 -2946 -508 -2942
rect -452 -2946 -448 -2942
rect -428 -2946 -424 -2942
rect -192 -2946 -188 -2942
rect -154 -2946 -150 -2942
rect -94 -2946 -90 -2942
rect -70 -2946 -66 -2942
rect 166 -2946 170 -2942
rect 204 -2946 208 -2942
rect 264 -2946 268 -2942
rect 288 -2946 292 -2942
rect -1552 -2954 -1548 -2950
rect -1518 -2954 -1514 -2950
rect -1466 -2954 -1462 -2950
rect -1406 -2954 -1402 -2950
rect -1368 -2954 -1364 -2950
rect -1227 -2954 -1223 -2950
rect -1193 -2954 -1189 -2950
rect -1141 -2954 -1137 -2950
rect -1081 -2954 -1077 -2950
rect -1043 -2954 -1039 -2950
rect -928 -2954 -924 -2950
rect -894 -2954 -890 -2950
rect -842 -2954 -838 -2950
rect -782 -2954 -778 -2950
rect -744 -2954 -740 -2950
rect -570 -2954 -566 -2950
rect -536 -2954 -532 -2950
rect -484 -2954 -480 -2950
rect -424 -2954 -420 -2950
rect -386 -2954 -382 -2950
rect -212 -2954 -208 -2950
rect -178 -2954 -174 -2950
rect -126 -2954 -122 -2950
rect -66 -2954 -62 -2950
rect -28 -2954 -24 -2950
rect 146 -2954 150 -2950
rect 180 -2954 184 -2950
rect 232 -2954 236 -2950
rect 292 -2954 296 -2950
rect 330 -2954 334 -2950
rect -1508 -2961 -1504 -2957
rect -1476 -2961 -1472 -2957
rect -1424 -2961 -1420 -2957
rect -1392 -2961 -1388 -2957
rect -1183 -2961 -1179 -2957
rect -1151 -2961 -1147 -2957
rect -1099 -2961 -1095 -2957
rect -1067 -2961 -1063 -2957
rect -884 -2961 -880 -2957
rect -852 -2961 -848 -2957
rect -800 -2961 -796 -2957
rect -768 -2961 -764 -2957
rect -526 -2961 -522 -2957
rect -494 -2961 -490 -2957
rect -442 -2961 -438 -2957
rect -410 -2961 -406 -2957
rect -168 -2961 -164 -2957
rect -136 -2961 -132 -2957
rect -84 -2961 -80 -2957
rect -52 -2961 -48 -2957
rect 190 -2961 194 -2957
rect 222 -2961 226 -2957
rect 274 -2961 278 -2957
rect 306 -2961 310 -2957
rect -1548 -2968 -1544 -2964
rect -1434 -2968 -1430 -2964
rect -1382 -2968 -1378 -2964
rect -1223 -2968 -1219 -2964
rect -1109 -2968 -1105 -2964
rect -1057 -2968 -1053 -2964
rect -924 -2968 -920 -2964
rect -810 -2968 -806 -2964
rect -758 -2968 -754 -2964
rect -566 -2968 -562 -2964
rect -452 -2968 -448 -2964
rect -400 -2968 -396 -2964
rect -208 -2968 -204 -2964
rect -94 -2968 -90 -2964
rect -42 -2968 -38 -2964
rect 150 -2968 154 -2964
rect 264 -2968 268 -2964
rect 316 -2968 320 -2964
rect -1490 -2975 -1486 -2971
rect -1452 -2975 -1448 -2971
rect -1165 -2975 -1161 -2971
rect -1127 -2975 -1123 -2971
rect -866 -2975 -862 -2971
rect -828 -2975 -824 -2971
rect -508 -2975 -504 -2971
rect -470 -2975 -466 -2971
rect -150 -2975 -146 -2971
rect -112 -2975 -108 -2971
rect 208 -2975 212 -2971
rect 246 -2975 250 -2971
rect -1532 -3117 -1528 -3113
rect -1494 -3117 -1490 -3113
rect -1434 -3117 -1430 -3113
rect -1410 -3117 -1406 -3113
rect -1207 -3117 -1203 -3113
rect -1169 -3117 -1165 -3113
rect -1109 -3117 -1105 -3113
rect -1085 -3117 -1081 -3113
rect -908 -3117 -904 -3113
rect -870 -3117 -866 -3113
rect -810 -3117 -806 -3113
rect -786 -3117 -782 -3113
rect -550 -3117 -546 -3113
rect -512 -3117 -508 -3113
rect -452 -3117 -448 -3113
rect -428 -3117 -424 -3113
rect -192 -3117 -188 -3113
rect -154 -3117 -150 -3113
rect -94 -3117 -90 -3113
rect -70 -3117 -66 -3113
rect 166 -3117 170 -3113
rect 204 -3117 208 -3113
rect 264 -3117 268 -3113
rect 288 -3117 292 -3113
rect 522 -3117 526 -3113
rect 560 -3117 564 -3113
rect 620 -3117 624 -3113
rect 644 -3117 648 -3113
rect 880 -3117 884 -3113
rect 918 -3117 922 -3113
rect 978 -3117 982 -3113
rect 1002 -3117 1006 -3113
rect 1238 -3117 1242 -3113
rect 1276 -3117 1280 -3113
rect 1336 -3117 1340 -3113
rect 1360 -3117 1364 -3113
rect -1552 -3125 -1548 -3121
rect -1518 -3125 -1514 -3121
rect -1466 -3125 -1462 -3121
rect -1406 -3125 -1402 -3121
rect -1368 -3125 -1364 -3121
rect -1227 -3125 -1223 -3121
rect -1193 -3125 -1189 -3121
rect -1141 -3125 -1137 -3121
rect -1081 -3125 -1077 -3121
rect -1043 -3125 -1039 -3121
rect -928 -3125 -924 -3121
rect -894 -3125 -890 -3121
rect -842 -3125 -838 -3121
rect -782 -3125 -778 -3121
rect -744 -3125 -740 -3121
rect -570 -3125 -566 -3121
rect -536 -3125 -532 -3121
rect -484 -3125 -480 -3121
rect -424 -3125 -420 -3121
rect -386 -3125 -382 -3121
rect -212 -3125 -208 -3121
rect -178 -3125 -174 -3121
rect -126 -3125 -122 -3121
rect -66 -3125 -62 -3121
rect -28 -3125 -24 -3121
rect 146 -3125 150 -3121
rect 180 -3125 184 -3121
rect 232 -3125 236 -3121
rect 292 -3125 296 -3121
rect 330 -3125 334 -3121
rect 502 -3125 506 -3121
rect 536 -3125 540 -3121
rect 588 -3125 592 -3121
rect 648 -3125 652 -3121
rect 686 -3125 690 -3121
rect 860 -3125 864 -3121
rect 894 -3125 898 -3121
rect 946 -3125 950 -3121
rect 1006 -3125 1010 -3121
rect 1044 -3125 1048 -3121
rect 1218 -3125 1222 -3121
rect 1252 -3125 1256 -3121
rect 1304 -3125 1308 -3121
rect 1364 -3125 1368 -3121
rect 1402 -3125 1406 -3121
rect -1508 -3132 -1504 -3128
rect -1476 -3132 -1472 -3128
rect -1424 -3132 -1420 -3128
rect -1392 -3132 -1388 -3128
rect -1183 -3132 -1179 -3128
rect -1151 -3132 -1147 -3128
rect -1099 -3132 -1095 -3128
rect -1067 -3132 -1063 -3128
rect -884 -3132 -880 -3128
rect -852 -3132 -848 -3128
rect -800 -3132 -796 -3128
rect -768 -3132 -764 -3128
rect -526 -3132 -522 -3128
rect -494 -3132 -490 -3128
rect -442 -3132 -438 -3128
rect -410 -3132 -406 -3128
rect -168 -3132 -164 -3128
rect -136 -3132 -132 -3128
rect -84 -3132 -80 -3128
rect -52 -3132 -48 -3128
rect 190 -3132 194 -3128
rect 222 -3132 226 -3128
rect 274 -3132 278 -3128
rect 306 -3132 310 -3128
rect 546 -3132 550 -3128
rect 578 -3132 582 -3128
rect 630 -3132 634 -3128
rect 662 -3132 666 -3128
rect 904 -3132 908 -3128
rect 936 -3132 940 -3128
rect 988 -3132 992 -3128
rect 1020 -3132 1024 -3128
rect 1262 -3132 1266 -3128
rect 1294 -3132 1298 -3128
rect 1346 -3132 1350 -3128
rect 1378 -3132 1382 -3128
rect -1548 -3139 -1544 -3135
rect -1434 -3139 -1430 -3135
rect -1382 -3139 -1378 -3135
rect -1223 -3139 -1219 -3135
rect -1109 -3139 -1105 -3135
rect -1057 -3139 -1053 -3135
rect -924 -3139 -920 -3135
rect -810 -3139 -806 -3135
rect -758 -3139 -754 -3135
rect -566 -3139 -562 -3135
rect -452 -3139 -448 -3135
rect -400 -3139 -396 -3135
rect -208 -3139 -204 -3135
rect -94 -3139 -90 -3135
rect -42 -3139 -38 -3135
rect 150 -3139 154 -3135
rect 264 -3139 268 -3135
rect 316 -3139 320 -3135
rect 506 -3139 510 -3135
rect 620 -3139 624 -3135
rect 672 -3139 676 -3135
rect 864 -3139 868 -3135
rect 978 -3139 982 -3135
rect 1030 -3139 1034 -3135
rect 1222 -3139 1226 -3135
rect 1336 -3139 1340 -3135
rect 1388 -3139 1392 -3135
rect -1490 -3146 -1486 -3142
rect -1452 -3146 -1448 -3142
rect -1165 -3146 -1161 -3142
rect -1127 -3146 -1123 -3142
rect -866 -3146 -862 -3142
rect -828 -3146 -824 -3142
rect -508 -3146 -504 -3142
rect -470 -3146 -466 -3142
rect -150 -3146 -146 -3142
rect -112 -3146 -108 -3142
rect 208 -3146 212 -3142
rect 246 -3146 250 -3142
rect 564 -3146 568 -3142
rect 602 -3146 606 -3142
rect 922 -3146 926 -3142
rect 960 -3146 964 -3142
rect 1280 -3146 1284 -3142
rect 1318 -3146 1322 -3142
rect -1532 -3288 -1528 -3284
rect -1494 -3288 -1490 -3284
rect -1434 -3288 -1430 -3284
rect -1410 -3288 -1406 -3284
rect -1207 -3288 -1203 -3284
rect -1169 -3288 -1165 -3284
rect -1109 -3288 -1105 -3284
rect -1085 -3288 -1081 -3284
rect -908 -3288 -904 -3284
rect -870 -3288 -866 -3284
rect -810 -3288 -806 -3284
rect -786 -3288 -782 -3284
rect -550 -3288 -546 -3284
rect -512 -3288 -508 -3284
rect -452 -3288 -448 -3284
rect -428 -3288 -424 -3284
rect -192 -3288 -188 -3284
rect -154 -3288 -150 -3284
rect -94 -3288 -90 -3284
rect -70 -3288 -66 -3284
rect 166 -3288 170 -3284
rect 204 -3288 208 -3284
rect 264 -3288 268 -3284
rect 288 -3288 292 -3284
rect 522 -3288 526 -3284
rect 560 -3288 564 -3284
rect 620 -3288 624 -3284
rect 644 -3288 648 -3284
rect 880 -3288 884 -3284
rect 918 -3288 922 -3284
rect 978 -3288 982 -3284
rect 1002 -3288 1006 -3284
rect 1238 -3288 1242 -3284
rect 1276 -3288 1280 -3284
rect 1336 -3288 1340 -3284
rect 1360 -3288 1364 -3284
rect -1552 -3296 -1548 -3292
rect -1518 -3296 -1514 -3292
rect -1466 -3296 -1462 -3292
rect -1406 -3296 -1402 -3292
rect -1368 -3296 -1364 -3292
rect -1227 -3296 -1223 -3292
rect -1193 -3296 -1189 -3292
rect -1141 -3296 -1137 -3292
rect -1081 -3296 -1077 -3292
rect -1043 -3296 -1039 -3292
rect -928 -3296 -924 -3292
rect -894 -3296 -890 -3292
rect -842 -3296 -838 -3292
rect -782 -3296 -778 -3292
rect -744 -3296 -740 -3292
rect -570 -3296 -566 -3292
rect -536 -3296 -532 -3292
rect -484 -3296 -480 -3292
rect -424 -3296 -420 -3292
rect -386 -3296 -382 -3292
rect -212 -3296 -208 -3292
rect -178 -3296 -174 -3292
rect -126 -3296 -122 -3292
rect -66 -3296 -62 -3292
rect -28 -3296 -24 -3292
rect 146 -3296 150 -3292
rect 180 -3296 184 -3292
rect 232 -3296 236 -3292
rect 292 -3296 296 -3292
rect 330 -3296 334 -3292
rect 502 -3296 506 -3292
rect 536 -3296 540 -3292
rect 588 -3296 592 -3292
rect 648 -3296 652 -3292
rect 686 -3296 690 -3292
rect 860 -3296 864 -3292
rect 894 -3296 898 -3292
rect 946 -3296 950 -3292
rect 1006 -3296 1010 -3292
rect 1044 -3296 1048 -3292
rect 1218 -3296 1222 -3292
rect 1252 -3296 1256 -3292
rect 1304 -3296 1308 -3292
rect 1364 -3296 1368 -3292
rect 1402 -3296 1406 -3292
rect -1508 -3303 -1504 -3299
rect -1476 -3303 -1472 -3299
rect -1424 -3303 -1420 -3299
rect -1392 -3303 -1388 -3299
rect -1183 -3303 -1179 -3299
rect -1151 -3303 -1147 -3299
rect -1099 -3303 -1095 -3299
rect -1067 -3303 -1063 -3299
rect -884 -3303 -880 -3299
rect -852 -3303 -848 -3299
rect -800 -3303 -796 -3299
rect -768 -3303 -764 -3299
rect -526 -3303 -522 -3299
rect -494 -3303 -490 -3299
rect -442 -3303 -438 -3299
rect -410 -3303 -406 -3299
rect -168 -3303 -164 -3299
rect -136 -3303 -132 -3299
rect -84 -3303 -80 -3299
rect -52 -3303 -48 -3299
rect 190 -3303 194 -3299
rect 222 -3303 226 -3299
rect 274 -3303 278 -3299
rect 306 -3303 310 -3299
rect 546 -3303 550 -3299
rect 578 -3303 582 -3299
rect 630 -3303 634 -3299
rect 662 -3303 666 -3299
rect 904 -3303 908 -3299
rect 936 -3303 940 -3299
rect 988 -3303 992 -3299
rect 1020 -3303 1024 -3299
rect 1262 -3303 1266 -3299
rect 1294 -3303 1298 -3299
rect 1346 -3303 1350 -3299
rect 1378 -3303 1382 -3299
rect -1548 -3310 -1544 -3306
rect -1434 -3310 -1430 -3306
rect -1382 -3310 -1378 -3306
rect -1223 -3310 -1219 -3306
rect -1109 -3310 -1105 -3306
rect -1057 -3310 -1053 -3306
rect -924 -3310 -920 -3306
rect -810 -3310 -806 -3306
rect -758 -3310 -754 -3306
rect -566 -3310 -562 -3306
rect -452 -3310 -448 -3306
rect -400 -3310 -396 -3306
rect -208 -3310 -204 -3306
rect -94 -3310 -90 -3306
rect -42 -3310 -38 -3306
rect 150 -3310 154 -3306
rect 264 -3310 268 -3306
rect 316 -3310 320 -3306
rect 506 -3310 510 -3306
rect 620 -3310 624 -3306
rect 672 -3310 676 -3306
rect 864 -3310 868 -3306
rect 978 -3310 982 -3306
rect 1030 -3310 1034 -3306
rect 1222 -3310 1226 -3306
rect 1336 -3310 1340 -3306
rect 1388 -3310 1392 -3306
rect -1490 -3317 -1486 -3313
rect -1452 -3317 -1448 -3313
rect -1165 -3317 -1161 -3313
rect -1127 -3317 -1123 -3313
rect -866 -3317 -862 -3313
rect -828 -3317 -824 -3313
rect -508 -3317 -504 -3313
rect -470 -3317 -466 -3313
rect -150 -3317 -146 -3313
rect -112 -3317 -108 -3313
rect 208 -3317 212 -3313
rect 246 -3317 250 -3313
rect 564 -3317 568 -3313
rect 602 -3317 606 -3313
rect 922 -3317 926 -3313
rect 960 -3317 964 -3313
rect 1280 -3317 1284 -3313
rect 1318 -3317 1322 -3313
rect -1308 -3383 -1304 -3379
rect -934 -3383 -930 -3379
rect -576 -3383 -572 -3379
rect -218 -3383 -214 -3379
rect 140 -3383 144 -3379
rect 496 -3383 500 -3379
rect 854 -3383 858 -3379
rect 1212 -3383 1216 -3379
rect -1297 -3391 -1293 -3387
rect -923 -3391 -919 -3387
rect -565 -3391 -561 -3387
rect -207 -3391 -203 -3387
rect 151 -3391 155 -3387
rect 507 -3391 511 -3387
rect 865 -3391 869 -3387
rect 1223 -3391 1227 -3387
rect -924 -3529 -920 -3525
rect -858 -3529 -854 -3525
rect -824 -3529 -820 -3525
rect -780 -3529 -776 -3525
rect -746 -3529 -742 -3525
rect -566 -3529 -562 -3525
rect -500 -3529 -496 -3525
rect -466 -3529 -462 -3525
rect -422 -3529 -418 -3525
rect -388 -3529 -384 -3525
rect -208 -3529 -204 -3525
rect -142 -3529 -138 -3525
rect -108 -3529 -104 -3525
rect -64 -3529 -60 -3525
rect -30 -3529 -26 -3525
rect 150 -3529 154 -3525
rect 216 -3529 220 -3525
rect 250 -3529 254 -3525
rect 294 -3529 298 -3525
rect 328 -3529 332 -3525
rect 506 -3529 510 -3525
rect 572 -3529 576 -3525
rect 606 -3529 610 -3525
rect 650 -3529 654 -3525
rect 684 -3529 688 -3525
rect 864 -3529 868 -3525
rect 930 -3529 934 -3525
rect 964 -3529 968 -3525
rect 1008 -3529 1012 -3525
rect 1042 -3529 1046 -3525
rect 1222 -3529 1226 -3525
rect 1288 -3529 1292 -3525
rect 1322 -3529 1326 -3525
rect 1366 -3529 1370 -3525
rect 1400 -3529 1404 -3525
rect -882 -3536 -878 -3532
rect -524 -3536 -520 -3532
rect -166 -3536 -162 -3532
rect 192 -3536 196 -3532
rect 548 -3536 552 -3532
rect 906 -3536 910 -3532
rect 1264 -3536 1268 -3532
rect -848 -3543 -844 -3539
rect -706 -3543 -702 -3539
rect -490 -3543 -486 -3539
rect -348 -3543 -344 -3539
rect -132 -3543 -128 -3539
rect 10 -3543 14 -3539
rect 226 -3543 230 -3539
rect 368 -3543 372 -3539
rect 582 -3543 586 -3539
rect 724 -3543 728 -3539
rect 940 -3543 944 -3539
rect 1082 -3543 1086 -3539
rect 1298 -3543 1302 -3539
rect 1440 -3543 1444 -3539
rect -928 -3550 -924 -3546
rect -898 -3550 -894 -3546
rect -780 -3550 -776 -3546
rect -570 -3550 -566 -3546
rect -540 -3550 -536 -3546
rect -422 -3550 -418 -3546
rect -212 -3550 -208 -3546
rect -182 -3550 -178 -3546
rect -64 -3550 -60 -3546
rect 146 -3550 150 -3546
rect 176 -3550 180 -3546
rect 294 -3550 298 -3546
rect 502 -3550 506 -3546
rect 532 -3550 536 -3546
rect 650 -3550 654 -3546
rect 860 -3550 864 -3546
rect 890 -3550 894 -3546
rect 1008 -3550 1012 -3546
rect 1218 -3550 1222 -3546
rect 1248 -3550 1252 -3546
rect 1366 -3550 1370 -3546
rect -1173 -3559 -1169 -3555
rect -902 -3558 -898 -3554
rect -804 -3558 -800 -3554
rect -544 -3558 -540 -3554
rect -446 -3558 -442 -3554
rect -186 -3558 -182 -3554
rect -88 -3558 -84 -3554
rect 172 -3558 176 -3554
rect 270 -3558 274 -3554
rect 528 -3558 532 -3554
rect 626 -3558 630 -3554
rect 886 -3558 890 -3554
rect 984 -3558 988 -3554
rect 1244 -3558 1248 -3554
rect 1342 -3558 1346 -3554
rect -1223 -3566 -1219 -3562
rect -1183 -3566 -1179 -3562
rect -1163 -3566 -1159 -3562
rect -924 -3565 -920 -3561
rect -776 -3565 -772 -3561
rect -566 -3565 -562 -3561
rect -418 -3565 -414 -3561
rect -208 -3565 -204 -3561
rect -60 -3565 -56 -3561
rect 150 -3565 154 -3561
rect 298 -3565 302 -3561
rect 506 -3565 510 -3561
rect 654 -3565 658 -3561
rect 864 -3565 868 -3561
rect 1012 -3565 1016 -3561
rect 1222 -3565 1226 -3561
rect 1370 -3565 1374 -3561
rect -1227 -3573 -1223 -3569
rect -1197 -3573 -1193 -3569
rect -1149 -3573 -1145 -3569
rect -902 -3572 -898 -3568
rect -794 -3572 -790 -3568
rect -760 -3572 -756 -3568
rect -544 -3572 -540 -3568
rect -436 -3572 -432 -3568
rect -402 -3572 -398 -3568
rect -186 -3572 -182 -3568
rect -78 -3572 -74 -3568
rect -44 -3572 -40 -3568
rect 172 -3572 176 -3568
rect 280 -3572 284 -3568
rect 314 -3572 318 -3568
rect 528 -3572 532 -3568
rect 636 -3572 640 -3568
rect 670 -3572 674 -3568
rect 886 -3572 890 -3568
rect 994 -3572 998 -3568
rect 1028 -3572 1032 -3568
rect 1244 -3572 1248 -3568
rect 1352 -3572 1356 -3568
rect 1386 -3572 1390 -3568
rect -928 -3579 -924 -3575
rect -872 -3579 -868 -3575
rect -838 -3579 -834 -3575
rect -570 -3579 -566 -3575
rect -514 -3579 -510 -3575
rect -480 -3579 -476 -3575
rect -212 -3579 -208 -3575
rect -156 -3579 -152 -3575
rect -122 -3579 -118 -3575
rect 146 -3579 150 -3575
rect 202 -3579 206 -3575
rect 236 -3579 240 -3575
rect 502 -3579 506 -3575
rect 558 -3579 562 -3575
rect 592 -3579 596 -3575
rect 860 -3579 864 -3575
rect 916 -3579 920 -3575
rect 950 -3579 954 -3575
rect 1218 -3579 1222 -3575
rect 1274 -3579 1278 -3575
rect 1308 -3579 1312 -3575
rect -1795 -3688 -1791 -3684
rect -1757 -3688 -1753 -3684
rect -1697 -3688 -1693 -3684
rect -1673 -3688 -1669 -3684
rect -1532 -3688 -1528 -3684
rect -1494 -3688 -1490 -3684
rect -1434 -3688 -1430 -3684
rect -1410 -3688 -1406 -3684
rect -1207 -3688 -1203 -3684
rect -1169 -3688 -1165 -3684
rect -1109 -3688 -1105 -3684
rect -1085 -3688 -1081 -3684
rect -907 -3688 -903 -3684
rect -869 -3688 -865 -3684
rect -809 -3688 -805 -3684
rect -785 -3688 -781 -3684
rect -550 -3688 -546 -3684
rect -512 -3688 -508 -3684
rect -452 -3688 -448 -3684
rect -428 -3688 -424 -3684
rect -192 -3688 -188 -3684
rect -154 -3688 -150 -3684
rect -94 -3688 -90 -3684
rect -70 -3688 -66 -3684
rect -1815 -3696 -1811 -3692
rect -1781 -3696 -1777 -3692
rect -1729 -3696 -1725 -3692
rect -1669 -3696 -1665 -3692
rect -1631 -3696 -1627 -3692
rect -1552 -3696 -1548 -3692
rect -1518 -3696 -1514 -3692
rect -1466 -3696 -1462 -3692
rect -1406 -3696 -1402 -3692
rect -1368 -3696 -1364 -3692
rect -1227 -3696 -1223 -3692
rect -1193 -3696 -1189 -3692
rect -1141 -3696 -1137 -3692
rect -1081 -3696 -1077 -3692
rect -1043 -3696 -1039 -3692
rect -927 -3696 -923 -3692
rect -893 -3696 -889 -3692
rect -841 -3696 -837 -3692
rect -781 -3696 -777 -3692
rect -743 -3696 -739 -3692
rect -570 -3696 -566 -3692
rect -536 -3696 -532 -3692
rect -484 -3696 -480 -3692
rect -424 -3696 -420 -3692
rect -386 -3696 -382 -3692
rect -212 -3696 -208 -3692
rect -178 -3696 -174 -3692
rect -126 -3696 -122 -3692
rect -66 -3696 -62 -3692
rect -28 -3696 -24 -3692
rect -1771 -3703 -1767 -3699
rect -1739 -3703 -1735 -3699
rect -1687 -3703 -1683 -3699
rect -1655 -3703 -1651 -3699
rect -1508 -3703 -1504 -3699
rect -1476 -3703 -1472 -3699
rect -1424 -3703 -1420 -3699
rect -1392 -3703 -1388 -3699
rect -1183 -3703 -1179 -3699
rect -1151 -3703 -1147 -3699
rect -1099 -3703 -1095 -3699
rect -1067 -3703 -1063 -3699
rect -883 -3703 -879 -3699
rect -851 -3703 -847 -3699
rect -799 -3703 -795 -3699
rect -767 -3703 -763 -3699
rect -526 -3703 -522 -3699
rect -494 -3703 -490 -3699
rect -442 -3703 -438 -3699
rect -410 -3703 -406 -3699
rect -168 -3703 -164 -3699
rect -136 -3703 -132 -3699
rect -84 -3703 -80 -3699
rect -52 -3703 -48 -3699
rect -1811 -3710 -1807 -3706
rect -1697 -3710 -1693 -3706
rect -1645 -3710 -1641 -3706
rect -1548 -3710 -1544 -3706
rect -1434 -3710 -1430 -3706
rect -1382 -3710 -1378 -3706
rect -1223 -3710 -1219 -3706
rect -1109 -3710 -1105 -3706
rect -1057 -3710 -1053 -3706
rect -923 -3710 -919 -3706
rect -809 -3710 -805 -3706
rect -757 -3710 -753 -3706
rect -566 -3710 -562 -3706
rect -452 -3710 -448 -3706
rect -400 -3710 -396 -3706
rect -208 -3710 -204 -3706
rect -94 -3710 -90 -3706
rect -42 -3710 -38 -3706
rect -1753 -3717 -1749 -3713
rect -1715 -3717 -1711 -3713
rect -1490 -3717 -1486 -3713
rect -1452 -3717 -1448 -3713
rect -1165 -3717 -1161 -3713
rect -1127 -3717 -1123 -3713
rect -865 -3717 -861 -3713
rect -827 -3717 -823 -3713
rect -508 -3717 -504 -3713
rect -470 -3717 -466 -3713
rect -150 -3717 -146 -3713
rect -112 -3717 -108 -3713
rect -1532 -3859 -1528 -3855
rect -1494 -3859 -1490 -3855
rect -1434 -3859 -1430 -3855
rect -1410 -3859 -1406 -3855
rect -1207 -3859 -1203 -3855
rect -1169 -3859 -1165 -3855
rect -1109 -3859 -1105 -3855
rect -1085 -3859 -1081 -3855
rect -907 -3859 -903 -3855
rect -869 -3859 -865 -3855
rect -809 -3859 -805 -3855
rect -785 -3859 -781 -3855
rect -550 -3859 -546 -3855
rect -512 -3859 -508 -3855
rect -452 -3859 -448 -3855
rect -428 -3859 -424 -3855
rect -192 -3859 -188 -3855
rect -154 -3859 -150 -3855
rect -94 -3859 -90 -3855
rect -70 -3859 -66 -3855
rect 166 -3859 170 -3855
rect 204 -3859 208 -3855
rect 264 -3859 268 -3855
rect 288 -3859 292 -3855
rect 522 -3859 526 -3855
rect 560 -3859 564 -3855
rect 620 -3859 624 -3855
rect 644 -3859 648 -3855
rect 880 -3859 884 -3855
rect 918 -3859 922 -3855
rect 978 -3859 982 -3855
rect 1002 -3859 1006 -3855
rect 1238 -3859 1242 -3855
rect 1276 -3859 1280 -3855
rect 1336 -3859 1340 -3855
rect 1360 -3859 1364 -3855
rect -1552 -3867 -1548 -3863
rect -1518 -3867 -1514 -3863
rect -1466 -3867 -1462 -3863
rect -1406 -3867 -1402 -3863
rect -1368 -3867 -1364 -3863
rect -1227 -3867 -1223 -3863
rect -1193 -3867 -1189 -3863
rect -1141 -3867 -1137 -3863
rect -1081 -3867 -1077 -3863
rect -1043 -3867 -1039 -3863
rect -927 -3867 -923 -3863
rect -893 -3867 -889 -3863
rect -841 -3867 -837 -3863
rect -781 -3867 -777 -3863
rect -743 -3867 -739 -3863
rect -570 -3867 -566 -3863
rect -536 -3867 -532 -3863
rect -484 -3867 -480 -3863
rect -424 -3867 -420 -3863
rect -386 -3867 -382 -3863
rect -212 -3867 -208 -3863
rect -178 -3867 -174 -3863
rect -126 -3867 -122 -3863
rect -66 -3867 -62 -3863
rect -28 -3867 -24 -3863
rect 146 -3867 150 -3863
rect 180 -3867 184 -3863
rect 232 -3867 236 -3863
rect 292 -3867 296 -3863
rect 330 -3867 334 -3863
rect 502 -3867 506 -3863
rect 536 -3867 540 -3863
rect 588 -3867 592 -3863
rect 648 -3867 652 -3863
rect 686 -3867 690 -3863
rect 860 -3867 864 -3863
rect 894 -3867 898 -3863
rect 946 -3867 950 -3863
rect 1006 -3867 1010 -3863
rect 1044 -3867 1048 -3863
rect 1218 -3867 1222 -3863
rect 1252 -3867 1256 -3863
rect 1304 -3867 1308 -3863
rect 1364 -3867 1368 -3863
rect 1402 -3867 1406 -3863
rect -1508 -3874 -1504 -3870
rect -1476 -3874 -1472 -3870
rect -1424 -3874 -1420 -3870
rect -1392 -3874 -1388 -3870
rect -1183 -3874 -1179 -3870
rect -1151 -3874 -1147 -3870
rect -1099 -3874 -1095 -3870
rect -1067 -3874 -1063 -3870
rect -883 -3874 -879 -3870
rect -851 -3874 -847 -3870
rect -799 -3874 -795 -3870
rect -767 -3874 -763 -3870
rect -526 -3874 -522 -3870
rect -494 -3874 -490 -3870
rect -442 -3874 -438 -3870
rect -410 -3874 -406 -3870
rect -168 -3874 -164 -3870
rect -136 -3874 -132 -3870
rect -84 -3874 -80 -3870
rect -52 -3874 -48 -3870
rect 190 -3874 194 -3870
rect 222 -3874 226 -3870
rect 274 -3874 278 -3870
rect 306 -3874 310 -3870
rect 546 -3874 550 -3870
rect 578 -3874 582 -3870
rect 630 -3874 634 -3870
rect 662 -3874 666 -3870
rect 904 -3874 908 -3870
rect 936 -3874 940 -3870
rect 988 -3874 992 -3870
rect 1020 -3874 1024 -3870
rect 1262 -3874 1266 -3870
rect 1294 -3874 1298 -3870
rect 1346 -3874 1350 -3870
rect 1378 -3874 1382 -3870
rect -1548 -3881 -1544 -3877
rect -1434 -3881 -1430 -3877
rect -1382 -3881 -1378 -3877
rect -1223 -3881 -1219 -3877
rect -1109 -3881 -1105 -3877
rect -1057 -3881 -1053 -3877
rect -923 -3881 -919 -3877
rect -809 -3881 -805 -3877
rect -757 -3881 -753 -3877
rect -566 -3881 -562 -3877
rect -452 -3881 -448 -3877
rect -400 -3881 -396 -3877
rect -208 -3881 -204 -3877
rect -94 -3881 -90 -3877
rect -42 -3881 -38 -3877
rect 150 -3881 154 -3877
rect 264 -3881 268 -3877
rect 316 -3881 320 -3877
rect 506 -3881 510 -3877
rect 620 -3881 624 -3877
rect 672 -3881 676 -3877
rect 864 -3881 868 -3877
rect 978 -3881 982 -3877
rect 1030 -3881 1034 -3877
rect 1222 -3881 1226 -3877
rect 1336 -3881 1340 -3877
rect 1388 -3881 1392 -3877
rect -1490 -3888 -1486 -3884
rect -1452 -3888 -1448 -3884
rect -1165 -3888 -1161 -3884
rect -1127 -3888 -1123 -3884
rect -865 -3888 -861 -3884
rect -827 -3888 -823 -3884
rect -508 -3888 -504 -3884
rect -470 -3888 -466 -3884
rect -150 -3888 -146 -3884
rect -112 -3888 -108 -3884
rect 208 -3888 212 -3884
rect 246 -3888 250 -3884
rect 564 -3888 568 -3884
rect 602 -3888 606 -3884
rect 922 -3888 926 -3884
rect 960 -3888 964 -3884
rect 1280 -3888 1284 -3884
rect 1318 -3888 1322 -3884
rect -1532 -4034 -1528 -4030
rect -1494 -4034 -1490 -4030
rect -1434 -4034 -1430 -4030
rect -1410 -4034 -1406 -4030
rect -1207 -4034 -1203 -4030
rect -1169 -4034 -1165 -4030
rect -1109 -4034 -1105 -4030
rect -1085 -4034 -1081 -4030
rect -908 -4034 -904 -4030
rect -870 -4034 -866 -4030
rect -810 -4034 -806 -4030
rect -786 -4034 -782 -4030
rect -550 -4034 -546 -4030
rect -512 -4034 -508 -4030
rect -452 -4034 -448 -4030
rect -428 -4034 -424 -4030
rect -192 -4034 -188 -4030
rect -154 -4034 -150 -4030
rect -94 -4034 -90 -4030
rect -70 -4034 -66 -4030
rect 166 -4034 170 -4030
rect 204 -4034 208 -4030
rect 264 -4034 268 -4030
rect 288 -4034 292 -4030
rect 522 -4034 526 -4030
rect 560 -4034 564 -4030
rect 620 -4034 624 -4030
rect 644 -4034 648 -4030
rect 880 -4034 884 -4030
rect 918 -4034 922 -4030
rect 978 -4034 982 -4030
rect 1002 -4034 1006 -4030
rect 1238 -4034 1242 -4030
rect 1276 -4034 1280 -4030
rect 1336 -4034 1340 -4030
rect 1360 -4034 1364 -4030
rect -1552 -4042 -1548 -4038
rect -1518 -4042 -1514 -4038
rect -1466 -4042 -1462 -4038
rect -1406 -4042 -1402 -4038
rect -1368 -4042 -1364 -4038
rect -1227 -4042 -1223 -4038
rect -1193 -4042 -1189 -4038
rect -1141 -4042 -1137 -4038
rect -1081 -4042 -1077 -4038
rect -1043 -4042 -1039 -4038
rect -928 -4042 -924 -4038
rect -894 -4042 -890 -4038
rect -842 -4042 -838 -4038
rect -782 -4042 -778 -4038
rect -744 -4042 -740 -4038
rect -570 -4042 -566 -4038
rect -536 -4042 -532 -4038
rect -484 -4042 -480 -4038
rect -424 -4042 -420 -4038
rect -386 -4042 -382 -4038
rect -212 -4042 -208 -4038
rect -178 -4042 -174 -4038
rect -126 -4042 -122 -4038
rect -66 -4042 -62 -4038
rect -28 -4042 -24 -4038
rect 146 -4042 150 -4038
rect 180 -4042 184 -4038
rect 232 -4042 236 -4038
rect 292 -4042 296 -4038
rect 330 -4042 334 -4038
rect 502 -4042 506 -4038
rect 536 -4042 540 -4038
rect 588 -4042 592 -4038
rect 648 -4042 652 -4038
rect 686 -4042 690 -4038
rect 860 -4042 864 -4038
rect 894 -4042 898 -4038
rect 946 -4042 950 -4038
rect 1006 -4042 1010 -4038
rect 1044 -4042 1048 -4038
rect 1218 -4042 1222 -4038
rect 1252 -4042 1256 -4038
rect 1304 -4042 1308 -4038
rect 1364 -4042 1368 -4038
rect 1402 -4042 1406 -4038
rect -1508 -4049 -1504 -4045
rect -1476 -4049 -1472 -4045
rect -1424 -4049 -1420 -4045
rect -1392 -4049 -1388 -4045
rect -1183 -4049 -1179 -4045
rect -1151 -4049 -1147 -4045
rect -1099 -4049 -1095 -4045
rect -1067 -4049 -1063 -4045
rect -884 -4049 -880 -4045
rect -852 -4049 -848 -4045
rect -800 -4049 -796 -4045
rect -768 -4049 -764 -4045
rect -526 -4049 -522 -4045
rect -494 -4049 -490 -4045
rect -442 -4049 -438 -4045
rect -410 -4049 -406 -4045
rect -168 -4049 -164 -4045
rect -136 -4049 -132 -4045
rect -84 -4049 -80 -4045
rect -52 -4049 -48 -4045
rect 190 -4049 194 -4045
rect 222 -4049 226 -4045
rect 274 -4049 278 -4045
rect 306 -4049 310 -4045
rect 546 -4049 550 -4045
rect 578 -4049 582 -4045
rect 630 -4049 634 -4045
rect 662 -4049 666 -4045
rect 904 -4049 908 -4045
rect 936 -4049 940 -4045
rect 988 -4049 992 -4045
rect 1020 -4049 1024 -4045
rect 1262 -4049 1266 -4045
rect 1294 -4049 1298 -4045
rect 1346 -4049 1350 -4045
rect 1378 -4049 1382 -4045
rect -1548 -4056 -1544 -4052
rect -1434 -4056 -1430 -4052
rect -1382 -4056 -1378 -4052
rect -1223 -4056 -1219 -4052
rect -1109 -4056 -1105 -4052
rect -1057 -4056 -1053 -4052
rect -924 -4056 -920 -4052
rect -810 -4056 -806 -4052
rect -758 -4056 -754 -4052
rect -566 -4056 -562 -4052
rect -452 -4056 -448 -4052
rect -400 -4056 -396 -4052
rect -208 -4056 -204 -4052
rect -94 -4056 -90 -4052
rect -42 -4056 -38 -4052
rect 150 -4056 154 -4052
rect 264 -4056 268 -4052
rect 316 -4056 320 -4052
rect 506 -4056 510 -4052
rect 620 -4056 624 -4052
rect 672 -4056 676 -4052
rect 864 -4056 868 -4052
rect 978 -4056 982 -4052
rect 1030 -4056 1034 -4052
rect 1222 -4056 1226 -4052
rect 1336 -4056 1340 -4052
rect 1388 -4056 1392 -4052
rect -1490 -4063 -1486 -4059
rect -1452 -4063 -1448 -4059
rect -1165 -4063 -1161 -4059
rect -1127 -4063 -1123 -4059
rect -866 -4063 -862 -4059
rect -828 -4063 -824 -4059
rect -508 -4063 -504 -4059
rect -470 -4063 -466 -4059
rect -150 -4063 -146 -4059
rect -112 -4063 -108 -4059
rect 208 -4063 212 -4059
rect 246 -4063 250 -4059
rect 564 -4063 568 -4059
rect 602 -4063 606 -4059
rect 922 -4063 926 -4059
rect 960 -4063 964 -4059
rect 1280 -4063 1284 -4059
rect 1318 -4063 1322 -4059
rect -1308 -4133 -1304 -4129
rect -934 -4133 -930 -4129
rect -576 -4133 -572 -4129
rect -218 -4133 -214 -4129
rect 140 -4133 144 -4129
rect 496 -4133 500 -4129
rect 854 -4133 858 -4129
rect 1212 -4133 1216 -4129
rect -1297 -4141 -1293 -4137
rect -923 -4141 -919 -4137
rect -565 -4141 -561 -4137
rect -207 -4141 -203 -4137
rect 151 -4141 155 -4137
rect 507 -4141 511 -4137
rect 865 -4141 869 -4137
rect 1223 -4141 1227 -4137
rect -924 -4279 -920 -4275
rect -858 -4279 -854 -4275
rect -824 -4279 -820 -4275
rect -780 -4279 -776 -4275
rect -746 -4279 -742 -4275
rect -566 -4279 -562 -4275
rect -500 -4279 -496 -4275
rect -466 -4279 -462 -4275
rect -422 -4279 -418 -4275
rect -388 -4279 -384 -4275
rect -208 -4279 -204 -4275
rect -142 -4279 -138 -4275
rect -108 -4279 -104 -4275
rect -64 -4279 -60 -4275
rect -30 -4279 -26 -4275
rect 150 -4279 154 -4275
rect 216 -4279 220 -4275
rect 250 -4279 254 -4275
rect 294 -4279 298 -4275
rect 328 -4279 332 -4275
rect 506 -4279 510 -4275
rect 572 -4279 576 -4275
rect 606 -4279 610 -4275
rect 650 -4279 654 -4275
rect 684 -4279 688 -4275
rect 864 -4279 868 -4275
rect 930 -4279 934 -4275
rect 964 -4279 968 -4275
rect 1008 -4279 1012 -4275
rect 1042 -4279 1046 -4275
rect 1222 -4279 1226 -4275
rect 1288 -4279 1292 -4275
rect 1322 -4279 1326 -4275
rect 1366 -4279 1370 -4275
rect 1400 -4279 1404 -4275
rect -882 -4286 -878 -4282
rect -524 -4286 -520 -4282
rect -166 -4286 -162 -4282
rect 192 -4286 196 -4282
rect 548 -4286 552 -4282
rect 906 -4286 910 -4282
rect 1264 -4286 1268 -4282
rect -848 -4293 -844 -4289
rect -706 -4293 -702 -4289
rect -490 -4293 -486 -4289
rect -348 -4293 -344 -4289
rect -132 -4293 -128 -4289
rect 10 -4293 14 -4289
rect 226 -4293 230 -4289
rect 368 -4293 372 -4289
rect 582 -4293 586 -4289
rect 724 -4293 728 -4289
rect 940 -4293 944 -4289
rect 1082 -4293 1086 -4289
rect 1298 -4293 1302 -4289
rect 1440 -4293 1444 -4289
rect -928 -4300 -924 -4296
rect -898 -4300 -894 -4296
rect -780 -4300 -776 -4296
rect -570 -4300 -566 -4296
rect -540 -4300 -536 -4296
rect -422 -4300 -418 -4296
rect -212 -4300 -208 -4296
rect -182 -4300 -178 -4296
rect -64 -4300 -60 -4296
rect 146 -4300 150 -4296
rect 176 -4300 180 -4296
rect 294 -4300 298 -4296
rect 502 -4300 506 -4296
rect 532 -4300 536 -4296
rect 650 -4300 654 -4296
rect 860 -4300 864 -4296
rect 890 -4300 894 -4296
rect 1008 -4300 1012 -4296
rect 1218 -4300 1222 -4296
rect 1248 -4300 1252 -4296
rect 1366 -4300 1370 -4296
rect -1173 -4309 -1169 -4305
rect -902 -4308 -898 -4304
rect -804 -4308 -800 -4304
rect -544 -4308 -540 -4304
rect -446 -4308 -442 -4304
rect -186 -4308 -182 -4304
rect -88 -4308 -84 -4304
rect 172 -4308 176 -4304
rect 270 -4308 274 -4304
rect 528 -4308 532 -4304
rect 626 -4308 630 -4304
rect 886 -4308 890 -4304
rect 984 -4308 988 -4304
rect 1244 -4308 1248 -4304
rect 1342 -4308 1346 -4304
rect -1223 -4316 -1219 -4312
rect -1183 -4316 -1179 -4312
rect -1163 -4316 -1159 -4312
rect -924 -4315 -920 -4311
rect -776 -4315 -772 -4311
rect -566 -4315 -562 -4311
rect -418 -4315 -414 -4311
rect -208 -4315 -204 -4311
rect -60 -4315 -56 -4311
rect 150 -4315 154 -4311
rect 298 -4315 302 -4311
rect 506 -4315 510 -4311
rect 654 -4315 658 -4311
rect 864 -4315 868 -4311
rect 1012 -4315 1016 -4311
rect 1222 -4315 1226 -4311
rect 1370 -4315 1374 -4311
rect -1227 -4323 -1223 -4319
rect -1197 -4323 -1193 -4319
rect -1149 -4323 -1145 -4319
rect -902 -4322 -898 -4318
rect -794 -4322 -790 -4318
rect -760 -4322 -756 -4318
rect -544 -4322 -540 -4318
rect -436 -4322 -432 -4318
rect -402 -4322 -398 -4318
rect -186 -4322 -182 -4318
rect -78 -4322 -74 -4318
rect -44 -4322 -40 -4318
rect 172 -4322 176 -4318
rect 280 -4322 284 -4318
rect 314 -4322 318 -4318
rect 528 -4322 532 -4318
rect 636 -4322 640 -4318
rect 670 -4322 674 -4318
rect 886 -4322 890 -4318
rect 994 -4322 998 -4318
rect 1028 -4322 1032 -4318
rect 1244 -4322 1248 -4318
rect 1352 -4322 1356 -4318
rect 1386 -4322 1390 -4318
rect -928 -4329 -924 -4325
rect -872 -4329 -868 -4325
rect -838 -4329 -834 -4325
rect -570 -4329 -566 -4325
rect -514 -4329 -510 -4325
rect -480 -4329 -476 -4325
rect -212 -4329 -208 -4325
rect -156 -4329 -152 -4325
rect -122 -4329 -118 -4325
rect 146 -4329 150 -4325
rect 202 -4329 206 -4325
rect 236 -4329 240 -4325
rect 502 -4329 506 -4325
rect 558 -4329 562 -4325
rect 592 -4329 596 -4325
rect 860 -4329 864 -4325
rect 916 -4329 920 -4325
rect 950 -4329 954 -4325
rect 1218 -4329 1222 -4325
rect 1274 -4329 1278 -4325
rect 1308 -4329 1312 -4325
rect -1787 -4431 -1783 -4427
rect -1749 -4431 -1745 -4427
rect -1689 -4431 -1685 -4427
rect -1665 -4431 -1661 -4427
rect -1524 -4431 -1520 -4427
rect -1486 -4431 -1482 -4427
rect -1426 -4431 -1422 -4427
rect -1402 -4431 -1398 -4427
rect -1207 -4431 -1203 -4427
rect -1169 -4431 -1165 -4427
rect -1109 -4431 -1105 -4427
rect -1085 -4431 -1081 -4427
rect -908 -4431 -904 -4427
rect -870 -4431 -866 -4427
rect -810 -4431 -806 -4427
rect -786 -4431 -782 -4427
rect -550 -4431 -546 -4427
rect -512 -4431 -508 -4427
rect -452 -4431 -448 -4427
rect -428 -4431 -424 -4427
rect -1807 -4439 -1803 -4435
rect -1773 -4439 -1769 -4435
rect -1721 -4439 -1717 -4435
rect -1661 -4439 -1657 -4435
rect -1623 -4439 -1619 -4435
rect -1544 -4439 -1540 -4435
rect -1510 -4439 -1506 -4435
rect -1458 -4439 -1454 -4435
rect -1398 -4439 -1394 -4435
rect -1360 -4439 -1356 -4435
rect -1227 -4439 -1223 -4435
rect -1193 -4439 -1189 -4435
rect -1141 -4439 -1137 -4435
rect -1081 -4439 -1077 -4435
rect -1043 -4439 -1039 -4435
rect -928 -4439 -924 -4435
rect -894 -4439 -890 -4435
rect -842 -4439 -838 -4435
rect -782 -4439 -778 -4435
rect -744 -4439 -740 -4435
rect -570 -4439 -566 -4435
rect -536 -4439 -532 -4435
rect -484 -4439 -480 -4435
rect -424 -4439 -420 -4435
rect -386 -4439 -382 -4435
rect -1763 -4446 -1759 -4442
rect -1731 -4446 -1727 -4442
rect -1679 -4446 -1675 -4442
rect -1647 -4446 -1643 -4442
rect -1500 -4446 -1496 -4442
rect -1468 -4446 -1464 -4442
rect -1416 -4446 -1412 -4442
rect -1384 -4446 -1380 -4442
rect -1183 -4446 -1179 -4442
rect -1151 -4446 -1147 -4442
rect -1099 -4446 -1095 -4442
rect -1067 -4446 -1063 -4442
rect -884 -4446 -880 -4442
rect -852 -4446 -848 -4442
rect -800 -4446 -796 -4442
rect -768 -4446 -764 -4442
rect -526 -4446 -522 -4442
rect -494 -4446 -490 -4442
rect -442 -4446 -438 -4442
rect -410 -4446 -406 -4442
rect -1803 -4453 -1799 -4449
rect -1689 -4453 -1685 -4449
rect -1637 -4453 -1633 -4449
rect -1540 -4453 -1536 -4449
rect -1426 -4453 -1422 -4449
rect -1374 -4453 -1370 -4449
rect -1223 -4453 -1219 -4449
rect -1109 -4453 -1105 -4449
rect -1057 -4453 -1053 -4449
rect -924 -4453 -920 -4449
rect -810 -4453 -806 -4449
rect -758 -4453 -754 -4449
rect -566 -4453 -562 -4449
rect -452 -4453 -448 -4449
rect -400 -4453 -396 -4449
rect -1745 -4460 -1741 -4456
rect -1707 -4460 -1703 -4456
rect -1482 -4460 -1478 -4456
rect -1444 -4460 -1440 -4456
rect -1165 -4460 -1161 -4456
rect -1127 -4460 -1123 -4456
rect -866 -4460 -862 -4456
rect -828 -4460 -824 -4456
rect -508 -4460 -504 -4456
rect -470 -4460 -466 -4456
rect -1787 -4602 -1783 -4598
rect -1749 -4602 -1745 -4598
rect -1689 -4602 -1685 -4598
rect -1665 -4602 -1661 -4598
rect -1524 -4602 -1520 -4598
rect -1486 -4602 -1482 -4598
rect -1426 -4602 -1422 -4598
rect -1402 -4602 -1398 -4598
rect -1207 -4602 -1203 -4598
rect -1169 -4602 -1165 -4598
rect -1109 -4602 -1105 -4598
rect -1085 -4602 -1081 -4598
rect -908 -4602 -904 -4598
rect -870 -4602 -866 -4598
rect -810 -4602 -806 -4598
rect -786 -4602 -782 -4598
rect -550 -4602 -546 -4598
rect -512 -4602 -508 -4598
rect -452 -4602 -448 -4598
rect -428 -4602 -424 -4598
rect -192 -4602 -188 -4598
rect -154 -4602 -150 -4598
rect -94 -4602 -90 -4598
rect -70 -4602 -66 -4598
rect 166 -4602 170 -4598
rect 204 -4602 208 -4598
rect 264 -4602 268 -4598
rect 288 -4602 292 -4598
rect 522 -4602 526 -4598
rect 560 -4602 564 -4598
rect 620 -4602 624 -4598
rect 644 -4602 648 -4598
rect 880 -4602 884 -4598
rect 918 -4602 922 -4598
rect 978 -4602 982 -4598
rect 1002 -4602 1006 -4598
rect 1238 -4602 1242 -4598
rect 1276 -4602 1280 -4598
rect 1336 -4602 1340 -4598
rect 1360 -4602 1364 -4598
rect -1807 -4610 -1803 -4606
rect -1773 -4610 -1769 -4606
rect -1721 -4610 -1717 -4606
rect -1661 -4610 -1657 -4606
rect -1623 -4610 -1619 -4606
rect -1544 -4610 -1540 -4606
rect -1510 -4610 -1506 -4606
rect -1458 -4610 -1454 -4606
rect -1398 -4610 -1394 -4606
rect -1360 -4610 -1356 -4606
rect -1227 -4610 -1223 -4606
rect -1193 -4610 -1189 -4606
rect -1141 -4610 -1137 -4606
rect -1081 -4610 -1077 -4606
rect -1043 -4610 -1039 -4606
rect -928 -4610 -924 -4606
rect -894 -4610 -890 -4606
rect -842 -4610 -838 -4606
rect -782 -4610 -778 -4606
rect -744 -4610 -740 -4606
rect -570 -4610 -566 -4606
rect -536 -4610 -532 -4606
rect -484 -4610 -480 -4606
rect -424 -4610 -420 -4606
rect -386 -4610 -382 -4606
rect -212 -4610 -208 -4606
rect -178 -4610 -174 -4606
rect -126 -4610 -122 -4606
rect -66 -4610 -62 -4606
rect -28 -4610 -24 -4606
rect 146 -4610 150 -4606
rect 180 -4610 184 -4606
rect 232 -4610 236 -4606
rect 292 -4610 296 -4606
rect 330 -4610 334 -4606
rect 502 -4610 506 -4606
rect 536 -4610 540 -4606
rect 588 -4610 592 -4606
rect 648 -4610 652 -4606
rect 686 -4610 690 -4606
rect 860 -4610 864 -4606
rect 894 -4610 898 -4606
rect 946 -4610 950 -4606
rect 1006 -4610 1010 -4606
rect 1044 -4610 1048 -4606
rect 1218 -4610 1222 -4606
rect 1252 -4610 1256 -4606
rect 1304 -4610 1308 -4606
rect 1364 -4610 1368 -4606
rect 1402 -4610 1406 -4606
rect -1763 -4617 -1759 -4613
rect -1731 -4617 -1727 -4613
rect -1679 -4617 -1675 -4613
rect -1647 -4617 -1643 -4613
rect -1500 -4617 -1496 -4613
rect -1468 -4617 -1464 -4613
rect -1416 -4617 -1412 -4613
rect -1384 -4617 -1380 -4613
rect -1183 -4617 -1179 -4613
rect -1151 -4617 -1147 -4613
rect -1099 -4617 -1095 -4613
rect -1067 -4617 -1063 -4613
rect -884 -4617 -880 -4613
rect -852 -4617 -848 -4613
rect -800 -4617 -796 -4613
rect -768 -4617 -764 -4613
rect -526 -4617 -522 -4613
rect -494 -4617 -490 -4613
rect -442 -4617 -438 -4613
rect -410 -4617 -406 -4613
rect -168 -4617 -164 -4613
rect -136 -4617 -132 -4613
rect -84 -4617 -80 -4613
rect -52 -4617 -48 -4613
rect 190 -4617 194 -4613
rect 222 -4617 226 -4613
rect 274 -4617 278 -4613
rect 306 -4617 310 -4613
rect 546 -4617 550 -4613
rect 578 -4617 582 -4613
rect 630 -4617 634 -4613
rect 662 -4617 666 -4613
rect 904 -4617 908 -4613
rect 936 -4617 940 -4613
rect 988 -4617 992 -4613
rect 1020 -4617 1024 -4613
rect 1262 -4617 1266 -4613
rect 1294 -4617 1298 -4613
rect 1346 -4617 1350 -4613
rect 1378 -4617 1382 -4613
rect -1803 -4624 -1799 -4620
rect -1689 -4624 -1685 -4620
rect -1637 -4624 -1633 -4620
rect -1540 -4624 -1536 -4620
rect -1426 -4624 -1422 -4620
rect -1374 -4624 -1370 -4620
rect -1223 -4624 -1219 -4620
rect -1109 -4624 -1105 -4620
rect -1057 -4624 -1053 -4620
rect -924 -4624 -920 -4620
rect -810 -4624 -806 -4620
rect -758 -4624 -754 -4620
rect -566 -4624 -562 -4620
rect -452 -4624 -448 -4620
rect -400 -4624 -396 -4620
rect -208 -4624 -204 -4620
rect -94 -4624 -90 -4620
rect -42 -4624 -38 -4620
rect 150 -4624 154 -4620
rect 264 -4624 268 -4620
rect 316 -4624 320 -4620
rect 506 -4624 510 -4620
rect 620 -4624 624 -4620
rect 672 -4624 676 -4620
rect 864 -4624 868 -4620
rect 978 -4624 982 -4620
rect 1030 -4624 1034 -4620
rect 1222 -4624 1226 -4620
rect 1336 -4624 1340 -4620
rect 1388 -4624 1392 -4620
rect -1745 -4631 -1741 -4627
rect -1707 -4631 -1703 -4627
rect -1482 -4631 -1478 -4627
rect -1444 -4631 -1440 -4627
rect -1165 -4631 -1161 -4627
rect -1127 -4631 -1123 -4627
rect -866 -4631 -862 -4627
rect -828 -4631 -824 -4627
rect -508 -4631 -504 -4627
rect -470 -4631 -466 -4627
rect -150 -4631 -146 -4627
rect -112 -4631 -108 -4627
rect 208 -4631 212 -4627
rect 246 -4631 250 -4627
rect 564 -4631 568 -4627
rect 602 -4631 606 -4627
rect 922 -4631 926 -4627
rect 960 -4631 964 -4627
rect 1280 -4631 1284 -4627
rect 1318 -4631 1322 -4627
rect -1524 -4773 -1520 -4769
rect -1486 -4773 -1482 -4769
rect -1426 -4773 -1422 -4769
rect -1402 -4773 -1398 -4769
rect -1207 -4773 -1203 -4769
rect -1169 -4773 -1165 -4769
rect -1109 -4773 -1105 -4769
rect -1085 -4773 -1081 -4769
rect -908 -4773 -904 -4769
rect -870 -4773 -866 -4769
rect -810 -4773 -806 -4769
rect -786 -4773 -782 -4769
rect -550 -4773 -546 -4769
rect -512 -4773 -508 -4769
rect -452 -4773 -448 -4769
rect -428 -4773 -424 -4769
rect -192 -4773 -188 -4769
rect -154 -4773 -150 -4769
rect -94 -4773 -90 -4769
rect -70 -4773 -66 -4769
rect 166 -4773 170 -4769
rect 204 -4773 208 -4769
rect 264 -4773 268 -4769
rect 288 -4773 292 -4769
rect 522 -4773 526 -4769
rect 560 -4773 564 -4769
rect 620 -4773 624 -4769
rect 644 -4773 648 -4769
rect 880 -4773 884 -4769
rect 918 -4773 922 -4769
rect 978 -4773 982 -4769
rect 1002 -4773 1006 -4769
rect 1238 -4773 1242 -4769
rect 1276 -4773 1280 -4769
rect 1336 -4773 1340 -4769
rect 1360 -4773 1364 -4769
rect -1544 -4781 -1540 -4777
rect -1510 -4781 -1506 -4777
rect -1458 -4781 -1454 -4777
rect -1398 -4781 -1394 -4777
rect -1360 -4781 -1356 -4777
rect -1227 -4781 -1223 -4777
rect -1193 -4781 -1189 -4777
rect -1141 -4781 -1137 -4777
rect -1081 -4781 -1077 -4777
rect -1043 -4781 -1039 -4777
rect -928 -4781 -924 -4777
rect -894 -4781 -890 -4777
rect -842 -4781 -838 -4777
rect -782 -4781 -778 -4777
rect -744 -4781 -740 -4777
rect -570 -4781 -566 -4777
rect -536 -4781 -532 -4777
rect -484 -4781 -480 -4777
rect -424 -4781 -420 -4777
rect -386 -4781 -382 -4777
rect -212 -4781 -208 -4777
rect -178 -4781 -174 -4777
rect -126 -4781 -122 -4777
rect -66 -4781 -62 -4777
rect -28 -4781 -24 -4777
rect 146 -4781 150 -4777
rect 180 -4781 184 -4777
rect 232 -4781 236 -4777
rect 292 -4781 296 -4777
rect 330 -4781 334 -4777
rect 502 -4781 506 -4777
rect 536 -4781 540 -4777
rect 588 -4781 592 -4777
rect 648 -4781 652 -4777
rect 686 -4781 690 -4777
rect 860 -4781 864 -4777
rect 894 -4781 898 -4777
rect 946 -4781 950 -4777
rect 1006 -4781 1010 -4777
rect 1044 -4781 1048 -4777
rect 1218 -4781 1222 -4777
rect 1252 -4781 1256 -4777
rect 1304 -4781 1308 -4777
rect 1364 -4781 1368 -4777
rect 1402 -4781 1406 -4777
rect -1500 -4788 -1496 -4784
rect -1468 -4788 -1464 -4784
rect -1416 -4788 -1412 -4784
rect -1384 -4788 -1380 -4784
rect -1183 -4788 -1179 -4784
rect -1151 -4788 -1147 -4784
rect -1099 -4788 -1095 -4784
rect -1067 -4788 -1063 -4784
rect -884 -4788 -880 -4784
rect -852 -4788 -848 -4784
rect -800 -4788 -796 -4784
rect -768 -4788 -764 -4784
rect -526 -4788 -522 -4784
rect -494 -4788 -490 -4784
rect -442 -4788 -438 -4784
rect -410 -4788 -406 -4784
rect -168 -4788 -164 -4784
rect -136 -4788 -132 -4784
rect -84 -4788 -80 -4784
rect -52 -4788 -48 -4784
rect 190 -4788 194 -4784
rect 222 -4788 226 -4784
rect 274 -4788 278 -4784
rect 306 -4788 310 -4784
rect 546 -4788 550 -4784
rect 578 -4788 582 -4784
rect 630 -4788 634 -4784
rect 662 -4788 666 -4784
rect 904 -4788 908 -4784
rect 936 -4788 940 -4784
rect 988 -4788 992 -4784
rect 1020 -4788 1024 -4784
rect 1262 -4788 1266 -4784
rect 1294 -4788 1298 -4784
rect 1346 -4788 1350 -4784
rect 1378 -4788 1382 -4784
rect -1540 -4795 -1536 -4791
rect -1426 -4795 -1422 -4791
rect -1374 -4795 -1370 -4791
rect -1223 -4795 -1219 -4791
rect -1109 -4795 -1105 -4791
rect -1057 -4795 -1053 -4791
rect -924 -4795 -920 -4791
rect -810 -4795 -806 -4791
rect -758 -4795 -754 -4791
rect -566 -4795 -562 -4791
rect -452 -4795 -448 -4791
rect -400 -4795 -396 -4791
rect -208 -4795 -204 -4791
rect -94 -4795 -90 -4791
rect -42 -4795 -38 -4791
rect 150 -4795 154 -4791
rect 264 -4795 268 -4791
rect 316 -4795 320 -4791
rect 506 -4795 510 -4791
rect 620 -4795 624 -4791
rect 672 -4795 676 -4791
rect 864 -4795 868 -4791
rect 978 -4795 982 -4791
rect 1030 -4795 1034 -4791
rect 1222 -4795 1226 -4791
rect 1336 -4795 1340 -4791
rect 1388 -4795 1392 -4791
rect -1482 -4802 -1478 -4798
rect -1444 -4802 -1440 -4798
rect -1165 -4802 -1161 -4798
rect -1127 -4802 -1123 -4798
rect -866 -4802 -862 -4798
rect -828 -4802 -824 -4798
rect -508 -4802 -504 -4798
rect -470 -4802 -466 -4798
rect -150 -4802 -146 -4798
rect -112 -4802 -108 -4798
rect 208 -4802 212 -4798
rect 246 -4802 250 -4798
rect 564 -4802 568 -4798
rect 602 -4802 606 -4798
rect 922 -4802 926 -4798
rect 960 -4802 964 -4798
rect 1280 -4802 1284 -4798
rect 1318 -4802 1322 -4798
rect -1308 -4872 -1304 -4868
rect -934 -4872 -930 -4868
rect -576 -4872 -572 -4868
rect -218 -4872 -214 -4868
rect 140 -4872 144 -4868
rect 854 -4872 858 -4868
rect 1212 -4872 1216 -4868
rect -1297 -4880 -1293 -4876
rect -923 -4880 -919 -4876
rect -565 -4880 -561 -4876
rect -207 -4880 -203 -4876
rect 151 -4880 155 -4876
rect 507 -4880 511 -4876
rect 865 -4880 869 -4876
rect 1223 -4880 1227 -4876
rect -924 -5018 -920 -5014
rect -858 -5018 -854 -5014
rect -824 -5018 -820 -5014
rect -780 -5018 -776 -5014
rect -746 -5018 -742 -5014
rect -566 -5018 -562 -5014
rect -500 -5018 -496 -5014
rect -466 -5018 -462 -5014
rect -422 -5018 -418 -5014
rect -388 -5018 -384 -5014
rect -208 -5018 -204 -5014
rect -142 -5018 -138 -5014
rect -108 -5018 -104 -5014
rect -64 -5018 -60 -5014
rect -30 -5018 -26 -5014
rect 150 -5018 154 -5014
rect 216 -5018 220 -5014
rect 250 -5018 254 -5014
rect 294 -5018 298 -5014
rect 328 -5018 332 -5014
rect 506 -5018 510 -5014
rect 572 -5018 576 -5014
rect 606 -5018 610 -5014
rect 650 -5018 654 -5014
rect 684 -5018 688 -5014
rect 864 -5018 868 -5014
rect 930 -5018 934 -5014
rect 964 -5018 968 -5014
rect 1008 -5018 1012 -5014
rect 1042 -5018 1046 -5014
rect 1222 -5018 1226 -5014
rect 1288 -5018 1292 -5014
rect 1322 -5018 1326 -5014
rect 1366 -5018 1370 -5014
rect 1400 -5018 1404 -5014
rect -882 -5025 -878 -5021
rect -524 -5025 -520 -5021
rect -166 -5025 -162 -5021
rect 192 -5025 196 -5021
rect 548 -5025 552 -5021
rect 906 -5025 910 -5021
rect 1264 -5025 1268 -5021
rect -848 -5032 -844 -5028
rect -706 -5032 -702 -5028
rect -490 -5032 -486 -5028
rect -348 -5032 -344 -5028
rect -132 -5032 -128 -5028
rect 10 -5032 14 -5028
rect 226 -5032 230 -5028
rect 368 -5032 372 -5028
rect 582 -5032 586 -5028
rect 724 -5032 728 -5028
rect 940 -5032 944 -5028
rect 1082 -5032 1086 -5028
rect 1298 -5032 1302 -5028
rect 1440 -5032 1444 -5028
rect -928 -5039 -924 -5035
rect -898 -5039 -894 -5035
rect -780 -5039 -776 -5035
rect -570 -5039 -566 -5035
rect -540 -5039 -536 -5035
rect -422 -5039 -418 -5035
rect -212 -5039 -208 -5035
rect -182 -5039 -178 -5035
rect -64 -5039 -60 -5035
rect 146 -5039 150 -5035
rect 176 -5039 180 -5035
rect 294 -5039 298 -5035
rect 502 -5039 506 -5035
rect 532 -5039 536 -5035
rect 650 -5039 654 -5035
rect 860 -5039 864 -5035
rect 890 -5039 894 -5035
rect 1008 -5039 1012 -5035
rect 1218 -5039 1222 -5035
rect 1248 -5039 1252 -5035
rect 1366 -5039 1370 -5035
rect -1173 -5048 -1169 -5044
rect -902 -5047 -898 -5043
rect -804 -5047 -800 -5043
rect -544 -5047 -540 -5043
rect -446 -5047 -442 -5043
rect -186 -5047 -182 -5043
rect -88 -5047 -84 -5043
rect 172 -5047 176 -5043
rect 270 -5047 274 -5043
rect 528 -5047 532 -5043
rect 626 -5047 630 -5043
rect 886 -5047 890 -5043
rect 984 -5047 988 -5043
rect 1244 -5047 1248 -5043
rect 1342 -5047 1346 -5043
rect -1223 -5055 -1219 -5051
rect -1183 -5055 -1179 -5051
rect -1163 -5055 -1159 -5051
rect -924 -5054 -920 -5050
rect -776 -5054 -772 -5050
rect -566 -5054 -562 -5050
rect -418 -5054 -414 -5050
rect -208 -5054 -204 -5050
rect -60 -5054 -56 -5050
rect 150 -5054 154 -5050
rect 298 -5054 302 -5050
rect 506 -5054 510 -5050
rect 654 -5054 658 -5050
rect 864 -5054 868 -5050
rect 1012 -5054 1016 -5050
rect 1222 -5054 1226 -5050
rect 1370 -5054 1374 -5050
rect -1227 -5062 -1223 -5058
rect -1197 -5062 -1193 -5058
rect -1149 -5062 -1145 -5058
rect -902 -5061 -898 -5057
rect -794 -5061 -790 -5057
rect -760 -5061 -756 -5057
rect -544 -5061 -540 -5057
rect -436 -5061 -432 -5057
rect -402 -5061 -398 -5057
rect -186 -5061 -182 -5057
rect -78 -5061 -74 -5057
rect -44 -5061 -40 -5057
rect 172 -5061 176 -5057
rect 280 -5061 284 -5057
rect 314 -5061 318 -5057
rect 528 -5061 532 -5057
rect 636 -5061 640 -5057
rect 670 -5061 674 -5057
rect 886 -5061 890 -5057
rect 994 -5061 998 -5057
rect 1028 -5061 1032 -5057
rect 1244 -5061 1248 -5057
rect 1352 -5061 1356 -5057
rect 1386 -5061 1390 -5057
rect -928 -5068 -924 -5064
rect -872 -5068 -868 -5064
rect -838 -5068 -834 -5064
rect -570 -5068 -566 -5064
rect -514 -5068 -510 -5064
rect -480 -5068 -476 -5064
rect -212 -5068 -208 -5064
rect -156 -5068 -152 -5064
rect -122 -5068 -118 -5064
rect 146 -5068 150 -5064
rect 202 -5068 206 -5064
rect 236 -5068 240 -5064
rect 502 -5068 506 -5064
rect 558 -5068 562 -5064
rect 592 -5068 596 -5064
rect 860 -5068 864 -5064
rect 916 -5068 920 -5064
rect 950 -5068 954 -5064
rect 1218 -5068 1222 -5064
rect 1274 -5068 1278 -5064
rect 1308 -5068 1312 -5064
rect -1783 -5166 -1779 -5162
rect -1745 -5166 -1741 -5162
rect -1685 -5166 -1681 -5162
rect -1661 -5166 -1657 -5162
rect -1520 -5166 -1516 -5162
rect -1482 -5166 -1478 -5162
rect -1422 -5166 -1418 -5162
rect -1398 -5166 -1394 -5162
rect -1207 -5166 -1203 -5162
rect -1169 -5166 -1165 -5162
rect -1109 -5166 -1105 -5162
rect -1085 -5166 -1081 -5162
rect -908 -5166 -904 -5162
rect -870 -5166 -866 -5162
rect -810 -5166 -806 -5162
rect -786 -5166 -782 -5162
rect -1803 -5174 -1799 -5170
rect -1769 -5174 -1765 -5170
rect -1717 -5174 -1713 -5170
rect -1657 -5174 -1653 -5170
rect -1619 -5174 -1615 -5170
rect -1540 -5174 -1536 -5170
rect -1506 -5174 -1502 -5170
rect -1454 -5174 -1450 -5170
rect -1394 -5174 -1390 -5170
rect -1356 -5174 -1352 -5170
rect -1227 -5174 -1223 -5170
rect -1193 -5174 -1189 -5170
rect -1141 -5174 -1137 -5170
rect -1081 -5174 -1077 -5170
rect -1043 -5174 -1039 -5170
rect -928 -5174 -924 -5170
rect -894 -5174 -890 -5170
rect -842 -5174 -838 -5170
rect -782 -5174 -778 -5170
rect -744 -5174 -740 -5170
rect -1759 -5181 -1755 -5177
rect -1727 -5181 -1723 -5177
rect -1675 -5181 -1671 -5177
rect -1643 -5181 -1639 -5177
rect -1496 -5181 -1492 -5177
rect -1464 -5181 -1460 -5177
rect -1412 -5181 -1408 -5177
rect -1380 -5181 -1376 -5177
rect -1183 -5181 -1179 -5177
rect -1151 -5181 -1147 -5177
rect -1099 -5181 -1095 -5177
rect -1067 -5181 -1063 -5177
rect -884 -5181 -880 -5177
rect -852 -5181 -848 -5177
rect -800 -5181 -796 -5177
rect -768 -5181 -764 -5177
rect -1799 -5188 -1795 -5184
rect -1685 -5188 -1681 -5184
rect -1633 -5188 -1629 -5184
rect -1536 -5188 -1532 -5184
rect -1422 -5188 -1418 -5184
rect -1370 -5188 -1366 -5184
rect -1223 -5188 -1219 -5184
rect -1109 -5188 -1105 -5184
rect -1057 -5188 -1053 -5184
rect -924 -5188 -920 -5184
rect -810 -5188 -806 -5184
rect -758 -5188 -754 -5184
rect -1741 -5195 -1737 -5191
rect -1703 -5195 -1699 -5191
rect -1478 -5195 -1474 -5191
rect -1440 -5195 -1436 -5191
rect -1165 -5195 -1161 -5191
rect -1127 -5195 -1123 -5191
rect -866 -5195 -862 -5191
rect -828 -5195 -824 -5191
rect -1783 -5337 -1779 -5333
rect -1745 -5337 -1741 -5333
rect -1685 -5337 -1681 -5333
rect -1661 -5337 -1657 -5333
rect -1520 -5337 -1516 -5333
rect -1482 -5337 -1478 -5333
rect -1422 -5337 -1418 -5333
rect -1398 -5337 -1394 -5333
rect -1207 -5337 -1203 -5333
rect -1169 -5337 -1165 -5333
rect -1109 -5337 -1105 -5333
rect -1085 -5337 -1081 -5333
rect -908 -5337 -904 -5333
rect -870 -5337 -866 -5333
rect -810 -5337 -806 -5333
rect -786 -5337 -782 -5333
rect -550 -5337 -546 -5333
rect -512 -5337 -508 -5333
rect -452 -5337 -448 -5333
rect -428 -5337 -424 -5333
rect -192 -5337 -188 -5333
rect -154 -5337 -150 -5333
rect -94 -5337 -90 -5333
rect -70 -5337 -66 -5333
rect 166 -5337 170 -5333
rect 204 -5337 208 -5333
rect 264 -5337 268 -5333
rect 288 -5337 292 -5333
rect 522 -5337 526 -5333
rect 560 -5337 564 -5333
rect 620 -5337 624 -5333
rect 644 -5337 648 -5333
rect 880 -5337 884 -5333
rect 918 -5337 922 -5333
rect 978 -5337 982 -5333
rect 1002 -5337 1006 -5333
rect 1238 -5337 1242 -5333
rect 1276 -5337 1280 -5333
rect 1336 -5337 1340 -5333
rect 1360 -5337 1364 -5333
rect -1803 -5345 -1799 -5341
rect -1769 -5345 -1765 -5341
rect -1717 -5345 -1713 -5341
rect -1657 -5345 -1653 -5341
rect -1619 -5345 -1615 -5341
rect -1540 -5345 -1536 -5341
rect -1506 -5345 -1502 -5341
rect -1454 -5345 -1450 -5341
rect -1394 -5345 -1390 -5341
rect -1356 -5345 -1352 -5341
rect -1227 -5345 -1223 -5341
rect -1193 -5345 -1189 -5341
rect -1141 -5345 -1137 -5341
rect -1081 -5345 -1077 -5341
rect -1043 -5345 -1039 -5341
rect -928 -5345 -924 -5341
rect -894 -5345 -890 -5341
rect -842 -5345 -838 -5341
rect -782 -5345 -778 -5341
rect -744 -5345 -740 -5341
rect -570 -5345 -566 -5341
rect -536 -5345 -532 -5341
rect -484 -5345 -480 -5341
rect -424 -5345 -420 -5341
rect -386 -5345 -382 -5341
rect -212 -5345 -208 -5341
rect -178 -5345 -174 -5341
rect -126 -5345 -122 -5341
rect -66 -5345 -62 -5341
rect -28 -5345 -24 -5341
rect 146 -5345 150 -5341
rect 180 -5345 184 -5341
rect 232 -5345 236 -5341
rect 292 -5345 296 -5341
rect 330 -5345 334 -5341
rect 502 -5345 506 -5341
rect 536 -5345 540 -5341
rect 588 -5345 592 -5341
rect 648 -5345 652 -5341
rect 686 -5345 690 -5341
rect 860 -5345 864 -5341
rect 894 -5345 898 -5341
rect 946 -5345 950 -5341
rect 1006 -5345 1010 -5341
rect 1044 -5345 1048 -5341
rect 1218 -5345 1222 -5341
rect 1252 -5345 1256 -5341
rect 1304 -5345 1308 -5341
rect 1364 -5345 1368 -5341
rect 1402 -5345 1406 -5341
rect -1759 -5352 -1755 -5348
rect -1727 -5352 -1723 -5348
rect -1675 -5352 -1671 -5348
rect -1643 -5352 -1639 -5348
rect -1496 -5352 -1492 -5348
rect -1464 -5352 -1460 -5348
rect -1412 -5352 -1408 -5348
rect -1380 -5352 -1376 -5348
rect -1183 -5352 -1179 -5348
rect -1151 -5352 -1147 -5348
rect -1099 -5352 -1095 -5348
rect -1067 -5352 -1063 -5348
rect -884 -5352 -880 -5348
rect -852 -5352 -848 -5348
rect -800 -5352 -796 -5348
rect -768 -5352 -764 -5348
rect -526 -5352 -522 -5348
rect -494 -5352 -490 -5348
rect -442 -5352 -438 -5348
rect -410 -5352 -406 -5348
rect -168 -5352 -164 -5348
rect -136 -5352 -132 -5348
rect -84 -5352 -80 -5348
rect -52 -5352 -48 -5348
rect 190 -5352 194 -5348
rect 222 -5352 226 -5348
rect 274 -5352 278 -5348
rect 306 -5352 310 -5348
rect 546 -5352 550 -5348
rect 578 -5352 582 -5348
rect 630 -5352 634 -5348
rect 662 -5352 666 -5348
rect 904 -5352 908 -5348
rect 936 -5352 940 -5348
rect 988 -5352 992 -5348
rect 1020 -5352 1024 -5348
rect 1262 -5352 1266 -5348
rect 1294 -5352 1298 -5348
rect 1346 -5352 1350 -5348
rect 1378 -5352 1382 -5348
rect -1799 -5359 -1795 -5355
rect -1685 -5359 -1681 -5355
rect -1633 -5359 -1629 -5355
rect -1536 -5359 -1532 -5355
rect -1422 -5359 -1418 -5355
rect -1370 -5359 -1366 -5355
rect -1223 -5359 -1219 -5355
rect -1109 -5359 -1105 -5355
rect -1057 -5359 -1053 -5355
rect -924 -5359 -920 -5355
rect -810 -5359 -806 -5355
rect -758 -5359 -754 -5355
rect -566 -5359 -562 -5355
rect -452 -5359 -448 -5355
rect -400 -5359 -396 -5355
rect -208 -5359 -204 -5355
rect -94 -5359 -90 -5355
rect -42 -5359 -38 -5355
rect 150 -5359 154 -5355
rect 264 -5359 268 -5355
rect 316 -5359 320 -5355
rect 506 -5359 510 -5355
rect 620 -5359 624 -5355
rect 672 -5359 676 -5355
rect 864 -5359 868 -5355
rect 978 -5359 982 -5355
rect 1030 -5359 1034 -5355
rect 1222 -5359 1226 -5355
rect 1336 -5359 1340 -5355
rect 1388 -5359 1392 -5355
rect -1741 -5366 -1737 -5362
rect -1703 -5366 -1699 -5362
rect -1478 -5366 -1474 -5362
rect -1440 -5366 -1436 -5362
rect -1165 -5366 -1161 -5362
rect -1127 -5366 -1123 -5362
rect -866 -5366 -862 -5362
rect -828 -5366 -824 -5362
rect -508 -5366 -504 -5362
rect -470 -5366 -466 -5362
rect -150 -5366 -146 -5362
rect -112 -5366 -108 -5362
rect 208 -5366 212 -5362
rect 246 -5366 250 -5362
rect 564 -5366 568 -5362
rect 602 -5366 606 -5362
rect 922 -5366 926 -5362
rect 960 -5366 964 -5362
rect 1280 -5366 1284 -5362
rect 1318 -5366 1322 -5362
rect -1783 -5497 -1779 -5493
rect -1745 -5497 -1741 -5493
rect -1685 -5497 -1681 -5493
rect -1661 -5497 -1657 -5493
rect -1520 -5497 -1516 -5493
rect -1482 -5497 -1478 -5493
rect -1422 -5497 -1418 -5493
rect -1398 -5497 -1394 -5493
rect -1207 -5497 -1203 -5493
rect -1169 -5497 -1165 -5493
rect -1109 -5497 -1105 -5493
rect -1085 -5497 -1081 -5493
rect -908 -5497 -904 -5493
rect -870 -5497 -866 -5493
rect -810 -5497 -806 -5493
rect -786 -5497 -782 -5493
rect -550 -5497 -546 -5493
rect -512 -5497 -508 -5493
rect -452 -5497 -448 -5493
rect -428 -5497 -424 -5493
rect -192 -5497 -188 -5493
rect -154 -5497 -150 -5493
rect -94 -5497 -90 -5493
rect -70 -5497 -66 -5493
rect 166 -5497 170 -5493
rect 204 -5497 208 -5493
rect 264 -5497 268 -5493
rect 288 -5497 292 -5493
rect 522 -5497 526 -5493
rect 560 -5497 564 -5493
rect 620 -5497 624 -5493
rect 644 -5497 648 -5493
rect 880 -5497 884 -5493
rect 918 -5497 922 -5493
rect 978 -5497 982 -5493
rect 1002 -5497 1006 -5493
rect 1238 -5497 1242 -5493
rect 1276 -5497 1280 -5493
rect 1336 -5497 1340 -5493
rect 1360 -5497 1364 -5493
rect -1803 -5505 -1799 -5501
rect -1769 -5505 -1765 -5501
rect -1717 -5505 -1713 -5501
rect -1657 -5505 -1653 -5501
rect -1619 -5505 -1615 -5501
rect -1540 -5505 -1536 -5501
rect -1506 -5505 -1502 -5501
rect -1454 -5505 -1450 -5501
rect -1394 -5505 -1390 -5501
rect -1356 -5505 -1352 -5501
rect -1227 -5505 -1223 -5501
rect -1193 -5505 -1189 -5501
rect -1141 -5505 -1137 -5501
rect -1081 -5505 -1077 -5501
rect -1043 -5505 -1039 -5501
rect -928 -5505 -924 -5501
rect -894 -5505 -890 -5501
rect -842 -5505 -838 -5501
rect -782 -5505 -778 -5501
rect -744 -5505 -740 -5501
rect -570 -5505 -566 -5501
rect -536 -5505 -532 -5501
rect -484 -5505 -480 -5501
rect -424 -5505 -420 -5501
rect -386 -5505 -382 -5501
rect -212 -5505 -208 -5501
rect -178 -5505 -174 -5501
rect -126 -5505 -122 -5501
rect -66 -5505 -62 -5501
rect -28 -5505 -24 -5501
rect 146 -5505 150 -5501
rect 180 -5505 184 -5501
rect 232 -5505 236 -5501
rect 292 -5505 296 -5501
rect 330 -5505 334 -5501
rect 502 -5505 506 -5501
rect 536 -5505 540 -5501
rect 588 -5505 592 -5501
rect 648 -5505 652 -5501
rect 686 -5505 690 -5501
rect 860 -5505 864 -5501
rect 894 -5505 898 -5501
rect 946 -5505 950 -5501
rect 1006 -5505 1010 -5501
rect 1044 -5505 1048 -5501
rect 1218 -5505 1222 -5501
rect 1252 -5505 1256 -5501
rect 1304 -5505 1308 -5501
rect 1364 -5505 1368 -5501
rect 1402 -5505 1406 -5501
rect -1759 -5512 -1755 -5508
rect -1727 -5512 -1723 -5508
rect -1675 -5512 -1671 -5508
rect -1643 -5512 -1639 -5508
rect -1496 -5512 -1492 -5508
rect -1464 -5512 -1460 -5508
rect -1412 -5512 -1408 -5508
rect -1380 -5512 -1376 -5508
rect -1183 -5512 -1179 -5508
rect -1151 -5512 -1147 -5508
rect -1099 -5512 -1095 -5508
rect -1067 -5512 -1063 -5508
rect -884 -5512 -880 -5508
rect -852 -5512 -848 -5508
rect -800 -5512 -796 -5508
rect -768 -5512 -764 -5508
rect -526 -5512 -522 -5508
rect -494 -5512 -490 -5508
rect -442 -5512 -438 -5508
rect -410 -5512 -406 -5508
rect -168 -5512 -164 -5508
rect -136 -5512 -132 -5508
rect -84 -5512 -80 -5508
rect -52 -5512 -48 -5508
rect 190 -5512 194 -5508
rect 222 -5512 226 -5508
rect 274 -5512 278 -5508
rect 306 -5512 310 -5508
rect 546 -5512 550 -5508
rect 578 -5512 582 -5508
rect 630 -5512 634 -5508
rect 662 -5512 666 -5508
rect 904 -5512 908 -5508
rect 936 -5512 940 -5508
rect 988 -5512 992 -5508
rect 1020 -5512 1024 -5508
rect 1262 -5512 1266 -5508
rect 1294 -5512 1298 -5508
rect 1346 -5512 1350 -5508
rect 1378 -5512 1382 -5508
rect -1799 -5519 -1795 -5515
rect -1685 -5519 -1681 -5515
rect -1633 -5519 -1629 -5515
rect -1536 -5519 -1532 -5515
rect -1422 -5519 -1418 -5515
rect -1370 -5519 -1366 -5515
rect -1223 -5519 -1219 -5515
rect -1109 -5519 -1105 -5515
rect -1057 -5519 -1053 -5515
rect -924 -5519 -920 -5515
rect -810 -5519 -806 -5515
rect -758 -5519 -754 -5515
rect -566 -5519 -562 -5515
rect -452 -5519 -448 -5515
rect -400 -5519 -396 -5515
rect -208 -5519 -204 -5515
rect -94 -5519 -90 -5515
rect -42 -5519 -38 -5515
rect 150 -5519 154 -5515
rect 264 -5519 268 -5515
rect 316 -5519 320 -5515
rect 506 -5519 510 -5515
rect 620 -5519 624 -5515
rect 672 -5519 676 -5515
rect 864 -5519 868 -5515
rect 978 -5519 982 -5515
rect 1030 -5519 1034 -5515
rect 1222 -5519 1226 -5515
rect 1336 -5519 1340 -5515
rect 1388 -5519 1392 -5515
rect -1741 -5526 -1737 -5522
rect -1703 -5526 -1699 -5522
rect -1478 -5526 -1474 -5522
rect -1440 -5526 -1436 -5522
rect -1165 -5526 -1161 -5522
rect -1127 -5526 -1123 -5522
rect -866 -5526 -862 -5522
rect -828 -5526 -824 -5522
rect -508 -5526 -504 -5522
rect -470 -5526 -466 -5522
rect -150 -5526 -146 -5522
rect -112 -5526 -108 -5522
rect 208 -5526 212 -5522
rect 246 -5526 250 -5522
rect 564 -5526 568 -5522
rect 602 -5526 606 -5522
rect 922 -5526 926 -5522
rect 960 -5526 964 -5522
rect 1280 -5526 1284 -5522
rect 1318 -5526 1322 -5522
rect -1308 -5595 -1304 -5591
rect -934 -5595 -930 -5591
rect -576 -5595 -572 -5591
rect -218 -5595 -214 -5591
rect 140 -5595 144 -5591
rect 496 -5595 500 -5591
rect 854 -5595 858 -5591
rect 1212 -5595 1216 -5591
rect -1297 -5603 -1293 -5599
rect -923 -5603 -919 -5599
rect -565 -5603 -561 -5599
rect -207 -5603 -203 -5599
rect 151 -5603 155 -5599
rect 507 -5603 511 -5599
rect 865 -5603 869 -5599
rect 1223 -5603 1227 -5599
rect -924 -5741 -920 -5737
rect -858 -5741 -854 -5737
rect -824 -5741 -820 -5737
rect -780 -5741 -776 -5737
rect -746 -5741 -742 -5737
rect -566 -5741 -562 -5737
rect -500 -5741 -496 -5737
rect -466 -5741 -462 -5737
rect -422 -5741 -418 -5737
rect -388 -5741 -384 -5737
rect -208 -5741 -204 -5737
rect -142 -5741 -138 -5737
rect -108 -5741 -104 -5737
rect -64 -5741 -60 -5737
rect -30 -5741 -26 -5737
rect 150 -5741 154 -5737
rect 216 -5741 220 -5737
rect 250 -5741 254 -5737
rect 294 -5741 298 -5737
rect 328 -5741 332 -5737
rect 506 -5741 510 -5737
rect 572 -5741 576 -5737
rect 606 -5741 610 -5737
rect 650 -5741 654 -5737
rect 684 -5741 688 -5737
rect 864 -5741 868 -5737
rect 930 -5741 934 -5737
rect 964 -5741 968 -5737
rect 1008 -5741 1012 -5737
rect 1042 -5741 1046 -5737
rect 1222 -5741 1226 -5737
rect 1288 -5741 1292 -5737
rect 1322 -5741 1326 -5737
rect 1366 -5741 1370 -5737
rect 1400 -5741 1404 -5737
rect -882 -5748 -878 -5744
rect -524 -5748 -520 -5744
rect -166 -5748 -162 -5744
rect 192 -5748 196 -5744
rect 548 -5748 552 -5744
rect 906 -5748 910 -5744
rect 1264 -5748 1268 -5744
rect -848 -5755 -844 -5751
rect -706 -5755 -702 -5751
rect -490 -5755 -486 -5751
rect -348 -5755 -344 -5751
rect -132 -5755 -128 -5751
rect 10 -5755 14 -5751
rect 226 -5755 230 -5751
rect 368 -5755 372 -5751
rect 582 -5755 586 -5751
rect 724 -5755 728 -5751
rect 940 -5755 944 -5751
rect 1082 -5755 1086 -5751
rect 1298 -5755 1302 -5751
rect 1440 -5755 1444 -5751
rect -928 -5762 -924 -5758
rect -898 -5762 -894 -5758
rect -780 -5762 -776 -5758
rect -570 -5762 -566 -5758
rect -540 -5762 -536 -5758
rect -422 -5762 -418 -5758
rect -212 -5762 -208 -5758
rect -182 -5762 -178 -5758
rect -64 -5762 -60 -5758
rect 146 -5762 150 -5758
rect 176 -5762 180 -5758
rect 294 -5762 298 -5758
rect 502 -5762 506 -5758
rect 532 -5762 536 -5758
rect 650 -5762 654 -5758
rect 860 -5762 864 -5758
rect 890 -5762 894 -5758
rect 1008 -5762 1012 -5758
rect 1218 -5762 1222 -5758
rect 1248 -5762 1252 -5758
rect 1366 -5762 1370 -5758
rect -1173 -5771 -1169 -5767
rect -902 -5770 -898 -5766
rect -804 -5770 -800 -5766
rect -544 -5770 -540 -5766
rect -446 -5770 -442 -5766
rect -186 -5770 -182 -5766
rect -88 -5770 -84 -5766
rect 172 -5770 176 -5766
rect 270 -5770 274 -5766
rect 528 -5770 532 -5766
rect 626 -5770 630 -5766
rect 886 -5770 890 -5766
rect 984 -5770 988 -5766
rect 1244 -5770 1248 -5766
rect 1342 -5770 1346 -5766
rect -1223 -5778 -1219 -5774
rect -1183 -5778 -1179 -5774
rect -1163 -5778 -1159 -5774
rect -924 -5777 -920 -5773
rect -776 -5777 -772 -5773
rect -566 -5777 -562 -5773
rect -418 -5777 -414 -5773
rect -208 -5777 -204 -5773
rect -60 -5777 -56 -5773
rect 150 -5777 154 -5773
rect 298 -5777 302 -5773
rect 506 -5777 510 -5773
rect 654 -5777 658 -5773
rect 864 -5777 868 -5773
rect 1012 -5777 1016 -5773
rect 1222 -5777 1226 -5773
rect 1370 -5777 1374 -5773
rect -1227 -5785 -1223 -5781
rect -1197 -5785 -1193 -5781
rect -1149 -5785 -1145 -5781
rect -902 -5784 -898 -5780
rect -794 -5784 -790 -5780
rect -760 -5784 -756 -5780
rect -544 -5784 -540 -5780
rect -436 -5784 -432 -5780
rect -402 -5784 -398 -5780
rect -186 -5784 -182 -5780
rect -78 -5784 -74 -5780
rect -44 -5784 -40 -5780
rect 172 -5784 176 -5780
rect 280 -5784 284 -5780
rect 314 -5784 318 -5780
rect 528 -5784 532 -5780
rect 636 -5784 640 -5780
rect 670 -5784 674 -5780
rect 886 -5784 890 -5780
rect 994 -5784 998 -5780
rect 1028 -5784 1032 -5780
rect 1244 -5784 1248 -5780
rect 1352 -5784 1356 -5780
rect 1386 -5784 1390 -5780
rect -928 -5791 -924 -5787
rect -872 -5791 -868 -5787
rect -838 -5791 -834 -5787
rect -570 -5791 -566 -5787
rect -514 -5791 -510 -5787
rect -480 -5791 -476 -5787
rect -212 -5791 -208 -5787
rect -156 -5791 -152 -5787
rect -122 -5791 -118 -5787
rect 146 -5791 150 -5787
rect 202 -5791 206 -5787
rect 236 -5791 240 -5787
rect 502 -5791 506 -5787
rect 558 -5791 562 -5787
rect 592 -5791 596 -5787
rect 860 -5791 864 -5787
rect 916 -5791 920 -5787
rect 950 -5791 954 -5787
rect 1218 -5791 1222 -5787
rect 1274 -5791 1278 -5787
rect 1308 -5791 1312 -5787
rect -1207 -5893 -1203 -5889
rect -1169 -5893 -1165 -5889
rect -1109 -5893 -1105 -5889
rect -1085 -5893 -1081 -5889
rect -908 -5893 -904 -5889
rect -870 -5893 -866 -5889
rect -810 -5893 -806 -5889
rect -786 -5893 -782 -5889
rect -550 -5893 -546 -5889
rect -512 -5893 -508 -5889
rect -452 -5893 -448 -5889
rect -428 -5893 -424 -5889
rect -192 -5893 -188 -5889
rect -154 -5893 -150 -5889
rect -94 -5893 -90 -5889
rect -70 -5893 -66 -5889
rect 166 -5893 170 -5889
rect 204 -5893 208 -5889
rect 264 -5893 268 -5889
rect 288 -5893 292 -5889
rect 522 -5893 526 -5889
rect 560 -5893 564 -5889
rect 620 -5893 624 -5889
rect 644 -5893 648 -5889
rect 880 -5893 884 -5889
rect 918 -5893 922 -5889
rect 978 -5893 982 -5889
rect 1002 -5893 1006 -5889
rect 1238 -5893 1242 -5889
rect 1276 -5893 1280 -5889
rect 1336 -5893 1340 -5889
rect 1360 -5893 1364 -5889
rect 1582 -5893 1586 -5889
rect 1620 -5893 1624 -5889
rect 1680 -5893 1684 -5889
rect 1704 -5893 1708 -5889
rect -1227 -5901 -1223 -5897
rect -1193 -5901 -1189 -5897
rect -1141 -5901 -1137 -5897
rect -1081 -5901 -1077 -5897
rect -1043 -5901 -1039 -5897
rect -928 -5901 -924 -5897
rect -894 -5901 -890 -5897
rect -842 -5901 -838 -5897
rect -782 -5901 -778 -5897
rect -744 -5901 -740 -5897
rect -570 -5901 -566 -5897
rect -536 -5901 -532 -5897
rect -484 -5901 -480 -5897
rect -424 -5901 -420 -5897
rect -386 -5901 -382 -5897
rect -212 -5901 -208 -5897
rect -178 -5901 -174 -5897
rect -126 -5901 -122 -5897
rect -66 -5901 -62 -5897
rect -28 -5901 -24 -5897
rect 146 -5901 150 -5897
rect 180 -5901 184 -5897
rect 232 -5901 236 -5897
rect 292 -5901 296 -5897
rect 330 -5901 334 -5897
rect 502 -5901 506 -5897
rect 536 -5901 540 -5897
rect 588 -5901 592 -5897
rect 648 -5901 652 -5897
rect 686 -5901 690 -5897
rect 860 -5901 864 -5897
rect 894 -5901 898 -5897
rect 946 -5901 950 -5897
rect 1006 -5901 1010 -5897
rect 1044 -5901 1048 -5897
rect 1218 -5901 1222 -5897
rect 1252 -5901 1256 -5897
rect 1304 -5901 1308 -5897
rect 1364 -5901 1368 -5897
rect 1402 -5901 1406 -5897
rect 1562 -5901 1566 -5897
rect 1596 -5901 1600 -5897
rect 1648 -5901 1652 -5897
rect 1708 -5901 1712 -5897
rect 1746 -5901 1750 -5897
rect -1183 -5908 -1179 -5904
rect -1151 -5908 -1147 -5904
rect -1099 -5908 -1095 -5904
rect -1067 -5908 -1063 -5904
rect -884 -5908 -880 -5904
rect -852 -5908 -848 -5904
rect -800 -5908 -796 -5904
rect -768 -5908 -764 -5904
rect -526 -5908 -522 -5904
rect -494 -5908 -490 -5904
rect -442 -5908 -438 -5904
rect -410 -5908 -406 -5904
rect -168 -5908 -164 -5904
rect -136 -5908 -132 -5904
rect -84 -5908 -80 -5904
rect -52 -5908 -48 -5904
rect 190 -5908 194 -5904
rect 222 -5908 226 -5904
rect 274 -5908 278 -5904
rect 306 -5908 310 -5904
rect 546 -5908 550 -5904
rect 578 -5908 582 -5904
rect 630 -5908 634 -5904
rect 662 -5908 666 -5904
rect 904 -5908 908 -5904
rect 936 -5908 940 -5904
rect 988 -5908 992 -5904
rect 1020 -5908 1024 -5904
rect 1262 -5908 1266 -5904
rect 1294 -5908 1298 -5904
rect 1346 -5908 1350 -5904
rect 1378 -5908 1382 -5904
rect 1606 -5908 1610 -5904
rect 1638 -5908 1642 -5904
rect 1690 -5908 1694 -5904
rect 1722 -5908 1726 -5904
rect -1223 -5915 -1219 -5911
rect -1109 -5915 -1105 -5911
rect -1057 -5915 -1053 -5911
rect -924 -5915 -920 -5911
rect -810 -5915 -806 -5911
rect -758 -5915 -754 -5911
rect -566 -5915 -562 -5911
rect -452 -5915 -448 -5911
rect -400 -5915 -396 -5911
rect -208 -5915 -204 -5911
rect -94 -5915 -90 -5911
rect -42 -5915 -38 -5911
rect 150 -5915 154 -5911
rect 264 -5915 268 -5911
rect 316 -5915 320 -5911
rect 506 -5915 510 -5911
rect 620 -5915 624 -5911
rect 672 -5915 676 -5911
rect 864 -5915 868 -5911
rect 978 -5915 982 -5911
rect 1030 -5915 1034 -5911
rect 1222 -5915 1226 -5911
rect 1336 -5915 1340 -5911
rect 1388 -5915 1392 -5911
rect 1566 -5915 1570 -5911
rect 1680 -5915 1684 -5911
rect 1732 -5915 1736 -5911
rect -1165 -5922 -1161 -5918
rect -1127 -5922 -1123 -5918
rect -866 -5922 -862 -5918
rect -828 -5922 -824 -5918
rect -508 -5922 -504 -5918
rect -470 -5922 -466 -5918
rect -150 -5922 -146 -5918
rect -112 -5922 -108 -5918
rect 208 -5922 212 -5918
rect 246 -5922 250 -5918
rect 564 -5922 568 -5918
rect 602 -5922 606 -5918
rect 922 -5922 926 -5918
rect 960 -5922 964 -5918
rect 1280 -5922 1284 -5918
rect 1318 -5922 1322 -5918
rect 1624 -5922 1628 -5918
rect 1662 -5922 1666 -5918
<< labels >>
rlabel metal2 -1411 -1174 -1411 -1170 1 Y1
rlabel metal1 -1319 -748 -1315 -748 5 X0
rlabel metal2 -1411 -824 -1411 -820 1 Y0
rlabel metal1 -949 -748 -945 -748 5 X1
rlabel metal1 -591 -749 -587 -749 5 X2
rlabel metal1 -233 -748 -229 -748 5 X3
rlabel metal1 481 -748 485 -748 5 X5
rlabel metal1 839 -748 843 -748 5 X6
rlabel metal1 1197 -748 1201 -748 5 X7
rlabel metal1 125 -748 129 -748 5 X4
rlabel metal2 -2041 -3508 -2041 -3508 1 VDD!
rlabel metal2 1053 -1469 1053 -1465 1 Z1
rlabel metal2 -1234 -1088 -1234 -1084 1 CLK!
rlabel metal2 -939 -1088 -939 -1084 1 CLK!
rlabel metal2 -581 -1088 -581 -1084 1 CLK!
rlabel metal2 -223 -1088 -223 -1084 1 CLK!
rlabel metal2 135 -1088 135 -1084 1 CLK!
rlabel metal2 491 -1088 491 -1084 1 CLK!
rlabel metal2 849 -1088 849 -1084 1 CLK!
rlabel metal2 1053 -1066 1053 -1062 1 Z0
rlabel metal2 -1234 -1491 -1234 -1487 1 CLK!
rlabel metal2 -939 -1491 -939 -1487 1 CLK!
rlabel metal2 -581 -1491 -581 -1487 1 CLK!
rlabel metal2 -223 -1491 -223 -1487 1 CLK!
rlabel metal2 135 -1491 135 -1487 1 CLK!
rlabel metal2 491 -1491 491 -1487 1 CLK!
rlabel metal2 849 -1491 849 -1487 1 CLK!
rlabel metal2 1207 -1662 1207 -1658 1 CLK!
rlabel metal2 1207 -1833 1207 -1829 1 CLK!
rlabel metal2 849 -1662 849 -1658 1 CLK!
rlabel metal2 849 -1833 849 -1829 1 CLK!
rlabel metal2 491 -1833 491 -1829 1 CLK!
rlabel metal2 491 -1662 491 -1658 1 CLK!
rlabel metal2 135 -1662 135 -1658 1 CLK!
rlabel metal2 135 -1833 135 -1829 1 CLK!
rlabel metal2 -223 -1662 -223 -1658 1 CLK!
rlabel metal2 -223 -1833 -223 -1829 1 CLK!
rlabel metal2 -581 -1662 -581 -1658 1 CLK!
rlabel metal2 -581 -1833 -581 -1829 1 CLK!
rlabel metal2 -939 -1833 -939 -1829 1 CLK!
rlabel metal2 -939 -1662 -939 -1658 1 CLK!
rlabel metal2 -1234 -1662 -1234 -1658 1 CLK!
rlabel metal2 -1234 -1833 -1234 -1829 1 CLK!
rlabel metal2 -1563 -1833 -1563 -1829 1 CLK!
rlabel metal2 -1563 -2414 -1563 -2410 1 CLK!
rlabel metal2 -1563 -2585 -1563 -2581 1 CLK!
rlabel metal2 -1238 -2414 -1238 -2410 1 CLK!
rlabel metal2 -1238 -2585 -1238 -2581 1 CLK!
rlabel metal2 -939 -2585 -939 -2581 1 CLK!
rlabel metal2 -939 -2414 -939 -2410 1 CLK!
rlabel metal2 -581 -2414 -581 -2410 1 CLK!
rlabel metal2 -1238 -2243 -1238 -2239 1 CLK!
rlabel metal2 -939 -2243 -939 -2239 1 CLK!
rlabel metal2 -581 -2243 -581 -2239 1 CLK!
rlabel metal2 -223 -2243 -223 -2239 1 CLK!
rlabel metal2 135 -2243 135 -2239 1 CLK!
rlabel metal2 491 -2243 491 -2239 1 CLK!
rlabel metal2 1207 -2414 1207 -2410 1 CLK!
rlabel metal2 849 -2414 849 -2410 1 CLK!
rlabel metal2 491 -2414 491 -2410 1 CLK!
rlabel metal2 135 -2414 135 -2410 1 CLK!
rlabel metal2 -223 -2414 -223 -2410 1 CLK!
rlabel metal2 -581 -2585 -581 -2581 1 CLK!
rlabel metal2 -224 -2585 -224 -2581 1 CLK!
rlabel metal2 135 -2585 135 -2581 1 CLK!
rlabel metal2 491 -2585 491 -2581 1 CLK!
rlabel metal2 849 -2585 849 -2581 1 CLK!
rlabel metal2 1207 -2585 1207 -2581 1 CLK!
rlabel metal2 1207 -3310 1207 -3306 1 CLK!
rlabel metal2 849 -3310 849 -3306 1 CLK!
rlabel metal2 491 -3310 491 -3306 1 CLK!
rlabel metal2 135 -3310 135 -3306 1 CLK!
rlabel metal2 -223 -3310 -223 -3306 1 CLK!
rlabel metal2 -581 -3310 -581 -3306 1 CLK!
rlabel metal2 -939 -3310 -939 -3306 1 CLK!
rlabel metal2 -1238 -3310 -1238 -3306 1 CLK!
rlabel metal2 -1563 -3310 -1563 -3306 1 CLK!
rlabel metal2 -1563 -3139 -1563 -3135 1 CLK!
rlabel metal2 -1238 -3139 -1238 -3135 1 CLK!
rlabel metal2 -939 -3139 -939 -3135 1 CLK!
rlabel metal2 -581 -3139 -581 -3135 1 CLK!
rlabel metal2 -223 -3139 -223 -3135 1 CLK!
rlabel metal2 135 -3139 135 -3135 1 CLK!
rlabel metal2 491 -3139 491 -3135 1 CLK!
rlabel metal2 849 -3139 849 -3135 1 CLK!
rlabel metal2 1207 -3139 1207 -3135 1 CLK!
rlabel metal2 135 -2968 135 -2964 1 CLK!
rlabel metal2 -223 -2968 -223 -2964 1 CLK!
rlabel metal2 -581 -2968 -581 -2964 1 CLK!
rlabel metal2 -939 -2968 -939 -2964 1 CLK!
rlabel metal2 -1238 -2968 -1238 -2964 1 CLK!
rlabel metal2 -1563 -2968 -1563 -2964 1 CLK!
rlabel metal2 -1826 -3710 -1826 -3706 1 CLK!
rlabel metal2 -1563 -3710 -1563 -3706 1 CLK!
rlabel metal2 -1563 -3881 -1563 -3877 1 CLK!
rlabel metal2 -1238 -3881 -1238 -3877 1 CLK!
rlabel metal2 -1563 -4056 -1563 -4052 1 CLK!
rlabel metal2 -1238 -4056 -1238 -4052 1 CLK!
rlabel metal2 -1238 -3710 -1238 -3706 1 CLK!
rlabel metal2 -938 -3710 -938 -3706 1 CLK!
rlabel metal2 -938 -3881 -938 -3877 1 CLK!
rlabel metal2 -939 -4056 -939 -4052 1 CLK!
rlabel metal2 -581 -4056 -581 -4052 1 CLK!
rlabel metal2 -581 -3881 -581 -3877 1 CLK!
rlabel metal2 -581 -3710 -581 -3706 1 CLK!
rlabel metal2 -223 -3710 -223 -3706 1 CLK!
rlabel metal2 -223 -3881 -223 -3877 1 CLK!
rlabel metal2 -223 -4056 -223 -4052 1 CLK!
rlabel metal2 135 -4056 135 -4052 1 CLK!
rlabel metal2 135 -3881 135 -3877 1 CLK!
rlabel metal2 491 -3881 491 -3877 1 CLK!
rlabel metal2 491 -4056 491 -4052 1 CLK!
rlabel metal2 849 -4056 849 -4052 1 CLK!
rlabel metal2 849 -3881 849 -3877 1 CLK!
rlabel metal2 1207 -3881 1207 -3877 1 CLK!
rlabel metal2 1207 -4056 1207 -4052 1 CLK!
rlabel metal2 -1818 -4453 -1818 -4449 1 CLK!
rlabel metal2 -1818 -4624 -1818 -4620 1 CLK!
rlabel metal2 -1555 -4624 -1555 -4620 1 CLK!
rlabel metal2 -1555 -4453 -1555 -4449 1 CLK!
rlabel metal2 -1555 -4795 -1555 -4791 1 CLK!
rlabel metal2 -1238 -4795 -1238 -4791 1 CLK!
rlabel metal2 -1238 -4624 -1238 -4620 1 CLK!
rlabel metal2 -1238 -4453 -1238 -4449 1 CLK!
rlabel metal2 -939 -4453 -939 -4449 1 CLK!
rlabel metal2 -939 -4624 -939 -4620 1 CLK!
rlabel metal2 -939 -4795 -939 -4791 1 CLK!
rlabel metal2 -581 -4795 -581 -4791 1 CLK!
rlabel metal2 -581 -4624 -581 -4620 1 CLK!
rlabel metal2 -581 -4453 -581 -4449 1 CLK!
rlabel metal2 -223 -4624 -223 -4620 1 CLK!
rlabel metal2 -223 -4795 -223 -4791 1 CLK!
rlabel metal2 135 -4795 135 -4791 1 CLK!
rlabel metal2 135 -4624 135 -4620 1 CLK!
rlabel metal2 491 -4624 491 -4620 1 CLK!
rlabel metal2 491 -4795 491 -4791 1 CLK!
rlabel metal2 849 -4795 849 -4791 1 CLK!
rlabel metal2 849 -4624 849 -4620 1 CLK!
rlabel metal2 1207 -4624 1207 -4620 1 CLK!
rlabel metal2 1207 -4795 1207 -4791 1 CLK!
rlabel metal2 -1814 -5519 -1814 -5515 1 CLK!
rlabel metal2 -1814 -5359 -1814 -5355 1 CLK!
rlabel metal2 -1814 -5188 -1814 -5184 1 CLK!
rlabel metal2 -1551 -5188 -1551 -5184 1 CLK!
rlabel metal2 -1551 -5359 -1551 -5355 1 CLK!
rlabel metal2 -1551 -5519 -1551 -5515 1 CLK!
rlabel metal2 -1238 -5519 -1238 -5515 1 CLK!
rlabel metal2 -1238 -5359 -1238 -5355 1 CLK!
rlabel metal2 -1238 -5188 -1238 -5184 1 CLK!
rlabel metal2 -939 -5188 -939 -5184 1 CLK!
rlabel metal2 -939 -5359 -939 -5355 1 CLK!
rlabel metal2 -939 -5519 -939 -5515 1 CLK!
rlabel metal2 -581 -5519 -581 -5515 1 CLK!
rlabel metal2 -581 -5359 -581 -5355 1 CLK!
rlabel metal2 -223 -5519 -223 -5515 1 CLK!
rlabel metal2 -223 -5359 -223 -5355 1 CLK!
rlabel metal2 135 -5359 135 -5355 1 CLK!
rlabel metal2 135 -5519 135 -5515 1 CLK!
rlabel metal2 491 -5519 491 -5515 1 CLK!
rlabel metal2 491 -5359 491 -5355 1 CLK!
rlabel metal2 849 -5359 849 -5355 1 CLK!
rlabel metal2 849 -5519 849 -5515 1 CLK!
rlabel metal2 1207 -5519 1207 -5515 1 CLK!
rlabel metal2 1207 -5359 1207 -5355 1 CLK!
rlabel metal2 -1238 -5915 -1238 -5911 1 CLK!
rlabel metal2 -939 -5915 -939 -5911 1 CLK!
rlabel metal2 -581 -5915 -581 -5911 1 CLK!
rlabel metal2 -223 -5915 -223 -5911 1 CLK!
rlabel metal2 135 -5915 135 -5911 1 CLK!
rlabel metal2 491 -5915 491 -5911 1 CLK!
rlabel metal2 849 -5915 849 -5911 1 CLK!
rlabel metal2 1207 -5915 1207 -5911 1 CLK!
rlabel metal2 1551 -5915 1551 -5911 1 CLK!
rlabel metal2 -1563 -1819 -1563 -1815 1 Y2
rlabel metal2 -1563 -2400 -1563 -2396 1 Y3
rlabel metal2 -1563 -2954 -1563 -2950 1 Y4
rlabel metal2 -1826 -3696 -1826 -3692 1 Y5
rlabel metal2 -1818 -4439 -1818 -4435 1 Y6
rlabel metal2 -1814 -5174 -1814 -5170 1 Y7
rlabel metal2 695 -2221 695 -2217 1 Z2
rlabel metal2 339 -2946 339 -2942 1 Z3
rlabel metal2 -19 -3688 -19 -3684 1 Z4
rlabel metal2 -377 -4431 -377 -4427 1 Z5
rlabel metal2 -735 -5166 -735 -5162 1 Z6
rlabel metal2 -1034 -5893 -1034 -5889 1 Z7
rlabel metal2 -735 -5893 -735 -5889 1 Z8
rlabel metal2 -377 -5893 -377 -5889 1 Z9
rlabel metal2 -19 -5893 -19 -5889 1 Z10
rlabel metal2 339 -5893 339 -5889 1 Z11
rlabel metal2 695 -5893 695 -5889 1 Z12
rlabel metal2 1053 -5893 1053 -5889 1 Z13
rlabel metal2 1411 -5893 1411 -5889 1 Z14
rlabel metal2 1755 -5893 1755 -5889 1 Z15
rlabel metal2 1818 -3600 1818 -3600 1 GND!
<< end >>
