magic
tech scmos
timestamp 1612988216
<< ntransistor >>
rect 3 -14 5 -10
rect 11 -14 13 -10
<< ptransistor >>
rect 3 14 5 23
rect 11 14 13 23
<< ndiffusion >>
rect 2 -14 3 -10
rect 5 -14 6 -10
rect 10 -14 11 -10
rect 13 -14 14 -10
<< pdiffusion >>
rect 2 14 3 23
rect 5 14 11 23
rect 13 14 14 23
<< ndcontact >>
rect -2 -14 2 -10
rect 6 -14 10 -10
rect 14 -14 18 -10
<< pdcontact >>
rect -2 14 2 23
rect 14 14 18 23
<< psubstratepcontact >>
rect -2 -22 2 -18
rect 14 -22 18 -18
<< nsubstratencontact >>
rect -2 27 2 31
rect 14 27 18 31
<< polysilicon >>
rect 3 23 5 25
rect 11 23 13 25
rect 3 11 5 14
rect 3 -10 5 7
rect 11 4 13 14
rect 11 -10 13 0
rect 3 -16 5 -14
rect 11 -16 13 -14
<< polycontact >>
rect 1 7 5 11
rect 9 0 13 4
<< metal1 >>
rect 2 27 14 31
rect -2 23 2 27
rect -2 7 1 11
rect 18 6 22 23
rect -2 0 9 4
rect 18 2 26 6
rect 18 -3 22 2
rect 6 -7 22 -3
rect 6 -10 10 -7
rect -2 -18 2 -14
rect 14 -18 18 -14
rect 2 -22 14 -18
<< labels >>
rlabel metal1 -2 7 -2 11 3 a
rlabel metal1 -2 0 -2 4 3 b
rlabel metal1 8 29 8 29 5 VDD!
rlabel metal1 8 -20 8 -20 1 GND!
rlabel metal1 26 2 26 6 7 out
<< end >>
