magic
tech scmos
timestamp 1615598126
<< ntransistor >>
rect 3 -25 5 -21
rect 11 -25 13 -21
<< ptransistor >>
rect 3 31 5 40
rect 11 31 13 40
<< ndiffusion >>
rect 2 -25 3 -21
rect 5 -25 6 -21
rect 10 -25 11 -21
rect 13 -25 14 -21
<< pdiffusion >>
rect 2 31 3 40
rect 5 31 11 40
rect 13 31 14 40
<< ndcontact >>
rect -2 -25 2 -21
rect 6 -25 10 -21
rect 14 -25 18 -21
<< pdcontact >>
rect -2 31 2 40
rect 14 31 18 40
<< psubstratepcontact >>
rect -2 -33 2 -29
rect 14 -33 18 -29
<< nsubstratencontact >>
rect -2 44 2 48
<< polysilicon >>
rect 3 40 5 42
rect 11 40 13 42
rect 3 11 5 31
rect 3 -21 5 7
rect 11 4 13 31
rect 11 -21 13 0
rect 3 -27 5 -25
rect 11 -27 13 -25
<< polycontact >>
rect 1 7 5 11
rect 9 0 13 4
<< metal1 >>
rect -6 44 -2 48
rect 2 44 22 48
rect -2 40 2 44
rect -2 7 1 11
rect -2 0 9 4
rect 18 -14 22 40
rect 6 -18 22 -14
rect 6 -21 10 -18
rect -2 -29 2 -25
rect 14 -29 18 -25
rect -6 -33 -2 -29
rect 2 -33 14 -29
rect 18 -33 22 -29
<< labels >>
rlabel metal1 8 46 8 46 5 VDD!
rlabel metal1 -2 7 -2 11 3 A
rlabel metal1 -2 0 -2 4 3 B
rlabel metal1 22 7 22 11 7 OUT
rlabel metal1 8 -31 8 -31 1 GND!
<< end >>
