magic
tech scmos
timestamp 1612915487
<< ntransistor >>
rect 5 -25 7 -21
<< ptransistor >>
rect 5 -9 7 0
<< ndiffusion >>
rect 4 -25 5 -21
rect 7 -25 8 -21
<< pdiffusion >>
rect 4 -9 5 0
rect 7 -9 8 0
<< ndcontact >>
rect 0 -25 4 -21
rect 8 -25 12 -21
<< pdcontact >>
rect 0 -9 4 0
rect 8 -9 12 0
<< psubstratepcontact >>
rect -4 -33 0 -29
rect 8 -33 12 -29
<< nsubstratencontact >>
rect -4 4 0 8
rect 8 4 12 8
<< polysilicon >>
rect 5 0 7 2
rect 5 -13 7 -9
rect 4 -17 7 -13
rect 5 -21 7 -17
rect 5 -27 7 -25
<< polycontact >>
rect 0 -17 4 -13
<< metal1 >>
rect 0 4 8 8
rect 0 0 4 4
rect 8 -13 12 -9
rect 8 -17 16 -13
rect 8 -21 12 -17
rect 0 -29 4 -25
rect 0 -33 8 -29
<< labels >>
rlabel polycontact 0 -17 0 -13 3 in
rlabel metal1 16 -17 16 -13 7 out
rlabel metal1 4 6 4 6 5 VDD!
rlabel metal1 4 -31 4 -31 1 GND!
<< end >>
