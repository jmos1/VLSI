magic
tech scmos
timestamp 1612987764
<< ntransistor >>
rect -60 2 -58 6
rect -37 2 -35 6
rect -9 2 -7 6
rect -1 2 1 6
rect 7 2 9 6
rect 15 2 17 6
<< ptransistor >>
rect -60 32 -58 41
rect -37 32 -35 41
rect -9 32 -7 41
rect -1 32 1 41
rect 7 32 9 41
rect 15 32 17 41
<< ndiffusion >>
rect -61 2 -60 6
rect -58 2 -57 6
rect -38 2 -37 6
rect -35 2 -34 6
rect -10 2 -9 6
rect -7 2 -1 6
rect 1 2 2 6
rect 6 2 7 6
rect 9 2 15 6
rect 17 2 18 6
<< pdiffusion >>
rect -61 32 -60 41
rect -58 32 -57 41
rect -38 32 -37 41
rect -35 32 -34 41
rect -10 32 -9 41
rect -7 32 -1 41
rect 1 32 2 41
rect 6 32 7 41
rect 9 32 15 41
rect 17 32 18 41
<< ndcontact >>
rect -65 2 -61 6
rect -57 2 -53 6
rect -42 2 -38 6
rect -34 2 -30 6
rect -14 2 -10 6
rect 2 2 6 6
rect 18 2 22 6
<< pdcontact >>
rect -65 32 -61 41
rect -57 32 -53 41
rect -42 32 -38 41
rect -34 32 -30 41
rect -14 32 -10 41
rect 2 32 6 41
rect 18 32 22 41
<< psubstratepcontact >>
rect -65 -10 -61 -6
rect -42 -10 -38 -6
rect -14 -10 -10 -6
rect 18 -10 22 -6
<< nsubstratencontact >>
rect -65 54 -61 58
rect -42 54 -38 58
rect -14 54 -10 58
rect 18 54 22 58
<< polysilicon >>
rect -60 51 17 53
rect -60 41 -58 51
rect -19 46 1 48
rect -37 41 -35 43
rect -60 24 -58 32
rect -61 20 -58 24
rect -60 6 -58 20
rect -37 17 -35 32
rect -38 13 -35 17
rect -37 6 -35 13
rect -60 0 -58 2
rect -37 -1 -35 2
rect -19 -1 -17 46
rect -9 41 -7 43
rect -1 41 1 46
rect 7 41 9 43
rect 15 41 17 51
rect -9 29 -7 32
rect -1 30 1 32
rect -9 19 -7 25
rect 7 24 9 32
rect 15 29 17 32
rect 15 27 25 29
rect 7 22 17 24
rect -9 17 9 19
rect -9 6 -7 8
rect -1 6 1 8
rect 7 6 9 17
rect 15 6 17 18
rect -9 -1 -7 2
rect -37 -3 -7 -1
rect -1 -3 1 2
rect 7 0 9 2
rect 15 0 17 2
rect 23 -3 25 27
rect -1 -5 25 -3
<< polycontact >>
rect -65 20 -61 24
rect 13 18 17 22
<< metal1 >>
rect -69 54 -65 58
rect -61 54 -42 58
rect -38 54 -14 58
rect -10 54 18 58
rect 22 54 26 58
rect -65 41 -61 54
rect -42 41 -38 54
rect -14 41 -10 54
rect 18 41 22 54
rect -57 6 -53 32
rect -34 22 -30 32
rect 2 29 6 32
rect 2 25 24 29
rect -34 18 13 22
rect 20 21 24 25
rect -34 6 -30 18
rect 20 17 29 21
rect 20 13 24 17
rect 2 9 24 13
rect 2 6 6 9
rect -65 -6 -61 2
rect -42 -6 -38 2
rect -14 -6 -10 2
rect 18 -6 22 2
rect -69 -10 -65 -6
rect -61 -10 -42 -6
rect -38 -10 -14 -6
rect -10 -10 18 -6
rect 22 -10 26 -6
<< m2contact >>
rect -53 25 -49 29
<< pm12contact >>
rect -11 25 -7 29
rect -42 13 -38 17
<< metal2 >>
rect -49 25 -11 29
rect -65 13 -42 17
<< labels >>
rlabel polycontact -65 20 -65 24 3 a
rlabel metal2 -65 13 -65 17 3 b
rlabel metal1 29 17 29 21 7 out
rlabel metal1 -20 56 -20 56 5 VDD!
rlabel metal1 -22 -8 -22 -8 1 GND!
<< end >>
