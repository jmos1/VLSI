magic
tech scmos
timestamp 1615598037
<< ntransistor >>
rect 55 23 57 27
rect 63 23 65 27
<< ptransistor >>
rect 55 79 57 88
rect 63 79 65 88
<< ndiffusion >>
rect 54 23 55 27
rect 57 23 63 27
rect 65 23 66 27
<< pdiffusion >>
rect 54 79 55 88
rect 57 79 58 88
rect 62 79 63 88
rect 65 79 66 88
<< ndcontact >>
rect 50 23 54 27
rect 66 23 70 27
<< pdcontact >>
rect 50 79 54 88
rect 58 79 62 88
rect 66 79 70 88
<< psubstratepcontact >>
rect 50 15 54 19
<< nsubstratencontact >>
rect 50 92 54 96
rect 66 92 70 96
<< polysilicon >>
rect 55 88 57 90
rect 63 88 65 90
rect 55 27 57 79
rect 63 52 65 79
rect 63 27 65 48
rect 55 21 57 23
rect 63 21 65 23
<< polycontact >>
rect 51 55 55 59
rect 61 48 65 52
<< metal1 >>
rect 46 92 50 96
rect 54 92 66 96
rect 70 92 74 96
rect 50 88 54 92
rect 66 88 70 92
rect 58 59 62 79
rect 46 55 51 59
rect 58 55 74 59
rect 46 48 61 52
rect 70 23 74 55
rect 50 19 54 23
rect 46 15 50 19
rect 54 15 74 19
<< labels >>
rlabel metal1 60 17 60 17 1 GND!
rlabel metal1 46 55 46 59 3 A
rlabel metal1 46 48 46 52 3 B
rlabel metal1 74 48 74 52 7 OUT
rlabel metal1 60 94 60 94 5 VDD!
<< end >>
