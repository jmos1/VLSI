magic
tech scmos
timestamp 1613140719
<< ntransistor >>
rect -121 -21 -119 -17
rect -91 -21 -89 -17
rect -61 -21 -59 -17
rect -53 -21 -51 -17
rect -19 -21 -17 -17
rect -11 -21 -9 -17
rect 20 -21 22 -17
rect 28 -21 30 -17
rect 58 -21 60 -17
rect 66 -21 68 -17
rect 106 -21 108 -17
rect 114 -21 116 -17
rect 148 -21 150 -17
rect 156 -21 158 -17
rect 187 -21 189 -17
rect 195 -21 197 -17
rect 225 -21 227 -17
rect 233 -21 235 -17
<< ptransistor >>
rect -121 7 -119 16
rect -91 7 -89 16
rect -61 7 -59 16
rect -53 7 -51 16
rect -19 7 -17 16
rect -11 7 -9 16
rect 20 7 22 16
rect 28 7 30 16
rect 58 7 60 16
rect 66 7 68 16
rect 106 7 108 16
rect 114 7 116 16
rect 148 7 150 16
rect 156 7 158 16
rect 187 7 189 16
rect 195 7 197 16
rect 225 7 227 16
rect 233 7 235 16
<< ndiffusion >>
rect -122 -21 -121 -17
rect -119 -21 -118 -17
rect -92 -21 -91 -17
rect -89 -21 -88 -17
rect -62 -21 -61 -17
rect -59 -21 -53 -17
rect -51 -21 -50 -17
rect -20 -21 -19 -17
rect -17 -21 -11 -17
rect -9 -21 -8 -17
rect 19 -21 20 -17
rect 22 -21 28 -17
rect 30 -21 31 -17
rect 57 -21 58 -17
rect 60 -21 66 -17
rect 68 -21 69 -17
rect 105 -21 106 -17
rect 108 -21 114 -17
rect 116 -21 117 -17
rect 147 -21 148 -17
rect 150 -21 156 -17
rect 158 -21 159 -17
rect 186 -21 187 -17
rect 189 -21 195 -17
rect 197 -21 198 -17
rect 224 -21 225 -17
rect 227 -21 233 -17
rect 235 -21 236 -17
<< pdiffusion >>
rect -122 7 -121 16
rect -119 7 -118 16
rect -92 7 -91 16
rect -89 7 -88 16
rect -62 7 -61 16
rect -59 7 -58 16
rect -54 7 -53 16
rect -51 7 -50 16
rect -20 7 -19 16
rect -17 7 -16 16
rect -12 7 -11 16
rect -9 7 -8 16
rect 19 7 20 16
rect 22 7 23 16
rect 27 7 28 16
rect 30 7 31 16
rect 57 7 58 16
rect 60 7 61 16
rect 65 7 66 16
rect 68 7 69 16
rect 105 7 106 16
rect 108 7 109 16
rect 113 7 114 16
rect 116 7 117 16
rect 147 7 148 16
rect 150 7 151 16
rect 155 7 156 16
rect 158 7 159 16
rect 186 7 187 16
rect 189 7 190 16
rect 194 7 195 16
rect 197 7 198 16
rect 224 7 225 16
rect 227 7 228 16
rect 232 7 233 16
rect 235 7 236 16
<< ndcontact >>
rect -126 -21 -122 -17
rect -118 -21 -114 -17
rect -96 -21 -92 -17
rect -88 -21 -84 -17
rect -66 -21 -62 -17
rect -50 -21 -46 -17
rect -24 -21 -20 -17
rect -8 -21 -4 -17
rect 15 -21 19 -17
rect 31 -21 35 -17
rect 53 -21 57 -17
rect 69 -21 73 -17
rect 101 -21 105 -17
rect 117 -21 121 -17
rect 143 -21 147 -17
rect 159 -21 163 -17
rect 182 -21 186 -17
rect 198 -21 202 -17
rect 220 -21 224 -17
rect 236 -21 240 -17
<< pdcontact >>
rect -126 7 -122 16
rect -118 7 -114 16
rect -96 7 -92 16
rect -88 7 -84 16
rect -66 7 -62 16
rect -58 7 -54 16
rect -50 7 -46 16
rect -24 7 -20 16
rect -16 7 -12 16
rect -8 7 -4 16
rect 15 7 19 16
rect 23 7 27 16
rect 31 7 35 16
rect 53 7 57 16
rect 61 7 65 16
rect 69 7 73 16
rect 101 7 105 16
rect 109 7 113 16
rect 117 7 121 16
rect 143 7 147 16
rect 151 7 155 16
rect 159 7 163 16
rect 182 7 186 16
rect 190 7 194 16
rect 198 7 202 16
rect 220 7 224 16
rect 228 7 232 16
rect 236 7 240 16
<< psubstratepcontact >>
rect -126 -34 -122 -30
rect -96 -34 -92 -30
rect -66 -34 -62 -30
rect -24 -34 -20 -30
rect 15 -34 19 -30
rect 53 -34 57 -30
rect 101 -34 105 -30
rect 143 -34 147 -30
rect 182 -34 186 -30
rect 220 -34 224 -30
<< nsubstratencontact >>
rect -126 20 -122 24
rect -96 20 -92 24
rect -66 20 -62 24
rect -50 20 -46 24
rect -24 20 -20 24
rect -8 20 -4 24
rect 15 20 19 24
rect 31 20 35 24
rect 53 20 57 24
rect 69 20 73 24
rect 101 20 105 24
rect 117 20 121 24
rect 143 20 147 24
rect 159 20 163 24
rect 182 20 186 24
rect 198 20 202 24
rect 220 20 224 24
rect 236 20 240 24
<< polysilicon >>
rect -121 16 -119 18
rect -91 16 -89 18
rect -61 16 -59 18
rect -53 16 -51 18
rect -19 16 -17 18
rect -11 16 -9 18
rect 20 16 22 18
rect 28 16 30 18
rect 58 16 60 18
rect 66 16 68 18
rect 106 16 108 18
rect 114 16 116 18
rect 148 16 150 18
rect 156 16 158 18
rect 187 16 189 18
rect 195 16 197 18
rect 225 16 227 18
rect 233 16 235 18
rect -121 -10 -119 7
rect -91 3 -89 7
rect -92 -1 -89 3
rect -122 -14 -119 -10
rect -121 -17 -119 -14
rect -91 -17 -89 -1
rect -61 -17 -59 7
rect -53 -10 -51 7
rect -53 -17 -51 -14
rect -19 -17 -17 7
rect -11 -10 -9 7
rect -11 -17 -9 -14
rect 20 -17 22 7
rect 28 -10 30 7
rect 58 -3 60 7
rect 28 -17 30 -14
rect 58 -17 60 -7
rect 66 -10 68 7
rect 66 -17 68 -14
rect 106 -17 108 7
rect 114 -10 116 7
rect 114 -17 116 -14
rect 148 -17 150 7
rect 156 -10 158 7
rect 156 -17 158 -14
rect 187 -17 189 7
rect 195 -10 197 7
rect 225 -3 227 7
rect 195 -17 197 -14
rect 225 -17 227 -7
rect 233 -10 235 7
rect 233 -17 235 -14
rect -121 -23 -119 -21
rect -91 -23 -89 -21
rect -61 -23 -59 -21
rect -53 -23 -51 -21
rect -19 -23 -17 -21
rect -11 -23 -9 -21
rect 20 -23 22 -21
rect 28 -23 30 -21
rect 58 -23 60 -21
rect 66 -23 68 -21
rect 106 -23 108 -21
rect 114 -23 116 -21
rect 148 -23 150 -21
rect 156 -23 158 -21
rect 187 -23 189 -21
rect 195 -23 197 -21
rect 225 -23 227 -21
rect 233 -23 235 -21
<< polycontact >>
rect -65 0 -61 4
<< metal1 >>
rect -130 20 -126 24
rect -122 20 -96 24
rect -92 20 -66 24
rect -62 20 -50 24
rect -46 20 -24 24
rect -20 20 -8 24
rect -4 20 15 24
rect 19 20 31 24
rect 35 20 53 24
rect 57 20 69 24
rect 73 20 101 24
rect 105 20 117 24
rect 121 20 143 24
rect 147 20 159 24
rect 163 20 182 24
rect 186 20 198 24
rect 202 20 220 24
rect 224 20 236 24
rect 240 20 247 24
rect -126 16 -122 20
rect -96 16 -92 20
rect -66 16 -62 20
rect -50 16 -46 20
rect -24 16 -20 20
rect -8 16 -4 20
rect 15 16 19 20
rect 31 16 35 20
rect 53 16 57 20
rect 69 16 73 20
rect 101 16 105 20
rect 117 16 121 20
rect 143 16 147 20
rect 159 16 163 20
rect 182 16 186 20
rect 198 16 202 20
rect 220 16 224 20
rect 236 16 240 20
rect -118 -10 -114 7
rect -88 4 -84 7
rect -58 4 -54 7
rect -16 4 -12 7
rect 23 4 27 7
rect 61 4 65 7
rect 109 4 113 7
rect 151 4 155 7
rect 190 4 194 7
rect 228 4 232 7
rect -88 0 -65 4
rect -58 0 -42 4
rect -16 0 0 4
rect 23 0 39 4
rect 61 0 73 4
rect 109 0 125 4
rect 151 0 167 4
rect 190 0 206 4
rect 228 0 240 4
rect 244 0 248 4
rect -118 -14 -100 -10
rect -118 -17 -114 -14
rect -88 -17 -84 0
rect -46 -3 -42 0
rect -46 -21 -42 -7
rect -4 -10 0 0
rect 35 -10 39 0
rect 73 -3 77 0
rect 121 -3 125 0
rect 73 -7 90 -3
rect -4 -21 0 -14
rect 35 -21 39 -14
rect 73 -21 77 -7
rect 121 -21 125 -7
rect 163 -10 167 0
rect 202 -10 206 0
rect 163 -21 167 -14
rect 202 -21 206 -14
rect 240 -21 244 0
rect -126 -30 -122 -21
rect -96 -30 -92 -21
rect -66 -30 -62 -21
rect -24 -30 -20 -21
rect 15 -30 19 -21
rect 53 -30 57 -21
rect 101 -30 105 -21
rect 143 -30 147 -21
rect 182 -30 186 -21
rect 220 -30 224 -21
rect -130 -34 -126 -30
rect -122 -34 -96 -30
rect -92 -34 -66 -30
rect -62 -34 -24 -30
rect -20 -34 15 -30
rect 19 -34 53 -30
rect 57 -34 101 -30
rect 105 -34 143 -30
rect 147 -34 182 -30
rect 186 -34 220 -30
rect 224 -34 246 -30
<< m2contact >>
rect 73 0 77 4
rect 240 0 244 4
rect 35 -14 39 -10
rect 202 -14 206 -10
<< pm12contact >>
rect -96 -1 -92 3
rect -23 0 -19 4
rect 16 0 20 4
rect 102 0 106 4
rect 144 0 148 4
rect 183 0 187 4
rect -126 -14 -122 -10
rect -100 -14 -96 -10
rect -46 -7 -42 -3
rect -55 -14 -51 -10
rect 56 -7 60 -3
rect 90 -7 94 -3
rect 121 -7 125 -3
rect -13 -14 -9 -10
rect -4 -14 0 -10
rect 26 -14 30 -10
rect 64 -14 68 -10
rect 112 -14 116 -10
rect 223 -7 227 -3
rect 154 -14 158 -10
rect 163 -14 167 -10
rect 193 -14 197 -10
rect 231 -14 235 -10
<< metal2 >>
rect -96 -3 -92 -1
rect -56 0 -23 4
rect 20 0 73 4
rect 83 0 102 4
rect 111 0 144 4
rect 187 0 240 4
rect -56 -3 -52 0
rect -137 -7 -52 -3
rect -42 -7 56 -3
rect 83 -10 87 0
rect 111 -3 115 0
rect 94 -7 115 -3
rect 125 -7 223 -3
rect -137 -14 -126 -10
rect -96 -14 -55 -10
rect -51 -14 -13 -10
rect 0 -14 26 -10
rect 39 -14 64 -10
rect 68 -14 87 -10
rect 91 -14 112 -10
rect 116 -14 154 -10
rect 167 -14 193 -10
rect 206 -14 231 -10
rect 235 -14 248 -10
rect -133 -22 -129 -14
rect 91 -22 95 -14
rect -133 -26 95 -22
<< labels >>
rlabel metal2 -137 -7 -137 -3 3 D
rlabel metal2 -137 -14 -137 -10 3 CLK
rlabel metal2 248 -14 248 -10 7 QNOT
rlabel metal1 248 0 248 4 7 Q
rlabel metal1 80 -33 80 -33 1 GND!
rlabel metal1 82 23 82 23 5 VDD!
<< end >>
