magic
tech scmos
timestamp 1612988274
<< ntransistor >>
rect -3 -9 -1 -5
rect 5 -9 7 -5
rect 24 -9 26 -5
<< ptransistor >>
rect -3 19 -1 28
rect 5 19 7 28
rect 24 19 26 28
<< ndiffusion >>
rect -4 -9 -3 -5
rect -1 -9 0 -5
rect 4 -9 5 -5
rect 7 -9 8 -5
rect 23 -9 24 -5
rect 26 -9 27 -5
<< pdiffusion >>
rect -4 19 -3 28
rect -1 19 5 28
rect 7 19 8 28
rect 23 19 24 28
rect 26 19 27 28
<< ndcontact >>
rect -8 -9 -4 -5
rect 0 -9 4 -5
rect 8 -9 12 -5
rect 19 -9 23 -5
rect 27 -9 31 -5
<< pdcontact >>
rect -8 19 -4 28
rect 8 19 12 28
rect 19 19 23 28
rect 27 19 31 28
<< psubstratepcontact >>
rect -8 -17 -4 -13
rect 8 -17 12 -13
rect 19 -17 23 -13
<< nsubstratencontact >>
rect -8 32 -4 36
rect 19 32 23 36
<< polysilicon >>
rect -3 28 -1 30
rect 5 28 7 30
rect 24 28 26 30
rect -3 16 -1 19
rect -3 -5 -1 12
rect 5 9 7 19
rect 24 11 26 19
rect 23 7 26 11
rect 5 -5 7 5
rect 24 -5 26 7
rect -3 -11 -1 -9
rect 5 -11 7 -9
rect 24 -11 26 -9
<< polycontact >>
rect -5 12 -1 16
rect 3 5 7 9
rect 19 7 23 11
<< metal1 >>
rect -12 32 -8 36
rect -4 32 19 36
rect 23 32 35 36
rect -8 28 -4 32
rect 19 28 23 32
rect -12 12 -5 16
rect 12 11 16 28
rect 27 11 31 19
rect -12 5 3 9
rect 12 7 19 11
rect 27 7 35 11
rect 12 2 16 7
rect 0 -2 16 2
rect 0 -5 4 -2
rect 27 -5 31 7
rect -8 -13 -4 -9
rect 8 -13 12 -9
rect 19 -13 23 -9
rect -12 -17 -8 -13
rect -4 -17 8 -13
rect 12 -17 19 -13
rect 23 -17 35 -13
<< labels >>
rlabel metal1 35 7 35 11 7 out
rlabel psubstratepcontact 10 -15 10 -15 1 GND!
rlabel metal1 -12 12 -12 16 3 a
rlabel metal1 -12 5 -12 9 3 b
rlabel metal1 10 34 10 34 5 VDD!
<< end >>
