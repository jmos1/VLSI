magic
tech scmos
timestamp 1619535334
<< polysilicon >>
rect -1332 -1038 -1330 -1036
rect -1324 -1038 -1322 -1036
rect -1314 -1038 -1312 -1036
rect -931 -1038 -929 -1036
rect -923 -1038 -921 -1036
rect -913 -1038 -911 -1036
rect -572 -1038 -570 -1036
rect -564 -1038 -562 -1036
rect -554 -1038 -552 -1036
rect -214 -1038 -212 -1036
rect -206 -1038 -204 -1036
rect -196 -1038 -194 -1036
rect 214 -1038 216 -1036
rect 222 -1038 224 -1036
rect 232 -1038 234 -1036
rect 570 -1038 572 -1036
rect 578 -1038 580 -1036
rect 588 -1038 590 -1036
rect 968 -1038 970 -1036
rect 976 -1038 978 -1036
rect 986 -1038 988 -1036
rect 1326 -1038 1328 -1036
rect 1334 -1038 1336 -1036
rect 1344 -1038 1346 -1036
rect -1332 -1114 -1330 -1046
rect -1324 -1070 -1322 -1046
rect -1324 -1114 -1322 -1074
rect -1314 -1114 -1312 -1046
rect -931 -1114 -929 -1046
rect -923 -1070 -921 -1046
rect -923 -1114 -921 -1074
rect -913 -1114 -911 -1046
rect -572 -1114 -570 -1046
rect -564 -1070 -562 -1046
rect -564 -1114 -562 -1074
rect -554 -1114 -552 -1046
rect -214 -1114 -212 -1046
rect -206 -1070 -204 -1046
rect -206 -1114 -204 -1074
rect -196 -1114 -194 -1046
rect 214 -1114 216 -1046
rect 222 -1070 224 -1046
rect 222 -1114 224 -1074
rect 232 -1114 234 -1046
rect 570 -1114 572 -1046
rect 578 -1070 580 -1046
rect 578 -1114 580 -1074
rect 588 -1114 590 -1046
rect 968 -1114 970 -1046
rect 976 -1070 978 -1046
rect 976 -1114 978 -1074
rect 986 -1114 988 -1046
rect 1326 -1114 1328 -1046
rect 1334 -1070 1336 -1046
rect 1334 -1114 1336 -1074
rect 1344 -1114 1346 -1046
rect -1332 -1120 -1330 -1118
rect -1324 -1120 -1322 -1118
rect -1314 -1120 -1312 -1118
rect -931 -1120 -929 -1118
rect -923 -1120 -921 -1118
rect -913 -1120 -911 -1118
rect -572 -1120 -570 -1118
rect -564 -1120 -562 -1118
rect -554 -1120 -552 -1118
rect -214 -1120 -212 -1118
rect -206 -1120 -204 -1118
rect -196 -1120 -194 -1118
rect 214 -1120 216 -1118
rect 222 -1120 224 -1118
rect 232 -1120 234 -1118
rect 570 -1120 572 -1118
rect 578 -1120 580 -1118
rect 588 -1120 590 -1118
rect 968 -1120 970 -1118
rect 976 -1120 978 -1118
rect 986 -1120 988 -1118
rect 1326 -1120 1328 -1118
rect 1334 -1120 1336 -1118
rect 1344 -1120 1346 -1118
rect -1255 -1152 -1253 -1150
rect -1245 -1152 -1243 -1150
rect -1229 -1152 -1227 -1150
rect -1221 -1152 -1219 -1150
rect -1205 -1152 -1203 -1150
rect -1197 -1152 -1195 -1150
rect -1187 -1152 -1185 -1150
rect -1179 -1152 -1177 -1150
rect -1163 -1152 -1161 -1150
rect -1155 -1152 -1153 -1150
rect -1145 -1152 -1143 -1150
rect -1137 -1152 -1135 -1150
rect -1121 -1152 -1119 -1150
rect -1113 -1152 -1111 -1150
rect -1103 -1152 -1101 -1150
rect -1095 -1152 -1093 -1150
rect -1079 -1152 -1077 -1150
rect -1071 -1152 -1069 -1150
rect -930 -1152 -928 -1150
rect -920 -1152 -918 -1150
rect -904 -1152 -902 -1150
rect -896 -1152 -894 -1150
rect -880 -1152 -878 -1150
rect -872 -1152 -870 -1150
rect -862 -1152 -860 -1150
rect -854 -1152 -852 -1150
rect -838 -1152 -836 -1150
rect -830 -1152 -828 -1150
rect -820 -1152 -818 -1150
rect -812 -1152 -810 -1150
rect -796 -1152 -794 -1150
rect -788 -1152 -786 -1150
rect -778 -1152 -776 -1150
rect -770 -1152 -768 -1150
rect -754 -1152 -752 -1150
rect -746 -1152 -744 -1150
rect -572 -1152 -570 -1150
rect -562 -1152 -560 -1150
rect -546 -1152 -544 -1150
rect -538 -1152 -536 -1150
rect -522 -1152 -520 -1150
rect -514 -1152 -512 -1150
rect -504 -1152 -502 -1150
rect -496 -1152 -494 -1150
rect -480 -1152 -478 -1150
rect -472 -1152 -470 -1150
rect -462 -1152 -460 -1150
rect -454 -1152 -452 -1150
rect -438 -1152 -436 -1150
rect -430 -1152 -428 -1150
rect -420 -1152 -418 -1150
rect -412 -1152 -410 -1150
rect -396 -1152 -394 -1150
rect -388 -1152 -386 -1150
rect -214 -1152 -212 -1150
rect -204 -1152 -202 -1150
rect -188 -1152 -186 -1150
rect -180 -1152 -178 -1150
rect -164 -1152 -162 -1150
rect -156 -1152 -154 -1150
rect -146 -1152 -144 -1150
rect -138 -1152 -136 -1150
rect -122 -1152 -120 -1150
rect -114 -1152 -112 -1150
rect -104 -1152 -102 -1150
rect -96 -1152 -94 -1150
rect -80 -1152 -78 -1150
rect -72 -1152 -70 -1150
rect -62 -1152 -60 -1150
rect -54 -1152 -52 -1150
rect -38 -1152 -36 -1150
rect -30 -1152 -28 -1150
rect 214 -1152 216 -1150
rect 224 -1152 226 -1150
rect 240 -1152 242 -1150
rect 248 -1152 250 -1150
rect 264 -1152 266 -1150
rect 272 -1152 274 -1150
rect 282 -1152 284 -1150
rect 290 -1152 292 -1150
rect 306 -1152 308 -1150
rect 314 -1152 316 -1150
rect 324 -1152 326 -1150
rect 332 -1152 334 -1150
rect 348 -1152 350 -1150
rect 356 -1152 358 -1150
rect 366 -1152 368 -1150
rect 374 -1152 376 -1150
rect 390 -1152 392 -1150
rect 398 -1152 400 -1150
rect 570 -1152 572 -1150
rect 580 -1152 582 -1150
rect 596 -1152 598 -1150
rect 604 -1152 606 -1150
rect 620 -1152 622 -1150
rect 628 -1152 630 -1150
rect 638 -1152 640 -1150
rect 646 -1152 648 -1150
rect 662 -1152 664 -1150
rect 670 -1152 672 -1150
rect 680 -1152 682 -1150
rect 688 -1152 690 -1150
rect 704 -1152 706 -1150
rect 712 -1152 714 -1150
rect 722 -1152 724 -1150
rect 730 -1152 732 -1150
rect 746 -1152 748 -1150
rect 754 -1152 756 -1150
rect 968 -1152 970 -1150
rect 978 -1152 980 -1150
rect 994 -1152 996 -1150
rect 1002 -1152 1004 -1150
rect 1018 -1152 1020 -1150
rect 1026 -1152 1028 -1150
rect 1036 -1152 1038 -1150
rect 1044 -1152 1046 -1150
rect 1060 -1152 1062 -1150
rect 1068 -1152 1070 -1150
rect 1078 -1152 1080 -1150
rect 1086 -1152 1088 -1150
rect 1102 -1152 1104 -1150
rect 1110 -1152 1112 -1150
rect 1120 -1152 1122 -1150
rect 1128 -1152 1130 -1150
rect 1144 -1152 1146 -1150
rect 1152 -1152 1154 -1150
rect -1255 -1228 -1253 -1160
rect -1245 -1228 -1243 -1160
rect -1229 -1228 -1227 -1160
rect -1221 -1228 -1219 -1160
rect -1205 -1228 -1203 -1160
rect -1197 -1228 -1195 -1160
rect -1187 -1228 -1185 -1160
rect -1179 -1228 -1177 -1160
rect -1163 -1228 -1161 -1160
rect -1155 -1193 -1153 -1160
rect -1145 -1193 -1143 -1160
rect -1155 -1195 -1143 -1193
rect -1155 -1228 -1153 -1195
rect -1145 -1228 -1143 -1195
rect -1137 -1228 -1135 -1160
rect -1121 -1228 -1119 -1160
rect -1113 -1228 -1111 -1160
rect -1103 -1228 -1101 -1160
rect -1095 -1228 -1093 -1160
rect -1079 -1228 -1077 -1160
rect -1071 -1228 -1069 -1160
rect -930 -1228 -928 -1160
rect -920 -1228 -918 -1160
rect -904 -1228 -902 -1160
rect -896 -1228 -894 -1160
rect -880 -1228 -878 -1160
rect -872 -1228 -870 -1160
rect -862 -1228 -860 -1160
rect -854 -1228 -852 -1160
rect -838 -1228 -836 -1160
rect -830 -1193 -828 -1160
rect -820 -1193 -818 -1160
rect -830 -1195 -818 -1193
rect -830 -1228 -828 -1195
rect -820 -1228 -818 -1195
rect -812 -1228 -810 -1160
rect -796 -1228 -794 -1160
rect -788 -1228 -786 -1160
rect -778 -1228 -776 -1160
rect -770 -1228 -768 -1160
rect -754 -1228 -752 -1160
rect -746 -1228 -744 -1160
rect -572 -1228 -570 -1160
rect -562 -1228 -560 -1160
rect -546 -1228 -544 -1160
rect -538 -1228 -536 -1160
rect -522 -1228 -520 -1160
rect -514 -1228 -512 -1160
rect -504 -1228 -502 -1160
rect -496 -1228 -494 -1160
rect -480 -1228 -478 -1160
rect -472 -1193 -470 -1160
rect -462 -1193 -460 -1160
rect -472 -1195 -460 -1193
rect -472 -1228 -470 -1195
rect -462 -1228 -460 -1195
rect -454 -1228 -452 -1160
rect -438 -1228 -436 -1160
rect -430 -1228 -428 -1160
rect -420 -1228 -418 -1160
rect -412 -1228 -410 -1160
rect -396 -1228 -394 -1160
rect -388 -1228 -386 -1160
rect -214 -1228 -212 -1160
rect -204 -1228 -202 -1160
rect -188 -1228 -186 -1160
rect -180 -1228 -178 -1160
rect -164 -1228 -162 -1160
rect -156 -1228 -154 -1160
rect -146 -1228 -144 -1160
rect -138 -1228 -136 -1160
rect -122 -1228 -120 -1160
rect -114 -1193 -112 -1160
rect -104 -1193 -102 -1160
rect -114 -1195 -102 -1193
rect -114 -1228 -112 -1195
rect -104 -1228 -102 -1195
rect -96 -1228 -94 -1160
rect -80 -1228 -78 -1160
rect -72 -1228 -70 -1160
rect -62 -1228 -60 -1160
rect -54 -1228 -52 -1160
rect -38 -1228 -36 -1160
rect -30 -1228 -28 -1160
rect 214 -1228 216 -1160
rect 224 -1228 226 -1160
rect 240 -1228 242 -1160
rect 248 -1228 250 -1160
rect 264 -1228 266 -1160
rect 272 -1228 274 -1160
rect 282 -1228 284 -1160
rect 290 -1228 292 -1160
rect 306 -1228 308 -1160
rect 314 -1193 316 -1160
rect 324 -1193 326 -1160
rect 314 -1195 326 -1193
rect 314 -1228 316 -1195
rect 324 -1228 326 -1195
rect 332 -1228 334 -1160
rect 348 -1228 350 -1160
rect 356 -1228 358 -1160
rect 366 -1228 368 -1160
rect 374 -1228 376 -1160
rect 390 -1228 392 -1160
rect 398 -1228 400 -1160
rect 570 -1228 572 -1160
rect 580 -1228 582 -1160
rect 596 -1228 598 -1160
rect 604 -1228 606 -1160
rect 620 -1228 622 -1160
rect 628 -1228 630 -1160
rect 638 -1228 640 -1160
rect 646 -1228 648 -1160
rect 662 -1228 664 -1160
rect 670 -1193 672 -1160
rect 680 -1193 682 -1160
rect 670 -1195 682 -1193
rect 670 -1228 672 -1195
rect 680 -1228 682 -1195
rect 688 -1228 690 -1160
rect 704 -1228 706 -1160
rect 712 -1228 714 -1160
rect 722 -1228 724 -1160
rect 730 -1228 732 -1160
rect 746 -1228 748 -1160
rect 754 -1228 756 -1160
rect 968 -1228 970 -1160
rect 978 -1228 980 -1160
rect 994 -1228 996 -1160
rect 1002 -1228 1004 -1160
rect 1018 -1228 1020 -1160
rect 1026 -1228 1028 -1160
rect 1036 -1228 1038 -1160
rect 1044 -1228 1046 -1160
rect 1060 -1228 1062 -1160
rect 1068 -1193 1070 -1160
rect 1078 -1193 1080 -1160
rect 1068 -1195 1080 -1193
rect 1068 -1228 1070 -1195
rect 1078 -1228 1080 -1195
rect 1086 -1228 1088 -1160
rect 1102 -1228 1104 -1160
rect 1110 -1228 1112 -1160
rect 1120 -1228 1122 -1160
rect 1128 -1228 1130 -1160
rect 1144 -1228 1146 -1160
rect 1152 -1228 1154 -1160
rect -1255 -1234 -1253 -1232
rect -1245 -1234 -1243 -1232
rect -1229 -1234 -1227 -1232
rect -1221 -1234 -1219 -1232
rect -1205 -1234 -1203 -1232
rect -1197 -1234 -1195 -1232
rect -1187 -1234 -1185 -1232
rect -1179 -1234 -1177 -1232
rect -1163 -1234 -1161 -1232
rect -1155 -1234 -1153 -1232
rect -1145 -1234 -1143 -1232
rect -1137 -1234 -1135 -1232
rect -1121 -1234 -1119 -1232
rect -1113 -1234 -1111 -1232
rect -1103 -1234 -1101 -1232
rect -1095 -1234 -1093 -1232
rect -1079 -1234 -1077 -1232
rect -1071 -1234 -1069 -1232
rect -930 -1234 -928 -1232
rect -920 -1234 -918 -1232
rect -904 -1234 -902 -1232
rect -896 -1234 -894 -1232
rect -880 -1234 -878 -1232
rect -872 -1234 -870 -1232
rect -862 -1234 -860 -1232
rect -854 -1234 -852 -1232
rect -838 -1234 -836 -1232
rect -830 -1234 -828 -1232
rect -820 -1234 -818 -1232
rect -812 -1234 -810 -1232
rect -796 -1234 -794 -1232
rect -788 -1234 -786 -1232
rect -778 -1234 -776 -1232
rect -770 -1234 -768 -1232
rect -754 -1234 -752 -1232
rect -746 -1234 -744 -1232
rect -572 -1234 -570 -1232
rect -562 -1234 -560 -1232
rect -546 -1234 -544 -1232
rect -538 -1234 -536 -1232
rect -522 -1234 -520 -1232
rect -514 -1234 -512 -1232
rect -504 -1234 -502 -1232
rect -496 -1234 -494 -1232
rect -480 -1234 -478 -1232
rect -472 -1234 -470 -1232
rect -462 -1234 -460 -1232
rect -454 -1234 -452 -1232
rect -438 -1234 -436 -1232
rect -430 -1234 -428 -1232
rect -420 -1234 -418 -1232
rect -412 -1234 -410 -1232
rect -396 -1234 -394 -1232
rect -388 -1234 -386 -1232
rect -214 -1234 -212 -1232
rect -204 -1234 -202 -1232
rect -188 -1234 -186 -1232
rect -180 -1234 -178 -1232
rect -164 -1234 -162 -1232
rect -156 -1234 -154 -1232
rect -146 -1234 -144 -1232
rect -138 -1234 -136 -1232
rect -122 -1234 -120 -1232
rect -114 -1234 -112 -1232
rect -104 -1234 -102 -1232
rect -96 -1234 -94 -1232
rect -80 -1234 -78 -1232
rect -72 -1234 -70 -1232
rect -62 -1234 -60 -1232
rect -54 -1234 -52 -1232
rect -38 -1234 -36 -1232
rect -30 -1234 -28 -1232
rect 214 -1234 216 -1232
rect 224 -1234 226 -1232
rect 240 -1234 242 -1232
rect 248 -1234 250 -1232
rect 264 -1234 266 -1232
rect 272 -1234 274 -1232
rect 282 -1234 284 -1232
rect 290 -1234 292 -1232
rect 306 -1234 308 -1232
rect 314 -1234 316 -1232
rect 324 -1234 326 -1232
rect 332 -1234 334 -1232
rect 348 -1234 350 -1232
rect 356 -1234 358 -1232
rect 366 -1234 368 -1232
rect 374 -1234 376 -1232
rect 390 -1234 392 -1232
rect 398 -1234 400 -1232
rect 570 -1234 572 -1232
rect 580 -1234 582 -1232
rect 596 -1234 598 -1232
rect 604 -1234 606 -1232
rect 620 -1234 622 -1232
rect 628 -1234 630 -1232
rect 638 -1234 640 -1232
rect 646 -1234 648 -1232
rect 662 -1234 664 -1232
rect 670 -1234 672 -1232
rect 680 -1234 682 -1232
rect 688 -1234 690 -1232
rect 704 -1234 706 -1232
rect 712 -1234 714 -1232
rect 722 -1234 724 -1232
rect 730 -1234 732 -1232
rect 746 -1234 748 -1232
rect 754 -1234 756 -1232
rect 968 -1234 970 -1232
rect 978 -1234 980 -1232
rect 994 -1234 996 -1232
rect 1002 -1234 1004 -1232
rect 1018 -1234 1020 -1232
rect 1026 -1234 1028 -1232
rect 1036 -1234 1038 -1232
rect 1044 -1234 1046 -1232
rect 1060 -1234 1062 -1232
rect 1068 -1234 1070 -1232
rect 1078 -1234 1080 -1232
rect 1086 -1234 1088 -1232
rect 1102 -1234 1104 -1232
rect 1110 -1234 1112 -1232
rect 1120 -1234 1122 -1232
rect 1128 -1234 1130 -1232
rect 1144 -1234 1146 -1232
rect 1152 -1234 1154 -1232
rect -1334 -1268 -1332 -1266
rect -1326 -1268 -1324 -1266
rect -1316 -1268 -1314 -1266
rect -930 -1268 -928 -1266
rect -922 -1268 -920 -1266
rect -912 -1268 -910 -1266
rect -572 -1268 -570 -1266
rect -564 -1268 -562 -1266
rect -554 -1268 -552 -1266
rect -214 -1268 -212 -1266
rect -206 -1268 -204 -1266
rect -196 -1268 -194 -1266
rect 214 -1268 216 -1266
rect 222 -1268 224 -1266
rect 232 -1268 234 -1266
rect 570 -1268 572 -1266
rect 578 -1268 580 -1266
rect 588 -1268 590 -1266
rect 968 -1268 970 -1266
rect 976 -1268 978 -1266
rect 986 -1268 988 -1266
rect 1326 -1268 1328 -1266
rect 1334 -1268 1336 -1266
rect 1344 -1268 1346 -1266
rect -1334 -1344 -1332 -1276
rect -1326 -1300 -1324 -1276
rect -1326 -1344 -1324 -1304
rect -1316 -1344 -1314 -1276
rect -930 -1344 -928 -1276
rect -922 -1300 -920 -1276
rect -922 -1344 -920 -1304
rect -912 -1344 -910 -1276
rect -572 -1344 -570 -1276
rect -564 -1300 -562 -1276
rect -564 -1344 -562 -1304
rect -554 -1344 -552 -1276
rect -214 -1344 -212 -1276
rect -206 -1300 -204 -1276
rect -206 -1344 -204 -1304
rect -196 -1344 -194 -1276
rect 214 -1344 216 -1276
rect 222 -1300 224 -1276
rect 222 -1344 224 -1304
rect 232 -1344 234 -1276
rect 570 -1344 572 -1276
rect 578 -1300 580 -1276
rect 578 -1344 580 -1304
rect 588 -1344 590 -1276
rect 968 -1344 970 -1276
rect 976 -1300 978 -1276
rect 976 -1344 978 -1304
rect 986 -1344 988 -1276
rect 1326 -1344 1328 -1276
rect 1334 -1300 1336 -1276
rect 1334 -1344 1336 -1304
rect 1344 -1344 1346 -1276
rect -1334 -1350 -1332 -1348
rect -1326 -1350 -1324 -1348
rect -1316 -1350 -1314 -1348
rect -930 -1350 -928 -1348
rect -922 -1350 -920 -1348
rect -912 -1350 -910 -1348
rect -572 -1350 -570 -1348
rect -564 -1350 -562 -1348
rect -554 -1350 -552 -1348
rect -214 -1350 -212 -1348
rect -206 -1350 -204 -1348
rect -196 -1350 -194 -1348
rect 214 -1350 216 -1348
rect 222 -1350 224 -1348
rect 232 -1350 234 -1348
rect 570 -1350 572 -1348
rect 578 -1350 580 -1348
rect 588 -1350 590 -1348
rect 968 -1350 970 -1348
rect 976 -1350 978 -1348
rect 986 -1350 988 -1348
rect 1326 -1350 1328 -1348
rect 1334 -1350 1336 -1348
rect 1344 -1350 1346 -1348
rect -1255 -1382 -1253 -1380
rect -1245 -1382 -1243 -1380
rect -1229 -1382 -1227 -1380
rect -1219 -1382 -1217 -1380
rect -1211 -1382 -1209 -1380
rect -1201 -1382 -1199 -1380
rect -1185 -1382 -1183 -1380
rect -1177 -1382 -1175 -1380
rect -1167 -1382 -1165 -1380
rect -930 -1382 -928 -1380
rect -920 -1382 -918 -1380
rect -904 -1382 -902 -1380
rect -894 -1382 -892 -1380
rect -878 -1382 -876 -1380
rect -868 -1382 -866 -1380
rect -860 -1382 -858 -1380
rect -850 -1382 -848 -1380
rect -834 -1382 -832 -1380
rect -826 -1382 -824 -1380
rect -816 -1382 -814 -1380
rect -800 -1382 -798 -1380
rect -790 -1382 -788 -1380
rect -782 -1382 -780 -1380
rect -772 -1382 -770 -1380
rect -756 -1382 -754 -1380
rect -748 -1382 -746 -1380
rect -732 -1382 -730 -1380
rect -716 -1382 -714 -1380
rect -708 -1382 -706 -1380
rect -698 -1382 -696 -1380
rect -572 -1382 -570 -1380
rect -562 -1382 -560 -1380
rect -546 -1382 -544 -1380
rect -536 -1382 -534 -1380
rect -520 -1382 -518 -1380
rect -510 -1382 -508 -1380
rect -502 -1382 -500 -1380
rect -492 -1382 -490 -1380
rect -476 -1382 -474 -1380
rect -468 -1382 -466 -1380
rect -458 -1382 -456 -1380
rect -442 -1382 -440 -1380
rect -432 -1382 -430 -1380
rect -424 -1382 -422 -1380
rect -414 -1382 -412 -1380
rect -398 -1382 -396 -1380
rect -390 -1382 -388 -1380
rect -374 -1382 -372 -1380
rect -358 -1382 -356 -1380
rect -350 -1382 -348 -1380
rect -340 -1382 -338 -1380
rect -214 -1382 -212 -1380
rect -204 -1382 -202 -1380
rect -188 -1382 -186 -1380
rect -178 -1382 -176 -1380
rect -162 -1382 -160 -1380
rect -152 -1382 -150 -1380
rect -144 -1382 -142 -1380
rect -134 -1382 -132 -1380
rect -118 -1382 -116 -1380
rect -110 -1382 -108 -1380
rect -100 -1382 -98 -1380
rect -84 -1382 -82 -1380
rect -74 -1382 -72 -1380
rect -66 -1382 -64 -1380
rect -56 -1382 -54 -1380
rect -40 -1382 -38 -1380
rect -32 -1382 -30 -1380
rect -16 -1382 -14 -1380
rect 0 -1382 2 -1380
rect 8 -1382 10 -1380
rect 18 -1382 20 -1380
rect 214 -1382 216 -1380
rect 224 -1382 226 -1380
rect 240 -1382 242 -1380
rect 250 -1382 252 -1380
rect 266 -1382 268 -1380
rect 276 -1382 278 -1380
rect 284 -1382 286 -1380
rect 294 -1382 296 -1380
rect 310 -1382 312 -1380
rect 318 -1382 320 -1380
rect 328 -1382 330 -1380
rect 344 -1382 346 -1380
rect 354 -1382 356 -1380
rect 362 -1382 364 -1380
rect 372 -1382 374 -1380
rect 388 -1382 390 -1380
rect 396 -1382 398 -1380
rect 412 -1382 414 -1380
rect 428 -1382 430 -1380
rect 436 -1382 438 -1380
rect 446 -1382 448 -1380
rect 570 -1382 572 -1380
rect 580 -1382 582 -1380
rect 596 -1382 598 -1380
rect 606 -1382 608 -1380
rect 622 -1382 624 -1380
rect 632 -1382 634 -1380
rect 640 -1382 642 -1380
rect 650 -1382 652 -1380
rect 666 -1382 668 -1380
rect 674 -1382 676 -1380
rect 684 -1382 686 -1380
rect 700 -1382 702 -1380
rect 710 -1382 712 -1380
rect 718 -1382 720 -1380
rect 728 -1382 730 -1380
rect 744 -1382 746 -1380
rect 752 -1382 754 -1380
rect 768 -1382 770 -1380
rect 784 -1382 786 -1380
rect 792 -1382 794 -1380
rect 802 -1382 804 -1380
rect 968 -1382 970 -1380
rect 978 -1382 980 -1380
rect 994 -1382 996 -1380
rect 1004 -1382 1006 -1380
rect 1020 -1382 1022 -1380
rect 1030 -1382 1032 -1380
rect 1038 -1382 1040 -1380
rect 1048 -1382 1050 -1380
rect 1064 -1382 1066 -1380
rect 1072 -1382 1074 -1380
rect 1082 -1382 1084 -1380
rect 1098 -1382 1100 -1380
rect 1108 -1382 1110 -1380
rect 1116 -1382 1118 -1380
rect 1126 -1382 1128 -1380
rect 1142 -1382 1144 -1380
rect 1150 -1382 1152 -1380
rect 1166 -1382 1168 -1380
rect 1182 -1382 1184 -1380
rect 1190 -1382 1192 -1380
rect 1200 -1382 1202 -1380
rect 1326 -1382 1328 -1380
rect 1336 -1382 1338 -1380
rect 1352 -1382 1354 -1380
rect 1362 -1382 1364 -1380
rect 1370 -1382 1372 -1380
rect 1380 -1382 1382 -1380
rect 1396 -1382 1398 -1380
rect 1404 -1382 1406 -1380
rect 1414 -1382 1416 -1380
rect -1255 -1458 -1253 -1390
rect -1245 -1458 -1243 -1390
rect -1229 -1458 -1227 -1390
rect -1219 -1458 -1217 -1390
rect -1211 -1458 -1209 -1390
rect -1201 -1458 -1199 -1390
rect -1185 -1458 -1183 -1390
rect -1177 -1458 -1175 -1390
rect -1167 -1458 -1165 -1390
rect -930 -1458 -928 -1390
rect -920 -1458 -918 -1390
rect -904 -1458 -902 -1390
rect -894 -1458 -892 -1390
rect -878 -1458 -876 -1390
rect -868 -1458 -866 -1390
rect -860 -1458 -858 -1390
rect -850 -1458 -848 -1390
rect -834 -1458 -832 -1390
rect -826 -1458 -824 -1390
rect -816 -1458 -814 -1390
rect -800 -1458 -798 -1390
rect -790 -1458 -788 -1390
rect -782 -1458 -780 -1390
rect -772 -1458 -770 -1390
rect -756 -1458 -754 -1390
rect -748 -1458 -746 -1390
rect -732 -1458 -730 -1390
rect -716 -1458 -714 -1390
rect -708 -1458 -706 -1390
rect -698 -1458 -696 -1390
rect -572 -1458 -570 -1390
rect -562 -1458 -560 -1390
rect -546 -1458 -544 -1390
rect -536 -1458 -534 -1390
rect -520 -1458 -518 -1390
rect -510 -1458 -508 -1390
rect -502 -1458 -500 -1390
rect -492 -1458 -490 -1390
rect -476 -1458 -474 -1390
rect -468 -1458 -466 -1390
rect -458 -1458 -456 -1390
rect -442 -1458 -440 -1390
rect -432 -1458 -430 -1390
rect -424 -1458 -422 -1390
rect -414 -1458 -412 -1390
rect -398 -1458 -396 -1390
rect -390 -1458 -388 -1390
rect -374 -1458 -372 -1390
rect -358 -1458 -356 -1390
rect -350 -1458 -348 -1390
rect -340 -1458 -338 -1390
rect -214 -1458 -212 -1390
rect -204 -1458 -202 -1390
rect -188 -1458 -186 -1390
rect -178 -1458 -176 -1390
rect -162 -1458 -160 -1390
rect -152 -1458 -150 -1390
rect -144 -1458 -142 -1390
rect -134 -1458 -132 -1390
rect -118 -1458 -116 -1390
rect -110 -1458 -108 -1390
rect -100 -1458 -98 -1390
rect -84 -1458 -82 -1390
rect -74 -1458 -72 -1390
rect -66 -1458 -64 -1390
rect -56 -1458 -54 -1390
rect -40 -1458 -38 -1390
rect -32 -1458 -30 -1390
rect -16 -1458 -14 -1390
rect 0 -1458 2 -1390
rect 8 -1458 10 -1390
rect 18 -1458 20 -1390
rect 214 -1458 216 -1390
rect 224 -1458 226 -1390
rect 240 -1458 242 -1390
rect 250 -1458 252 -1390
rect 266 -1458 268 -1390
rect 276 -1458 278 -1390
rect 284 -1458 286 -1390
rect 294 -1458 296 -1390
rect 310 -1458 312 -1390
rect 318 -1458 320 -1390
rect 328 -1458 330 -1390
rect 344 -1458 346 -1390
rect 354 -1458 356 -1390
rect 362 -1458 364 -1390
rect 372 -1458 374 -1390
rect 388 -1458 390 -1390
rect 396 -1458 398 -1390
rect 412 -1458 414 -1390
rect 428 -1458 430 -1390
rect 436 -1458 438 -1390
rect 446 -1458 448 -1390
rect 570 -1458 572 -1390
rect 580 -1458 582 -1390
rect 596 -1458 598 -1390
rect 606 -1458 608 -1390
rect 622 -1458 624 -1390
rect 632 -1458 634 -1390
rect 640 -1458 642 -1390
rect 650 -1458 652 -1390
rect 666 -1458 668 -1390
rect 674 -1458 676 -1390
rect 684 -1458 686 -1390
rect 700 -1458 702 -1390
rect 710 -1458 712 -1390
rect 718 -1458 720 -1390
rect 728 -1458 730 -1390
rect 744 -1458 746 -1390
rect 752 -1458 754 -1390
rect 768 -1458 770 -1390
rect 784 -1458 786 -1390
rect 792 -1458 794 -1390
rect 802 -1458 804 -1390
rect 968 -1458 970 -1390
rect 978 -1458 980 -1390
rect 994 -1458 996 -1390
rect 1004 -1458 1006 -1390
rect 1020 -1458 1022 -1390
rect 1030 -1458 1032 -1390
rect 1038 -1458 1040 -1390
rect 1048 -1458 1050 -1390
rect 1064 -1458 1066 -1390
rect 1072 -1458 1074 -1390
rect 1082 -1458 1084 -1390
rect 1098 -1458 1100 -1390
rect 1108 -1458 1110 -1390
rect 1116 -1458 1118 -1390
rect 1126 -1458 1128 -1390
rect 1142 -1458 1144 -1390
rect 1150 -1458 1152 -1390
rect 1166 -1458 1168 -1390
rect 1182 -1458 1184 -1390
rect 1190 -1458 1192 -1390
rect 1200 -1458 1202 -1390
rect 1326 -1458 1328 -1390
rect 1336 -1458 1338 -1390
rect 1352 -1458 1354 -1390
rect 1362 -1458 1364 -1390
rect 1370 -1458 1372 -1390
rect 1380 -1458 1382 -1390
rect 1396 -1458 1398 -1390
rect 1404 -1458 1406 -1390
rect 1414 -1458 1416 -1390
rect -1255 -1464 -1253 -1462
rect -1245 -1464 -1243 -1462
rect -1229 -1464 -1227 -1462
rect -1219 -1464 -1217 -1462
rect -1211 -1464 -1209 -1462
rect -1201 -1464 -1199 -1462
rect -1185 -1464 -1183 -1462
rect -1177 -1464 -1175 -1462
rect -1167 -1464 -1165 -1462
rect -930 -1464 -928 -1462
rect -920 -1464 -918 -1462
rect -904 -1464 -902 -1462
rect -894 -1464 -892 -1462
rect -878 -1464 -876 -1462
rect -868 -1464 -866 -1462
rect -860 -1464 -858 -1462
rect -850 -1464 -848 -1462
rect -834 -1464 -832 -1462
rect -826 -1464 -824 -1462
rect -816 -1464 -814 -1462
rect -800 -1464 -798 -1462
rect -790 -1464 -788 -1462
rect -782 -1464 -780 -1462
rect -772 -1464 -770 -1462
rect -756 -1464 -754 -1462
rect -748 -1464 -746 -1462
rect -732 -1464 -730 -1462
rect -716 -1464 -714 -1462
rect -708 -1464 -706 -1462
rect -698 -1464 -696 -1462
rect -572 -1464 -570 -1462
rect -562 -1464 -560 -1462
rect -546 -1464 -544 -1462
rect -536 -1464 -534 -1462
rect -520 -1464 -518 -1462
rect -510 -1464 -508 -1462
rect -502 -1464 -500 -1462
rect -492 -1464 -490 -1462
rect -476 -1464 -474 -1462
rect -468 -1464 -466 -1462
rect -458 -1464 -456 -1462
rect -442 -1464 -440 -1462
rect -432 -1464 -430 -1462
rect -424 -1464 -422 -1462
rect -414 -1464 -412 -1462
rect -398 -1464 -396 -1462
rect -390 -1464 -388 -1462
rect -374 -1464 -372 -1462
rect -358 -1464 -356 -1462
rect -350 -1464 -348 -1462
rect -340 -1464 -338 -1462
rect -214 -1464 -212 -1462
rect -204 -1464 -202 -1462
rect -188 -1464 -186 -1462
rect -178 -1464 -176 -1462
rect -162 -1464 -160 -1462
rect -152 -1464 -150 -1462
rect -144 -1464 -142 -1462
rect -134 -1464 -132 -1462
rect -118 -1464 -116 -1462
rect -110 -1464 -108 -1462
rect -100 -1464 -98 -1462
rect -84 -1464 -82 -1462
rect -74 -1464 -72 -1462
rect -66 -1464 -64 -1462
rect -56 -1464 -54 -1462
rect -40 -1464 -38 -1462
rect -32 -1464 -30 -1462
rect -16 -1464 -14 -1462
rect 0 -1464 2 -1462
rect 8 -1464 10 -1462
rect 18 -1464 20 -1462
rect 214 -1464 216 -1462
rect 224 -1464 226 -1462
rect 240 -1464 242 -1462
rect 250 -1464 252 -1462
rect 266 -1464 268 -1462
rect 276 -1464 278 -1462
rect 284 -1464 286 -1462
rect 294 -1464 296 -1462
rect 310 -1464 312 -1462
rect 318 -1464 320 -1462
rect 328 -1464 330 -1462
rect 344 -1464 346 -1462
rect 354 -1464 356 -1462
rect 362 -1464 364 -1462
rect 372 -1464 374 -1462
rect 388 -1464 390 -1462
rect 396 -1464 398 -1462
rect 412 -1464 414 -1462
rect 428 -1464 430 -1462
rect 436 -1464 438 -1462
rect 446 -1464 448 -1462
rect 570 -1464 572 -1462
rect 580 -1464 582 -1462
rect 596 -1464 598 -1462
rect 606 -1464 608 -1462
rect 622 -1464 624 -1462
rect 632 -1464 634 -1462
rect 640 -1464 642 -1462
rect 650 -1464 652 -1462
rect 666 -1464 668 -1462
rect 674 -1464 676 -1462
rect 684 -1464 686 -1462
rect 700 -1464 702 -1462
rect 710 -1464 712 -1462
rect 718 -1464 720 -1462
rect 728 -1464 730 -1462
rect 744 -1464 746 -1462
rect 752 -1464 754 -1462
rect 768 -1464 770 -1462
rect 784 -1464 786 -1462
rect 792 -1464 794 -1462
rect 802 -1464 804 -1462
rect 968 -1464 970 -1462
rect 978 -1464 980 -1462
rect 994 -1464 996 -1462
rect 1004 -1464 1006 -1462
rect 1020 -1464 1022 -1462
rect 1030 -1464 1032 -1462
rect 1038 -1464 1040 -1462
rect 1048 -1464 1050 -1462
rect 1064 -1464 1066 -1462
rect 1072 -1464 1074 -1462
rect 1082 -1464 1084 -1462
rect 1098 -1464 1100 -1462
rect 1108 -1464 1110 -1462
rect 1116 -1464 1118 -1462
rect 1126 -1464 1128 -1462
rect 1142 -1464 1144 -1462
rect 1150 -1464 1152 -1462
rect 1166 -1464 1168 -1462
rect 1182 -1464 1184 -1462
rect 1190 -1464 1192 -1462
rect 1200 -1464 1202 -1462
rect 1326 -1464 1328 -1462
rect 1336 -1464 1338 -1462
rect 1352 -1464 1354 -1462
rect 1362 -1464 1364 -1462
rect 1370 -1464 1372 -1462
rect 1380 -1464 1382 -1462
rect 1396 -1464 1398 -1462
rect 1404 -1464 1406 -1462
rect 1414 -1464 1416 -1462
rect -1255 -1505 -1253 -1503
rect -1245 -1505 -1243 -1503
rect -1229 -1505 -1227 -1503
rect -1221 -1505 -1219 -1503
rect -1205 -1505 -1203 -1503
rect -1197 -1505 -1195 -1503
rect -1187 -1505 -1185 -1503
rect -1179 -1505 -1177 -1503
rect -1163 -1505 -1161 -1503
rect -1155 -1505 -1153 -1503
rect -1145 -1505 -1143 -1503
rect -1137 -1505 -1135 -1503
rect -1121 -1505 -1119 -1503
rect -1113 -1505 -1111 -1503
rect -1103 -1505 -1101 -1503
rect -1095 -1505 -1093 -1503
rect -1079 -1505 -1077 -1503
rect -1071 -1505 -1069 -1503
rect -930 -1505 -928 -1503
rect -920 -1505 -918 -1503
rect -904 -1505 -902 -1503
rect -896 -1505 -894 -1503
rect -880 -1505 -878 -1503
rect -872 -1505 -870 -1503
rect -862 -1505 -860 -1503
rect -854 -1505 -852 -1503
rect -838 -1505 -836 -1503
rect -830 -1505 -828 -1503
rect -820 -1505 -818 -1503
rect -812 -1505 -810 -1503
rect -796 -1505 -794 -1503
rect -788 -1505 -786 -1503
rect -778 -1505 -776 -1503
rect -770 -1505 -768 -1503
rect -754 -1505 -752 -1503
rect -746 -1505 -744 -1503
rect -572 -1505 -570 -1503
rect -562 -1505 -560 -1503
rect -546 -1505 -544 -1503
rect -538 -1505 -536 -1503
rect -522 -1505 -520 -1503
rect -514 -1505 -512 -1503
rect -504 -1505 -502 -1503
rect -496 -1505 -494 -1503
rect -480 -1505 -478 -1503
rect -472 -1505 -470 -1503
rect -462 -1505 -460 -1503
rect -454 -1505 -452 -1503
rect -438 -1505 -436 -1503
rect -430 -1505 -428 -1503
rect -420 -1505 -418 -1503
rect -412 -1505 -410 -1503
rect -396 -1505 -394 -1503
rect -388 -1505 -386 -1503
rect -214 -1505 -212 -1503
rect -204 -1505 -202 -1503
rect -188 -1505 -186 -1503
rect -180 -1505 -178 -1503
rect -164 -1505 -162 -1503
rect -156 -1505 -154 -1503
rect -146 -1505 -144 -1503
rect -138 -1505 -136 -1503
rect -122 -1505 -120 -1503
rect -114 -1505 -112 -1503
rect -104 -1505 -102 -1503
rect -96 -1505 -94 -1503
rect -80 -1505 -78 -1503
rect -72 -1505 -70 -1503
rect -62 -1505 -60 -1503
rect -54 -1505 -52 -1503
rect -38 -1505 -36 -1503
rect -30 -1505 -28 -1503
rect 214 -1505 216 -1503
rect 224 -1505 226 -1503
rect 240 -1505 242 -1503
rect 248 -1505 250 -1503
rect 264 -1505 266 -1503
rect 272 -1505 274 -1503
rect 282 -1505 284 -1503
rect 290 -1505 292 -1503
rect 306 -1505 308 -1503
rect 314 -1505 316 -1503
rect 324 -1505 326 -1503
rect 332 -1505 334 -1503
rect 348 -1505 350 -1503
rect 356 -1505 358 -1503
rect 366 -1505 368 -1503
rect 374 -1505 376 -1503
rect 390 -1505 392 -1503
rect 398 -1505 400 -1503
rect 570 -1505 572 -1503
rect 580 -1505 582 -1503
rect 596 -1505 598 -1503
rect 604 -1505 606 -1503
rect 620 -1505 622 -1503
rect 628 -1505 630 -1503
rect 638 -1505 640 -1503
rect 646 -1505 648 -1503
rect 662 -1505 664 -1503
rect 670 -1505 672 -1503
rect 680 -1505 682 -1503
rect 688 -1505 690 -1503
rect 704 -1505 706 -1503
rect 712 -1505 714 -1503
rect 722 -1505 724 -1503
rect 730 -1505 732 -1503
rect 746 -1505 748 -1503
rect 754 -1505 756 -1503
rect 968 -1505 970 -1503
rect 978 -1505 980 -1503
rect 994 -1505 996 -1503
rect 1002 -1505 1004 -1503
rect 1018 -1505 1020 -1503
rect 1026 -1505 1028 -1503
rect 1036 -1505 1038 -1503
rect 1044 -1505 1046 -1503
rect 1060 -1505 1062 -1503
rect 1068 -1505 1070 -1503
rect 1078 -1505 1080 -1503
rect 1086 -1505 1088 -1503
rect 1102 -1505 1104 -1503
rect 1110 -1505 1112 -1503
rect 1120 -1505 1122 -1503
rect 1128 -1505 1130 -1503
rect 1144 -1505 1146 -1503
rect 1152 -1505 1154 -1503
rect -1255 -1581 -1253 -1513
rect -1245 -1581 -1243 -1513
rect -1229 -1581 -1227 -1513
rect -1221 -1581 -1219 -1513
rect -1205 -1581 -1203 -1513
rect -1197 -1581 -1195 -1513
rect -1187 -1581 -1185 -1513
rect -1179 -1581 -1177 -1513
rect -1163 -1581 -1161 -1513
rect -1155 -1546 -1153 -1513
rect -1145 -1546 -1143 -1513
rect -1155 -1548 -1143 -1546
rect -1155 -1581 -1153 -1548
rect -1145 -1581 -1143 -1548
rect -1137 -1581 -1135 -1513
rect -1121 -1581 -1119 -1513
rect -1113 -1581 -1111 -1513
rect -1103 -1581 -1101 -1513
rect -1095 -1581 -1093 -1513
rect -1079 -1581 -1077 -1513
rect -1071 -1581 -1069 -1513
rect -930 -1581 -928 -1513
rect -920 -1581 -918 -1513
rect -904 -1581 -902 -1513
rect -896 -1581 -894 -1513
rect -880 -1581 -878 -1513
rect -872 -1581 -870 -1513
rect -862 -1581 -860 -1513
rect -854 -1581 -852 -1513
rect -838 -1581 -836 -1513
rect -830 -1546 -828 -1513
rect -820 -1546 -818 -1513
rect -830 -1548 -818 -1546
rect -830 -1581 -828 -1548
rect -820 -1581 -818 -1548
rect -812 -1581 -810 -1513
rect -796 -1581 -794 -1513
rect -788 -1581 -786 -1513
rect -778 -1581 -776 -1513
rect -770 -1581 -768 -1513
rect -754 -1581 -752 -1513
rect -746 -1581 -744 -1513
rect -572 -1581 -570 -1513
rect -562 -1581 -560 -1513
rect -546 -1581 -544 -1513
rect -538 -1581 -536 -1513
rect -522 -1581 -520 -1513
rect -514 -1581 -512 -1513
rect -504 -1581 -502 -1513
rect -496 -1581 -494 -1513
rect -480 -1581 -478 -1513
rect -472 -1546 -470 -1513
rect -462 -1546 -460 -1513
rect -472 -1548 -460 -1546
rect -472 -1581 -470 -1548
rect -462 -1581 -460 -1548
rect -454 -1581 -452 -1513
rect -438 -1581 -436 -1513
rect -430 -1581 -428 -1513
rect -420 -1581 -418 -1513
rect -412 -1581 -410 -1513
rect -396 -1581 -394 -1513
rect -388 -1581 -386 -1513
rect -214 -1581 -212 -1513
rect -204 -1581 -202 -1513
rect -188 -1581 -186 -1513
rect -180 -1581 -178 -1513
rect -164 -1581 -162 -1513
rect -156 -1581 -154 -1513
rect -146 -1581 -144 -1513
rect -138 -1581 -136 -1513
rect -122 -1581 -120 -1513
rect -114 -1546 -112 -1513
rect -104 -1546 -102 -1513
rect -114 -1548 -102 -1546
rect -114 -1581 -112 -1548
rect -104 -1581 -102 -1548
rect -96 -1581 -94 -1513
rect -80 -1581 -78 -1513
rect -72 -1581 -70 -1513
rect -62 -1581 -60 -1513
rect -54 -1581 -52 -1513
rect -38 -1581 -36 -1513
rect -30 -1581 -28 -1513
rect 214 -1581 216 -1513
rect 224 -1581 226 -1513
rect 240 -1581 242 -1513
rect 248 -1581 250 -1513
rect 264 -1581 266 -1513
rect 272 -1581 274 -1513
rect 282 -1581 284 -1513
rect 290 -1581 292 -1513
rect 306 -1581 308 -1513
rect 314 -1546 316 -1513
rect 324 -1546 326 -1513
rect 314 -1548 326 -1546
rect 314 -1581 316 -1548
rect 324 -1581 326 -1548
rect 332 -1581 334 -1513
rect 348 -1581 350 -1513
rect 356 -1581 358 -1513
rect 366 -1581 368 -1513
rect 374 -1581 376 -1513
rect 390 -1581 392 -1513
rect 398 -1581 400 -1513
rect 570 -1581 572 -1513
rect 580 -1581 582 -1513
rect 596 -1581 598 -1513
rect 604 -1581 606 -1513
rect 620 -1581 622 -1513
rect 628 -1581 630 -1513
rect 638 -1581 640 -1513
rect 646 -1581 648 -1513
rect 662 -1581 664 -1513
rect 670 -1546 672 -1513
rect 680 -1546 682 -1513
rect 670 -1548 682 -1546
rect 670 -1581 672 -1548
rect 680 -1581 682 -1548
rect 688 -1581 690 -1513
rect 704 -1581 706 -1513
rect 712 -1581 714 -1513
rect 722 -1581 724 -1513
rect 730 -1581 732 -1513
rect 746 -1581 748 -1513
rect 754 -1581 756 -1513
rect 968 -1581 970 -1513
rect 978 -1581 980 -1513
rect 994 -1581 996 -1513
rect 1002 -1581 1004 -1513
rect 1018 -1581 1020 -1513
rect 1026 -1581 1028 -1513
rect 1036 -1581 1038 -1513
rect 1044 -1581 1046 -1513
rect 1060 -1581 1062 -1513
rect 1068 -1546 1070 -1513
rect 1078 -1546 1080 -1513
rect 1068 -1548 1080 -1546
rect 1068 -1581 1070 -1548
rect 1078 -1581 1080 -1548
rect 1086 -1581 1088 -1513
rect 1102 -1581 1104 -1513
rect 1110 -1581 1112 -1513
rect 1120 -1581 1122 -1513
rect 1128 -1581 1130 -1513
rect 1144 -1581 1146 -1513
rect 1152 -1581 1154 -1513
rect -1255 -1587 -1253 -1585
rect -1245 -1587 -1243 -1585
rect -1229 -1587 -1227 -1585
rect -1221 -1587 -1219 -1585
rect -1205 -1587 -1203 -1585
rect -1197 -1587 -1195 -1585
rect -1187 -1587 -1185 -1585
rect -1179 -1587 -1177 -1585
rect -1163 -1587 -1161 -1585
rect -1155 -1587 -1153 -1585
rect -1145 -1587 -1143 -1585
rect -1137 -1587 -1135 -1585
rect -1121 -1587 -1119 -1585
rect -1113 -1587 -1111 -1585
rect -1103 -1587 -1101 -1585
rect -1095 -1587 -1093 -1585
rect -1079 -1587 -1077 -1585
rect -1071 -1587 -1069 -1585
rect -930 -1587 -928 -1585
rect -920 -1587 -918 -1585
rect -904 -1587 -902 -1585
rect -896 -1587 -894 -1585
rect -880 -1587 -878 -1585
rect -872 -1587 -870 -1585
rect -862 -1587 -860 -1585
rect -854 -1587 -852 -1585
rect -838 -1587 -836 -1585
rect -830 -1587 -828 -1585
rect -820 -1587 -818 -1585
rect -812 -1587 -810 -1585
rect -796 -1587 -794 -1585
rect -788 -1587 -786 -1585
rect -778 -1587 -776 -1585
rect -770 -1587 -768 -1585
rect -754 -1587 -752 -1585
rect -746 -1587 -744 -1585
rect -572 -1587 -570 -1585
rect -562 -1587 -560 -1585
rect -546 -1587 -544 -1585
rect -538 -1587 -536 -1585
rect -522 -1587 -520 -1585
rect -514 -1587 -512 -1585
rect -504 -1587 -502 -1585
rect -496 -1587 -494 -1585
rect -480 -1587 -478 -1585
rect -472 -1587 -470 -1585
rect -462 -1587 -460 -1585
rect -454 -1587 -452 -1585
rect -438 -1587 -436 -1585
rect -430 -1587 -428 -1585
rect -420 -1587 -418 -1585
rect -412 -1587 -410 -1585
rect -396 -1587 -394 -1585
rect -388 -1587 -386 -1585
rect -214 -1587 -212 -1585
rect -204 -1587 -202 -1585
rect -188 -1587 -186 -1585
rect -180 -1587 -178 -1585
rect -164 -1587 -162 -1585
rect -156 -1587 -154 -1585
rect -146 -1587 -144 -1585
rect -138 -1587 -136 -1585
rect -122 -1587 -120 -1585
rect -114 -1587 -112 -1585
rect -104 -1587 -102 -1585
rect -96 -1587 -94 -1585
rect -80 -1587 -78 -1585
rect -72 -1587 -70 -1585
rect -62 -1587 -60 -1585
rect -54 -1587 -52 -1585
rect -38 -1587 -36 -1585
rect -30 -1587 -28 -1585
rect 214 -1587 216 -1585
rect 224 -1587 226 -1585
rect 240 -1587 242 -1585
rect 248 -1587 250 -1585
rect 264 -1587 266 -1585
rect 272 -1587 274 -1585
rect 282 -1587 284 -1585
rect 290 -1587 292 -1585
rect 306 -1587 308 -1585
rect 314 -1587 316 -1585
rect 324 -1587 326 -1585
rect 332 -1587 334 -1585
rect 348 -1587 350 -1585
rect 356 -1587 358 -1585
rect 366 -1587 368 -1585
rect 374 -1587 376 -1585
rect 390 -1587 392 -1585
rect 398 -1587 400 -1585
rect 570 -1587 572 -1585
rect 580 -1587 582 -1585
rect 596 -1587 598 -1585
rect 604 -1587 606 -1585
rect 620 -1587 622 -1585
rect 628 -1587 630 -1585
rect 638 -1587 640 -1585
rect 646 -1587 648 -1585
rect 662 -1587 664 -1585
rect 670 -1587 672 -1585
rect 680 -1587 682 -1585
rect 688 -1587 690 -1585
rect 704 -1587 706 -1585
rect 712 -1587 714 -1585
rect 722 -1587 724 -1585
rect 730 -1587 732 -1585
rect 746 -1587 748 -1585
rect 754 -1587 756 -1585
rect 968 -1587 970 -1585
rect 978 -1587 980 -1585
rect 994 -1587 996 -1585
rect 1002 -1587 1004 -1585
rect 1018 -1587 1020 -1585
rect 1026 -1587 1028 -1585
rect 1036 -1587 1038 -1585
rect 1044 -1587 1046 -1585
rect 1060 -1587 1062 -1585
rect 1068 -1587 1070 -1585
rect 1078 -1587 1080 -1585
rect 1086 -1587 1088 -1585
rect 1102 -1587 1104 -1585
rect 1110 -1587 1112 -1585
rect 1120 -1587 1122 -1585
rect 1128 -1587 1130 -1585
rect 1144 -1587 1146 -1585
rect 1152 -1587 1154 -1585
rect -1255 -1626 -1253 -1624
rect -1245 -1626 -1243 -1624
rect -1229 -1626 -1227 -1624
rect -1221 -1626 -1219 -1624
rect -1205 -1626 -1203 -1624
rect -1197 -1626 -1195 -1624
rect -1187 -1626 -1185 -1624
rect -1179 -1626 -1177 -1624
rect -1163 -1626 -1161 -1624
rect -1155 -1626 -1153 -1624
rect -1145 -1626 -1143 -1624
rect -1137 -1626 -1135 -1624
rect -1121 -1626 -1119 -1624
rect -1113 -1626 -1111 -1624
rect -1103 -1626 -1101 -1624
rect -1095 -1626 -1093 -1624
rect -1079 -1626 -1077 -1624
rect -1071 -1626 -1069 -1624
rect -930 -1626 -928 -1624
rect -920 -1626 -918 -1624
rect -904 -1626 -902 -1624
rect -896 -1626 -894 -1624
rect -880 -1626 -878 -1624
rect -872 -1626 -870 -1624
rect -862 -1626 -860 -1624
rect -854 -1626 -852 -1624
rect -838 -1626 -836 -1624
rect -830 -1626 -828 -1624
rect -820 -1626 -818 -1624
rect -812 -1626 -810 -1624
rect -796 -1626 -794 -1624
rect -788 -1626 -786 -1624
rect -778 -1626 -776 -1624
rect -770 -1626 -768 -1624
rect -754 -1626 -752 -1624
rect -746 -1626 -744 -1624
rect -572 -1626 -570 -1624
rect -562 -1626 -560 -1624
rect -546 -1626 -544 -1624
rect -538 -1626 -536 -1624
rect -522 -1626 -520 -1624
rect -514 -1626 -512 -1624
rect -504 -1626 -502 -1624
rect -496 -1626 -494 -1624
rect -480 -1626 -478 -1624
rect -472 -1626 -470 -1624
rect -462 -1626 -460 -1624
rect -454 -1626 -452 -1624
rect -438 -1626 -436 -1624
rect -430 -1626 -428 -1624
rect -420 -1626 -418 -1624
rect -412 -1626 -410 -1624
rect -396 -1626 -394 -1624
rect -388 -1626 -386 -1624
rect -214 -1626 -212 -1624
rect -204 -1626 -202 -1624
rect -188 -1626 -186 -1624
rect -180 -1626 -178 -1624
rect -164 -1626 -162 -1624
rect -156 -1626 -154 -1624
rect -146 -1626 -144 -1624
rect -138 -1626 -136 -1624
rect -122 -1626 -120 -1624
rect -114 -1626 -112 -1624
rect -104 -1626 -102 -1624
rect -96 -1626 -94 -1624
rect -80 -1626 -78 -1624
rect -72 -1626 -70 -1624
rect -62 -1626 -60 -1624
rect -54 -1626 -52 -1624
rect -38 -1626 -36 -1624
rect -30 -1626 -28 -1624
rect 214 -1626 216 -1624
rect 224 -1626 226 -1624
rect 240 -1626 242 -1624
rect 248 -1626 250 -1624
rect 264 -1626 266 -1624
rect 272 -1626 274 -1624
rect 282 -1626 284 -1624
rect 290 -1626 292 -1624
rect 306 -1626 308 -1624
rect 314 -1626 316 -1624
rect 324 -1626 326 -1624
rect 332 -1626 334 -1624
rect 348 -1626 350 -1624
rect 356 -1626 358 -1624
rect 366 -1626 368 -1624
rect 374 -1626 376 -1624
rect 390 -1626 392 -1624
rect 398 -1626 400 -1624
rect 570 -1626 572 -1624
rect 580 -1626 582 -1624
rect 596 -1626 598 -1624
rect 604 -1626 606 -1624
rect 620 -1626 622 -1624
rect 628 -1626 630 -1624
rect 638 -1626 640 -1624
rect 646 -1626 648 -1624
rect 662 -1626 664 -1624
rect 670 -1626 672 -1624
rect 680 -1626 682 -1624
rect 688 -1626 690 -1624
rect 704 -1626 706 -1624
rect 712 -1626 714 -1624
rect 722 -1626 724 -1624
rect 730 -1626 732 -1624
rect 746 -1626 748 -1624
rect 754 -1626 756 -1624
rect 968 -1626 970 -1624
rect 978 -1626 980 -1624
rect 994 -1626 996 -1624
rect 1002 -1626 1004 -1624
rect 1018 -1626 1020 -1624
rect 1026 -1626 1028 -1624
rect 1036 -1626 1038 -1624
rect 1044 -1626 1046 -1624
rect 1060 -1626 1062 -1624
rect 1068 -1626 1070 -1624
rect 1078 -1626 1080 -1624
rect 1086 -1626 1088 -1624
rect 1102 -1626 1104 -1624
rect 1110 -1626 1112 -1624
rect 1120 -1626 1122 -1624
rect 1128 -1626 1130 -1624
rect 1144 -1626 1146 -1624
rect 1152 -1626 1154 -1624
rect 1326 -1626 1328 -1624
rect 1336 -1626 1338 -1624
rect 1352 -1626 1354 -1624
rect 1360 -1626 1362 -1624
rect 1376 -1626 1378 -1624
rect 1384 -1626 1386 -1624
rect 1394 -1626 1396 -1624
rect 1402 -1626 1404 -1624
rect 1418 -1626 1420 -1624
rect 1426 -1626 1428 -1624
rect 1436 -1626 1438 -1624
rect 1444 -1626 1446 -1624
rect 1460 -1626 1462 -1624
rect 1468 -1626 1470 -1624
rect 1478 -1626 1480 -1624
rect 1486 -1626 1488 -1624
rect 1502 -1626 1504 -1624
rect 1510 -1626 1512 -1624
rect -1255 -1702 -1253 -1634
rect -1245 -1702 -1243 -1634
rect -1229 -1702 -1227 -1634
rect -1221 -1702 -1219 -1634
rect -1205 -1702 -1203 -1634
rect -1197 -1702 -1195 -1634
rect -1187 -1702 -1185 -1634
rect -1179 -1702 -1177 -1634
rect -1163 -1702 -1161 -1634
rect -1155 -1667 -1153 -1634
rect -1145 -1667 -1143 -1634
rect -1155 -1669 -1143 -1667
rect -1155 -1702 -1153 -1669
rect -1145 -1702 -1143 -1669
rect -1137 -1702 -1135 -1634
rect -1121 -1702 -1119 -1634
rect -1113 -1702 -1111 -1634
rect -1103 -1702 -1101 -1634
rect -1095 -1702 -1093 -1634
rect -1079 -1702 -1077 -1634
rect -1071 -1702 -1069 -1634
rect -930 -1702 -928 -1634
rect -920 -1702 -918 -1634
rect -904 -1702 -902 -1634
rect -896 -1702 -894 -1634
rect -880 -1702 -878 -1634
rect -872 -1702 -870 -1634
rect -862 -1702 -860 -1634
rect -854 -1702 -852 -1634
rect -838 -1702 -836 -1634
rect -830 -1667 -828 -1634
rect -820 -1667 -818 -1634
rect -830 -1669 -818 -1667
rect -830 -1702 -828 -1669
rect -820 -1702 -818 -1669
rect -812 -1702 -810 -1634
rect -796 -1702 -794 -1634
rect -788 -1702 -786 -1634
rect -778 -1702 -776 -1634
rect -770 -1702 -768 -1634
rect -754 -1702 -752 -1634
rect -746 -1702 -744 -1634
rect -572 -1702 -570 -1634
rect -562 -1702 -560 -1634
rect -546 -1702 -544 -1634
rect -538 -1702 -536 -1634
rect -522 -1702 -520 -1634
rect -514 -1702 -512 -1634
rect -504 -1702 -502 -1634
rect -496 -1702 -494 -1634
rect -480 -1702 -478 -1634
rect -472 -1667 -470 -1634
rect -462 -1667 -460 -1634
rect -472 -1669 -460 -1667
rect -472 -1702 -470 -1669
rect -462 -1702 -460 -1669
rect -454 -1702 -452 -1634
rect -438 -1702 -436 -1634
rect -430 -1702 -428 -1634
rect -420 -1702 -418 -1634
rect -412 -1702 -410 -1634
rect -396 -1702 -394 -1634
rect -388 -1702 -386 -1634
rect -214 -1702 -212 -1634
rect -204 -1702 -202 -1634
rect -188 -1702 -186 -1634
rect -180 -1702 -178 -1634
rect -164 -1702 -162 -1634
rect -156 -1702 -154 -1634
rect -146 -1702 -144 -1634
rect -138 -1702 -136 -1634
rect -122 -1702 -120 -1634
rect -114 -1667 -112 -1634
rect -104 -1667 -102 -1634
rect -114 -1669 -102 -1667
rect -114 -1702 -112 -1669
rect -104 -1702 -102 -1669
rect -96 -1702 -94 -1634
rect -80 -1702 -78 -1634
rect -72 -1702 -70 -1634
rect -62 -1702 -60 -1634
rect -54 -1702 -52 -1634
rect -38 -1702 -36 -1634
rect -30 -1702 -28 -1634
rect 214 -1702 216 -1634
rect 224 -1702 226 -1634
rect 240 -1702 242 -1634
rect 248 -1702 250 -1634
rect 264 -1702 266 -1634
rect 272 -1702 274 -1634
rect 282 -1702 284 -1634
rect 290 -1702 292 -1634
rect 306 -1702 308 -1634
rect 314 -1667 316 -1634
rect 324 -1667 326 -1634
rect 314 -1669 326 -1667
rect 314 -1702 316 -1669
rect 324 -1702 326 -1669
rect 332 -1702 334 -1634
rect 348 -1702 350 -1634
rect 356 -1702 358 -1634
rect 366 -1702 368 -1634
rect 374 -1702 376 -1634
rect 390 -1702 392 -1634
rect 398 -1702 400 -1634
rect 570 -1702 572 -1634
rect 580 -1702 582 -1634
rect 596 -1702 598 -1634
rect 604 -1702 606 -1634
rect 620 -1702 622 -1634
rect 628 -1702 630 -1634
rect 638 -1702 640 -1634
rect 646 -1702 648 -1634
rect 662 -1702 664 -1634
rect 670 -1667 672 -1634
rect 680 -1667 682 -1634
rect 670 -1669 682 -1667
rect 670 -1702 672 -1669
rect 680 -1702 682 -1669
rect 688 -1702 690 -1634
rect 704 -1702 706 -1634
rect 712 -1702 714 -1634
rect 722 -1702 724 -1634
rect 730 -1702 732 -1634
rect 746 -1702 748 -1634
rect 754 -1702 756 -1634
rect 968 -1702 970 -1634
rect 978 -1702 980 -1634
rect 994 -1702 996 -1634
rect 1002 -1702 1004 -1634
rect 1018 -1702 1020 -1634
rect 1026 -1702 1028 -1634
rect 1036 -1702 1038 -1634
rect 1044 -1702 1046 -1634
rect 1060 -1702 1062 -1634
rect 1068 -1667 1070 -1634
rect 1078 -1667 1080 -1634
rect 1068 -1669 1080 -1667
rect 1068 -1702 1070 -1669
rect 1078 -1702 1080 -1669
rect 1086 -1702 1088 -1634
rect 1102 -1702 1104 -1634
rect 1110 -1702 1112 -1634
rect 1120 -1702 1122 -1634
rect 1128 -1702 1130 -1634
rect 1144 -1702 1146 -1634
rect 1152 -1702 1154 -1634
rect 1326 -1702 1328 -1634
rect 1336 -1702 1338 -1634
rect 1352 -1702 1354 -1634
rect 1360 -1702 1362 -1634
rect 1376 -1702 1378 -1634
rect 1384 -1702 1386 -1634
rect 1394 -1702 1396 -1634
rect 1402 -1702 1404 -1634
rect 1418 -1702 1420 -1634
rect 1426 -1667 1428 -1634
rect 1436 -1667 1438 -1634
rect 1426 -1669 1438 -1667
rect 1426 -1702 1428 -1669
rect 1436 -1702 1438 -1669
rect 1444 -1702 1446 -1634
rect 1460 -1702 1462 -1634
rect 1468 -1702 1470 -1634
rect 1478 -1702 1480 -1634
rect 1486 -1702 1488 -1634
rect 1502 -1702 1504 -1634
rect 1510 -1702 1512 -1634
rect -1255 -1708 -1253 -1706
rect -1245 -1708 -1243 -1706
rect -1229 -1708 -1227 -1706
rect -1221 -1708 -1219 -1706
rect -1205 -1708 -1203 -1706
rect -1197 -1708 -1195 -1706
rect -1187 -1708 -1185 -1706
rect -1179 -1708 -1177 -1706
rect -1163 -1708 -1161 -1706
rect -1155 -1708 -1153 -1706
rect -1145 -1708 -1143 -1706
rect -1137 -1708 -1135 -1706
rect -1121 -1708 -1119 -1706
rect -1113 -1708 -1111 -1706
rect -1103 -1708 -1101 -1706
rect -1095 -1708 -1093 -1706
rect -1079 -1708 -1077 -1706
rect -1071 -1708 -1069 -1706
rect -930 -1708 -928 -1706
rect -920 -1708 -918 -1706
rect -904 -1708 -902 -1706
rect -896 -1708 -894 -1706
rect -880 -1708 -878 -1706
rect -872 -1708 -870 -1706
rect -862 -1708 -860 -1706
rect -854 -1708 -852 -1706
rect -838 -1708 -836 -1706
rect -830 -1708 -828 -1706
rect -820 -1708 -818 -1706
rect -812 -1708 -810 -1706
rect -796 -1708 -794 -1706
rect -788 -1708 -786 -1706
rect -778 -1708 -776 -1706
rect -770 -1708 -768 -1706
rect -754 -1708 -752 -1706
rect -746 -1708 -744 -1706
rect -572 -1708 -570 -1706
rect -562 -1708 -560 -1706
rect -546 -1708 -544 -1706
rect -538 -1708 -536 -1706
rect -522 -1708 -520 -1706
rect -514 -1708 -512 -1706
rect -504 -1708 -502 -1706
rect -496 -1708 -494 -1706
rect -480 -1708 -478 -1706
rect -472 -1708 -470 -1706
rect -462 -1708 -460 -1706
rect -454 -1708 -452 -1706
rect -438 -1708 -436 -1706
rect -430 -1708 -428 -1706
rect -420 -1708 -418 -1706
rect -412 -1708 -410 -1706
rect -396 -1708 -394 -1706
rect -388 -1708 -386 -1706
rect -214 -1708 -212 -1706
rect -204 -1708 -202 -1706
rect -188 -1708 -186 -1706
rect -180 -1708 -178 -1706
rect -164 -1708 -162 -1706
rect -156 -1708 -154 -1706
rect -146 -1708 -144 -1706
rect -138 -1708 -136 -1706
rect -122 -1708 -120 -1706
rect -114 -1708 -112 -1706
rect -104 -1708 -102 -1706
rect -96 -1708 -94 -1706
rect -80 -1708 -78 -1706
rect -72 -1708 -70 -1706
rect -62 -1708 -60 -1706
rect -54 -1708 -52 -1706
rect -38 -1708 -36 -1706
rect -30 -1708 -28 -1706
rect 214 -1708 216 -1706
rect 224 -1708 226 -1706
rect 240 -1708 242 -1706
rect 248 -1708 250 -1706
rect 264 -1708 266 -1706
rect 272 -1708 274 -1706
rect 282 -1708 284 -1706
rect 290 -1708 292 -1706
rect 306 -1708 308 -1706
rect 314 -1708 316 -1706
rect 324 -1708 326 -1706
rect 332 -1708 334 -1706
rect 348 -1708 350 -1706
rect 356 -1708 358 -1706
rect 366 -1708 368 -1706
rect 374 -1708 376 -1706
rect 390 -1708 392 -1706
rect 398 -1708 400 -1706
rect 570 -1708 572 -1706
rect 580 -1708 582 -1706
rect 596 -1708 598 -1706
rect 604 -1708 606 -1706
rect 620 -1708 622 -1706
rect 628 -1708 630 -1706
rect 638 -1708 640 -1706
rect 646 -1708 648 -1706
rect 662 -1708 664 -1706
rect 670 -1708 672 -1706
rect 680 -1708 682 -1706
rect 688 -1708 690 -1706
rect 704 -1708 706 -1706
rect 712 -1708 714 -1706
rect 722 -1708 724 -1706
rect 730 -1708 732 -1706
rect 746 -1708 748 -1706
rect 754 -1708 756 -1706
rect 968 -1708 970 -1706
rect 978 -1708 980 -1706
rect 994 -1708 996 -1706
rect 1002 -1708 1004 -1706
rect 1018 -1708 1020 -1706
rect 1026 -1708 1028 -1706
rect 1036 -1708 1038 -1706
rect 1044 -1708 1046 -1706
rect 1060 -1708 1062 -1706
rect 1068 -1708 1070 -1706
rect 1078 -1708 1080 -1706
rect 1086 -1708 1088 -1706
rect 1102 -1708 1104 -1706
rect 1110 -1708 1112 -1706
rect 1120 -1708 1122 -1706
rect 1128 -1708 1130 -1706
rect 1144 -1708 1146 -1706
rect 1152 -1708 1154 -1706
rect 1326 -1708 1328 -1706
rect 1336 -1708 1338 -1706
rect 1352 -1708 1354 -1706
rect 1360 -1708 1362 -1706
rect 1376 -1708 1378 -1706
rect 1384 -1708 1386 -1706
rect 1394 -1708 1396 -1706
rect 1402 -1708 1404 -1706
rect 1418 -1708 1420 -1706
rect 1426 -1708 1428 -1706
rect 1436 -1708 1438 -1706
rect 1444 -1708 1446 -1706
rect 1460 -1708 1462 -1706
rect 1468 -1708 1470 -1706
rect 1478 -1708 1480 -1706
rect 1486 -1708 1488 -1706
rect 1502 -1708 1504 -1706
rect 1510 -1708 1512 -1706
rect -1255 -1747 -1253 -1745
rect -1245 -1747 -1243 -1745
rect -1229 -1747 -1227 -1745
rect -1221 -1747 -1219 -1745
rect -1205 -1747 -1203 -1745
rect -1197 -1747 -1195 -1745
rect -1187 -1747 -1185 -1745
rect -1179 -1747 -1177 -1745
rect -1163 -1747 -1161 -1745
rect -1155 -1747 -1153 -1745
rect -1145 -1747 -1143 -1745
rect -1137 -1747 -1135 -1745
rect -1121 -1747 -1119 -1745
rect -1113 -1747 -1111 -1745
rect -1103 -1747 -1101 -1745
rect -1095 -1747 -1093 -1745
rect -1079 -1747 -1077 -1745
rect -1071 -1747 -1069 -1745
rect -1024 -1747 -1022 -1745
rect -930 -1747 -928 -1745
rect -920 -1747 -918 -1745
rect -904 -1747 -902 -1745
rect -896 -1747 -894 -1745
rect -880 -1747 -878 -1745
rect -872 -1747 -870 -1745
rect -862 -1747 -860 -1745
rect -854 -1747 -852 -1745
rect -838 -1747 -836 -1745
rect -830 -1747 -828 -1745
rect -820 -1747 -818 -1745
rect -812 -1747 -810 -1745
rect -796 -1747 -794 -1745
rect -788 -1747 -786 -1745
rect -778 -1747 -776 -1745
rect -770 -1747 -768 -1745
rect -754 -1747 -752 -1745
rect -746 -1747 -744 -1745
rect -572 -1747 -570 -1745
rect -562 -1747 -560 -1745
rect -546 -1747 -544 -1745
rect -538 -1747 -536 -1745
rect -522 -1747 -520 -1745
rect -514 -1747 -512 -1745
rect -504 -1747 -502 -1745
rect -496 -1747 -494 -1745
rect -480 -1747 -478 -1745
rect -472 -1747 -470 -1745
rect -462 -1747 -460 -1745
rect -454 -1747 -452 -1745
rect -438 -1747 -436 -1745
rect -430 -1747 -428 -1745
rect -420 -1747 -418 -1745
rect -412 -1747 -410 -1745
rect -396 -1747 -394 -1745
rect -388 -1747 -386 -1745
rect -327 -1747 -325 -1745
rect -214 -1747 -212 -1745
rect -204 -1747 -202 -1745
rect -188 -1747 -186 -1745
rect -180 -1747 -178 -1745
rect -164 -1747 -162 -1745
rect -156 -1747 -154 -1745
rect -146 -1747 -144 -1745
rect -138 -1747 -136 -1745
rect -122 -1747 -120 -1745
rect -114 -1747 -112 -1745
rect -104 -1747 -102 -1745
rect -96 -1747 -94 -1745
rect -80 -1747 -78 -1745
rect -72 -1747 -70 -1745
rect -62 -1747 -60 -1745
rect -54 -1747 -52 -1745
rect -38 -1747 -36 -1745
rect -30 -1747 -28 -1745
rect 214 -1747 216 -1745
rect 224 -1747 226 -1745
rect 240 -1747 242 -1745
rect 248 -1747 250 -1745
rect 264 -1747 266 -1745
rect 272 -1747 274 -1745
rect 282 -1747 284 -1745
rect 290 -1747 292 -1745
rect 306 -1747 308 -1745
rect 314 -1747 316 -1745
rect 324 -1747 326 -1745
rect 332 -1747 334 -1745
rect 348 -1747 350 -1745
rect 356 -1747 358 -1745
rect 366 -1747 368 -1745
rect 374 -1747 376 -1745
rect 390 -1747 392 -1745
rect 398 -1747 400 -1745
rect 469 -1747 471 -1745
rect 570 -1747 572 -1745
rect 580 -1747 582 -1745
rect 596 -1747 598 -1745
rect 604 -1747 606 -1745
rect 620 -1747 622 -1745
rect 628 -1747 630 -1745
rect 638 -1747 640 -1745
rect 646 -1747 648 -1745
rect 662 -1747 664 -1745
rect 670 -1747 672 -1745
rect 680 -1747 682 -1745
rect 688 -1747 690 -1745
rect 704 -1747 706 -1745
rect 712 -1747 714 -1745
rect 722 -1747 724 -1745
rect 730 -1747 732 -1745
rect 746 -1747 748 -1745
rect 754 -1747 756 -1745
rect 968 -1747 970 -1745
rect 978 -1747 980 -1745
rect 994 -1747 996 -1745
rect 1002 -1747 1004 -1745
rect 1018 -1747 1020 -1745
rect 1026 -1747 1028 -1745
rect 1036 -1747 1038 -1745
rect 1044 -1747 1046 -1745
rect 1060 -1747 1062 -1745
rect 1068 -1747 1070 -1745
rect 1078 -1747 1080 -1745
rect 1086 -1747 1088 -1745
rect 1102 -1747 1104 -1745
rect 1110 -1747 1112 -1745
rect 1120 -1747 1122 -1745
rect 1128 -1747 1130 -1745
rect 1144 -1747 1146 -1745
rect 1152 -1747 1154 -1745
rect 1208 -1747 1210 -1745
rect 1326 -1747 1328 -1745
rect 1336 -1747 1338 -1745
rect 1352 -1747 1354 -1745
rect 1360 -1747 1362 -1745
rect 1376 -1747 1378 -1745
rect 1384 -1747 1386 -1745
rect 1394 -1747 1396 -1745
rect 1402 -1747 1404 -1745
rect 1418 -1747 1420 -1745
rect 1426 -1747 1428 -1745
rect 1436 -1747 1438 -1745
rect 1444 -1747 1446 -1745
rect 1460 -1747 1462 -1745
rect 1468 -1747 1470 -1745
rect 1478 -1747 1480 -1745
rect 1486 -1747 1488 -1745
rect 1502 -1747 1504 -1745
rect 1510 -1747 1512 -1745
rect -1255 -1823 -1253 -1755
rect -1245 -1823 -1243 -1755
rect -1229 -1823 -1227 -1755
rect -1221 -1823 -1219 -1755
rect -1205 -1823 -1203 -1755
rect -1197 -1823 -1195 -1755
rect -1187 -1823 -1185 -1755
rect -1179 -1823 -1177 -1755
rect -1163 -1823 -1161 -1755
rect -1155 -1788 -1153 -1755
rect -1145 -1788 -1143 -1755
rect -1155 -1790 -1143 -1788
rect -1155 -1823 -1153 -1790
rect -1145 -1823 -1143 -1790
rect -1137 -1823 -1135 -1755
rect -1121 -1823 -1119 -1755
rect -1113 -1823 -1111 -1755
rect -1103 -1823 -1101 -1755
rect -1095 -1823 -1093 -1755
rect -1079 -1823 -1077 -1755
rect -1071 -1823 -1069 -1755
rect -1024 -1823 -1022 -1755
rect -930 -1823 -928 -1755
rect -920 -1823 -918 -1755
rect -904 -1823 -902 -1755
rect -896 -1823 -894 -1755
rect -880 -1823 -878 -1755
rect -872 -1823 -870 -1755
rect -862 -1823 -860 -1755
rect -854 -1823 -852 -1755
rect -838 -1823 -836 -1755
rect -830 -1788 -828 -1755
rect -820 -1788 -818 -1755
rect -830 -1790 -818 -1788
rect -830 -1823 -828 -1790
rect -820 -1823 -818 -1790
rect -812 -1823 -810 -1755
rect -796 -1823 -794 -1755
rect -788 -1823 -786 -1755
rect -778 -1823 -776 -1755
rect -770 -1823 -768 -1755
rect -754 -1823 -752 -1755
rect -746 -1823 -744 -1755
rect -572 -1823 -570 -1755
rect -562 -1823 -560 -1755
rect -546 -1823 -544 -1755
rect -538 -1823 -536 -1755
rect -522 -1823 -520 -1755
rect -514 -1823 -512 -1755
rect -504 -1823 -502 -1755
rect -496 -1823 -494 -1755
rect -480 -1823 -478 -1755
rect -472 -1788 -470 -1755
rect -462 -1788 -460 -1755
rect -472 -1790 -460 -1788
rect -472 -1823 -470 -1790
rect -462 -1823 -460 -1790
rect -454 -1823 -452 -1755
rect -438 -1823 -436 -1755
rect -430 -1823 -428 -1755
rect -420 -1823 -418 -1755
rect -412 -1823 -410 -1755
rect -396 -1823 -394 -1755
rect -388 -1823 -386 -1755
rect -327 -1823 -325 -1755
rect -214 -1823 -212 -1755
rect -204 -1823 -202 -1755
rect -188 -1823 -186 -1755
rect -180 -1823 -178 -1755
rect -164 -1823 -162 -1755
rect -156 -1823 -154 -1755
rect -146 -1823 -144 -1755
rect -138 -1823 -136 -1755
rect -122 -1823 -120 -1755
rect -114 -1788 -112 -1755
rect -104 -1788 -102 -1755
rect -114 -1790 -102 -1788
rect -114 -1823 -112 -1790
rect -104 -1823 -102 -1790
rect -96 -1823 -94 -1755
rect -80 -1823 -78 -1755
rect -72 -1823 -70 -1755
rect -62 -1823 -60 -1755
rect -54 -1823 -52 -1755
rect -38 -1823 -36 -1755
rect -30 -1823 -28 -1755
rect 214 -1823 216 -1755
rect 224 -1823 226 -1755
rect 240 -1823 242 -1755
rect 248 -1823 250 -1755
rect 264 -1823 266 -1755
rect 272 -1823 274 -1755
rect 282 -1823 284 -1755
rect 290 -1823 292 -1755
rect 306 -1823 308 -1755
rect 314 -1788 316 -1755
rect 324 -1788 326 -1755
rect 314 -1790 326 -1788
rect 314 -1823 316 -1790
rect 324 -1823 326 -1790
rect 332 -1823 334 -1755
rect 348 -1823 350 -1755
rect 356 -1823 358 -1755
rect 366 -1823 368 -1755
rect 374 -1823 376 -1755
rect 390 -1823 392 -1755
rect 398 -1823 400 -1755
rect 469 -1823 471 -1755
rect 570 -1823 572 -1755
rect 580 -1823 582 -1755
rect 596 -1823 598 -1755
rect 604 -1823 606 -1755
rect 620 -1823 622 -1755
rect 628 -1823 630 -1755
rect 638 -1823 640 -1755
rect 646 -1823 648 -1755
rect 662 -1823 664 -1755
rect 670 -1788 672 -1755
rect 680 -1788 682 -1755
rect 670 -1790 682 -1788
rect 670 -1823 672 -1790
rect 680 -1823 682 -1790
rect 688 -1823 690 -1755
rect 704 -1823 706 -1755
rect 712 -1823 714 -1755
rect 722 -1823 724 -1755
rect 730 -1823 732 -1755
rect 746 -1823 748 -1755
rect 754 -1823 756 -1755
rect 968 -1823 970 -1755
rect 978 -1823 980 -1755
rect 994 -1823 996 -1755
rect 1002 -1823 1004 -1755
rect 1018 -1823 1020 -1755
rect 1026 -1823 1028 -1755
rect 1036 -1823 1038 -1755
rect 1044 -1823 1046 -1755
rect 1060 -1823 1062 -1755
rect 1068 -1788 1070 -1755
rect 1078 -1788 1080 -1755
rect 1068 -1790 1080 -1788
rect 1068 -1823 1070 -1790
rect 1078 -1823 1080 -1790
rect 1086 -1823 1088 -1755
rect 1102 -1823 1104 -1755
rect 1110 -1823 1112 -1755
rect 1120 -1823 1122 -1755
rect 1128 -1823 1130 -1755
rect 1144 -1823 1146 -1755
rect 1152 -1823 1154 -1755
rect 1208 -1823 1210 -1755
rect 1326 -1823 1328 -1755
rect 1336 -1823 1338 -1755
rect 1352 -1823 1354 -1755
rect 1360 -1823 1362 -1755
rect 1376 -1823 1378 -1755
rect 1384 -1823 1386 -1755
rect 1394 -1823 1396 -1755
rect 1402 -1823 1404 -1755
rect 1418 -1823 1420 -1755
rect 1426 -1788 1428 -1755
rect 1436 -1788 1438 -1755
rect 1426 -1790 1438 -1788
rect 1426 -1823 1428 -1790
rect 1436 -1823 1438 -1790
rect 1444 -1823 1446 -1755
rect 1460 -1823 1462 -1755
rect 1468 -1823 1470 -1755
rect 1478 -1823 1480 -1755
rect 1486 -1823 1488 -1755
rect 1502 -1823 1504 -1755
rect 1510 -1823 1512 -1755
rect -1255 -1829 -1253 -1827
rect -1245 -1829 -1243 -1827
rect -1229 -1829 -1227 -1827
rect -1221 -1829 -1219 -1827
rect -1205 -1829 -1203 -1827
rect -1197 -1829 -1195 -1827
rect -1187 -1829 -1185 -1827
rect -1179 -1829 -1177 -1827
rect -1163 -1829 -1161 -1827
rect -1155 -1829 -1153 -1827
rect -1145 -1829 -1143 -1827
rect -1137 -1829 -1135 -1827
rect -1121 -1829 -1119 -1827
rect -1113 -1829 -1111 -1827
rect -1103 -1829 -1101 -1827
rect -1095 -1829 -1093 -1827
rect -1079 -1829 -1077 -1827
rect -1071 -1829 -1069 -1827
rect -1024 -1829 -1022 -1827
rect -930 -1829 -928 -1827
rect -920 -1829 -918 -1827
rect -904 -1829 -902 -1827
rect -896 -1829 -894 -1827
rect -880 -1829 -878 -1827
rect -872 -1829 -870 -1827
rect -862 -1829 -860 -1827
rect -854 -1829 -852 -1827
rect -838 -1829 -836 -1827
rect -830 -1829 -828 -1827
rect -820 -1829 -818 -1827
rect -812 -1829 -810 -1827
rect -796 -1829 -794 -1827
rect -788 -1829 -786 -1827
rect -778 -1829 -776 -1827
rect -770 -1829 -768 -1827
rect -754 -1829 -752 -1827
rect -746 -1829 -744 -1827
rect -572 -1829 -570 -1827
rect -562 -1829 -560 -1827
rect -546 -1829 -544 -1827
rect -538 -1829 -536 -1827
rect -522 -1829 -520 -1827
rect -514 -1829 -512 -1827
rect -504 -1829 -502 -1827
rect -496 -1829 -494 -1827
rect -480 -1829 -478 -1827
rect -472 -1829 -470 -1827
rect -462 -1829 -460 -1827
rect -454 -1829 -452 -1827
rect -438 -1829 -436 -1827
rect -430 -1829 -428 -1827
rect -420 -1829 -418 -1827
rect -412 -1829 -410 -1827
rect -396 -1829 -394 -1827
rect -388 -1829 -386 -1827
rect -327 -1829 -325 -1827
rect -214 -1829 -212 -1827
rect -204 -1829 -202 -1827
rect -188 -1829 -186 -1827
rect -180 -1829 -178 -1827
rect -164 -1829 -162 -1827
rect -156 -1829 -154 -1827
rect -146 -1829 -144 -1827
rect -138 -1829 -136 -1827
rect -122 -1829 -120 -1827
rect -114 -1829 -112 -1827
rect -104 -1829 -102 -1827
rect -96 -1829 -94 -1827
rect -80 -1829 -78 -1827
rect -72 -1829 -70 -1827
rect -62 -1829 -60 -1827
rect -54 -1829 -52 -1827
rect -38 -1829 -36 -1827
rect -30 -1829 -28 -1827
rect 214 -1829 216 -1827
rect 224 -1829 226 -1827
rect 240 -1829 242 -1827
rect 248 -1829 250 -1827
rect 264 -1829 266 -1827
rect 272 -1829 274 -1827
rect 282 -1829 284 -1827
rect 290 -1829 292 -1827
rect 306 -1829 308 -1827
rect 314 -1829 316 -1827
rect 324 -1829 326 -1827
rect 332 -1829 334 -1827
rect 348 -1829 350 -1827
rect 356 -1829 358 -1827
rect 366 -1829 368 -1827
rect 374 -1829 376 -1827
rect 390 -1829 392 -1827
rect 398 -1829 400 -1827
rect 469 -1829 471 -1827
rect 570 -1829 572 -1827
rect 580 -1829 582 -1827
rect 596 -1829 598 -1827
rect 604 -1829 606 -1827
rect 620 -1829 622 -1827
rect 628 -1829 630 -1827
rect 638 -1829 640 -1827
rect 646 -1829 648 -1827
rect 662 -1829 664 -1827
rect 670 -1829 672 -1827
rect 680 -1829 682 -1827
rect 688 -1829 690 -1827
rect 704 -1829 706 -1827
rect 712 -1829 714 -1827
rect 722 -1829 724 -1827
rect 730 -1829 732 -1827
rect 746 -1829 748 -1827
rect 754 -1829 756 -1827
rect 968 -1829 970 -1827
rect 978 -1829 980 -1827
rect 994 -1829 996 -1827
rect 1002 -1829 1004 -1827
rect 1018 -1829 1020 -1827
rect 1026 -1829 1028 -1827
rect 1036 -1829 1038 -1827
rect 1044 -1829 1046 -1827
rect 1060 -1829 1062 -1827
rect 1068 -1829 1070 -1827
rect 1078 -1829 1080 -1827
rect 1086 -1829 1088 -1827
rect 1102 -1829 1104 -1827
rect 1110 -1829 1112 -1827
rect 1120 -1829 1122 -1827
rect 1128 -1829 1130 -1827
rect 1144 -1829 1146 -1827
rect 1152 -1829 1154 -1827
rect 1208 -1829 1210 -1827
rect 1326 -1829 1328 -1827
rect 1336 -1829 1338 -1827
rect 1352 -1829 1354 -1827
rect 1360 -1829 1362 -1827
rect 1376 -1829 1378 -1827
rect 1384 -1829 1386 -1827
rect 1394 -1829 1396 -1827
rect 1402 -1829 1404 -1827
rect 1418 -1829 1420 -1827
rect 1426 -1829 1428 -1827
rect 1436 -1829 1438 -1827
rect 1444 -1829 1446 -1827
rect 1460 -1829 1462 -1827
rect 1468 -1829 1470 -1827
rect 1478 -1829 1480 -1827
rect 1486 -1829 1488 -1827
rect 1502 -1829 1504 -1827
rect 1510 -1829 1512 -1827
rect -1255 -1862 -1253 -1860
rect -1245 -1862 -1243 -1860
rect -1229 -1862 -1227 -1860
rect -1221 -1862 -1219 -1860
rect -1205 -1862 -1203 -1860
rect -1197 -1862 -1195 -1860
rect -1187 -1862 -1185 -1860
rect -1179 -1862 -1177 -1860
rect -1163 -1862 -1161 -1860
rect -1155 -1862 -1153 -1860
rect -1145 -1862 -1143 -1860
rect -1137 -1862 -1135 -1860
rect -1121 -1862 -1119 -1860
rect -1113 -1862 -1111 -1860
rect -1103 -1862 -1101 -1860
rect -1095 -1862 -1093 -1860
rect -1079 -1862 -1077 -1860
rect -1071 -1862 -1069 -1860
rect -1024 -1862 -1022 -1860
rect -668 -1862 -666 -1860
rect -327 -1862 -325 -1860
rect 469 -1862 471 -1860
rect 846 -1862 848 -1860
rect 1208 -1862 1210 -1860
rect -1255 -1938 -1253 -1870
rect -1245 -1938 -1243 -1870
rect -1229 -1938 -1227 -1870
rect -1221 -1938 -1219 -1870
rect -1205 -1938 -1203 -1870
rect -1197 -1938 -1195 -1870
rect -1187 -1938 -1185 -1870
rect -1179 -1938 -1177 -1870
rect -1163 -1938 -1161 -1870
rect -1155 -1903 -1153 -1870
rect -1145 -1903 -1143 -1870
rect -1155 -1905 -1143 -1903
rect -1155 -1938 -1153 -1905
rect -1145 -1938 -1143 -1905
rect -1137 -1938 -1135 -1870
rect -1121 -1938 -1119 -1870
rect -1113 -1938 -1111 -1870
rect -1103 -1938 -1101 -1870
rect -1095 -1938 -1093 -1870
rect -1079 -1938 -1077 -1870
rect -1071 -1938 -1069 -1870
rect -1024 -1938 -1022 -1870
rect -668 -1934 -666 -1878
rect -327 -1938 -325 -1870
rect 469 -1938 471 -1870
rect 846 -1934 848 -1878
rect 1208 -1938 1210 -1870
rect -1255 -1944 -1253 -1942
rect -1245 -1944 -1243 -1942
rect -1229 -1944 -1227 -1942
rect -1221 -1944 -1219 -1942
rect -1205 -1944 -1203 -1942
rect -1197 -1944 -1195 -1942
rect -1187 -1944 -1185 -1942
rect -1179 -1944 -1177 -1942
rect -1163 -1944 -1161 -1942
rect -1155 -1944 -1153 -1942
rect -1145 -1944 -1143 -1942
rect -1137 -1944 -1135 -1942
rect -1121 -1944 -1119 -1942
rect -1113 -1944 -1111 -1942
rect -1103 -1944 -1101 -1942
rect -1095 -1944 -1093 -1942
rect -1079 -1944 -1077 -1942
rect -1071 -1944 -1069 -1942
rect -1024 -1944 -1022 -1942
rect -668 -1944 -666 -1942
rect -327 -1944 -325 -1942
rect 469 -1944 471 -1942
rect 846 -1944 848 -1942
rect 1208 -1944 1210 -1942
rect -1334 -1974 -1332 -1972
rect -1326 -1974 -1324 -1972
rect -1316 -1974 -1314 -1972
rect -930 -1974 -928 -1972
rect -922 -1974 -920 -1972
rect -912 -1974 -910 -1972
rect -572 -1974 -570 -1972
rect -564 -1974 -562 -1972
rect -554 -1974 -552 -1972
rect -214 -1974 -212 -1972
rect -206 -1974 -204 -1972
rect -196 -1974 -194 -1972
rect 214 -1974 216 -1972
rect 222 -1974 224 -1972
rect 232 -1974 234 -1972
rect 570 -1974 572 -1972
rect 578 -1974 580 -1972
rect 588 -1974 590 -1972
rect 968 -1974 970 -1972
rect 976 -1974 978 -1972
rect 986 -1974 988 -1972
rect 1326 -1974 1328 -1972
rect 1334 -1974 1336 -1972
rect 1344 -1974 1346 -1972
rect -1334 -2050 -1332 -1982
rect -1326 -2006 -1324 -1982
rect -1326 -2050 -1324 -2010
rect -1316 -2050 -1314 -1982
rect -930 -2050 -928 -1982
rect -922 -2006 -920 -1982
rect -922 -2050 -920 -2010
rect -912 -2050 -910 -1982
rect -572 -2050 -570 -1982
rect -564 -2006 -562 -1982
rect -564 -2050 -562 -2010
rect -554 -2050 -552 -1982
rect -214 -2050 -212 -1982
rect -206 -2006 -204 -1982
rect -206 -2050 -204 -2010
rect -196 -2050 -194 -1982
rect 214 -2050 216 -1982
rect 222 -2006 224 -1982
rect 222 -2050 224 -2010
rect 232 -2050 234 -1982
rect 570 -2050 572 -1982
rect 578 -2006 580 -1982
rect 578 -2050 580 -2010
rect 588 -2050 590 -1982
rect 968 -2050 970 -1982
rect 976 -2006 978 -1982
rect 976 -2050 978 -2010
rect 986 -2050 988 -1982
rect 1326 -2050 1328 -1982
rect 1334 -2006 1336 -1982
rect 1334 -2050 1336 -2010
rect 1344 -2050 1346 -1982
rect -1334 -2056 -1332 -2054
rect -1326 -2056 -1324 -2054
rect -1316 -2056 -1314 -2054
rect -930 -2056 -928 -2054
rect -922 -2056 -920 -2054
rect -912 -2056 -910 -2054
rect -572 -2056 -570 -2054
rect -564 -2056 -562 -2054
rect -554 -2056 -552 -2054
rect -214 -2056 -212 -2054
rect -206 -2056 -204 -2054
rect -196 -2056 -194 -2054
rect 214 -2056 216 -2054
rect 222 -2056 224 -2054
rect 232 -2056 234 -2054
rect 570 -2056 572 -2054
rect 578 -2056 580 -2054
rect 588 -2056 590 -2054
rect 968 -2056 970 -2054
rect 976 -2056 978 -2054
rect 986 -2056 988 -2054
rect 1326 -2056 1328 -2054
rect 1334 -2056 1336 -2054
rect 1344 -2056 1346 -2054
rect -1255 -2093 -1253 -2091
rect -1245 -2093 -1243 -2091
rect -1229 -2093 -1227 -2091
rect -1219 -2093 -1217 -2091
rect -1211 -2093 -1209 -2091
rect -1201 -2093 -1199 -2091
rect -1185 -2093 -1183 -2091
rect -1177 -2093 -1175 -2091
rect -1167 -2093 -1165 -2091
rect -930 -2093 -928 -2091
rect -920 -2093 -918 -2091
rect -904 -2093 -902 -2091
rect -894 -2093 -892 -2091
rect -878 -2093 -876 -2091
rect -868 -2093 -866 -2091
rect -860 -2093 -858 -2091
rect -850 -2093 -848 -2091
rect -834 -2093 -832 -2091
rect -826 -2093 -824 -2091
rect -816 -2093 -814 -2091
rect -800 -2093 -798 -2091
rect -790 -2093 -788 -2091
rect -782 -2093 -780 -2091
rect -772 -2093 -770 -2091
rect -756 -2093 -754 -2091
rect -748 -2093 -746 -2091
rect -732 -2093 -730 -2091
rect -716 -2093 -714 -2091
rect -708 -2093 -706 -2091
rect -698 -2093 -696 -2091
rect -572 -2093 -570 -2091
rect -562 -2093 -560 -2091
rect -546 -2093 -544 -2091
rect -536 -2093 -534 -2091
rect -520 -2093 -518 -2091
rect -510 -2093 -508 -2091
rect -502 -2093 -500 -2091
rect -492 -2093 -490 -2091
rect -476 -2093 -474 -2091
rect -468 -2093 -466 -2091
rect -458 -2093 -456 -2091
rect -442 -2093 -440 -2091
rect -432 -2093 -430 -2091
rect -424 -2093 -422 -2091
rect -414 -2093 -412 -2091
rect -398 -2093 -396 -2091
rect -390 -2093 -388 -2091
rect -374 -2093 -372 -2091
rect -358 -2093 -356 -2091
rect -350 -2093 -348 -2091
rect -340 -2093 -338 -2091
rect -214 -2093 -212 -2091
rect -204 -2093 -202 -2091
rect -188 -2093 -186 -2091
rect -178 -2093 -176 -2091
rect -162 -2093 -160 -2091
rect -152 -2093 -150 -2091
rect -144 -2093 -142 -2091
rect -134 -2093 -132 -2091
rect -118 -2093 -116 -2091
rect -110 -2093 -108 -2091
rect -100 -2093 -98 -2091
rect -84 -2093 -82 -2091
rect -74 -2093 -72 -2091
rect -66 -2093 -64 -2091
rect -56 -2093 -54 -2091
rect -40 -2093 -38 -2091
rect -32 -2093 -30 -2091
rect -16 -2093 -14 -2091
rect 0 -2093 2 -2091
rect 8 -2093 10 -2091
rect 18 -2093 20 -2091
rect 214 -2093 216 -2091
rect 224 -2093 226 -2091
rect 240 -2093 242 -2091
rect 250 -2093 252 -2091
rect 266 -2093 268 -2091
rect 276 -2093 278 -2091
rect 284 -2093 286 -2091
rect 294 -2093 296 -2091
rect 310 -2093 312 -2091
rect 318 -2093 320 -2091
rect 328 -2093 330 -2091
rect 344 -2093 346 -2091
rect 354 -2093 356 -2091
rect 362 -2093 364 -2091
rect 372 -2093 374 -2091
rect 388 -2093 390 -2091
rect 396 -2093 398 -2091
rect 412 -2093 414 -2091
rect 428 -2093 430 -2091
rect 436 -2093 438 -2091
rect 446 -2093 448 -2091
rect 570 -2093 572 -2091
rect 580 -2093 582 -2091
rect 596 -2093 598 -2091
rect 606 -2093 608 -2091
rect 622 -2093 624 -2091
rect 632 -2093 634 -2091
rect 640 -2093 642 -2091
rect 650 -2093 652 -2091
rect 666 -2093 668 -2091
rect 674 -2093 676 -2091
rect 684 -2093 686 -2091
rect 700 -2093 702 -2091
rect 710 -2093 712 -2091
rect 718 -2093 720 -2091
rect 728 -2093 730 -2091
rect 744 -2093 746 -2091
rect 752 -2093 754 -2091
rect 768 -2093 770 -2091
rect 784 -2093 786 -2091
rect 792 -2093 794 -2091
rect 802 -2093 804 -2091
rect 968 -2093 970 -2091
rect 978 -2093 980 -2091
rect 994 -2093 996 -2091
rect 1004 -2093 1006 -2091
rect 1020 -2093 1022 -2091
rect 1030 -2093 1032 -2091
rect 1038 -2093 1040 -2091
rect 1048 -2093 1050 -2091
rect 1064 -2093 1066 -2091
rect 1072 -2093 1074 -2091
rect 1082 -2093 1084 -2091
rect 1098 -2093 1100 -2091
rect 1108 -2093 1110 -2091
rect 1116 -2093 1118 -2091
rect 1126 -2093 1128 -2091
rect 1142 -2093 1144 -2091
rect 1150 -2093 1152 -2091
rect 1166 -2093 1168 -2091
rect 1182 -2093 1184 -2091
rect 1190 -2093 1192 -2091
rect 1200 -2093 1202 -2091
rect 1326 -2093 1328 -2091
rect 1336 -2093 1338 -2091
rect 1352 -2093 1354 -2091
rect 1362 -2093 1364 -2091
rect 1378 -2093 1380 -2091
rect 1388 -2093 1390 -2091
rect 1396 -2093 1398 -2091
rect 1406 -2093 1408 -2091
rect 1422 -2093 1424 -2091
rect 1430 -2093 1432 -2091
rect 1440 -2093 1442 -2091
rect 1456 -2093 1458 -2091
rect 1466 -2093 1468 -2091
rect 1474 -2093 1476 -2091
rect 1484 -2093 1486 -2091
rect 1500 -2093 1502 -2091
rect 1508 -2093 1510 -2091
rect 1524 -2093 1526 -2091
rect 1540 -2093 1542 -2091
rect 1548 -2093 1550 -2091
rect 1558 -2093 1560 -2091
rect -1255 -2169 -1253 -2101
rect -1245 -2169 -1243 -2101
rect -1229 -2169 -1227 -2101
rect -1219 -2169 -1217 -2101
rect -1211 -2169 -1209 -2101
rect -1201 -2169 -1199 -2101
rect -1185 -2169 -1183 -2101
rect -1177 -2169 -1175 -2101
rect -1167 -2169 -1165 -2101
rect -930 -2169 -928 -2101
rect -920 -2169 -918 -2101
rect -904 -2169 -902 -2101
rect -894 -2169 -892 -2101
rect -878 -2169 -876 -2101
rect -868 -2169 -866 -2101
rect -860 -2169 -858 -2101
rect -850 -2169 -848 -2101
rect -834 -2169 -832 -2101
rect -826 -2169 -824 -2101
rect -816 -2169 -814 -2101
rect -800 -2169 -798 -2101
rect -790 -2169 -788 -2101
rect -782 -2169 -780 -2101
rect -772 -2169 -770 -2101
rect -756 -2169 -754 -2101
rect -748 -2169 -746 -2101
rect -732 -2169 -730 -2101
rect -716 -2169 -714 -2101
rect -708 -2169 -706 -2101
rect -698 -2169 -696 -2101
rect -572 -2169 -570 -2101
rect -562 -2169 -560 -2101
rect -546 -2169 -544 -2101
rect -536 -2169 -534 -2101
rect -520 -2169 -518 -2101
rect -510 -2169 -508 -2101
rect -502 -2169 -500 -2101
rect -492 -2169 -490 -2101
rect -476 -2169 -474 -2101
rect -468 -2169 -466 -2101
rect -458 -2169 -456 -2101
rect -442 -2169 -440 -2101
rect -432 -2169 -430 -2101
rect -424 -2169 -422 -2101
rect -414 -2169 -412 -2101
rect -398 -2169 -396 -2101
rect -390 -2169 -388 -2101
rect -374 -2169 -372 -2101
rect -358 -2169 -356 -2101
rect -350 -2169 -348 -2101
rect -340 -2169 -338 -2101
rect -214 -2169 -212 -2101
rect -204 -2169 -202 -2101
rect -188 -2169 -186 -2101
rect -178 -2169 -176 -2101
rect -162 -2169 -160 -2101
rect -152 -2169 -150 -2101
rect -144 -2169 -142 -2101
rect -134 -2169 -132 -2101
rect -118 -2169 -116 -2101
rect -110 -2169 -108 -2101
rect -100 -2169 -98 -2101
rect -84 -2169 -82 -2101
rect -74 -2169 -72 -2101
rect -66 -2169 -64 -2101
rect -56 -2169 -54 -2101
rect -40 -2169 -38 -2101
rect -32 -2169 -30 -2101
rect -16 -2169 -14 -2101
rect 0 -2169 2 -2101
rect 8 -2169 10 -2101
rect 18 -2169 20 -2101
rect 214 -2169 216 -2101
rect 224 -2169 226 -2101
rect 240 -2169 242 -2101
rect 250 -2169 252 -2101
rect 266 -2169 268 -2101
rect 276 -2169 278 -2101
rect 284 -2169 286 -2101
rect 294 -2169 296 -2101
rect 310 -2169 312 -2101
rect 318 -2169 320 -2101
rect 328 -2169 330 -2101
rect 344 -2169 346 -2101
rect 354 -2169 356 -2101
rect 362 -2169 364 -2101
rect 372 -2169 374 -2101
rect 388 -2169 390 -2101
rect 396 -2169 398 -2101
rect 412 -2169 414 -2101
rect 428 -2169 430 -2101
rect 436 -2169 438 -2101
rect 446 -2169 448 -2101
rect 570 -2169 572 -2101
rect 580 -2169 582 -2101
rect 596 -2169 598 -2101
rect 606 -2169 608 -2101
rect 622 -2169 624 -2101
rect 632 -2169 634 -2101
rect 640 -2169 642 -2101
rect 650 -2169 652 -2101
rect 666 -2169 668 -2101
rect 674 -2169 676 -2101
rect 684 -2169 686 -2101
rect 700 -2169 702 -2101
rect 710 -2169 712 -2101
rect 718 -2169 720 -2101
rect 728 -2169 730 -2101
rect 744 -2169 746 -2101
rect 752 -2169 754 -2101
rect 768 -2169 770 -2101
rect 784 -2169 786 -2101
rect 792 -2169 794 -2101
rect 802 -2169 804 -2101
rect 968 -2169 970 -2101
rect 978 -2169 980 -2101
rect 994 -2169 996 -2101
rect 1004 -2169 1006 -2101
rect 1020 -2169 1022 -2101
rect 1030 -2169 1032 -2101
rect 1038 -2169 1040 -2101
rect 1048 -2169 1050 -2101
rect 1064 -2169 1066 -2101
rect 1072 -2169 1074 -2101
rect 1082 -2169 1084 -2101
rect 1098 -2169 1100 -2101
rect 1108 -2169 1110 -2101
rect 1116 -2169 1118 -2101
rect 1126 -2169 1128 -2101
rect 1142 -2169 1144 -2101
rect 1150 -2169 1152 -2101
rect 1166 -2169 1168 -2101
rect 1182 -2169 1184 -2101
rect 1190 -2169 1192 -2101
rect 1200 -2169 1202 -2101
rect 1326 -2169 1328 -2101
rect 1336 -2169 1338 -2101
rect 1352 -2169 1354 -2101
rect 1362 -2169 1364 -2101
rect 1378 -2169 1380 -2101
rect 1388 -2169 1390 -2101
rect 1396 -2169 1398 -2101
rect 1406 -2169 1408 -2101
rect 1422 -2169 1424 -2101
rect 1430 -2169 1432 -2101
rect 1440 -2169 1442 -2101
rect 1456 -2169 1458 -2101
rect 1466 -2169 1468 -2101
rect 1474 -2169 1476 -2101
rect 1484 -2169 1486 -2101
rect 1500 -2169 1502 -2101
rect 1508 -2169 1510 -2101
rect 1524 -2169 1526 -2101
rect 1540 -2169 1542 -2101
rect 1548 -2169 1550 -2101
rect 1558 -2169 1560 -2101
rect -1255 -2175 -1253 -2173
rect -1245 -2175 -1243 -2173
rect -1229 -2175 -1227 -2173
rect -1219 -2175 -1217 -2173
rect -1211 -2175 -1209 -2173
rect -1201 -2175 -1199 -2173
rect -1185 -2175 -1183 -2173
rect -1177 -2175 -1175 -2173
rect -1167 -2175 -1165 -2173
rect -930 -2175 -928 -2173
rect -920 -2175 -918 -2173
rect -904 -2175 -902 -2173
rect -894 -2175 -892 -2173
rect -878 -2175 -876 -2173
rect -868 -2175 -866 -2173
rect -860 -2175 -858 -2173
rect -850 -2175 -848 -2173
rect -834 -2175 -832 -2173
rect -826 -2175 -824 -2173
rect -816 -2175 -814 -2173
rect -800 -2175 -798 -2173
rect -790 -2175 -788 -2173
rect -782 -2175 -780 -2173
rect -772 -2175 -770 -2173
rect -756 -2175 -754 -2173
rect -748 -2175 -746 -2173
rect -732 -2175 -730 -2173
rect -716 -2175 -714 -2173
rect -708 -2175 -706 -2173
rect -698 -2175 -696 -2173
rect -572 -2175 -570 -2173
rect -562 -2175 -560 -2173
rect -546 -2175 -544 -2173
rect -536 -2175 -534 -2173
rect -520 -2175 -518 -2173
rect -510 -2175 -508 -2173
rect -502 -2175 -500 -2173
rect -492 -2175 -490 -2173
rect -476 -2175 -474 -2173
rect -468 -2175 -466 -2173
rect -458 -2175 -456 -2173
rect -442 -2175 -440 -2173
rect -432 -2175 -430 -2173
rect -424 -2175 -422 -2173
rect -414 -2175 -412 -2173
rect -398 -2175 -396 -2173
rect -390 -2175 -388 -2173
rect -374 -2175 -372 -2173
rect -358 -2175 -356 -2173
rect -350 -2175 -348 -2173
rect -340 -2175 -338 -2173
rect -214 -2175 -212 -2173
rect -204 -2175 -202 -2173
rect -188 -2175 -186 -2173
rect -178 -2175 -176 -2173
rect -162 -2175 -160 -2173
rect -152 -2175 -150 -2173
rect -144 -2175 -142 -2173
rect -134 -2175 -132 -2173
rect -118 -2175 -116 -2173
rect -110 -2175 -108 -2173
rect -100 -2175 -98 -2173
rect -84 -2175 -82 -2173
rect -74 -2175 -72 -2173
rect -66 -2175 -64 -2173
rect -56 -2175 -54 -2173
rect -40 -2175 -38 -2173
rect -32 -2175 -30 -2173
rect -16 -2175 -14 -2173
rect 0 -2175 2 -2173
rect 8 -2175 10 -2173
rect 18 -2175 20 -2173
rect 214 -2175 216 -2173
rect 224 -2175 226 -2173
rect 240 -2175 242 -2173
rect 250 -2175 252 -2173
rect 266 -2175 268 -2173
rect 276 -2175 278 -2173
rect 284 -2175 286 -2173
rect 294 -2175 296 -2173
rect 310 -2175 312 -2173
rect 318 -2175 320 -2173
rect 328 -2175 330 -2173
rect 344 -2175 346 -2173
rect 354 -2175 356 -2173
rect 362 -2175 364 -2173
rect 372 -2175 374 -2173
rect 388 -2175 390 -2173
rect 396 -2175 398 -2173
rect 412 -2175 414 -2173
rect 428 -2175 430 -2173
rect 436 -2175 438 -2173
rect 446 -2175 448 -2173
rect 570 -2175 572 -2173
rect 580 -2175 582 -2173
rect 596 -2175 598 -2173
rect 606 -2175 608 -2173
rect 622 -2175 624 -2173
rect 632 -2175 634 -2173
rect 640 -2175 642 -2173
rect 650 -2175 652 -2173
rect 666 -2175 668 -2173
rect 674 -2175 676 -2173
rect 684 -2175 686 -2173
rect 700 -2175 702 -2173
rect 710 -2175 712 -2173
rect 718 -2175 720 -2173
rect 728 -2175 730 -2173
rect 744 -2175 746 -2173
rect 752 -2175 754 -2173
rect 768 -2175 770 -2173
rect 784 -2175 786 -2173
rect 792 -2175 794 -2173
rect 802 -2175 804 -2173
rect 968 -2175 970 -2173
rect 978 -2175 980 -2173
rect 994 -2175 996 -2173
rect 1004 -2175 1006 -2173
rect 1020 -2175 1022 -2173
rect 1030 -2175 1032 -2173
rect 1038 -2175 1040 -2173
rect 1048 -2175 1050 -2173
rect 1064 -2175 1066 -2173
rect 1072 -2175 1074 -2173
rect 1082 -2175 1084 -2173
rect 1098 -2175 1100 -2173
rect 1108 -2175 1110 -2173
rect 1116 -2175 1118 -2173
rect 1126 -2175 1128 -2173
rect 1142 -2175 1144 -2173
rect 1150 -2175 1152 -2173
rect 1166 -2175 1168 -2173
rect 1182 -2175 1184 -2173
rect 1190 -2175 1192 -2173
rect 1200 -2175 1202 -2173
rect 1326 -2175 1328 -2173
rect 1336 -2175 1338 -2173
rect 1352 -2175 1354 -2173
rect 1362 -2175 1364 -2173
rect 1378 -2175 1380 -2173
rect 1388 -2175 1390 -2173
rect 1396 -2175 1398 -2173
rect 1406 -2175 1408 -2173
rect 1422 -2175 1424 -2173
rect 1430 -2175 1432 -2173
rect 1440 -2175 1442 -2173
rect 1456 -2175 1458 -2173
rect 1466 -2175 1468 -2173
rect 1474 -2175 1476 -2173
rect 1484 -2175 1486 -2173
rect 1500 -2175 1502 -2173
rect 1508 -2175 1510 -2173
rect 1524 -2175 1526 -2173
rect 1540 -2175 1542 -2173
rect 1548 -2175 1550 -2173
rect 1558 -2175 1560 -2173
rect -1259 -2237 -1257 -2235
rect -1249 -2237 -1247 -2235
rect -1233 -2237 -1231 -2235
rect -1225 -2237 -1223 -2235
rect -1209 -2237 -1207 -2235
rect -1201 -2237 -1199 -2235
rect -1191 -2237 -1189 -2235
rect -1183 -2237 -1181 -2235
rect -1167 -2237 -1165 -2235
rect -1159 -2237 -1157 -2235
rect -1149 -2237 -1147 -2235
rect -1141 -2237 -1139 -2235
rect -1125 -2237 -1123 -2235
rect -1117 -2237 -1115 -2235
rect -1107 -2237 -1105 -2235
rect -1099 -2237 -1097 -2235
rect -1083 -2237 -1081 -2235
rect -1075 -2237 -1073 -2235
rect -930 -2237 -928 -2235
rect -920 -2237 -918 -2235
rect -904 -2237 -902 -2235
rect -896 -2237 -894 -2235
rect -880 -2237 -878 -2235
rect -872 -2237 -870 -2235
rect -862 -2237 -860 -2235
rect -854 -2237 -852 -2235
rect -838 -2237 -836 -2235
rect -830 -2237 -828 -2235
rect -820 -2237 -818 -2235
rect -812 -2237 -810 -2235
rect -796 -2237 -794 -2235
rect -788 -2237 -786 -2235
rect -778 -2237 -776 -2235
rect -770 -2237 -768 -2235
rect -754 -2237 -752 -2235
rect -746 -2237 -744 -2235
rect -572 -2237 -570 -2235
rect -562 -2237 -560 -2235
rect -546 -2237 -544 -2235
rect -538 -2237 -536 -2235
rect -522 -2237 -520 -2235
rect -514 -2237 -512 -2235
rect -504 -2237 -502 -2235
rect -496 -2237 -494 -2235
rect -480 -2237 -478 -2235
rect -472 -2237 -470 -2235
rect -462 -2237 -460 -2235
rect -454 -2237 -452 -2235
rect -438 -2237 -436 -2235
rect -430 -2237 -428 -2235
rect -420 -2237 -418 -2235
rect -412 -2237 -410 -2235
rect -396 -2237 -394 -2235
rect -388 -2237 -386 -2235
rect -214 -2237 -212 -2235
rect -204 -2237 -202 -2235
rect -188 -2237 -186 -2235
rect -180 -2237 -178 -2235
rect -164 -2237 -162 -2235
rect -156 -2237 -154 -2235
rect -146 -2237 -144 -2235
rect -138 -2237 -136 -2235
rect -122 -2237 -120 -2235
rect -114 -2237 -112 -2235
rect -104 -2237 -102 -2235
rect -96 -2237 -94 -2235
rect -80 -2237 -78 -2235
rect -72 -2237 -70 -2235
rect -62 -2237 -60 -2235
rect -54 -2237 -52 -2235
rect -38 -2237 -36 -2235
rect -30 -2237 -28 -2235
rect 214 -2237 216 -2235
rect 224 -2237 226 -2235
rect 240 -2237 242 -2235
rect 248 -2237 250 -2235
rect 264 -2237 266 -2235
rect 272 -2237 274 -2235
rect 282 -2237 284 -2235
rect 290 -2237 292 -2235
rect 306 -2237 308 -2235
rect 314 -2237 316 -2235
rect 324 -2237 326 -2235
rect 332 -2237 334 -2235
rect 348 -2237 350 -2235
rect 356 -2237 358 -2235
rect 366 -2237 368 -2235
rect 374 -2237 376 -2235
rect 390 -2237 392 -2235
rect 398 -2237 400 -2235
rect 570 -2237 572 -2235
rect 580 -2237 582 -2235
rect 596 -2237 598 -2235
rect 604 -2237 606 -2235
rect 620 -2237 622 -2235
rect 628 -2237 630 -2235
rect 638 -2237 640 -2235
rect 646 -2237 648 -2235
rect 662 -2237 664 -2235
rect 670 -2237 672 -2235
rect 680 -2237 682 -2235
rect 688 -2237 690 -2235
rect 704 -2237 706 -2235
rect 712 -2237 714 -2235
rect 722 -2237 724 -2235
rect 730 -2237 732 -2235
rect 746 -2237 748 -2235
rect 754 -2237 756 -2235
rect -1259 -2313 -1257 -2245
rect -1249 -2313 -1247 -2245
rect -1233 -2313 -1231 -2245
rect -1225 -2313 -1223 -2245
rect -1209 -2313 -1207 -2245
rect -1201 -2313 -1199 -2245
rect -1191 -2313 -1189 -2245
rect -1183 -2313 -1181 -2245
rect -1167 -2313 -1165 -2245
rect -1159 -2278 -1157 -2245
rect -1149 -2278 -1147 -2245
rect -1159 -2280 -1147 -2278
rect -1159 -2313 -1157 -2280
rect -1149 -2313 -1147 -2280
rect -1141 -2313 -1139 -2245
rect -1125 -2313 -1123 -2245
rect -1117 -2313 -1115 -2245
rect -1107 -2313 -1105 -2245
rect -1099 -2313 -1097 -2245
rect -1083 -2313 -1081 -2245
rect -1075 -2313 -1073 -2245
rect -930 -2313 -928 -2245
rect -920 -2313 -918 -2245
rect -904 -2313 -902 -2245
rect -896 -2313 -894 -2245
rect -880 -2313 -878 -2245
rect -872 -2313 -870 -2245
rect -862 -2313 -860 -2245
rect -854 -2313 -852 -2245
rect -838 -2313 -836 -2245
rect -830 -2278 -828 -2245
rect -820 -2278 -818 -2245
rect -830 -2280 -818 -2278
rect -830 -2313 -828 -2280
rect -820 -2313 -818 -2280
rect -812 -2313 -810 -2245
rect -796 -2313 -794 -2245
rect -788 -2313 -786 -2245
rect -778 -2313 -776 -2245
rect -770 -2313 -768 -2245
rect -754 -2313 -752 -2245
rect -746 -2313 -744 -2245
rect -572 -2313 -570 -2245
rect -562 -2313 -560 -2245
rect -546 -2313 -544 -2245
rect -538 -2313 -536 -2245
rect -522 -2313 -520 -2245
rect -514 -2313 -512 -2245
rect -504 -2313 -502 -2245
rect -496 -2313 -494 -2245
rect -480 -2313 -478 -2245
rect -472 -2278 -470 -2245
rect -462 -2278 -460 -2245
rect -472 -2280 -460 -2278
rect -472 -2313 -470 -2280
rect -462 -2313 -460 -2280
rect -454 -2313 -452 -2245
rect -438 -2313 -436 -2245
rect -430 -2313 -428 -2245
rect -420 -2313 -418 -2245
rect -412 -2313 -410 -2245
rect -396 -2313 -394 -2245
rect -388 -2313 -386 -2245
rect -214 -2313 -212 -2245
rect -204 -2313 -202 -2245
rect -188 -2313 -186 -2245
rect -180 -2313 -178 -2245
rect -164 -2313 -162 -2245
rect -156 -2313 -154 -2245
rect -146 -2313 -144 -2245
rect -138 -2313 -136 -2245
rect -122 -2313 -120 -2245
rect -114 -2278 -112 -2245
rect -104 -2278 -102 -2245
rect -114 -2280 -102 -2278
rect -114 -2313 -112 -2280
rect -104 -2313 -102 -2280
rect -96 -2313 -94 -2245
rect -80 -2313 -78 -2245
rect -72 -2313 -70 -2245
rect -62 -2313 -60 -2245
rect -54 -2313 -52 -2245
rect -38 -2313 -36 -2245
rect -30 -2313 -28 -2245
rect 214 -2313 216 -2245
rect 224 -2313 226 -2245
rect 240 -2313 242 -2245
rect 248 -2313 250 -2245
rect 264 -2313 266 -2245
rect 272 -2313 274 -2245
rect 282 -2313 284 -2245
rect 290 -2313 292 -2245
rect 306 -2313 308 -2245
rect 314 -2278 316 -2245
rect 324 -2278 326 -2245
rect 314 -2280 326 -2278
rect 314 -2313 316 -2280
rect 324 -2313 326 -2280
rect 332 -2313 334 -2245
rect 348 -2313 350 -2245
rect 356 -2313 358 -2245
rect 366 -2313 368 -2245
rect 374 -2313 376 -2245
rect 390 -2313 392 -2245
rect 398 -2313 400 -2245
rect 570 -2313 572 -2245
rect 580 -2313 582 -2245
rect 596 -2313 598 -2245
rect 604 -2313 606 -2245
rect 620 -2313 622 -2245
rect 628 -2313 630 -2245
rect 638 -2313 640 -2245
rect 646 -2313 648 -2245
rect 662 -2313 664 -2245
rect 670 -2278 672 -2245
rect 680 -2278 682 -2245
rect 670 -2280 682 -2278
rect 670 -2313 672 -2280
rect 680 -2313 682 -2280
rect 688 -2313 690 -2245
rect 704 -2313 706 -2245
rect 712 -2313 714 -2245
rect 722 -2313 724 -2245
rect 730 -2313 732 -2245
rect 746 -2313 748 -2245
rect 754 -2313 756 -2245
rect -1259 -2319 -1257 -2317
rect -1249 -2319 -1247 -2317
rect -1233 -2319 -1231 -2317
rect -1225 -2319 -1223 -2317
rect -1209 -2319 -1207 -2317
rect -1201 -2319 -1199 -2317
rect -1191 -2319 -1189 -2317
rect -1183 -2319 -1181 -2317
rect -1167 -2319 -1165 -2317
rect -1159 -2319 -1157 -2317
rect -1149 -2319 -1147 -2317
rect -1141 -2319 -1139 -2317
rect -1125 -2319 -1123 -2317
rect -1117 -2319 -1115 -2317
rect -1107 -2319 -1105 -2317
rect -1099 -2319 -1097 -2317
rect -1083 -2319 -1081 -2317
rect -1075 -2319 -1073 -2317
rect -930 -2319 -928 -2317
rect -920 -2319 -918 -2317
rect -904 -2319 -902 -2317
rect -896 -2319 -894 -2317
rect -880 -2319 -878 -2317
rect -872 -2319 -870 -2317
rect -862 -2319 -860 -2317
rect -854 -2319 -852 -2317
rect -838 -2319 -836 -2317
rect -830 -2319 -828 -2317
rect -820 -2319 -818 -2317
rect -812 -2319 -810 -2317
rect -796 -2319 -794 -2317
rect -788 -2319 -786 -2317
rect -778 -2319 -776 -2317
rect -770 -2319 -768 -2317
rect -754 -2319 -752 -2317
rect -746 -2319 -744 -2317
rect -572 -2319 -570 -2317
rect -562 -2319 -560 -2317
rect -546 -2319 -544 -2317
rect -538 -2319 -536 -2317
rect -522 -2319 -520 -2317
rect -514 -2319 -512 -2317
rect -504 -2319 -502 -2317
rect -496 -2319 -494 -2317
rect -480 -2319 -478 -2317
rect -472 -2319 -470 -2317
rect -462 -2319 -460 -2317
rect -454 -2319 -452 -2317
rect -438 -2319 -436 -2317
rect -430 -2319 -428 -2317
rect -420 -2319 -418 -2317
rect -412 -2319 -410 -2317
rect -396 -2319 -394 -2317
rect -388 -2319 -386 -2317
rect -214 -2319 -212 -2317
rect -204 -2319 -202 -2317
rect -188 -2319 -186 -2317
rect -180 -2319 -178 -2317
rect -164 -2319 -162 -2317
rect -156 -2319 -154 -2317
rect -146 -2319 -144 -2317
rect -138 -2319 -136 -2317
rect -122 -2319 -120 -2317
rect -114 -2319 -112 -2317
rect -104 -2319 -102 -2317
rect -96 -2319 -94 -2317
rect -80 -2319 -78 -2317
rect -72 -2319 -70 -2317
rect -62 -2319 -60 -2317
rect -54 -2319 -52 -2317
rect -38 -2319 -36 -2317
rect -30 -2319 -28 -2317
rect 214 -2319 216 -2317
rect 224 -2319 226 -2317
rect 240 -2319 242 -2317
rect 248 -2319 250 -2317
rect 264 -2319 266 -2317
rect 272 -2319 274 -2317
rect 282 -2319 284 -2317
rect 290 -2319 292 -2317
rect 306 -2319 308 -2317
rect 314 -2319 316 -2317
rect 324 -2319 326 -2317
rect 332 -2319 334 -2317
rect 348 -2319 350 -2317
rect 356 -2319 358 -2317
rect 366 -2319 368 -2317
rect 374 -2319 376 -2317
rect 390 -2319 392 -2317
rect 398 -2319 400 -2317
rect 570 -2319 572 -2317
rect 580 -2319 582 -2317
rect 596 -2319 598 -2317
rect 604 -2319 606 -2317
rect 620 -2319 622 -2317
rect 628 -2319 630 -2317
rect 638 -2319 640 -2317
rect 646 -2319 648 -2317
rect 662 -2319 664 -2317
rect 670 -2319 672 -2317
rect 680 -2319 682 -2317
rect 688 -2319 690 -2317
rect 704 -2319 706 -2317
rect 712 -2319 714 -2317
rect 722 -2319 724 -2317
rect 730 -2319 732 -2317
rect 746 -2319 748 -2317
rect 754 -2319 756 -2317
rect -1259 -2368 -1257 -2366
rect -1249 -2368 -1247 -2366
rect -1233 -2368 -1231 -2366
rect -1225 -2368 -1223 -2366
rect -1209 -2368 -1207 -2366
rect -1201 -2368 -1199 -2366
rect -1191 -2368 -1189 -2366
rect -1183 -2368 -1181 -2366
rect -1167 -2368 -1165 -2366
rect -1159 -2368 -1157 -2366
rect -1149 -2368 -1147 -2366
rect -1141 -2368 -1139 -2366
rect -1125 -2368 -1123 -2366
rect -1117 -2368 -1115 -2366
rect -1107 -2368 -1105 -2366
rect -1099 -2368 -1097 -2366
rect -1083 -2368 -1081 -2366
rect -1075 -2368 -1073 -2366
rect -930 -2368 -928 -2366
rect -920 -2368 -918 -2366
rect -904 -2368 -902 -2366
rect -896 -2368 -894 -2366
rect -880 -2368 -878 -2366
rect -872 -2368 -870 -2366
rect -862 -2368 -860 -2366
rect -854 -2368 -852 -2366
rect -838 -2368 -836 -2366
rect -830 -2368 -828 -2366
rect -820 -2368 -818 -2366
rect -812 -2368 -810 -2366
rect -796 -2368 -794 -2366
rect -788 -2368 -786 -2366
rect -778 -2368 -776 -2366
rect -770 -2368 -768 -2366
rect -754 -2368 -752 -2366
rect -746 -2368 -744 -2366
rect -572 -2368 -570 -2366
rect -562 -2368 -560 -2366
rect -546 -2368 -544 -2366
rect -538 -2368 -536 -2366
rect -522 -2368 -520 -2366
rect -514 -2368 -512 -2366
rect -504 -2368 -502 -2366
rect -496 -2368 -494 -2366
rect -480 -2368 -478 -2366
rect -472 -2368 -470 -2366
rect -462 -2368 -460 -2366
rect -454 -2368 -452 -2366
rect -438 -2368 -436 -2366
rect -430 -2368 -428 -2366
rect -420 -2368 -418 -2366
rect -412 -2368 -410 -2366
rect -396 -2368 -394 -2366
rect -388 -2368 -386 -2366
rect -214 -2368 -212 -2366
rect -204 -2368 -202 -2366
rect -188 -2368 -186 -2366
rect -180 -2368 -178 -2366
rect -164 -2368 -162 -2366
rect -156 -2368 -154 -2366
rect -146 -2368 -144 -2366
rect -138 -2368 -136 -2366
rect -122 -2368 -120 -2366
rect -114 -2368 -112 -2366
rect -104 -2368 -102 -2366
rect -96 -2368 -94 -2366
rect -80 -2368 -78 -2366
rect -72 -2368 -70 -2366
rect -62 -2368 -60 -2366
rect -54 -2368 -52 -2366
rect -38 -2368 -36 -2366
rect -30 -2368 -28 -2366
rect 214 -2368 216 -2366
rect 224 -2368 226 -2366
rect 240 -2368 242 -2366
rect 248 -2368 250 -2366
rect 264 -2368 266 -2366
rect 272 -2368 274 -2366
rect 282 -2368 284 -2366
rect 290 -2368 292 -2366
rect 306 -2368 308 -2366
rect 314 -2368 316 -2366
rect 324 -2368 326 -2366
rect 332 -2368 334 -2366
rect 348 -2368 350 -2366
rect 356 -2368 358 -2366
rect 366 -2368 368 -2366
rect 374 -2368 376 -2366
rect 390 -2368 392 -2366
rect 398 -2368 400 -2366
rect 570 -2368 572 -2366
rect 580 -2368 582 -2366
rect 596 -2368 598 -2366
rect 604 -2368 606 -2366
rect 620 -2368 622 -2366
rect 628 -2368 630 -2366
rect 638 -2368 640 -2366
rect 646 -2368 648 -2366
rect 662 -2368 664 -2366
rect 670 -2368 672 -2366
rect 680 -2368 682 -2366
rect 688 -2368 690 -2366
rect 704 -2368 706 -2366
rect 712 -2368 714 -2366
rect 722 -2368 724 -2366
rect 730 -2368 732 -2366
rect 746 -2368 748 -2366
rect 754 -2368 756 -2366
rect 968 -2368 970 -2366
rect 978 -2368 980 -2366
rect 994 -2368 996 -2366
rect 1002 -2368 1004 -2366
rect 1018 -2368 1020 -2366
rect 1026 -2368 1028 -2366
rect 1036 -2368 1038 -2366
rect 1044 -2368 1046 -2366
rect 1060 -2368 1062 -2366
rect 1068 -2368 1070 -2366
rect 1078 -2368 1080 -2366
rect 1086 -2368 1088 -2366
rect 1102 -2368 1104 -2366
rect 1110 -2368 1112 -2366
rect 1120 -2368 1122 -2366
rect 1128 -2368 1130 -2366
rect 1144 -2368 1146 -2366
rect 1152 -2368 1154 -2366
rect 1326 -2368 1328 -2366
rect 1336 -2368 1338 -2366
rect 1352 -2368 1354 -2366
rect 1360 -2368 1362 -2366
rect 1376 -2368 1378 -2366
rect 1384 -2368 1386 -2366
rect 1394 -2368 1396 -2366
rect 1402 -2368 1404 -2366
rect 1418 -2368 1420 -2366
rect 1426 -2368 1428 -2366
rect 1436 -2368 1438 -2366
rect 1444 -2368 1446 -2366
rect 1460 -2368 1462 -2366
rect 1468 -2368 1470 -2366
rect 1478 -2368 1480 -2366
rect 1486 -2368 1488 -2366
rect 1502 -2368 1504 -2366
rect 1510 -2368 1512 -2366
rect -1259 -2444 -1257 -2376
rect -1249 -2444 -1247 -2376
rect -1233 -2444 -1231 -2376
rect -1225 -2444 -1223 -2376
rect -1209 -2444 -1207 -2376
rect -1201 -2444 -1199 -2376
rect -1191 -2444 -1189 -2376
rect -1183 -2444 -1181 -2376
rect -1167 -2444 -1165 -2376
rect -1159 -2409 -1157 -2376
rect -1149 -2409 -1147 -2376
rect -1159 -2411 -1147 -2409
rect -1159 -2444 -1157 -2411
rect -1149 -2444 -1147 -2411
rect -1141 -2444 -1139 -2376
rect -1125 -2444 -1123 -2376
rect -1117 -2444 -1115 -2376
rect -1107 -2444 -1105 -2376
rect -1099 -2444 -1097 -2376
rect -1083 -2444 -1081 -2376
rect -1075 -2444 -1073 -2376
rect -930 -2444 -928 -2376
rect -920 -2444 -918 -2376
rect -904 -2444 -902 -2376
rect -896 -2444 -894 -2376
rect -880 -2444 -878 -2376
rect -872 -2444 -870 -2376
rect -862 -2444 -860 -2376
rect -854 -2444 -852 -2376
rect -838 -2444 -836 -2376
rect -830 -2409 -828 -2376
rect -820 -2409 -818 -2376
rect -830 -2411 -818 -2409
rect -830 -2444 -828 -2411
rect -820 -2444 -818 -2411
rect -812 -2444 -810 -2376
rect -796 -2444 -794 -2376
rect -788 -2444 -786 -2376
rect -778 -2444 -776 -2376
rect -770 -2444 -768 -2376
rect -754 -2444 -752 -2376
rect -746 -2444 -744 -2376
rect -572 -2444 -570 -2376
rect -562 -2444 -560 -2376
rect -546 -2444 -544 -2376
rect -538 -2444 -536 -2376
rect -522 -2444 -520 -2376
rect -514 -2444 -512 -2376
rect -504 -2444 -502 -2376
rect -496 -2444 -494 -2376
rect -480 -2444 -478 -2376
rect -472 -2409 -470 -2376
rect -462 -2409 -460 -2376
rect -472 -2411 -460 -2409
rect -472 -2444 -470 -2411
rect -462 -2444 -460 -2411
rect -454 -2444 -452 -2376
rect -438 -2444 -436 -2376
rect -430 -2444 -428 -2376
rect -420 -2444 -418 -2376
rect -412 -2444 -410 -2376
rect -396 -2444 -394 -2376
rect -388 -2444 -386 -2376
rect -214 -2444 -212 -2376
rect -204 -2444 -202 -2376
rect -188 -2444 -186 -2376
rect -180 -2444 -178 -2376
rect -164 -2444 -162 -2376
rect -156 -2444 -154 -2376
rect -146 -2444 -144 -2376
rect -138 -2444 -136 -2376
rect -122 -2444 -120 -2376
rect -114 -2409 -112 -2376
rect -104 -2409 -102 -2376
rect -114 -2411 -102 -2409
rect -114 -2444 -112 -2411
rect -104 -2444 -102 -2411
rect -96 -2444 -94 -2376
rect -80 -2444 -78 -2376
rect -72 -2444 -70 -2376
rect -62 -2444 -60 -2376
rect -54 -2444 -52 -2376
rect -38 -2444 -36 -2376
rect -30 -2444 -28 -2376
rect 214 -2444 216 -2376
rect 224 -2444 226 -2376
rect 240 -2444 242 -2376
rect 248 -2444 250 -2376
rect 264 -2444 266 -2376
rect 272 -2444 274 -2376
rect 282 -2444 284 -2376
rect 290 -2444 292 -2376
rect 306 -2444 308 -2376
rect 314 -2409 316 -2376
rect 324 -2409 326 -2376
rect 314 -2411 326 -2409
rect 314 -2444 316 -2411
rect 324 -2444 326 -2411
rect 332 -2444 334 -2376
rect 348 -2444 350 -2376
rect 356 -2444 358 -2376
rect 366 -2444 368 -2376
rect 374 -2444 376 -2376
rect 390 -2444 392 -2376
rect 398 -2444 400 -2376
rect 570 -2444 572 -2376
rect 580 -2444 582 -2376
rect 596 -2444 598 -2376
rect 604 -2444 606 -2376
rect 620 -2444 622 -2376
rect 628 -2444 630 -2376
rect 638 -2444 640 -2376
rect 646 -2444 648 -2376
rect 662 -2444 664 -2376
rect 670 -2409 672 -2376
rect 680 -2409 682 -2376
rect 670 -2411 682 -2409
rect 670 -2444 672 -2411
rect 680 -2444 682 -2411
rect 688 -2444 690 -2376
rect 704 -2444 706 -2376
rect 712 -2444 714 -2376
rect 722 -2444 724 -2376
rect 730 -2444 732 -2376
rect 746 -2444 748 -2376
rect 754 -2444 756 -2376
rect 968 -2444 970 -2376
rect 978 -2444 980 -2376
rect 994 -2444 996 -2376
rect 1002 -2444 1004 -2376
rect 1018 -2444 1020 -2376
rect 1026 -2444 1028 -2376
rect 1036 -2444 1038 -2376
rect 1044 -2444 1046 -2376
rect 1060 -2444 1062 -2376
rect 1068 -2409 1070 -2376
rect 1078 -2409 1080 -2376
rect 1068 -2411 1080 -2409
rect 1068 -2444 1070 -2411
rect 1078 -2444 1080 -2411
rect 1086 -2444 1088 -2376
rect 1102 -2444 1104 -2376
rect 1110 -2444 1112 -2376
rect 1120 -2444 1122 -2376
rect 1128 -2444 1130 -2376
rect 1144 -2444 1146 -2376
rect 1152 -2444 1154 -2376
rect 1326 -2444 1328 -2376
rect 1336 -2444 1338 -2376
rect 1352 -2444 1354 -2376
rect 1360 -2444 1362 -2376
rect 1376 -2444 1378 -2376
rect 1384 -2444 1386 -2376
rect 1394 -2444 1396 -2376
rect 1402 -2444 1404 -2376
rect 1418 -2444 1420 -2376
rect 1426 -2409 1428 -2376
rect 1436 -2409 1438 -2376
rect 1426 -2411 1438 -2409
rect 1426 -2444 1428 -2411
rect 1436 -2444 1438 -2411
rect 1444 -2444 1446 -2376
rect 1460 -2444 1462 -2376
rect 1468 -2444 1470 -2376
rect 1478 -2444 1480 -2376
rect 1486 -2444 1488 -2376
rect 1502 -2444 1504 -2376
rect 1510 -2444 1512 -2376
rect -1259 -2450 -1257 -2448
rect -1249 -2450 -1247 -2448
rect -1233 -2450 -1231 -2448
rect -1225 -2450 -1223 -2448
rect -1209 -2450 -1207 -2448
rect -1201 -2450 -1199 -2448
rect -1191 -2450 -1189 -2448
rect -1183 -2450 -1181 -2448
rect -1167 -2450 -1165 -2448
rect -1159 -2450 -1157 -2448
rect -1149 -2450 -1147 -2448
rect -1141 -2450 -1139 -2448
rect -1125 -2450 -1123 -2448
rect -1117 -2450 -1115 -2448
rect -1107 -2450 -1105 -2448
rect -1099 -2450 -1097 -2448
rect -1083 -2450 -1081 -2448
rect -1075 -2450 -1073 -2448
rect -930 -2450 -928 -2448
rect -920 -2450 -918 -2448
rect -904 -2450 -902 -2448
rect -896 -2450 -894 -2448
rect -880 -2450 -878 -2448
rect -872 -2450 -870 -2448
rect -862 -2450 -860 -2448
rect -854 -2450 -852 -2448
rect -838 -2450 -836 -2448
rect -830 -2450 -828 -2448
rect -820 -2450 -818 -2448
rect -812 -2450 -810 -2448
rect -796 -2450 -794 -2448
rect -788 -2450 -786 -2448
rect -778 -2450 -776 -2448
rect -770 -2450 -768 -2448
rect -754 -2450 -752 -2448
rect -746 -2450 -744 -2448
rect -572 -2450 -570 -2448
rect -562 -2450 -560 -2448
rect -546 -2450 -544 -2448
rect -538 -2450 -536 -2448
rect -522 -2450 -520 -2448
rect -514 -2450 -512 -2448
rect -504 -2450 -502 -2448
rect -496 -2450 -494 -2448
rect -480 -2450 -478 -2448
rect -472 -2450 -470 -2448
rect -462 -2450 -460 -2448
rect -454 -2450 -452 -2448
rect -438 -2450 -436 -2448
rect -430 -2450 -428 -2448
rect -420 -2450 -418 -2448
rect -412 -2450 -410 -2448
rect -396 -2450 -394 -2448
rect -388 -2450 -386 -2448
rect -214 -2450 -212 -2448
rect -204 -2450 -202 -2448
rect -188 -2450 -186 -2448
rect -180 -2450 -178 -2448
rect -164 -2450 -162 -2448
rect -156 -2450 -154 -2448
rect -146 -2450 -144 -2448
rect -138 -2450 -136 -2448
rect -122 -2450 -120 -2448
rect -114 -2450 -112 -2448
rect -104 -2450 -102 -2448
rect -96 -2450 -94 -2448
rect -80 -2450 -78 -2448
rect -72 -2450 -70 -2448
rect -62 -2450 -60 -2448
rect -54 -2450 -52 -2448
rect -38 -2450 -36 -2448
rect -30 -2450 -28 -2448
rect 214 -2450 216 -2448
rect 224 -2450 226 -2448
rect 240 -2450 242 -2448
rect 248 -2450 250 -2448
rect 264 -2450 266 -2448
rect 272 -2450 274 -2448
rect 282 -2450 284 -2448
rect 290 -2450 292 -2448
rect 306 -2450 308 -2448
rect 314 -2450 316 -2448
rect 324 -2450 326 -2448
rect 332 -2450 334 -2448
rect 348 -2450 350 -2448
rect 356 -2450 358 -2448
rect 366 -2450 368 -2448
rect 374 -2450 376 -2448
rect 390 -2450 392 -2448
rect 398 -2450 400 -2448
rect 570 -2450 572 -2448
rect 580 -2450 582 -2448
rect 596 -2450 598 -2448
rect 604 -2450 606 -2448
rect 620 -2450 622 -2448
rect 628 -2450 630 -2448
rect 638 -2450 640 -2448
rect 646 -2450 648 -2448
rect 662 -2450 664 -2448
rect 670 -2450 672 -2448
rect 680 -2450 682 -2448
rect 688 -2450 690 -2448
rect 704 -2450 706 -2448
rect 712 -2450 714 -2448
rect 722 -2450 724 -2448
rect 730 -2450 732 -2448
rect 746 -2450 748 -2448
rect 754 -2450 756 -2448
rect 968 -2450 970 -2448
rect 978 -2450 980 -2448
rect 994 -2450 996 -2448
rect 1002 -2450 1004 -2448
rect 1018 -2450 1020 -2448
rect 1026 -2450 1028 -2448
rect 1036 -2450 1038 -2448
rect 1044 -2450 1046 -2448
rect 1060 -2450 1062 -2448
rect 1068 -2450 1070 -2448
rect 1078 -2450 1080 -2448
rect 1086 -2450 1088 -2448
rect 1102 -2450 1104 -2448
rect 1110 -2450 1112 -2448
rect 1120 -2450 1122 -2448
rect 1128 -2450 1130 -2448
rect 1144 -2450 1146 -2448
rect 1152 -2450 1154 -2448
rect 1326 -2450 1328 -2448
rect 1336 -2450 1338 -2448
rect 1352 -2450 1354 -2448
rect 1360 -2450 1362 -2448
rect 1376 -2450 1378 -2448
rect 1384 -2450 1386 -2448
rect 1394 -2450 1396 -2448
rect 1402 -2450 1404 -2448
rect 1418 -2450 1420 -2448
rect 1426 -2450 1428 -2448
rect 1436 -2450 1438 -2448
rect 1444 -2450 1446 -2448
rect 1460 -2450 1462 -2448
rect 1468 -2450 1470 -2448
rect 1478 -2450 1480 -2448
rect 1486 -2450 1488 -2448
rect 1502 -2450 1504 -2448
rect 1510 -2450 1512 -2448
rect -1259 -2499 -1257 -2497
rect -1249 -2499 -1247 -2497
rect -1233 -2499 -1231 -2497
rect -1225 -2499 -1223 -2497
rect -1209 -2499 -1207 -2497
rect -1201 -2499 -1199 -2497
rect -1191 -2499 -1189 -2497
rect -1183 -2499 -1181 -2497
rect -1167 -2499 -1165 -2497
rect -1159 -2499 -1157 -2497
rect -1149 -2499 -1147 -2497
rect -1141 -2499 -1139 -2497
rect -1125 -2499 -1123 -2497
rect -1117 -2499 -1115 -2497
rect -1107 -2499 -1105 -2497
rect -1099 -2499 -1097 -2497
rect -1083 -2499 -1081 -2497
rect -1075 -2499 -1073 -2497
rect -930 -2499 -928 -2497
rect -920 -2499 -918 -2497
rect -904 -2499 -902 -2497
rect -896 -2499 -894 -2497
rect -880 -2499 -878 -2497
rect -872 -2499 -870 -2497
rect -862 -2499 -860 -2497
rect -854 -2499 -852 -2497
rect -838 -2499 -836 -2497
rect -830 -2499 -828 -2497
rect -820 -2499 -818 -2497
rect -812 -2499 -810 -2497
rect -796 -2499 -794 -2497
rect -788 -2499 -786 -2497
rect -778 -2499 -776 -2497
rect -770 -2499 -768 -2497
rect -754 -2499 -752 -2497
rect -746 -2499 -744 -2497
rect -572 -2499 -570 -2497
rect -562 -2499 -560 -2497
rect -546 -2499 -544 -2497
rect -538 -2499 -536 -2497
rect -522 -2499 -520 -2497
rect -514 -2499 -512 -2497
rect -504 -2499 -502 -2497
rect -496 -2499 -494 -2497
rect -480 -2499 -478 -2497
rect -472 -2499 -470 -2497
rect -462 -2499 -460 -2497
rect -454 -2499 -452 -2497
rect -438 -2499 -436 -2497
rect -430 -2499 -428 -2497
rect -420 -2499 -418 -2497
rect -412 -2499 -410 -2497
rect -396 -2499 -394 -2497
rect -388 -2499 -386 -2497
rect -214 -2499 -212 -2497
rect -204 -2499 -202 -2497
rect -188 -2499 -186 -2497
rect -180 -2499 -178 -2497
rect -164 -2499 -162 -2497
rect -156 -2499 -154 -2497
rect -146 -2499 -144 -2497
rect -138 -2499 -136 -2497
rect -122 -2499 -120 -2497
rect -114 -2499 -112 -2497
rect -104 -2499 -102 -2497
rect -96 -2499 -94 -2497
rect -80 -2499 -78 -2497
rect -72 -2499 -70 -2497
rect -62 -2499 -60 -2497
rect -54 -2499 -52 -2497
rect -38 -2499 -36 -2497
rect -30 -2499 -28 -2497
rect 95 -2499 97 -2497
rect 214 -2499 216 -2497
rect 224 -2499 226 -2497
rect 240 -2499 242 -2497
rect 248 -2499 250 -2497
rect 264 -2499 266 -2497
rect 272 -2499 274 -2497
rect 282 -2499 284 -2497
rect 290 -2499 292 -2497
rect 306 -2499 308 -2497
rect 314 -2499 316 -2497
rect 324 -2499 326 -2497
rect 332 -2499 334 -2497
rect 348 -2499 350 -2497
rect 356 -2499 358 -2497
rect 366 -2499 368 -2497
rect 374 -2499 376 -2497
rect 390 -2499 392 -2497
rect 398 -2499 400 -2497
rect 570 -2499 572 -2497
rect 580 -2499 582 -2497
rect 596 -2499 598 -2497
rect 604 -2499 606 -2497
rect 620 -2499 622 -2497
rect 628 -2499 630 -2497
rect 638 -2499 640 -2497
rect 646 -2499 648 -2497
rect 662 -2499 664 -2497
rect 670 -2499 672 -2497
rect 680 -2499 682 -2497
rect 688 -2499 690 -2497
rect 704 -2499 706 -2497
rect 712 -2499 714 -2497
rect 722 -2499 724 -2497
rect 730 -2499 732 -2497
rect 746 -2499 748 -2497
rect 754 -2499 756 -2497
rect 968 -2499 970 -2497
rect 978 -2499 980 -2497
rect 994 -2499 996 -2497
rect 1002 -2499 1004 -2497
rect 1018 -2499 1020 -2497
rect 1026 -2499 1028 -2497
rect 1036 -2499 1038 -2497
rect 1044 -2499 1046 -2497
rect 1060 -2499 1062 -2497
rect 1068 -2499 1070 -2497
rect 1078 -2499 1080 -2497
rect 1086 -2499 1088 -2497
rect 1102 -2499 1104 -2497
rect 1110 -2499 1112 -2497
rect 1120 -2499 1122 -2497
rect 1128 -2499 1130 -2497
rect 1144 -2499 1146 -2497
rect 1152 -2499 1154 -2497
rect 1326 -2499 1328 -2497
rect 1336 -2499 1338 -2497
rect 1352 -2499 1354 -2497
rect 1360 -2499 1362 -2497
rect 1376 -2499 1378 -2497
rect 1384 -2499 1386 -2497
rect 1394 -2499 1396 -2497
rect 1402 -2499 1404 -2497
rect 1418 -2499 1420 -2497
rect 1426 -2499 1428 -2497
rect 1436 -2499 1438 -2497
rect 1444 -2499 1446 -2497
rect 1460 -2499 1462 -2497
rect 1468 -2499 1470 -2497
rect 1478 -2499 1480 -2497
rect 1486 -2499 1488 -2497
rect 1502 -2499 1504 -2497
rect 1510 -2499 1512 -2497
rect -1259 -2575 -1257 -2507
rect -1249 -2575 -1247 -2507
rect -1233 -2575 -1231 -2507
rect -1225 -2575 -1223 -2507
rect -1209 -2575 -1207 -2507
rect -1201 -2575 -1199 -2507
rect -1191 -2575 -1189 -2507
rect -1183 -2575 -1181 -2507
rect -1167 -2575 -1165 -2507
rect -1159 -2540 -1157 -2507
rect -1149 -2540 -1147 -2507
rect -1159 -2542 -1147 -2540
rect -1159 -2575 -1157 -2542
rect -1149 -2575 -1147 -2542
rect -1141 -2575 -1139 -2507
rect -1125 -2575 -1123 -2507
rect -1117 -2575 -1115 -2507
rect -1107 -2575 -1105 -2507
rect -1099 -2575 -1097 -2507
rect -1083 -2575 -1081 -2507
rect -1075 -2575 -1073 -2507
rect -930 -2575 -928 -2507
rect -920 -2575 -918 -2507
rect -904 -2575 -902 -2507
rect -896 -2575 -894 -2507
rect -880 -2575 -878 -2507
rect -872 -2575 -870 -2507
rect -862 -2575 -860 -2507
rect -854 -2575 -852 -2507
rect -838 -2575 -836 -2507
rect -830 -2540 -828 -2507
rect -820 -2540 -818 -2507
rect -830 -2542 -818 -2540
rect -830 -2575 -828 -2542
rect -820 -2575 -818 -2542
rect -812 -2575 -810 -2507
rect -796 -2575 -794 -2507
rect -788 -2575 -786 -2507
rect -778 -2575 -776 -2507
rect -770 -2575 -768 -2507
rect -754 -2575 -752 -2507
rect -746 -2575 -744 -2507
rect -572 -2575 -570 -2507
rect -562 -2575 -560 -2507
rect -546 -2575 -544 -2507
rect -538 -2575 -536 -2507
rect -522 -2575 -520 -2507
rect -514 -2575 -512 -2507
rect -504 -2575 -502 -2507
rect -496 -2575 -494 -2507
rect -480 -2575 -478 -2507
rect -472 -2540 -470 -2507
rect -462 -2540 -460 -2507
rect -472 -2542 -460 -2540
rect -472 -2575 -470 -2542
rect -462 -2575 -460 -2542
rect -454 -2575 -452 -2507
rect -438 -2575 -436 -2507
rect -430 -2575 -428 -2507
rect -420 -2575 -418 -2507
rect -412 -2575 -410 -2507
rect -396 -2575 -394 -2507
rect -388 -2575 -386 -2507
rect -214 -2575 -212 -2507
rect -204 -2575 -202 -2507
rect -188 -2575 -186 -2507
rect -180 -2575 -178 -2507
rect -164 -2575 -162 -2507
rect -156 -2575 -154 -2507
rect -146 -2575 -144 -2507
rect -138 -2575 -136 -2507
rect -122 -2575 -120 -2507
rect -114 -2540 -112 -2507
rect -104 -2540 -102 -2507
rect -114 -2542 -102 -2540
rect -114 -2575 -112 -2542
rect -104 -2575 -102 -2542
rect -96 -2575 -94 -2507
rect -80 -2575 -78 -2507
rect -72 -2575 -70 -2507
rect -62 -2575 -60 -2507
rect -54 -2575 -52 -2507
rect -38 -2575 -36 -2507
rect -30 -2575 -28 -2507
rect 95 -2563 97 -2531
rect 214 -2575 216 -2507
rect 224 -2575 226 -2507
rect 240 -2575 242 -2507
rect 248 -2575 250 -2507
rect 264 -2575 266 -2507
rect 272 -2575 274 -2507
rect 282 -2575 284 -2507
rect 290 -2575 292 -2507
rect 306 -2575 308 -2507
rect 314 -2540 316 -2507
rect 324 -2540 326 -2507
rect 314 -2542 326 -2540
rect 314 -2575 316 -2542
rect 324 -2575 326 -2542
rect 332 -2575 334 -2507
rect 348 -2575 350 -2507
rect 356 -2575 358 -2507
rect 366 -2575 368 -2507
rect 374 -2575 376 -2507
rect 390 -2575 392 -2507
rect 398 -2575 400 -2507
rect 570 -2575 572 -2507
rect 580 -2575 582 -2507
rect 596 -2575 598 -2507
rect 604 -2575 606 -2507
rect 620 -2575 622 -2507
rect 628 -2575 630 -2507
rect 638 -2575 640 -2507
rect 646 -2575 648 -2507
rect 662 -2575 664 -2507
rect 670 -2540 672 -2507
rect 680 -2540 682 -2507
rect 670 -2542 682 -2540
rect 670 -2575 672 -2542
rect 680 -2575 682 -2542
rect 688 -2575 690 -2507
rect 704 -2575 706 -2507
rect 712 -2575 714 -2507
rect 722 -2575 724 -2507
rect 730 -2575 732 -2507
rect 746 -2575 748 -2507
rect 754 -2575 756 -2507
rect 968 -2575 970 -2507
rect 978 -2575 980 -2507
rect 994 -2575 996 -2507
rect 1002 -2575 1004 -2507
rect 1018 -2575 1020 -2507
rect 1026 -2575 1028 -2507
rect 1036 -2575 1038 -2507
rect 1044 -2575 1046 -2507
rect 1060 -2575 1062 -2507
rect 1068 -2540 1070 -2507
rect 1078 -2540 1080 -2507
rect 1068 -2542 1080 -2540
rect 1068 -2575 1070 -2542
rect 1078 -2575 1080 -2542
rect 1086 -2575 1088 -2507
rect 1102 -2575 1104 -2507
rect 1110 -2575 1112 -2507
rect 1120 -2575 1122 -2507
rect 1128 -2575 1130 -2507
rect 1144 -2575 1146 -2507
rect 1152 -2575 1154 -2507
rect 1326 -2575 1328 -2507
rect 1336 -2575 1338 -2507
rect 1352 -2575 1354 -2507
rect 1360 -2575 1362 -2507
rect 1376 -2575 1378 -2507
rect 1384 -2575 1386 -2507
rect 1394 -2575 1396 -2507
rect 1402 -2575 1404 -2507
rect 1418 -2575 1420 -2507
rect 1426 -2540 1428 -2507
rect 1436 -2540 1438 -2507
rect 1426 -2542 1438 -2540
rect 1426 -2575 1428 -2542
rect 1436 -2575 1438 -2542
rect 1444 -2575 1446 -2507
rect 1460 -2575 1462 -2507
rect 1468 -2575 1470 -2507
rect 1478 -2575 1480 -2507
rect 1486 -2575 1488 -2507
rect 1502 -2575 1504 -2507
rect 1510 -2575 1512 -2507
rect -1259 -2581 -1257 -2579
rect -1249 -2581 -1247 -2579
rect -1233 -2581 -1231 -2579
rect -1225 -2581 -1223 -2579
rect -1209 -2581 -1207 -2579
rect -1201 -2581 -1199 -2579
rect -1191 -2581 -1189 -2579
rect -1183 -2581 -1181 -2579
rect -1167 -2581 -1165 -2579
rect -1159 -2581 -1157 -2579
rect -1149 -2581 -1147 -2579
rect -1141 -2581 -1139 -2579
rect -1125 -2581 -1123 -2579
rect -1117 -2581 -1115 -2579
rect -1107 -2581 -1105 -2579
rect -1099 -2581 -1097 -2579
rect -1083 -2581 -1081 -2579
rect -1075 -2581 -1073 -2579
rect -930 -2581 -928 -2579
rect -920 -2581 -918 -2579
rect -904 -2581 -902 -2579
rect -896 -2581 -894 -2579
rect -880 -2581 -878 -2579
rect -872 -2581 -870 -2579
rect -862 -2581 -860 -2579
rect -854 -2581 -852 -2579
rect -838 -2581 -836 -2579
rect -830 -2581 -828 -2579
rect -820 -2581 -818 -2579
rect -812 -2581 -810 -2579
rect -796 -2581 -794 -2579
rect -788 -2581 -786 -2579
rect -778 -2581 -776 -2579
rect -770 -2581 -768 -2579
rect -754 -2581 -752 -2579
rect -746 -2581 -744 -2579
rect -572 -2581 -570 -2579
rect -562 -2581 -560 -2579
rect -546 -2581 -544 -2579
rect -538 -2581 -536 -2579
rect -522 -2581 -520 -2579
rect -514 -2581 -512 -2579
rect -504 -2581 -502 -2579
rect -496 -2581 -494 -2579
rect -480 -2581 -478 -2579
rect -472 -2581 -470 -2579
rect -462 -2581 -460 -2579
rect -454 -2581 -452 -2579
rect -438 -2581 -436 -2579
rect -430 -2581 -428 -2579
rect -420 -2581 -418 -2579
rect -412 -2581 -410 -2579
rect -396 -2581 -394 -2579
rect -388 -2581 -386 -2579
rect -214 -2581 -212 -2579
rect -204 -2581 -202 -2579
rect -188 -2581 -186 -2579
rect -180 -2581 -178 -2579
rect -164 -2581 -162 -2579
rect -156 -2581 -154 -2579
rect -146 -2581 -144 -2579
rect -138 -2581 -136 -2579
rect -122 -2581 -120 -2579
rect -114 -2581 -112 -2579
rect -104 -2581 -102 -2579
rect -96 -2581 -94 -2579
rect -80 -2581 -78 -2579
rect -72 -2581 -70 -2579
rect -62 -2581 -60 -2579
rect -54 -2581 -52 -2579
rect -38 -2581 -36 -2579
rect -30 -2581 -28 -2579
rect 95 -2581 97 -2579
rect 214 -2581 216 -2579
rect 224 -2581 226 -2579
rect 240 -2581 242 -2579
rect 248 -2581 250 -2579
rect 264 -2581 266 -2579
rect 272 -2581 274 -2579
rect 282 -2581 284 -2579
rect 290 -2581 292 -2579
rect 306 -2581 308 -2579
rect 314 -2581 316 -2579
rect 324 -2581 326 -2579
rect 332 -2581 334 -2579
rect 348 -2581 350 -2579
rect 356 -2581 358 -2579
rect 366 -2581 368 -2579
rect 374 -2581 376 -2579
rect 390 -2581 392 -2579
rect 398 -2581 400 -2579
rect 570 -2581 572 -2579
rect 580 -2581 582 -2579
rect 596 -2581 598 -2579
rect 604 -2581 606 -2579
rect 620 -2581 622 -2579
rect 628 -2581 630 -2579
rect 638 -2581 640 -2579
rect 646 -2581 648 -2579
rect 662 -2581 664 -2579
rect 670 -2581 672 -2579
rect 680 -2581 682 -2579
rect 688 -2581 690 -2579
rect 704 -2581 706 -2579
rect 712 -2581 714 -2579
rect 722 -2581 724 -2579
rect 730 -2581 732 -2579
rect 746 -2581 748 -2579
rect 754 -2581 756 -2579
rect 968 -2581 970 -2579
rect 978 -2581 980 -2579
rect 994 -2581 996 -2579
rect 1002 -2581 1004 -2579
rect 1018 -2581 1020 -2579
rect 1026 -2581 1028 -2579
rect 1036 -2581 1038 -2579
rect 1044 -2581 1046 -2579
rect 1060 -2581 1062 -2579
rect 1068 -2581 1070 -2579
rect 1078 -2581 1080 -2579
rect 1086 -2581 1088 -2579
rect 1102 -2581 1104 -2579
rect 1110 -2581 1112 -2579
rect 1120 -2581 1122 -2579
rect 1128 -2581 1130 -2579
rect 1144 -2581 1146 -2579
rect 1152 -2581 1154 -2579
rect 1326 -2581 1328 -2579
rect 1336 -2581 1338 -2579
rect 1352 -2581 1354 -2579
rect 1360 -2581 1362 -2579
rect 1376 -2581 1378 -2579
rect 1384 -2581 1386 -2579
rect 1394 -2581 1396 -2579
rect 1402 -2581 1404 -2579
rect 1418 -2581 1420 -2579
rect 1426 -2581 1428 -2579
rect 1436 -2581 1438 -2579
rect 1444 -2581 1446 -2579
rect 1460 -2581 1462 -2579
rect 1468 -2581 1470 -2579
rect 1478 -2581 1480 -2579
rect 1486 -2581 1488 -2579
rect 1502 -2581 1504 -2579
rect 1510 -2581 1512 -2579
rect -1259 -2611 -1257 -2609
rect -1249 -2611 -1247 -2609
rect -1233 -2611 -1231 -2609
rect -1225 -2611 -1223 -2609
rect -1209 -2611 -1207 -2609
rect -1201 -2611 -1199 -2609
rect -1191 -2611 -1189 -2609
rect -1183 -2611 -1181 -2609
rect -1167 -2611 -1165 -2609
rect -1159 -2611 -1157 -2609
rect -1149 -2611 -1147 -2609
rect -1141 -2611 -1139 -2609
rect -1125 -2611 -1123 -2609
rect -1117 -2611 -1115 -2609
rect -1107 -2611 -1105 -2609
rect -1099 -2611 -1097 -2609
rect -1083 -2611 -1081 -2609
rect -1075 -2611 -1073 -2609
rect -930 -2611 -928 -2609
rect -920 -2611 -918 -2609
rect -904 -2611 -902 -2609
rect -896 -2611 -894 -2609
rect -880 -2611 -878 -2609
rect -872 -2611 -870 -2609
rect -862 -2611 -860 -2609
rect -854 -2611 -852 -2609
rect -838 -2611 -836 -2609
rect -830 -2611 -828 -2609
rect -820 -2611 -818 -2609
rect -812 -2611 -810 -2609
rect -796 -2611 -794 -2609
rect -788 -2611 -786 -2609
rect -778 -2611 -776 -2609
rect -770 -2611 -768 -2609
rect -754 -2611 -752 -2609
rect -746 -2611 -744 -2609
rect -1259 -2687 -1257 -2619
rect -1249 -2687 -1247 -2619
rect -1233 -2687 -1231 -2619
rect -1225 -2687 -1223 -2619
rect -1209 -2687 -1207 -2619
rect -1201 -2687 -1199 -2619
rect -1191 -2687 -1189 -2619
rect -1183 -2687 -1181 -2619
rect -1167 -2687 -1165 -2619
rect -1159 -2652 -1157 -2619
rect -1149 -2652 -1147 -2619
rect -1159 -2654 -1147 -2652
rect -1159 -2687 -1157 -2654
rect -1149 -2687 -1147 -2654
rect -1141 -2687 -1139 -2619
rect -1125 -2687 -1123 -2619
rect -1117 -2687 -1115 -2619
rect -1107 -2687 -1105 -2619
rect -1099 -2687 -1097 -2619
rect -1083 -2687 -1081 -2619
rect -1075 -2687 -1073 -2619
rect -930 -2687 -928 -2619
rect -920 -2687 -918 -2619
rect -904 -2687 -902 -2619
rect -896 -2687 -894 -2619
rect -880 -2687 -878 -2619
rect -872 -2687 -870 -2619
rect -862 -2687 -860 -2619
rect -854 -2687 -852 -2619
rect -838 -2687 -836 -2619
rect -830 -2652 -828 -2619
rect -820 -2652 -818 -2619
rect -830 -2654 -818 -2652
rect -830 -2687 -828 -2654
rect -820 -2687 -818 -2654
rect -812 -2687 -810 -2619
rect -796 -2687 -794 -2619
rect -788 -2687 -786 -2619
rect -778 -2687 -776 -2619
rect -770 -2687 -768 -2619
rect -754 -2687 -752 -2619
rect -746 -2687 -744 -2619
rect -1259 -2693 -1257 -2691
rect -1249 -2693 -1247 -2691
rect -1233 -2693 -1231 -2691
rect -1225 -2693 -1223 -2691
rect -1209 -2693 -1207 -2691
rect -1201 -2693 -1199 -2691
rect -1191 -2693 -1189 -2691
rect -1183 -2693 -1181 -2691
rect -1167 -2693 -1165 -2691
rect -1159 -2693 -1157 -2691
rect -1149 -2693 -1147 -2691
rect -1141 -2693 -1139 -2691
rect -1125 -2693 -1123 -2691
rect -1117 -2693 -1115 -2691
rect -1107 -2693 -1105 -2691
rect -1099 -2693 -1097 -2691
rect -1083 -2693 -1081 -2691
rect -1075 -2693 -1073 -2691
rect -930 -2693 -928 -2691
rect -920 -2693 -918 -2691
rect -904 -2693 -902 -2691
rect -896 -2693 -894 -2691
rect -880 -2693 -878 -2691
rect -872 -2693 -870 -2691
rect -862 -2693 -860 -2691
rect -854 -2693 -852 -2691
rect -838 -2693 -836 -2691
rect -830 -2693 -828 -2691
rect -820 -2693 -818 -2691
rect -812 -2693 -810 -2691
rect -796 -2693 -794 -2691
rect -788 -2693 -786 -2691
rect -778 -2693 -776 -2691
rect -770 -2693 -768 -2691
rect -754 -2693 -752 -2691
rect -746 -2693 -744 -2691
rect -1334 -2724 -1332 -2722
rect -1326 -2724 -1324 -2722
rect -1316 -2724 -1314 -2722
rect -930 -2724 -928 -2722
rect -922 -2724 -920 -2722
rect -912 -2724 -910 -2722
rect -572 -2724 -570 -2722
rect -564 -2724 -562 -2722
rect -554 -2724 -552 -2722
rect -214 -2724 -212 -2722
rect -206 -2724 -204 -2722
rect -196 -2724 -194 -2722
rect 214 -2724 216 -2722
rect 222 -2724 224 -2722
rect 232 -2724 234 -2722
rect 570 -2724 572 -2722
rect 578 -2724 580 -2722
rect 588 -2724 590 -2722
rect 968 -2724 970 -2722
rect 976 -2724 978 -2722
rect 986 -2724 988 -2722
rect 1326 -2724 1328 -2722
rect 1334 -2724 1336 -2722
rect 1344 -2724 1346 -2722
rect -1334 -2800 -1332 -2732
rect -1326 -2756 -1324 -2732
rect -1326 -2800 -1324 -2760
rect -1316 -2800 -1314 -2732
rect -930 -2800 -928 -2732
rect -922 -2756 -920 -2732
rect -922 -2800 -920 -2760
rect -912 -2800 -910 -2732
rect -572 -2800 -570 -2732
rect -564 -2756 -562 -2732
rect -564 -2800 -562 -2760
rect -554 -2800 -552 -2732
rect -214 -2800 -212 -2732
rect -206 -2756 -204 -2732
rect -206 -2800 -204 -2760
rect -196 -2800 -194 -2732
rect 214 -2800 216 -2732
rect 222 -2756 224 -2732
rect 222 -2800 224 -2760
rect 232 -2800 234 -2732
rect 570 -2800 572 -2732
rect 578 -2756 580 -2732
rect 578 -2800 580 -2760
rect 588 -2800 590 -2732
rect 968 -2800 970 -2732
rect 976 -2756 978 -2732
rect 976 -2800 978 -2760
rect 986 -2800 988 -2732
rect 1326 -2800 1328 -2732
rect 1334 -2756 1336 -2732
rect 1334 -2800 1336 -2760
rect 1344 -2800 1346 -2732
rect -1334 -2806 -1332 -2804
rect -1326 -2806 -1324 -2804
rect -1316 -2806 -1314 -2804
rect -930 -2806 -928 -2804
rect -922 -2806 -920 -2804
rect -912 -2806 -910 -2804
rect -572 -2806 -570 -2804
rect -564 -2806 -562 -2804
rect -554 -2806 -552 -2804
rect -214 -2806 -212 -2804
rect -206 -2806 -204 -2804
rect -196 -2806 -194 -2804
rect 214 -2806 216 -2804
rect 222 -2806 224 -2804
rect 232 -2806 234 -2804
rect 570 -2806 572 -2804
rect 578 -2806 580 -2804
rect 588 -2806 590 -2804
rect 968 -2806 970 -2804
rect 976 -2806 978 -2804
rect 986 -2806 988 -2804
rect 1326 -2806 1328 -2804
rect 1334 -2806 1336 -2804
rect 1344 -2806 1346 -2804
rect -1259 -2843 -1257 -2841
rect -1249 -2843 -1247 -2841
rect -1233 -2843 -1231 -2841
rect -1223 -2843 -1221 -2841
rect -1215 -2843 -1213 -2841
rect -1205 -2843 -1203 -2841
rect -1189 -2843 -1187 -2841
rect -1181 -2843 -1179 -2841
rect -1171 -2843 -1169 -2841
rect -930 -2843 -928 -2841
rect -920 -2843 -918 -2841
rect -904 -2843 -902 -2841
rect -894 -2843 -892 -2841
rect -878 -2843 -876 -2841
rect -868 -2843 -866 -2841
rect -860 -2843 -858 -2841
rect -850 -2843 -848 -2841
rect -834 -2843 -832 -2841
rect -826 -2843 -824 -2841
rect -816 -2843 -814 -2841
rect -800 -2843 -798 -2841
rect -790 -2843 -788 -2841
rect -782 -2843 -780 -2841
rect -772 -2843 -770 -2841
rect -756 -2843 -754 -2841
rect -748 -2843 -746 -2841
rect -732 -2843 -730 -2841
rect -716 -2843 -714 -2841
rect -708 -2843 -706 -2841
rect -698 -2843 -696 -2841
rect -572 -2843 -570 -2841
rect -562 -2843 -560 -2841
rect -546 -2843 -544 -2841
rect -536 -2843 -534 -2841
rect -520 -2843 -518 -2841
rect -510 -2843 -508 -2841
rect -502 -2843 -500 -2841
rect -492 -2843 -490 -2841
rect -476 -2843 -474 -2841
rect -468 -2843 -466 -2841
rect -458 -2843 -456 -2841
rect -442 -2843 -440 -2841
rect -432 -2843 -430 -2841
rect -424 -2843 -422 -2841
rect -414 -2843 -412 -2841
rect -398 -2843 -396 -2841
rect -390 -2843 -388 -2841
rect -374 -2843 -372 -2841
rect -358 -2843 -356 -2841
rect -350 -2843 -348 -2841
rect -340 -2843 -338 -2841
rect -214 -2843 -212 -2841
rect -204 -2843 -202 -2841
rect -188 -2843 -186 -2841
rect -178 -2843 -176 -2841
rect -162 -2843 -160 -2841
rect -152 -2843 -150 -2841
rect -144 -2843 -142 -2841
rect -134 -2843 -132 -2841
rect -118 -2843 -116 -2841
rect -110 -2843 -108 -2841
rect -100 -2843 -98 -2841
rect -84 -2843 -82 -2841
rect -74 -2843 -72 -2841
rect -66 -2843 -64 -2841
rect -56 -2843 -54 -2841
rect -40 -2843 -38 -2841
rect -32 -2843 -30 -2841
rect -16 -2843 -14 -2841
rect 0 -2843 2 -2841
rect 8 -2843 10 -2841
rect 18 -2843 20 -2841
rect 214 -2843 216 -2841
rect 224 -2843 226 -2841
rect 240 -2843 242 -2841
rect 250 -2843 252 -2841
rect 266 -2843 268 -2841
rect 276 -2843 278 -2841
rect 284 -2843 286 -2841
rect 294 -2843 296 -2841
rect 310 -2843 312 -2841
rect 318 -2843 320 -2841
rect 328 -2843 330 -2841
rect 344 -2843 346 -2841
rect 354 -2843 356 -2841
rect 362 -2843 364 -2841
rect 372 -2843 374 -2841
rect 388 -2843 390 -2841
rect 396 -2843 398 -2841
rect 412 -2843 414 -2841
rect 428 -2843 430 -2841
rect 436 -2843 438 -2841
rect 446 -2843 448 -2841
rect 570 -2843 572 -2841
rect 580 -2843 582 -2841
rect 596 -2843 598 -2841
rect 606 -2843 608 -2841
rect 622 -2843 624 -2841
rect 632 -2843 634 -2841
rect 640 -2843 642 -2841
rect 650 -2843 652 -2841
rect 666 -2843 668 -2841
rect 674 -2843 676 -2841
rect 684 -2843 686 -2841
rect 700 -2843 702 -2841
rect 710 -2843 712 -2841
rect 718 -2843 720 -2841
rect 728 -2843 730 -2841
rect 744 -2843 746 -2841
rect 752 -2843 754 -2841
rect 768 -2843 770 -2841
rect 784 -2843 786 -2841
rect 792 -2843 794 -2841
rect 802 -2843 804 -2841
rect 968 -2843 970 -2841
rect 978 -2843 980 -2841
rect 994 -2843 996 -2841
rect 1004 -2843 1006 -2841
rect 1020 -2843 1022 -2841
rect 1030 -2843 1032 -2841
rect 1038 -2843 1040 -2841
rect 1048 -2843 1050 -2841
rect 1064 -2843 1066 -2841
rect 1072 -2843 1074 -2841
rect 1082 -2843 1084 -2841
rect 1098 -2843 1100 -2841
rect 1108 -2843 1110 -2841
rect 1116 -2843 1118 -2841
rect 1126 -2843 1128 -2841
rect 1142 -2843 1144 -2841
rect 1150 -2843 1152 -2841
rect 1166 -2843 1168 -2841
rect 1182 -2843 1184 -2841
rect 1190 -2843 1192 -2841
rect 1200 -2843 1202 -2841
rect 1326 -2843 1328 -2841
rect 1336 -2843 1338 -2841
rect 1352 -2843 1354 -2841
rect 1362 -2843 1364 -2841
rect 1378 -2843 1380 -2841
rect 1388 -2843 1390 -2841
rect 1396 -2843 1398 -2841
rect 1406 -2843 1408 -2841
rect 1422 -2843 1424 -2841
rect 1430 -2843 1432 -2841
rect 1440 -2843 1442 -2841
rect 1456 -2843 1458 -2841
rect 1466 -2843 1468 -2841
rect 1474 -2843 1476 -2841
rect 1484 -2843 1486 -2841
rect 1500 -2843 1502 -2841
rect 1508 -2843 1510 -2841
rect 1524 -2843 1526 -2841
rect 1540 -2843 1542 -2841
rect 1548 -2843 1550 -2841
rect 1558 -2843 1560 -2841
rect -1259 -2919 -1257 -2851
rect -1249 -2919 -1247 -2851
rect -1233 -2919 -1231 -2851
rect -1223 -2919 -1221 -2851
rect -1215 -2919 -1213 -2851
rect -1205 -2919 -1203 -2851
rect -1189 -2919 -1187 -2851
rect -1181 -2919 -1179 -2851
rect -1171 -2919 -1169 -2851
rect -930 -2919 -928 -2851
rect -920 -2919 -918 -2851
rect -904 -2919 -902 -2851
rect -894 -2919 -892 -2851
rect -878 -2919 -876 -2851
rect -868 -2919 -866 -2851
rect -860 -2919 -858 -2851
rect -850 -2919 -848 -2851
rect -834 -2919 -832 -2851
rect -826 -2919 -824 -2851
rect -816 -2919 -814 -2851
rect -800 -2919 -798 -2851
rect -790 -2919 -788 -2851
rect -782 -2919 -780 -2851
rect -772 -2919 -770 -2851
rect -756 -2919 -754 -2851
rect -748 -2919 -746 -2851
rect -732 -2919 -730 -2851
rect -716 -2919 -714 -2851
rect -708 -2919 -706 -2851
rect -698 -2919 -696 -2851
rect -572 -2919 -570 -2851
rect -562 -2919 -560 -2851
rect -546 -2919 -544 -2851
rect -536 -2919 -534 -2851
rect -520 -2919 -518 -2851
rect -510 -2919 -508 -2851
rect -502 -2919 -500 -2851
rect -492 -2919 -490 -2851
rect -476 -2919 -474 -2851
rect -468 -2919 -466 -2851
rect -458 -2919 -456 -2851
rect -442 -2919 -440 -2851
rect -432 -2919 -430 -2851
rect -424 -2919 -422 -2851
rect -414 -2919 -412 -2851
rect -398 -2919 -396 -2851
rect -390 -2919 -388 -2851
rect -374 -2919 -372 -2851
rect -358 -2919 -356 -2851
rect -350 -2919 -348 -2851
rect -340 -2919 -338 -2851
rect -214 -2919 -212 -2851
rect -204 -2919 -202 -2851
rect -188 -2919 -186 -2851
rect -178 -2919 -176 -2851
rect -162 -2919 -160 -2851
rect -152 -2919 -150 -2851
rect -144 -2919 -142 -2851
rect -134 -2919 -132 -2851
rect -118 -2919 -116 -2851
rect -110 -2919 -108 -2851
rect -100 -2919 -98 -2851
rect -84 -2919 -82 -2851
rect -74 -2919 -72 -2851
rect -66 -2919 -64 -2851
rect -56 -2919 -54 -2851
rect -40 -2919 -38 -2851
rect -32 -2919 -30 -2851
rect -16 -2919 -14 -2851
rect 0 -2919 2 -2851
rect 8 -2919 10 -2851
rect 18 -2919 20 -2851
rect 214 -2919 216 -2851
rect 224 -2919 226 -2851
rect 240 -2919 242 -2851
rect 250 -2919 252 -2851
rect 266 -2919 268 -2851
rect 276 -2919 278 -2851
rect 284 -2919 286 -2851
rect 294 -2919 296 -2851
rect 310 -2919 312 -2851
rect 318 -2919 320 -2851
rect 328 -2919 330 -2851
rect 344 -2919 346 -2851
rect 354 -2919 356 -2851
rect 362 -2919 364 -2851
rect 372 -2919 374 -2851
rect 388 -2919 390 -2851
rect 396 -2919 398 -2851
rect 412 -2919 414 -2851
rect 428 -2919 430 -2851
rect 436 -2919 438 -2851
rect 446 -2919 448 -2851
rect 570 -2919 572 -2851
rect 580 -2919 582 -2851
rect 596 -2919 598 -2851
rect 606 -2919 608 -2851
rect 622 -2919 624 -2851
rect 632 -2919 634 -2851
rect 640 -2919 642 -2851
rect 650 -2919 652 -2851
rect 666 -2919 668 -2851
rect 674 -2919 676 -2851
rect 684 -2919 686 -2851
rect 700 -2919 702 -2851
rect 710 -2919 712 -2851
rect 718 -2919 720 -2851
rect 728 -2919 730 -2851
rect 744 -2919 746 -2851
rect 752 -2919 754 -2851
rect 768 -2919 770 -2851
rect 784 -2919 786 -2851
rect 792 -2919 794 -2851
rect 802 -2919 804 -2851
rect 968 -2919 970 -2851
rect 978 -2919 980 -2851
rect 994 -2919 996 -2851
rect 1004 -2919 1006 -2851
rect 1020 -2919 1022 -2851
rect 1030 -2919 1032 -2851
rect 1038 -2919 1040 -2851
rect 1048 -2919 1050 -2851
rect 1064 -2919 1066 -2851
rect 1072 -2919 1074 -2851
rect 1082 -2919 1084 -2851
rect 1098 -2919 1100 -2851
rect 1108 -2919 1110 -2851
rect 1116 -2919 1118 -2851
rect 1126 -2919 1128 -2851
rect 1142 -2919 1144 -2851
rect 1150 -2919 1152 -2851
rect 1166 -2919 1168 -2851
rect 1182 -2919 1184 -2851
rect 1190 -2919 1192 -2851
rect 1200 -2919 1202 -2851
rect 1326 -2919 1328 -2851
rect 1336 -2919 1338 -2851
rect 1352 -2919 1354 -2851
rect 1362 -2919 1364 -2851
rect 1378 -2919 1380 -2851
rect 1388 -2919 1390 -2851
rect 1396 -2919 1398 -2851
rect 1406 -2919 1408 -2851
rect 1422 -2919 1424 -2851
rect 1430 -2919 1432 -2851
rect 1440 -2919 1442 -2851
rect 1456 -2919 1458 -2851
rect 1466 -2919 1468 -2851
rect 1474 -2919 1476 -2851
rect 1484 -2919 1486 -2851
rect 1500 -2919 1502 -2851
rect 1508 -2919 1510 -2851
rect 1524 -2919 1526 -2851
rect 1540 -2919 1542 -2851
rect 1548 -2919 1550 -2851
rect 1558 -2919 1560 -2851
rect -1259 -2925 -1257 -2923
rect -1249 -2925 -1247 -2923
rect -1233 -2925 -1231 -2923
rect -1223 -2925 -1221 -2923
rect -1215 -2925 -1213 -2923
rect -1205 -2925 -1203 -2923
rect -1189 -2925 -1187 -2923
rect -1181 -2925 -1179 -2923
rect -1171 -2925 -1169 -2923
rect -930 -2925 -928 -2923
rect -920 -2925 -918 -2923
rect -904 -2925 -902 -2923
rect -894 -2925 -892 -2923
rect -878 -2925 -876 -2923
rect -868 -2925 -866 -2923
rect -860 -2925 -858 -2923
rect -850 -2925 -848 -2923
rect -834 -2925 -832 -2923
rect -826 -2925 -824 -2923
rect -816 -2925 -814 -2923
rect -800 -2925 -798 -2923
rect -790 -2925 -788 -2923
rect -782 -2925 -780 -2923
rect -772 -2925 -770 -2923
rect -756 -2925 -754 -2923
rect -748 -2925 -746 -2923
rect -732 -2925 -730 -2923
rect -716 -2925 -714 -2923
rect -708 -2925 -706 -2923
rect -698 -2925 -696 -2923
rect -572 -2925 -570 -2923
rect -562 -2925 -560 -2923
rect -546 -2925 -544 -2923
rect -536 -2925 -534 -2923
rect -520 -2925 -518 -2923
rect -510 -2925 -508 -2923
rect -502 -2925 -500 -2923
rect -492 -2925 -490 -2923
rect -476 -2925 -474 -2923
rect -468 -2925 -466 -2923
rect -458 -2925 -456 -2923
rect -442 -2925 -440 -2923
rect -432 -2925 -430 -2923
rect -424 -2925 -422 -2923
rect -414 -2925 -412 -2923
rect -398 -2925 -396 -2923
rect -390 -2925 -388 -2923
rect -374 -2925 -372 -2923
rect -358 -2925 -356 -2923
rect -350 -2925 -348 -2923
rect -340 -2925 -338 -2923
rect -214 -2925 -212 -2923
rect -204 -2925 -202 -2923
rect -188 -2925 -186 -2923
rect -178 -2925 -176 -2923
rect -162 -2925 -160 -2923
rect -152 -2925 -150 -2923
rect -144 -2925 -142 -2923
rect -134 -2925 -132 -2923
rect -118 -2925 -116 -2923
rect -110 -2925 -108 -2923
rect -100 -2925 -98 -2923
rect -84 -2925 -82 -2923
rect -74 -2925 -72 -2923
rect -66 -2925 -64 -2923
rect -56 -2925 -54 -2923
rect -40 -2925 -38 -2923
rect -32 -2925 -30 -2923
rect -16 -2925 -14 -2923
rect 0 -2925 2 -2923
rect 8 -2925 10 -2923
rect 18 -2925 20 -2923
rect 214 -2925 216 -2923
rect 224 -2925 226 -2923
rect 240 -2925 242 -2923
rect 250 -2925 252 -2923
rect 266 -2925 268 -2923
rect 276 -2925 278 -2923
rect 284 -2925 286 -2923
rect 294 -2925 296 -2923
rect 310 -2925 312 -2923
rect 318 -2925 320 -2923
rect 328 -2925 330 -2923
rect 344 -2925 346 -2923
rect 354 -2925 356 -2923
rect 362 -2925 364 -2923
rect 372 -2925 374 -2923
rect 388 -2925 390 -2923
rect 396 -2925 398 -2923
rect 412 -2925 414 -2923
rect 428 -2925 430 -2923
rect 436 -2925 438 -2923
rect 446 -2925 448 -2923
rect 570 -2925 572 -2923
rect 580 -2925 582 -2923
rect 596 -2925 598 -2923
rect 606 -2925 608 -2923
rect 622 -2925 624 -2923
rect 632 -2925 634 -2923
rect 640 -2925 642 -2923
rect 650 -2925 652 -2923
rect 666 -2925 668 -2923
rect 674 -2925 676 -2923
rect 684 -2925 686 -2923
rect 700 -2925 702 -2923
rect 710 -2925 712 -2923
rect 718 -2925 720 -2923
rect 728 -2925 730 -2923
rect 744 -2925 746 -2923
rect 752 -2925 754 -2923
rect 768 -2925 770 -2923
rect 784 -2925 786 -2923
rect 792 -2925 794 -2923
rect 802 -2925 804 -2923
rect 968 -2925 970 -2923
rect 978 -2925 980 -2923
rect 994 -2925 996 -2923
rect 1004 -2925 1006 -2923
rect 1020 -2925 1022 -2923
rect 1030 -2925 1032 -2923
rect 1038 -2925 1040 -2923
rect 1048 -2925 1050 -2923
rect 1064 -2925 1066 -2923
rect 1072 -2925 1074 -2923
rect 1082 -2925 1084 -2923
rect 1098 -2925 1100 -2923
rect 1108 -2925 1110 -2923
rect 1116 -2925 1118 -2923
rect 1126 -2925 1128 -2923
rect 1142 -2925 1144 -2923
rect 1150 -2925 1152 -2923
rect 1166 -2925 1168 -2923
rect 1182 -2925 1184 -2923
rect 1190 -2925 1192 -2923
rect 1200 -2925 1202 -2923
rect 1326 -2925 1328 -2923
rect 1336 -2925 1338 -2923
rect 1352 -2925 1354 -2923
rect 1362 -2925 1364 -2923
rect 1378 -2925 1380 -2923
rect 1388 -2925 1390 -2923
rect 1396 -2925 1398 -2923
rect 1406 -2925 1408 -2923
rect 1422 -2925 1424 -2923
rect 1430 -2925 1432 -2923
rect 1440 -2925 1442 -2923
rect 1456 -2925 1458 -2923
rect 1466 -2925 1468 -2923
rect 1474 -2925 1476 -2923
rect 1484 -2925 1486 -2923
rect 1500 -2925 1502 -2923
rect 1508 -2925 1510 -2923
rect 1524 -2925 1526 -2923
rect 1540 -2925 1542 -2923
rect 1548 -2925 1550 -2923
rect 1558 -2925 1560 -2923
rect -1259 -2962 -1257 -2960
rect -1249 -2962 -1247 -2960
rect -1233 -2962 -1231 -2960
rect -1225 -2962 -1223 -2960
rect -1209 -2962 -1207 -2960
rect -1201 -2962 -1199 -2960
rect -1191 -2962 -1189 -2960
rect -1183 -2962 -1181 -2960
rect -1167 -2962 -1165 -2960
rect -1159 -2962 -1157 -2960
rect -1149 -2962 -1147 -2960
rect -1141 -2962 -1139 -2960
rect -1125 -2962 -1123 -2960
rect -1117 -2962 -1115 -2960
rect -1107 -2962 -1105 -2960
rect -1099 -2962 -1097 -2960
rect -1083 -2962 -1081 -2960
rect -1075 -2962 -1073 -2960
rect -1021 -2962 -1019 -2960
rect -930 -2962 -928 -2960
rect -920 -2962 -918 -2960
rect -904 -2962 -902 -2960
rect -896 -2962 -894 -2960
rect -880 -2962 -878 -2960
rect -872 -2962 -870 -2960
rect -862 -2962 -860 -2960
rect -854 -2962 -852 -2960
rect -838 -2962 -836 -2960
rect -830 -2962 -828 -2960
rect -820 -2962 -818 -2960
rect -812 -2962 -810 -2960
rect -796 -2962 -794 -2960
rect -788 -2962 -786 -2960
rect -778 -2962 -776 -2960
rect -770 -2962 -768 -2960
rect -754 -2962 -752 -2960
rect -746 -2962 -744 -2960
rect -667 -2962 -665 -2960
rect -572 -2962 -570 -2960
rect -562 -2962 -560 -2960
rect -546 -2962 -544 -2960
rect -538 -2962 -536 -2960
rect -522 -2962 -520 -2960
rect -514 -2962 -512 -2960
rect -504 -2962 -502 -2960
rect -496 -2962 -494 -2960
rect -480 -2962 -478 -2960
rect -472 -2962 -470 -2960
rect -462 -2962 -460 -2960
rect -454 -2962 -452 -2960
rect -438 -2962 -436 -2960
rect -430 -2962 -428 -2960
rect -420 -2962 -418 -2960
rect -412 -2962 -410 -2960
rect -396 -2962 -394 -2960
rect -388 -2962 -386 -2960
rect -324 -2962 -322 -2960
rect -214 -2962 -212 -2960
rect -204 -2962 -202 -2960
rect -188 -2962 -186 -2960
rect -180 -2962 -178 -2960
rect -164 -2962 -162 -2960
rect -156 -2962 -154 -2960
rect -146 -2962 -144 -2960
rect -138 -2962 -136 -2960
rect -122 -2962 -120 -2960
rect -114 -2962 -112 -2960
rect -104 -2962 -102 -2960
rect -96 -2962 -94 -2960
rect -80 -2962 -78 -2960
rect -72 -2962 -70 -2960
rect -62 -2962 -60 -2960
rect -54 -2962 -52 -2960
rect -38 -2962 -36 -2960
rect -30 -2962 -28 -2960
rect 214 -2962 216 -2960
rect 224 -2962 226 -2960
rect 240 -2962 242 -2960
rect 248 -2962 250 -2960
rect 264 -2962 266 -2960
rect 272 -2962 274 -2960
rect 282 -2962 284 -2960
rect 290 -2962 292 -2960
rect 306 -2962 308 -2960
rect 314 -2962 316 -2960
rect 324 -2962 326 -2960
rect 332 -2962 334 -2960
rect 348 -2962 350 -2960
rect 356 -2962 358 -2960
rect 366 -2962 368 -2960
rect 374 -2962 376 -2960
rect 390 -2962 392 -2960
rect 398 -2962 400 -2960
rect 477 -2962 479 -2960
rect 846 -2962 848 -2960
rect 1204 -2962 1206 -2960
rect -1259 -3038 -1257 -2970
rect -1249 -3038 -1247 -2970
rect -1233 -3038 -1231 -2970
rect -1225 -3038 -1223 -2970
rect -1209 -3038 -1207 -2970
rect -1201 -3038 -1199 -2970
rect -1191 -3038 -1189 -2970
rect -1183 -3038 -1181 -2970
rect -1167 -3038 -1165 -2970
rect -1159 -3003 -1157 -2970
rect -1149 -3003 -1147 -2970
rect -1159 -3005 -1147 -3003
rect -1159 -3038 -1157 -3005
rect -1149 -3038 -1147 -3005
rect -1141 -3038 -1139 -2970
rect -1125 -3038 -1123 -2970
rect -1117 -3038 -1115 -2970
rect -1107 -3038 -1105 -2970
rect -1099 -3038 -1097 -2970
rect -1083 -3038 -1081 -2970
rect -1075 -3038 -1073 -2970
rect -1021 -3038 -1019 -2970
rect -930 -3038 -928 -2970
rect -920 -3038 -918 -2970
rect -904 -3038 -902 -2970
rect -896 -3038 -894 -2970
rect -880 -3038 -878 -2970
rect -872 -3038 -870 -2970
rect -862 -3038 -860 -2970
rect -854 -3038 -852 -2970
rect -838 -3038 -836 -2970
rect -830 -3003 -828 -2970
rect -820 -3003 -818 -2970
rect -830 -3005 -818 -3003
rect -830 -3038 -828 -3005
rect -820 -3038 -818 -3005
rect -812 -3038 -810 -2970
rect -796 -3038 -794 -2970
rect -788 -3038 -786 -2970
rect -778 -3038 -776 -2970
rect -770 -3038 -768 -2970
rect -754 -3038 -752 -2970
rect -746 -3038 -744 -2970
rect -667 -3034 -665 -2978
rect -572 -3038 -570 -2970
rect -562 -3038 -560 -2970
rect -546 -3038 -544 -2970
rect -538 -3038 -536 -2970
rect -522 -3038 -520 -2970
rect -514 -3038 -512 -2970
rect -504 -3038 -502 -2970
rect -496 -3038 -494 -2970
rect -480 -3038 -478 -2970
rect -472 -3003 -470 -2970
rect -462 -3003 -460 -2970
rect -472 -3005 -460 -3003
rect -472 -3038 -470 -3005
rect -462 -3038 -460 -3005
rect -454 -3038 -452 -2970
rect -438 -3038 -436 -2970
rect -430 -3038 -428 -2970
rect -420 -3038 -418 -2970
rect -412 -3038 -410 -2970
rect -396 -3038 -394 -2970
rect -388 -3038 -386 -2970
rect -324 -3038 -322 -2970
rect -214 -3038 -212 -2970
rect -204 -3038 -202 -2970
rect -188 -3038 -186 -2970
rect -180 -3038 -178 -2970
rect -164 -3038 -162 -2970
rect -156 -3038 -154 -2970
rect -146 -3038 -144 -2970
rect -138 -3038 -136 -2970
rect -122 -3038 -120 -2970
rect -114 -3003 -112 -2970
rect -104 -3003 -102 -2970
rect -114 -3005 -102 -3003
rect -114 -3038 -112 -3005
rect -104 -3038 -102 -3005
rect -96 -3038 -94 -2970
rect -80 -3038 -78 -2970
rect -72 -3038 -70 -2970
rect -62 -3038 -60 -2970
rect -54 -3038 -52 -2970
rect -38 -3038 -36 -2970
rect -30 -3038 -28 -2970
rect 214 -3038 216 -2970
rect 224 -3038 226 -2970
rect 240 -3038 242 -2970
rect 248 -3038 250 -2970
rect 264 -3038 266 -2970
rect 272 -3038 274 -2970
rect 282 -3038 284 -2970
rect 290 -3038 292 -2970
rect 306 -3038 308 -2970
rect 314 -3003 316 -2970
rect 324 -3003 326 -2970
rect 314 -3005 326 -3003
rect 314 -3038 316 -3005
rect 324 -3038 326 -3005
rect 332 -3038 334 -2970
rect 348 -3038 350 -2970
rect 356 -3038 358 -2970
rect 366 -3038 368 -2970
rect 374 -3038 376 -2970
rect 390 -3038 392 -2970
rect 398 -3038 400 -2970
rect 477 -3038 479 -2970
rect 846 -3034 848 -2978
rect 1204 -3038 1206 -2970
rect -1259 -3044 -1257 -3042
rect -1249 -3044 -1247 -3042
rect -1233 -3044 -1231 -3042
rect -1225 -3044 -1223 -3042
rect -1209 -3044 -1207 -3042
rect -1201 -3044 -1199 -3042
rect -1191 -3044 -1189 -3042
rect -1183 -3044 -1181 -3042
rect -1167 -3044 -1165 -3042
rect -1159 -3044 -1157 -3042
rect -1149 -3044 -1147 -3042
rect -1141 -3044 -1139 -3042
rect -1125 -3044 -1123 -3042
rect -1117 -3044 -1115 -3042
rect -1107 -3044 -1105 -3042
rect -1099 -3044 -1097 -3042
rect -1083 -3044 -1081 -3042
rect -1075 -3044 -1073 -3042
rect -1021 -3044 -1019 -3042
rect -930 -3044 -928 -3042
rect -920 -3044 -918 -3042
rect -904 -3044 -902 -3042
rect -896 -3044 -894 -3042
rect -880 -3044 -878 -3042
rect -872 -3044 -870 -3042
rect -862 -3044 -860 -3042
rect -854 -3044 -852 -3042
rect -838 -3044 -836 -3042
rect -830 -3044 -828 -3042
rect -820 -3044 -818 -3042
rect -812 -3044 -810 -3042
rect -796 -3044 -794 -3042
rect -788 -3044 -786 -3042
rect -778 -3044 -776 -3042
rect -770 -3044 -768 -3042
rect -754 -3044 -752 -3042
rect -746 -3044 -744 -3042
rect -667 -3044 -665 -3042
rect -572 -3044 -570 -3042
rect -562 -3044 -560 -3042
rect -546 -3044 -544 -3042
rect -538 -3044 -536 -3042
rect -522 -3044 -520 -3042
rect -514 -3044 -512 -3042
rect -504 -3044 -502 -3042
rect -496 -3044 -494 -3042
rect -480 -3044 -478 -3042
rect -472 -3044 -470 -3042
rect -462 -3044 -460 -3042
rect -454 -3044 -452 -3042
rect -438 -3044 -436 -3042
rect -430 -3044 -428 -3042
rect -420 -3044 -418 -3042
rect -412 -3044 -410 -3042
rect -396 -3044 -394 -3042
rect -388 -3044 -386 -3042
rect -324 -3044 -322 -3042
rect -214 -3044 -212 -3042
rect -204 -3044 -202 -3042
rect -188 -3044 -186 -3042
rect -180 -3044 -178 -3042
rect -164 -3044 -162 -3042
rect -156 -3044 -154 -3042
rect -146 -3044 -144 -3042
rect -138 -3044 -136 -3042
rect -122 -3044 -120 -3042
rect -114 -3044 -112 -3042
rect -104 -3044 -102 -3042
rect -96 -3044 -94 -3042
rect -80 -3044 -78 -3042
rect -72 -3044 -70 -3042
rect -62 -3044 -60 -3042
rect -54 -3044 -52 -3042
rect -38 -3044 -36 -3042
rect -30 -3044 -28 -3042
rect 214 -3044 216 -3042
rect 224 -3044 226 -3042
rect 240 -3044 242 -3042
rect 248 -3044 250 -3042
rect 264 -3044 266 -3042
rect 272 -3044 274 -3042
rect 282 -3044 284 -3042
rect 290 -3044 292 -3042
rect 306 -3044 308 -3042
rect 314 -3044 316 -3042
rect 324 -3044 326 -3042
rect 332 -3044 334 -3042
rect 348 -3044 350 -3042
rect 356 -3044 358 -3042
rect 366 -3044 368 -3042
rect 374 -3044 376 -3042
rect 390 -3044 392 -3042
rect 398 -3044 400 -3042
rect 477 -3044 479 -3042
rect 846 -3044 848 -3042
rect 1204 -3044 1206 -3042
rect -1259 -3078 -1257 -3076
rect -1249 -3078 -1247 -3076
rect -1233 -3078 -1231 -3076
rect -1225 -3078 -1223 -3076
rect -1209 -3078 -1207 -3076
rect -1201 -3078 -1199 -3076
rect -1191 -3078 -1189 -3076
rect -1183 -3078 -1181 -3076
rect -1167 -3078 -1165 -3076
rect -1159 -3078 -1157 -3076
rect -1149 -3078 -1147 -3076
rect -1141 -3078 -1139 -3076
rect -1125 -3078 -1123 -3076
rect -1117 -3078 -1115 -3076
rect -1107 -3078 -1105 -3076
rect -1099 -3078 -1097 -3076
rect -1083 -3078 -1081 -3076
rect -1075 -3078 -1073 -3076
rect -1021 -3078 -1019 -3076
rect -930 -3078 -928 -3076
rect -920 -3078 -918 -3076
rect -904 -3078 -902 -3076
rect -896 -3078 -894 -3076
rect -880 -3078 -878 -3076
rect -872 -3078 -870 -3076
rect -862 -3078 -860 -3076
rect -854 -3078 -852 -3076
rect -838 -3078 -836 -3076
rect -830 -3078 -828 -3076
rect -820 -3078 -818 -3076
rect -812 -3078 -810 -3076
rect -796 -3078 -794 -3076
rect -788 -3078 -786 -3076
rect -778 -3078 -776 -3076
rect -770 -3078 -768 -3076
rect -754 -3078 -752 -3076
rect -746 -3078 -744 -3076
rect -572 -3078 -570 -3076
rect -562 -3078 -560 -3076
rect -546 -3078 -544 -3076
rect -538 -3078 -536 -3076
rect -522 -3078 -520 -3076
rect -514 -3078 -512 -3076
rect -504 -3078 -502 -3076
rect -496 -3078 -494 -3076
rect -480 -3078 -478 -3076
rect -472 -3078 -470 -3076
rect -462 -3078 -460 -3076
rect -454 -3078 -452 -3076
rect -438 -3078 -436 -3076
rect -430 -3078 -428 -3076
rect -420 -3078 -418 -3076
rect -412 -3078 -410 -3076
rect -396 -3078 -394 -3076
rect -388 -3078 -386 -3076
rect -324 -3078 -322 -3076
rect -214 -3078 -212 -3076
rect -204 -3078 -202 -3076
rect -188 -3078 -186 -3076
rect -180 -3078 -178 -3076
rect -164 -3078 -162 -3076
rect -156 -3078 -154 -3076
rect -146 -3078 -144 -3076
rect -138 -3078 -136 -3076
rect -122 -3078 -120 -3076
rect -114 -3078 -112 -3076
rect -104 -3078 -102 -3076
rect -96 -3078 -94 -3076
rect -80 -3078 -78 -3076
rect -72 -3078 -70 -3076
rect -62 -3078 -60 -3076
rect -54 -3078 -52 -3076
rect -38 -3078 -36 -3076
rect -30 -3078 -28 -3076
rect 214 -3078 216 -3076
rect 224 -3078 226 -3076
rect 240 -3078 242 -3076
rect 248 -3078 250 -3076
rect 264 -3078 266 -3076
rect 272 -3078 274 -3076
rect 282 -3078 284 -3076
rect 290 -3078 292 -3076
rect 306 -3078 308 -3076
rect 314 -3078 316 -3076
rect 324 -3078 326 -3076
rect 332 -3078 334 -3076
rect 348 -3078 350 -3076
rect 356 -3078 358 -3076
rect 366 -3078 368 -3076
rect 374 -3078 376 -3076
rect 390 -3078 392 -3076
rect 398 -3078 400 -3076
rect 477 -3078 479 -3076
rect 570 -3078 572 -3076
rect 580 -3078 582 -3076
rect 596 -3078 598 -3076
rect 604 -3078 606 -3076
rect 620 -3078 622 -3076
rect 628 -3078 630 -3076
rect 638 -3078 640 -3076
rect 646 -3078 648 -3076
rect 662 -3078 664 -3076
rect 670 -3078 672 -3076
rect 680 -3078 682 -3076
rect 688 -3078 690 -3076
rect 704 -3078 706 -3076
rect 712 -3078 714 -3076
rect 722 -3078 724 -3076
rect 730 -3078 732 -3076
rect 746 -3078 748 -3076
rect 754 -3078 756 -3076
rect 968 -3078 970 -3076
rect 978 -3078 980 -3076
rect 994 -3078 996 -3076
rect 1002 -3078 1004 -3076
rect 1018 -3078 1020 -3076
rect 1026 -3078 1028 -3076
rect 1036 -3078 1038 -3076
rect 1044 -3078 1046 -3076
rect 1060 -3078 1062 -3076
rect 1068 -3078 1070 -3076
rect 1078 -3078 1080 -3076
rect 1086 -3078 1088 -3076
rect 1102 -3078 1104 -3076
rect 1110 -3078 1112 -3076
rect 1120 -3078 1122 -3076
rect 1128 -3078 1130 -3076
rect 1144 -3078 1146 -3076
rect 1152 -3078 1154 -3076
rect 1204 -3078 1206 -3076
rect 1326 -3078 1328 -3076
rect 1336 -3078 1338 -3076
rect 1352 -3078 1354 -3076
rect 1360 -3078 1362 -3076
rect 1376 -3078 1378 -3076
rect 1384 -3078 1386 -3076
rect 1394 -3078 1396 -3076
rect 1402 -3078 1404 -3076
rect 1418 -3078 1420 -3076
rect 1426 -3078 1428 -3076
rect 1436 -3078 1438 -3076
rect 1444 -3078 1446 -3076
rect 1460 -3078 1462 -3076
rect 1468 -3078 1470 -3076
rect 1478 -3078 1480 -3076
rect 1486 -3078 1488 -3076
rect 1502 -3078 1504 -3076
rect 1510 -3078 1512 -3076
rect -1259 -3154 -1257 -3086
rect -1249 -3154 -1247 -3086
rect -1233 -3154 -1231 -3086
rect -1225 -3154 -1223 -3086
rect -1209 -3154 -1207 -3086
rect -1201 -3154 -1199 -3086
rect -1191 -3154 -1189 -3086
rect -1183 -3154 -1181 -3086
rect -1167 -3154 -1165 -3086
rect -1159 -3119 -1157 -3086
rect -1149 -3119 -1147 -3086
rect -1159 -3121 -1147 -3119
rect -1159 -3154 -1157 -3121
rect -1149 -3154 -1147 -3121
rect -1141 -3154 -1139 -3086
rect -1125 -3154 -1123 -3086
rect -1117 -3154 -1115 -3086
rect -1107 -3154 -1105 -3086
rect -1099 -3154 -1097 -3086
rect -1083 -3154 -1081 -3086
rect -1075 -3154 -1073 -3086
rect -1021 -3154 -1019 -3086
rect -930 -3154 -928 -3086
rect -920 -3154 -918 -3086
rect -904 -3154 -902 -3086
rect -896 -3154 -894 -3086
rect -880 -3154 -878 -3086
rect -872 -3154 -870 -3086
rect -862 -3154 -860 -3086
rect -854 -3154 -852 -3086
rect -838 -3154 -836 -3086
rect -830 -3119 -828 -3086
rect -820 -3119 -818 -3086
rect -830 -3121 -818 -3119
rect -830 -3154 -828 -3121
rect -820 -3154 -818 -3121
rect -812 -3154 -810 -3086
rect -796 -3154 -794 -3086
rect -788 -3154 -786 -3086
rect -778 -3154 -776 -3086
rect -770 -3154 -768 -3086
rect -754 -3154 -752 -3086
rect -746 -3154 -744 -3086
rect -572 -3154 -570 -3086
rect -562 -3154 -560 -3086
rect -546 -3154 -544 -3086
rect -538 -3154 -536 -3086
rect -522 -3154 -520 -3086
rect -514 -3154 -512 -3086
rect -504 -3154 -502 -3086
rect -496 -3154 -494 -3086
rect -480 -3154 -478 -3086
rect -472 -3119 -470 -3086
rect -462 -3119 -460 -3086
rect -472 -3121 -460 -3119
rect -472 -3154 -470 -3121
rect -462 -3154 -460 -3121
rect -454 -3154 -452 -3086
rect -438 -3154 -436 -3086
rect -430 -3154 -428 -3086
rect -420 -3154 -418 -3086
rect -412 -3154 -410 -3086
rect -396 -3154 -394 -3086
rect -388 -3154 -386 -3086
rect -324 -3154 -322 -3086
rect -214 -3154 -212 -3086
rect -204 -3154 -202 -3086
rect -188 -3154 -186 -3086
rect -180 -3154 -178 -3086
rect -164 -3154 -162 -3086
rect -156 -3154 -154 -3086
rect -146 -3154 -144 -3086
rect -138 -3154 -136 -3086
rect -122 -3154 -120 -3086
rect -114 -3119 -112 -3086
rect -104 -3119 -102 -3086
rect -114 -3121 -102 -3119
rect -114 -3154 -112 -3121
rect -104 -3154 -102 -3121
rect -96 -3154 -94 -3086
rect -80 -3154 -78 -3086
rect -72 -3154 -70 -3086
rect -62 -3154 -60 -3086
rect -54 -3154 -52 -3086
rect -38 -3154 -36 -3086
rect -30 -3154 -28 -3086
rect 214 -3154 216 -3086
rect 224 -3154 226 -3086
rect 240 -3154 242 -3086
rect 248 -3154 250 -3086
rect 264 -3154 266 -3086
rect 272 -3154 274 -3086
rect 282 -3154 284 -3086
rect 290 -3154 292 -3086
rect 306 -3154 308 -3086
rect 314 -3119 316 -3086
rect 324 -3119 326 -3086
rect 314 -3121 326 -3119
rect 314 -3154 316 -3121
rect 324 -3154 326 -3121
rect 332 -3154 334 -3086
rect 348 -3154 350 -3086
rect 356 -3154 358 -3086
rect 366 -3154 368 -3086
rect 374 -3154 376 -3086
rect 390 -3154 392 -3086
rect 398 -3154 400 -3086
rect 477 -3154 479 -3086
rect 570 -3154 572 -3086
rect 580 -3154 582 -3086
rect 596 -3154 598 -3086
rect 604 -3154 606 -3086
rect 620 -3154 622 -3086
rect 628 -3154 630 -3086
rect 638 -3154 640 -3086
rect 646 -3154 648 -3086
rect 662 -3154 664 -3086
rect 670 -3119 672 -3086
rect 680 -3119 682 -3086
rect 670 -3121 682 -3119
rect 670 -3154 672 -3121
rect 680 -3154 682 -3121
rect 688 -3154 690 -3086
rect 704 -3154 706 -3086
rect 712 -3154 714 -3086
rect 722 -3154 724 -3086
rect 730 -3154 732 -3086
rect 746 -3154 748 -3086
rect 754 -3154 756 -3086
rect 968 -3154 970 -3086
rect 978 -3154 980 -3086
rect 994 -3154 996 -3086
rect 1002 -3154 1004 -3086
rect 1018 -3154 1020 -3086
rect 1026 -3154 1028 -3086
rect 1036 -3154 1038 -3086
rect 1044 -3154 1046 -3086
rect 1060 -3154 1062 -3086
rect 1068 -3119 1070 -3086
rect 1078 -3119 1080 -3086
rect 1068 -3121 1080 -3119
rect 1068 -3154 1070 -3121
rect 1078 -3154 1080 -3121
rect 1086 -3154 1088 -3086
rect 1102 -3154 1104 -3086
rect 1110 -3154 1112 -3086
rect 1120 -3154 1122 -3086
rect 1128 -3154 1130 -3086
rect 1144 -3154 1146 -3086
rect 1152 -3154 1154 -3086
rect 1204 -3154 1206 -3086
rect 1326 -3154 1328 -3086
rect 1336 -3154 1338 -3086
rect 1352 -3154 1354 -3086
rect 1360 -3154 1362 -3086
rect 1376 -3154 1378 -3086
rect 1384 -3154 1386 -3086
rect 1394 -3154 1396 -3086
rect 1402 -3154 1404 -3086
rect 1418 -3154 1420 -3086
rect 1426 -3119 1428 -3086
rect 1436 -3119 1438 -3086
rect 1426 -3121 1438 -3119
rect 1426 -3154 1428 -3121
rect 1436 -3154 1438 -3121
rect 1444 -3154 1446 -3086
rect 1460 -3154 1462 -3086
rect 1468 -3154 1470 -3086
rect 1478 -3154 1480 -3086
rect 1486 -3154 1488 -3086
rect 1502 -3154 1504 -3086
rect 1510 -3154 1512 -3086
rect -1259 -3160 -1257 -3158
rect -1249 -3160 -1247 -3158
rect -1233 -3160 -1231 -3158
rect -1225 -3160 -1223 -3158
rect -1209 -3160 -1207 -3158
rect -1201 -3160 -1199 -3158
rect -1191 -3160 -1189 -3158
rect -1183 -3160 -1181 -3158
rect -1167 -3160 -1165 -3158
rect -1159 -3160 -1157 -3158
rect -1149 -3160 -1147 -3158
rect -1141 -3160 -1139 -3158
rect -1125 -3160 -1123 -3158
rect -1117 -3160 -1115 -3158
rect -1107 -3160 -1105 -3158
rect -1099 -3160 -1097 -3158
rect -1083 -3160 -1081 -3158
rect -1075 -3160 -1073 -3158
rect -1021 -3160 -1019 -3158
rect -930 -3160 -928 -3158
rect -920 -3160 -918 -3158
rect -904 -3160 -902 -3158
rect -896 -3160 -894 -3158
rect -880 -3160 -878 -3158
rect -872 -3160 -870 -3158
rect -862 -3160 -860 -3158
rect -854 -3160 -852 -3158
rect -838 -3160 -836 -3158
rect -830 -3160 -828 -3158
rect -820 -3160 -818 -3158
rect -812 -3160 -810 -3158
rect -796 -3160 -794 -3158
rect -788 -3160 -786 -3158
rect -778 -3160 -776 -3158
rect -770 -3160 -768 -3158
rect -754 -3160 -752 -3158
rect -746 -3160 -744 -3158
rect -572 -3160 -570 -3158
rect -562 -3160 -560 -3158
rect -546 -3160 -544 -3158
rect -538 -3160 -536 -3158
rect -522 -3160 -520 -3158
rect -514 -3160 -512 -3158
rect -504 -3160 -502 -3158
rect -496 -3160 -494 -3158
rect -480 -3160 -478 -3158
rect -472 -3160 -470 -3158
rect -462 -3160 -460 -3158
rect -454 -3160 -452 -3158
rect -438 -3160 -436 -3158
rect -430 -3160 -428 -3158
rect -420 -3160 -418 -3158
rect -412 -3160 -410 -3158
rect -396 -3160 -394 -3158
rect -388 -3160 -386 -3158
rect -324 -3160 -322 -3158
rect -214 -3160 -212 -3158
rect -204 -3160 -202 -3158
rect -188 -3160 -186 -3158
rect -180 -3160 -178 -3158
rect -164 -3160 -162 -3158
rect -156 -3160 -154 -3158
rect -146 -3160 -144 -3158
rect -138 -3160 -136 -3158
rect -122 -3160 -120 -3158
rect -114 -3160 -112 -3158
rect -104 -3160 -102 -3158
rect -96 -3160 -94 -3158
rect -80 -3160 -78 -3158
rect -72 -3160 -70 -3158
rect -62 -3160 -60 -3158
rect -54 -3160 -52 -3158
rect -38 -3160 -36 -3158
rect -30 -3160 -28 -3158
rect 214 -3160 216 -3158
rect 224 -3160 226 -3158
rect 240 -3160 242 -3158
rect 248 -3160 250 -3158
rect 264 -3160 266 -3158
rect 272 -3160 274 -3158
rect 282 -3160 284 -3158
rect 290 -3160 292 -3158
rect 306 -3160 308 -3158
rect 314 -3160 316 -3158
rect 324 -3160 326 -3158
rect 332 -3160 334 -3158
rect 348 -3160 350 -3158
rect 356 -3160 358 -3158
rect 366 -3160 368 -3158
rect 374 -3160 376 -3158
rect 390 -3160 392 -3158
rect 398 -3160 400 -3158
rect 477 -3160 479 -3158
rect 570 -3160 572 -3158
rect 580 -3160 582 -3158
rect 596 -3160 598 -3158
rect 604 -3160 606 -3158
rect 620 -3160 622 -3158
rect 628 -3160 630 -3158
rect 638 -3160 640 -3158
rect 646 -3160 648 -3158
rect 662 -3160 664 -3158
rect 670 -3160 672 -3158
rect 680 -3160 682 -3158
rect 688 -3160 690 -3158
rect 704 -3160 706 -3158
rect 712 -3160 714 -3158
rect 722 -3160 724 -3158
rect 730 -3160 732 -3158
rect 746 -3160 748 -3158
rect 754 -3160 756 -3158
rect 968 -3160 970 -3158
rect 978 -3160 980 -3158
rect 994 -3160 996 -3158
rect 1002 -3160 1004 -3158
rect 1018 -3160 1020 -3158
rect 1026 -3160 1028 -3158
rect 1036 -3160 1038 -3158
rect 1044 -3160 1046 -3158
rect 1060 -3160 1062 -3158
rect 1068 -3160 1070 -3158
rect 1078 -3160 1080 -3158
rect 1086 -3160 1088 -3158
rect 1102 -3160 1104 -3158
rect 1110 -3160 1112 -3158
rect 1120 -3160 1122 -3158
rect 1128 -3160 1130 -3158
rect 1144 -3160 1146 -3158
rect 1152 -3160 1154 -3158
rect 1204 -3160 1206 -3158
rect 1326 -3160 1328 -3158
rect 1336 -3160 1338 -3158
rect 1352 -3160 1354 -3158
rect 1360 -3160 1362 -3158
rect 1376 -3160 1378 -3158
rect 1384 -3160 1386 -3158
rect 1394 -3160 1396 -3158
rect 1402 -3160 1404 -3158
rect 1418 -3160 1420 -3158
rect 1426 -3160 1428 -3158
rect 1436 -3160 1438 -3158
rect 1444 -3160 1446 -3158
rect 1460 -3160 1462 -3158
rect 1468 -3160 1470 -3158
rect 1478 -3160 1480 -3158
rect 1486 -3160 1488 -3158
rect 1502 -3160 1504 -3158
rect 1510 -3160 1512 -3158
rect -1259 -3199 -1257 -3197
rect -1249 -3199 -1247 -3197
rect -1233 -3199 -1231 -3197
rect -1225 -3199 -1223 -3197
rect -1209 -3199 -1207 -3197
rect -1201 -3199 -1199 -3197
rect -1191 -3199 -1189 -3197
rect -1183 -3199 -1181 -3197
rect -1167 -3199 -1165 -3197
rect -1159 -3199 -1157 -3197
rect -1149 -3199 -1147 -3197
rect -1141 -3199 -1139 -3197
rect -1125 -3199 -1123 -3197
rect -1117 -3199 -1115 -3197
rect -1107 -3199 -1105 -3197
rect -1099 -3199 -1097 -3197
rect -1083 -3199 -1081 -3197
rect -1075 -3199 -1073 -3197
rect -930 -3199 -928 -3197
rect -920 -3199 -918 -3197
rect -904 -3199 -902 -3197
rect -896 -3199 -894 -3197
rect -880 -3199 -878 -3197
rect -872 -3199 -870 -3197
rect -862 -3199 -860 -3197
rect -854 -3199 -852 -3197
rect -838 -3199 -836 -3197
rect -830 -3199 -828 -3197
rect -820 -3199 -818 -3197
rect -812 -3199 -810 -3197
rect -796 -3199 -794 -3197
rect -788 -3199 -786 -3197
rect -778 -3199 -776 -3197
rect -770 -3199 -768 -3197
rect -754 -3199 -752 -3197
rect -746 -3199 -744 -3197
rect -572 -3199 -570 -3197
rect -562 -3199 -560 -3197
rect -546 -3199 -544 -3197
rect -538 -3199 -536 -3197
rect -522 -3199 -520 -3197
rect -514 -3199 -512 -3197
rect -504 -3199 -502 -3197
rect -496 -3199 -494 -3197
rect -480 -3199 -478 -3197
rect -472 -3199 -470 -3197
rect -462 -3199 -460 -3197
rect -454 -3199 -452 -3197
rect -438 -3199 -436 -3197
rect -430 -3199 -428 -3197
rect -420 -3199 -418 -3197
rect -412 -3199 -410 -3197
rect -396 -3199 -394 -3197
rect -388 -3199 -386 -3197
rect -214 -3199 -212 -3197
rect -204 -3199 -202 -3197
rect -188 -3199 -186 -3197
rect -180 -3199 -178 -3197
rect -164 -3199 -162 -3197
rect -156 -3199 -154 -3197
rect -146 -3199 -144 -3197
rect -138 -3199 -136 -3197
rect -122 -3199 -120 -3197
rect -114 -3199 -112 -3197
rect -104 -3199 -102 -3197
rect -96 -3199 -94 -3197
rect -80 -3199 -78 -3197
rect -72 -3199 -70 -3197
rect -62 -3199 -60 -3197
rect -54 -3199 -52 -3197
rect -38 -3199 -36 -3197
rect -30 -3199 -28 -3197
rect 214 -3199 216 -3197
rect 224 -3199 226 -3197
rect 240 -3199 242 -3197
rect 248 -3199 250 -3197
rect 264 -3199 266 -3197
rect 272 -3199 274 -3197
rect 282 -3199 284 -3197
rect 290 -3199 292 -3197
rect 306 -3199 308 -3197
rect 314 -3199 316 -3197
rect 324 -3199 326 -3197
rect 332 -3199 334 -3197
rect 348 -3199 350 -3197
rect 356 -3199 358 -3197
rect 366 -3199 368 -3197
rect 374 -3199 376 -3197
rect 390 -3199 392 -3197
rect 398 -3199 400 -3197
rect 570 -3199 572 -3197
rect 580 -3199 582 -3197
rect 596 -3199 598 -3197
rect 604 -3199 606 -3197
rect 620 -3199 622 -3197
rect 628 -3199 630 -3197
rect 638 -3199 640 -3197
rect 646 -3199 648 -3197
rect 662 -3199 664 -3197
rect 670 -3199 672 -3197
rect 680 -3199 682 -3197
rect 688 -3199 690 -3197
rect 704 -3199 706 -3197
rect 712 -3199 714 -3197
rect 722 -3199 724 -3197
rect 730 -3199 732 -3197
rect 746 -3199 748 -3197
rect 754 -3199 756 -3197
rect 968 -3199 970 -3197
rect 978 -3199 980 -3197
rect 994 -3199 996 -3197
rect 1002 -3199 1004 -3197
rect 1018 -3199 1020 -3197
rect 1026 -3199 1028 -3197
rect 1036 -3199 1038 -3197
rect 1044 -3199 1046 -3197
rect 1060 -3199 1062 -3197
rect 1068 -3199 1070 -3197
rect 1078 -3199 1080 -3197
rect 1086 -3199 1088 -3197
rect 1102 -3199 1104 -3197
rect 1110 -3199 1112 -3197
rect 1120 -3199 1122 -3197
rect 1128 -3199 1130 -3197
rect 1144 -3199 1146 -3197
rect 1152 -3199 1154 -3197
rect 1326 -3199 1328 -3197
rect 1336 -3199 1338 -3197
rect 1352 -3199 1354 -3197
rect 1360 -3199 1362 -3197
rect 1376 -3199 1378 -3197
rect 1384 -3199 1386 -3197
rect 1394 -3199 1396 -3197
rect 1402 -3199 1404 -3197
rect 1418 -3199 1420 -3197
rect 1426 -3199 1428 -3197
rect 1436 -3199 1438 -3197
rect 1444 -3199 1446 -3197
rect 1460 -3199 1462 -3197
rect 1468 -3199 1470 -3197
rect 1478 -3199 1480 -3197
rect 1486 -3199 1488 -3197
rect 1502 -3199 1504 -3197
rect 1510 -3199 1512 -3197
rect -1259 -3275 -1257 -3207
rect -1249 -3275 -1247 -3207
rect -1233 -3275 -1231 -3207
rect -1225 -3275 -1223 -3207
rect -1209 -3275 -1207 -3207
rect -1201 -3275 -1199 -3207
rect -1191 -3275 -1189 -3207
rect -1183 -3275 -1181 -3207
rect -1167 -3275 -1165 -3207
rect -1159 -3240 -1157 -3207
rect -1149 -3240 -1147 -3207
rect -1159 -3242 -1147 -3240
rect -1159 -3275 -1157 -3242
rect -1149 -3275 -1147 -3242
rect -1141 -3275 -1139 -3207
rect -1125 -3275 -1123 -3207
rect -1117 -3275 -1115 -3207
rect -1107 -3275 -1105 -3207
rect -1099 -3275 -1097 -3207
rect -1083 -3275 -1081 -3207
rect -1075 -3275 -1073 -3207
rect -930 -3275 -928 -3207
rect -920 -3275 -918 -3207
rect -904 -3275 -902 -3207
rect -896 -3275 -894 -3207
rect -880 -3275 -878 -3207
rect -872 -3275 -870 -3207
rect -862 -3275 -860 -3207
rect -854 -3275 -852 -3207
rect -838 -3275 -836 -3207
rect -830 -3240 -828 -3207
rect -820 -3240 -818 -3207
rect -830 -3242 -818 -3240
rect -830 -3275 -828 -3242
rect -820 -3275 -818 -3242
rect -812 -3275 -810 -3207
rect -796 -3275 -794 -3207
rect -788 -3275 -786 -3207
rect -778 -3275 -776 -3207
rect -770 -3275 -768 -3207
rect -754 -3275 -752 -3207
rect -746 -3275 -744 -3207
rect -572 -3275 -570 -3207
rect -562 -3275 -560 -3207
rect -546 -3275 -544 -3207
rect -538 -3275 -536 -3207
rect -522 -3275 -520 -3207
rect -514 -3275 -512 -3207
rect -504 -3275 -502 -3207
rect -496 -3275 -494 -3207
rect -480 -3275 -478 -3207
rect -472 -3240 -470 -3207
rect -462 -3240 -460 -3207
rect -472 -3242 -460 -3240
rect -472 -3275 -470 -3242
rect -462 -3275 -460 -3242
rect -454 -3275 -452 -3207
rect -438 -3275 -436 -3207
rect -430 -3275 -428 -3207
rect -420 -3275 -418 -3207
rect -412 -3275 -410 -3207
rect -396 -3275 -394 -3207
rect -388 -3275 -386 -3207
rect -214 -3275 -212 -3207
rect -204 -3275 -202 -3207
rect -188 -3275 -186 -3207
rect -180 -3275 -178 -3207
rect -164 -3275 -162 -3207
rect -156 -3275 -154 -3207
rect -146 -3275 -144 -3207
rect -138 -3275 -136 -3207
rect -122 -3275 -120 -3207
rect -114 -3240 -112 -3207
rect -104 -3240 -102 -3207
rect -114 -3242 -102 -3240
rect -114 -3275 -112 -3242
rect -104 -3275 -102 -3242
rect -96 -3275 -94 -3207
rect -80 -3275 -78 -3207
rect -72 -3275 -70 -3207
rect -62 -3275 -60 -3207
rect -54 -3275 -52 -3207
rect -38 -3275 -36 -3207
rect -30 -3275 -28 -3207
rect 214 -3275 216 -3207
rect 224 -3275 226 -3207
rect 240 -3275 242 -3207
rect 248 -3275 250 -3207
rect 264 -3275 266 -3207
rect 272 -3275 274 -3207
rect 282 -3275 284 -3207
rect 290 -3275 292 -3207
rect 306 -3275 308 -3207
rect 314 -3240 316 -3207
rect 324 -3240 326 -3207
rect 314 -3242 326 -3240
rect 314 -3275 316 -3242
rect 324 -3275 326 -3242
rect 332 -3275 334 -3207
rect 348 -3275 350 -3207
rect 356 -3275 358 -3207
rect 366 -3275 368 -3207
rect 374 -3275 376 -3207
rect 390 -3275 392 -3207
rect 398 -3275 400 -3207
rect 570 -3275 572 -3207
rect 580 -3275 582 -3207
rect 596 -3275 598 -3207
rect 604 -3275 606 -3207
rect 620 -3275 622 -3207
rect 628 -3275 630 -3207
rect 638 -3275 640 -3207
rect 646 -3275 648 -3207
rect 662 -3275 664 -3207
rect 670 -3240 672 -3207
rect 680 -3240 682 -3207
rect 670 -3242 682 -3240
rect 670 -3275 672 -3242
rect 680 -3275 682 -3242
rect 688 -3275 690 -3207
rect 704 -3275 706 -3207
rect 712 -3275 714 -3207
rect 722 -3275 724 -3207
rect 730 -3275 732 -3207
rect 746 -3275 748 -3207
rect 754 -3275 756 -3207
rect 968 -3275 970 -3207
rect 978 -3275 980 -3207
rect 994 -3275 996 -3207
rect 1002 -3275 1004 -3207
rect 1018 -3275 1020 -3207
rect 1026 -3275 1028 -3207
rect 1036 -3275 1038 -3207
rect 1044 -3275 1046 -3207
rect 1060 -3275 1062 -3207
rect 1068 -3240 1070 -3207
rect 1078 -3240 1080 -3207
rect 1068 -3242 1080 -3240
rect 1068 -3275 1070 -3242
rect 1078 -3275 1080 -3242
rect 1086 -3275 1088 -3207
rect 1102 -3275 1104 -3207
rect 1110 -3275 1112 -3207
rect 1120 -3275 1122 -3207
rect 1128 -3275 1130 -3207
rect 1144 -3275 1146 -3207
rect 1152 -3275 1154 -3207
rect 1326 -3275 1328 -3207
rect 1336 -3275 1338 -3207
rect 1352 -3275 1354 -3207
rect 1360 -3275 1362 -3207
rect 1376 -3275 1378 -3207
rect 1384 -3275 1386 -3207
rect 1394 -3275 1396 -3207
rect 1402 -3275 1404 -3207
rect 1418 -3275 1420 -3207
rect 1426 -3240 1428 -3207
rect 1436 -3240 1438 -3207
rect 1426 -3242 1438 -3240
rect 1426 -3275 1428 -3242
rect 1436 -3275 1438 -3242
rect 1444 -3275 1446 -3207
rect 1460 -3275 1462 -3207
rect 1468 -3275 1470 -3207
rect 1478 -3275 1480 -3207
rect 1486 -3275 1488 -3207
rect 1502 -3275 1504 -3207
rect 1510 -3275 1512 -3207
rect -1259 -3281 -1257 -3279
rect -1249 -3281 -1247 -3279
rect -1233 -3281 -1231 -3279
rect -1225 -3281 -1223 -3279
rect -1209 -3281 -1207 -3279
rect -1201 -3281 -1199 -3279
rect -1191 -3281 -1189 -3279
rect -1183 -3281 -1181 -3279
rect -1167 -3281 -1165 -3279
rect -1159 -3281 -1157 -3279
rect -1149 -3281 -1147 -3279
rect -1141 -3281 -1139 -3279
rect -1125 -3281 -1123 -3279
rect -1117 -3281 -1115 -3279
rect -1107 -3281 -1105 -3279
rect -1099 -3281 -1097 -3279
rect -1083 -3281 -1081 -3279
rect -1075 -3281 -1073 -3279
rect -930 -3281 -928 -3279
rect -920 -3281 -918 -3279
rect -904 -3281 -902 -3279
rect -896 -3281 -894 -3279
rect -880 -3281 -878 -3279
rect -872 -3281 -870 -3279
rect -862 -3281 -860 -3279
rect -854 -3281 -852 -3279
rect -838 -3281 -836 -3279
rect -830 -3281 -828 -3279
rect -820 -3281 -818 -3279
rect -812 -3281 -810 -3279
rect -796 -3281 -794 -3279
rect -788 -3281 -786 -3279
rect -778 -3281 -776 -3279
rect -770 -3281 -768 -3279
rect -754 -3281 -752 -3279
rect -746 -3281 -744 -3279
rect -572 -3281 -570 -3279
rect -562 -3281 -560 -3279
rect -546 -3281 -544 -3279
rect -538 -3281 -536 -3279
rect -522 -3281 -520 -3279
rect -514 -3281 -512 -3279
rect -504 -3281 -502 -3279
rect -496 -3281 -494 -3279
rect -480 -3281 -478 -3279
rect -472 -3281 -470 -3279
rect -462 -3281 -460 -3279
rect -454 -3281 -452 -3279
rect -438 -3281 -436 -3279
rect -430 -3281 -428 -3279
rect -420 -3281 -418 -3279
rect -412 -3281 -410 -3279
rect -396 -3281 -394 -3279
rect -388 -3281 -386 -3279
rect -214 -3281 -212 -3279
rect -204 -3281 -202 -3279
rect -188 -3281 -186 -3279
rect -180 -3281 -178 -3279
rect -164 -3281 -162 -3279
rect -156 -3281 -154 -3279
rect -146 -3281 -144 -3279
rect -138 -3281 -136 -3279
rect -122 -3281 -120 -3279
rect -114 -3281 -112 -3279
rect -104 -3281 -102 -3279
rect -96 -3281 -94 -3279
rect -80 -3281 -78 -3279
rect -72 -3281 -70 -3279
rect -62 -3281 -60 -3279
rect -54 -3281 -52 -3279
rect -38 -3281 -36 -3279
rect -30 -3281 -28 -3279
rect 214 -3281 216 -3279
rect 224 -3281 226 -3279
rect 240 -3281 242 -3279
rect 248 -3281 250 -3279
rect 264 -3281 266 -3279
rect 272 -3281 274 -3279
rect 282 -3281 284 -3279
rect 290 -3281 292 -3279
rect 306 -3281 308 -3279
rect 314 -3281 316 -3279
rect 324 -3281 326 -3279
rect 332 -3281 334 -3279
rect 348 -3281 350 -3279
rect 356 -3281 358 -3279
rect 366 -3281 368 -3279
rect 374 -3281 376 -3279
rect 390 -3281 392 -3279
rect 398 -3281 400 -3279
rect 570 -3281 572 -3279
rect 580 -3281 582 -3279
rect 596 -3281 598 -3279
rect 604 -3281 606 -3279
rect 620 -3281 622 -3279
rect 628 -3281 630 -3279
rect 638 -3281 640 -3279
rect 646 -3281 648 -3279
rect 662 -3281 664 -3279
rect 670 -3281 672 -3279
rect 680 -3281 682 -3279
rect 688 -3281 690 -3279
rect 704 -3281 706 -3279
rect 712 -3281 714 -3279
rect 722 -3281 724 -3279
rect 730 -3281 732 -3279
rect 746 -3281 748 -3279
rect 754 -3281 756 -3279
rect 968 -3281 970 -3279
rect 978 -3281 980 -3279
rect 994 -3281 996 -3279
rect 1002 -3281 1004 -3279
rect 1018 -3281 1020 -3279
rect 1026 -3281 1028 -3279
rect 1036 -3281 1038 -3279
rect 1044 -3281 1046 -3279
rect 1060 -3281 1062 -3279
rect 1068 -3281 1070 -3279
rect 1078 -3281 1080 -3279
rect 1086 -3281 1088 -3279
rect 1102 -3281 1104 -3279
rect 1110 -3281 1112 -3279
rect 1120 -3281 1122 -3279
rect 1128 -3281 1130 -3279
rect 1144 -3281 1146 -3279
rect 1152 -3281 1154 -3279
rect 1326 -3281 1328 -3279
rect 1336 -3281 1338 -3279
rect 1352 -3281 1354 -3279
rect 1360 -3281 1362 -3279
rect 1376 -3281 1378 -3279
rect 1384 -3281 1386 -3279
rect 1394 -3281 1396 -3279
rect 1402 -3281 1404 -3279
rect 1418 -3281 1420 -3279
rect 1426 -3281 1428 -3279
rect 1436 -3281 1438 -3279
rect 1444 -3281 1446 -3279
rect 1460 -3281 1462 -3279
rect 1468 -3281 1470 -3279
rect 1478 -3281 1480 -3279
rect 1486 -3281 1488 -3279
rect 1502 -3281 1504 -3279
rect 1510 -3281 1512 -3279
rect -1259 -3313 -1257 -3311
rect -1249 -3313 -1247 -3311
rect -1233 -3313 -1231 -3311
rect -1225 -3313 -1223 -3311
rect -1209 -3313 -1207 -3311
rect -1201 -3313 -1199 -3311
rect -1191 -3313 -1189 -3311
rect -1183 -3313 -1181 -3311
rect -1167 -3313 -1165 -3311
rect -1159 -3313 -1157 -3311
rect -1149 -3313 -1147 -3311
rect -1141 -3313 -1139 -3311
rect -1125 -3313 -1123 -3311
rect -1117 -3313 -1115 -3311
rect -1107 -3313 -1105 -3311
rect -1099 -3313 -1097 -3311
rect -1083 -3313 -1081 -3311
rect -1075 -3313 -1073 -3311
rect -930 -3313 -928 -3311
rect -920 -3313 -918 -3311
rect -904 -3313 -902 -3311
rect -896 -3313 -894 -3311
rect -880 -3313 -878 -3311
rect -872 -3313 -870 -3311
rect -862 -3313 -860 -3311
rect -854 -3313 -852 -3311
rect -838 -3313 -836 -3311
rect -830 -3313 -828 -3311
rect -820 -3313 -818 -3311
rect -812 -3313 -810 -3311
rect -796 -3313 -794 -3311
rect -788 -3313 -786 -3311
rect -778 -3313 -776 -3311
rect -770 -3313 -768 -3311
rect -754 -3313 -752 -3311
rect -746 -3313 -744 -3311
rect -572 -3313 -570 -3311
rect -562 -3313 -560 -3311
rect -546 -3313 -544 -3311
rect -538 -3313 -536 -3311
rect -522 -3313 -520 -3311
rect -514 -3313 -512 -3311
rect -504 -3313 -502 -3311
rect -496 -3313 -494 -3311
rect -480 -3313 -478 -3311
rect -472 -3313 -470 -3311
rect -462 -3313 -460 -3311
rect -454 -3313 -452 -3311
rect -438 -3313 -436 -3311
rect -430 -3313 -428 -3311
rect -420 -3313 -418 -3311
rect -412 -3313 -410 -3311
rect -396 -3313 -394 -3311
rect -388 -3313 -386 -3311
rect -1259 -3389 -1257 -3321
rect -1249 -3389 -1247 -3321
rect -1233 -3389 -1231 -3321
rect -1225 -3389 -1223 -3321
rect -1209 -3389 -1207 -3321
rect -1201 -3389 -1199 -3321
rect -1191 -3389 -1189 -3321
rect -1183 -3389 -1181 -3321
rect -1167 -3389 -1165 -3321
rect -1159 -3354 -1157 -3321
rect -1149 -3354 -1147 -3321
rect -1159 -3356 -1147 -3354
rect -1159 -3389 -1157 -3356
rect -1149 -3389 -1147 -3356
rect -1141 -3389 -1139 -3321
rect -1125 -3389 -1123 -3321
rect -1117 -3389 -1115 -3321
rect -1107 -3389 -1105 -3321
rect -1099 -3389 -1097 -3321
rect -1083 -3389 -1081 -3321
rect -1075 -3389 -1073 -3321
rect -930 -3389 -928 -3321
rect -920 -3389 -918 -3321
rect -904 -3389 -902 -3321
rect -896 -3389 -894 -3321
rect -880 -3389 -878 -3321
rect -872 -3389 -870 -3321
rect -862 -3389 -860 -3321
rect -854 -3389 -852 -3321
rect -838 -3389 -836 -3321
rect -830 -3354 -828 -3321
rect -820 -3354 -818 -3321
rect -830 -3356 -818 -3354
rect -830 -3389 -828 -3356
rect -820 -3389 -818 -3356
rect -812 -3389 -810 -3321
rect -796 -3389 -794 -3321
rect -788 -3389 -786 -3321
rect -778 -3389 -776 -3321
rect -770 -3389 -768 -3321
rect -754 -3389 -752 -3321
rect -746 -3389 -744 -3321
rect -572 -3389 -570 -3321
rect -562 -3389 -560 -3321
rect -546 -3389 -544 -3321
rect -538 -3389 -536 -3321
rect -522 -3389 -520 -3321
rect -514 -3389 -512 -3321
rect -504 -3389 -502 -3321
rect -496 -3389 -494 -3321
rect -480 -3389 -478 -3321
rect -472 -3354 -470 -3321
rect -462 -3354 -460 -3321
rect -472 -3356 -460 -3354
rect -472 -3389 -470 -3356
rect -462 -3389 -460 -3356
rect -454 -3389 -452 -3321
rect -438 -3389 -436 -3321
rect -430 -3389 -428 -3321
rect -420 -3389 -418 -3321
rect -412 -3389 -410 -3321
rect -396 -3389 -394 -3321
rect -388 -3389 -386 -3321
rect -1259 -3395 -1257 -3393
rect -1249 -3395 -1247 -3393
rect -1233 -3395 -1231 -3393
rect -1225 -3395 -1223 -3393
rect -1209 -3395 -1207 -3393
rect -1201 -3395 -1199 -3393
rect -1191 -3395 -1189 -3393
rect -1183 -3395 -1181 -3393
rect -1167 -3395 -1165 -3393
rect -1159 -3395 -1157 -3393
rect -1149 -3395 -1147 -3393
rect -1141 -3395 -1139 -3393
rect -1125 -3395 -1123 -3393
rect -1117 -3395 -1115 -3393
rect -1107 -3395 -1105 -3393
rect -1099 -3395 -1097 -3393
rect -1083 -3395 -1081 -3393
rect -1075 -3395 -1073 -3393
rect -930 -3395 -928 -3393
rect -920 -3395 -918 -3393
rect -904 -3395 -902 -3393
rect -896 -3395 -894 -3393
rect -880 -3395 -878 -3393
rect -872 -3395 -870 -3393
rect -862 -3395 -860 -3393
rect -854 -3395 -852 -3393
rect -838 -3395 -836 -3393
rect -830 -3395 -828 -3393
rect -820 -3395 -818 -3393
rect -812 -3395 -810 -3393
rect -796 -3395 -794 -3393
rect -788 -3395 -786 -3393
rect -778 -3395 -776 -3393
rect -770 -3395 -768 -3393
rect -754 -3395 -752 -3393
rect -746 -3395 -744 -3393
rect -572 -3395 -570 -3393
rect -562 -3395 -560 -3393
rect -546 -3395 -544 -3393
rect -538 -3395 -536 -3393
rect -522 -3395 -520 -3393
rect -514 -3395 -512 -3393
rect -504 -3395 -502 -3393
rect -496 -3395 -494 -3393
rect -480 -3395 -478 -3393
rect -472 -3395 -470 -3393
rect -462 -3395 -460 -3393
rect -454 -3395 -452 -3393
rect -438 -3395 -436 -3393
rect -430 -3395 -428 -3393
rect -420 -3395 -418 -3393
rect -412 -3395 -410 -3393
rect -396 -3395 -394 -3393
rect -388 -3395 -386 -3393
rect -1334 -3430 -1332 -3428
rect -1326 -3430 -1324 -3428
rect -1316 -3430 -1314 -3428
rect -930 -3430 -928 -3428
rect -922 -3430 -920 -3428
rect -912 -3430 -910 -3428
rect -572 -3430 -570 -3428
rect -564 -3430 -562 -3428
rect -554 -3430 -552 -3428
rect -214 -3430 -212 -3428
rect -206 -3430 -204 -3428
rect -196 -3430 -194 -3428
rect 214 -3430 216 -3428
rect 222 -3430 224 -3428
rect 232 -3430 234 -3428
rect 570 -3430 572 -3428
rect 578 -3430 580 -3428
rect 588 -3430 590 -3428
rect 968 -3430 970 -3428
rect 976 -3430 978 -3428
rect 986 -3430 988 -3428
rect 1326 -3430 1328 -3428
rect 1334 -3430 1336 -3428
rect 1344 -3430 1346 -3428
rect -1334 -3506 -1332 -3438
rect -1326 -3462 -1324 -3438
rect -1326 -3506 -1324 -3466
rect -1316 -3506 -1314 -3438
rect -930 -3506 -928 -3438
rect -922 -3462 -920 -3438
rect -922 -3506 -920 -3466
rect -912 -3506 -910 -3438
rect -572 -3506 -570 -3438
rect -564 -3462 -562 -3438
rect -564 -3506 -562 -3466
rect -554 -3506 -552 -3438
rect -214 -3506 -212 -3438
rect -206 -3462 -204 -3438
rect -206 -3506 -204 -3466
rect -196 -3506 -194 -3438
rect 214 -3506 216 -3438
rect 222 -3462 224 -3438
rect 222 -3506 224 -3466
rect 232 -3506 234 -3438
rect 570 -3506 572 -3438
rect 578 -3462 580 -3438
rect 578 -3506 580 -3466
rect 588 -3506 590 -3438
rect 968 -3506 970 -3438
rect 976 -3462 978 -3438
rect 976 -3506 978 -3466
rect 986 -3506 988 -3438
rect 1326 -3506 1328 -3438
rect 1334 -3462 1336 -3438
rect 1334 -3506 1336 -3466
rect 1344 -3506 1346 -3438
rect -1334 -3512 -1332 -3510
rect -1326 -3512 -1324 -3510
rect -1316 -3512 -1314 -3510
rect -930 -3512 -928 -3510
rect -922 -3512 -920 -3510
rect -912 -3512 -910 -3510
rect -572 -3512 -570 -3510
rect -564 -3512 -562 -3510
rect -554 -3512 -552 -3510
rect -214 -3512 -212 -3510
rect -206 -3512 -204 -3510
rect -196 -3512 -194 -3510
rect 214 -3512 216 -3510
rect 222 -3512 224 -3510
rect 232 -3512 234 -3510
rect 570 -3512 572 -3510
rect 578 -3512 580 -3510
rect 588 -3512 590 -3510
rect 968 -3512 970 -3510
rect 976 -3512 978 -3510
rect 986 -3512 988 -3510
rect 1326 -3512 1328 -3510
rect 1334 -3512 1336 -3510
rect 1344 -3512 1346 -3510
rect -1259 -3554 -1257 -3552
rect -1249 -3554 -1247 -3552
rect -1233 -3554 -1231 -3552
rect -1223 -3554 -1221 -3552
rect -1215 -3554 -1213 -3552
rect -1205 -3554 -1203 -3552
rect -1189 -3554 -1187 -3552
rect -1181 -3554 -1179 -3552
rect -1171 -3554 -1169 -3552
rect -930 -3554 -928 -3552
rect -920 -3554 -918 -3552
rect -904 -3554 -902 -3552
rect -894 -3554 -892 -3552
rect -878 -3554 -876 -3552
rect -868 -3554 -866 -3552
rect -860 -3554 -858 -3552
rect -850 -3554 -848 -3552
rect -834 -3554 -832 -3552
rect -826 -3554 -824 -3552
rect -816 -3554 -814 -3552
rect -800 -3554 -798 -3552
rect -790 -3554 -788 -3552
rect -782 -3554 -780 -3552
rect -772 -3554 -770 -3552
rect -756 -3554 -754 -3552
rect -748 -3554 -746 -3552
rect -732 -3554 -730 -3552
rect -716 -3554 -714 -3552
rect -708 -3554 -706 -3552
rect -698 -3554 -696 -3552
rect -572 -3554 -570 -3552
rect -562 -3554 -560 -3552
rect -546 -3554 -544 -3552
rect -536 -3554 -534 -3552
rect -520 -3554 -518 -3552
rect -510 -3554 -508 -3552
rect -502 -3554 -500 -3552
rect -492 -3554 -490 -3552
rect -476 -3554 -474 -3552
rect -468 -3554 -466 -3552
rect -458 -3554 -456 -3552
rect -442 -3554 -440 -3552
rect -432 -3554 -430 -3552
rect -424 -3554 -422 -3552
rect -414 -3554 -412 -3552
rect -398 -3554 -396 -3552
rect -390 -3554 -388 -3552
rect -374 -3554 -372 -3552
rect -358 -3554 -356 -3552
rect -350 -3554 -348 -3552
rect -340 -3554 -338 -3552
rect -214 -3554 -212 -3552
rect -204 -3554 -202 -3552
rect -188 -3554 -186 -3552
rect -178 -3554 -176 -3552
rect -162 -3554 -160 -3552
rect -152 -3554 -150 -3552
rect -144 -3554 -142 -3552
rect -134 -3554 -132 -3552
rect -118 -3554 -116 -3552
rect -110 -3554 -108 -3552
rect -100 -3554 -98 -3552
rect -84 -3554 -82 -3552
rect -74 -3554 -72 -3552
rect -66 -3554 -64 -3552
rect -56 -3554 -54 -3552
rect -40 -3554 -38 -3552
rect -32 -3554 -30 -3552
rect -16 -3554 -14 -3552
rect 0 -3554 2 -3552
rect 8 -3554 10 -3552
rect 18 -3554 20 -3552
rect 214 -3554 216 -3552
rect 224 -3554 226 -3552
rect 240 -3554 242 -3552
rect 250 -3554 252 -3552
rect 266 -3554 268 -3552
rect 276 -3554 278 -3552
rect 284 -3554 286 -3552
rect 294 -3554 296 -3552
rect 310 -3554 312 -3552
rect 318 -3554 320 -3552
rect 328 -3554 330 -3552
rect 344 -3554 346 -3552
rect 354 -3554 356 -3552
rect 362 -3554 364 -3552
rect 372 -3554 374 -3552
rect 388 -3554 390 -3552
rect 396 -3554 398 -3552
rect 412 -3554 414 -3552
rect 428 -3554 430 -3552
rect 436 -3554 438 -3552
rect 446 -3554 448 -3552
rect 570 -3554 572 -3552
rect 580 -3554 582 -3552
rect 596 -3554 598 -3552
rect 606 -3554 608 -3552
rect 622 -3554 624 -3552
rect 632 -3554 634 -3552
rect 640 -3554 642 -3552
rect 650 -3554 652 -3552
rect 666 -3554 668 -3552
rect 674 -3554 676 -3552
rect 684 -3554 686 -3552
rect 700 -3554 702 -3552
rect 710 -3554 712 -3552
rect 718 -3554 720 -3552
rect 728 -3554 730 -3552
rect 744 -3554 746 -3552
rect 752 -3554 754 -3552
rect 768 -3554 770 -3552
rect 784 -3554 786 -3552
rect 792 -3554 794 -3552
rect 802 -3554 804 -3552
rect 968 -3554 970 -3552
rect 978 -3554 980 -3552
rect 994 -3554 996 -3552
rect 1004 -3554 1006 -3552
rect 1020 -3554 1022 -3552
rect 1030 -3554 1032 -3552
rect 1038 -3554 1040 -3552
rect 1048 -3554 1050 -3552
rect 1064 -3554 1066 -3552
rect 1072 -3554 1074 -3552
rect 1082 -3554 1084 -3552
rect 1098 -3554 1100 -3552
rect 1108 -3554 1110 -3552
rect 1116 -3554 1118 -3552
rect 1126 -3554 1128 -3552
rect 1142 -3554 1144 -3552
rect 1150 -3554 1152 -3552
rect 1166 -3554 1168 -3552
rect 1182 -3554 1184 -3552
rect 1190 -3554 1192 -3552
rect 1200 -3554 1202 -3552
rect 1326 -3554 1328 -3552
rect 1336 -3554 1338 -3552
rect 1352 -3554 1354 -3552
rect 1362 -3554 1364 -3552
rect 1378 -3554 1380 -3552
rect 1388 -3554 1390 -3552
rect 1396 -3554 1398 -3552
rect 1406 -3554 1408 -3552
rect 1422 -3554 1424 -3552
rect 1430 -3554 1432 -3552
rect 1440 -3554 1442 -3552
rect 1456 -3554 1458 -3552
rect 1466 -3554 1468 -3552
rect 1474 -3554 1476 -3552
rect 1484 -3554 1486 -3552
rect 1500 -3554 1502 -3552
rect 1508 -3554 1510 -3552
rect 1524 -3554 1526 -3552
rect 1540 -3554 1542 -3552
rect 1548 -3554 1550 -3552
rect 1558 -3554 1560 -3552
rect -1259 -3630 -1257 -3562
rect -1249 -3630 -1247 -3562
rect -1233 -3630 -1231 -3562
rect -1223 -3630 -1221 -3562
rect -1215 -3630 -1213 -3562
rect -1205 -3630 -1203 -3562
rect -1189 -3630 -1187 -3562
rect -1181 -3630 -1179 -3562
rect -1171 -3630 -1169 -3562
rect -930 -3630 -928 -3562
rect -920 -3630 -918 -3562
rect -904 -3630 -902 -3562
rect -894 -3630 -892 -3562
rect -878 -3630 -876 -3562
rect -868 -3630 -866 -3562
rect -860 -3630 -858 -3562
rect -850 -3630 -848 -3562
rect -834 -3630 -832 -3562
rect -826 -3630 -824 -3562
rect -816 -3630 -814 -3562
rect -800 -3630 -798 -3562
rect -790 -3630 -788 -3562
rect -782 -3630 -780 -3562
rect -772 -3630 -770 -3562
rect -756 -3630 -754 -3562
rect -748 -3630 -746 -3562
rect -732 -3630 -730 -3562
rect -716 -3630 -714 -3562
rect -708 -3630 -706 -3562
rect -698 -3630 -696 -3562
rect -572 -3630 -570 -3562
rect -562 -3630 -560 -3562
rect -546 -3630 -544 -3562
rect -536 -3630 -534 -3562
rect -520 -3630 -518 -3562
rect -510 -3630 -508 -3562
rect -502 -3630 -500 -3562
rect -492 -3630 -490 -3562
rect -476 -3630 -474 -3562
rect -468 -3630 -466 -3562
rect -458 -3630 -456 -3562
rect -442 -3630 -440 -3562
rect -432 -3630 -430 -3562
rect -424 -3630 -422 -3562
rect -414 -3630 -412 -3562
rect -398 -3630 -396 -3562
rect -390 -3630 -388 -3562
rect -374 -3630 -372 -3562
rect -358 -3630 -356 -3562
rect -350 -3630 -348 -3562
rect -340 -3630 -338 -3562
rect -214 -3630 -212 -3562
rect -204 -3630 -202 -3562
rect -188 -3630 -186 -3562
rect -178 -3630 -176 -3562
rect -162 -3630 -160 -3562
rect -152 -3630 -150 -3562
rect -144 -3630 -142 -3562
rect -134 -3630 -132 -3562
rect -118 -3630 -116 -3562
rect -110 -3630 -108 -3562
rect -100 -3630 -98 -3562
rect -84 -3630 -82 -3562
rect -74 -3630 -72 -3562
rect -66 -3630 -64 -3562
rect -56 -3630 -54 -3562
rect -40 -3630 -38 -3562
rect -32 -3630 -30 -3562
rect -16 -3630 -14 -3562
rect 0 -3630 2 -3562
rect 8 -3630 10 -3562
rect 18 -3630 20 -3562
rect 214 -3630 216 -3562
rect 224 -3630 226 -3562
rect 240 -3630 242 -3562
rect 250 -3630 252 -3562
rect 266 -3630 268 -3562
rect 276 -3630 278 -3562
rect 284 -3630 286 -3562
rect 294 -3630 296 -3562
rect 310 -3630 312 -3562
rect 318 -3630 320 -3562
rect 328 -3630 330 -3562
rect 344 -3630 346 -3562
rect 354 -3630 356 -3562
rect 362 -3630 364 -3562
rect 372 -3630 374 -3562
rect 388 -3630 390 -3562
rect 396 -3630 398 -3562
rect 412 -3630 414 -3562
rect 428 -3630 430 -3562
rect 436 -3630 438 -3562
rect 446 -3630 448 -3562
rect 570 -3630 572 -3562
rect 580 -3630 582 -3562
rect 596 -3630 598 -3562
rect 606 -3630 608 -3562
rect 622 -3630 624 -3562
rect 632 -3630 634 -3562
rect 640 -3630 642 -3562
rect 650 -3630 652 -3562
rect 666 -3630 668 -3562
rect 674 -3630 676 -3562
rect 684 -3630 686 -3562
rect 700 -3630 702 -3562
rect 710 -3630 712 -3562
rect 718 -3630 720 -3562
rect 728 -3630 730 -3562
rect 744 -3630 746 -3562
rect 752 -3630 754 -3562
rect 768 -3630 770 -3562
rect 784 -3630 786 -3562
rect 792 -3630 794 -3562
rect 802 -3630 804 -3562
rect 968 -3630 970 -3562
rect 978 -3630 980 -3562
rect 994 -3630 996 -3562
rect 1004 -3630 1006 -3562
rect 1020 -3630 1022 -3562
rect 1030 -3630 1032 -3562
rect 1038 -3630 1040 -3562
rect 1048 -3630 1050 -3562
rect 1064 -3630 1066 -3562
rect 1072 -3630 1074 -3562
rect 1082 -3630 1084 -3562
rect 1098 -3630 1100 -3562
rect 1108 -3630 1110 -3562
rect 1116 -3630 1118 -3562
rect 1126 -3630 1128 -3562
rect 1142 -3630 1144 -3562
rect 1150 -3630 1152 -3562
rect 1166 -3630 1168 -3562
rect 1182 -3630 1184 -3562
rect 1190 -3630 1192 -3562
rect 1200 -3630 1202 -3562
rect 1326 -3630 1328 -3562
rect 1336 -3630 1338 -3562
rect 1352 -3630 1354 -3562
rect 1362 -3630 1364 -3562
rect 1378 -3630 1380 -3562
rect 1388 -3630 1390 -3562
rect 1396 -3630 1398 -3562
rect 1406 -3630 1408 -3562
rect 1422 -3630 1424 -3562
rect 1430 -3630 1432 -3562
rect 1440 -3630 1442 -3562
rect 1456 -3630 1458 -3562
rect 1466 -3630 1468 -3562
rect 1474 -3630 1476 -3562
rect 1484 -3630 1486 -3562
rect 1500 -3630 1502 -3562
rect 1508 -3630 1510 -3562
rect 1524 -3630 1526 -3562
rect 1540 -3630 1542 -3562
rect 1548 -3630 1550 -3562
rect 1558 -3630 1560 -3562
rect -1259 -3636 -1257 -3634
rect -1249 -3636 -1247 -3634
rect -1233 -3636 -1231 -3634
rect -1223 -3636 -1221 -3634
rect -1215 -3636 -1213 -3634
rect -1205 -3636 -1203 -3634
rect -1189 -3636 -1187 -3634
rect -1181 -3636 -1179 -3634
rect -1171 -3636 -1169 -3634
rect -930 -3636 -928 -3634
rect -920 -3636 -918 -3634
rect -904 -3636 -902 -3634
rect -894 -3636 -892 -3634
rect -878 -3636 -876 -3634
rect -868 -3636 -866 -3634
rect -860 -3636 -858 -3634
rect -850 -3636 -848 -3634
rect -834 -3636 -832 -3634
rect -826 -3636 -824 -3634
rect -816 -3636 -814 -3634
rect -800 -3636 -798 -3634
rect -790 -3636 -788 -3634
rect -782 -3636 -780 -3634
rect -772 -3636 -770 -3634
rect -756 -3636 -754 -3634
rect -748 -3636 -746 -3634
rect -732 -3636 -730 -3634
rect -716 -3636 -714 -3634
rect -708 -3636 -706 -3634
rect -698 -3636 -696 -3634
rect -572 -3636 -570 -3634
rect -562 -3636 -560 -3634
rect -546 -3636 -544 -3634
rect -536 -3636 -534 -3634
rect -520 -3636 -518 -3634
rect -510 -3636 -508 -3634
rect -502 -3636 -500 -3634
rect -492 -3636 -490 -3634
rect -476 -3636 -474 -3634
rect -468 -3636 -466 -3634
rect -458 -3636 -456 -3634
rect -442 -3636 -440 -3634
rect -432 -3636 -430 -3634
rect -424 -3636 -422 -3634
rect -414 -3636 -412 -3634
rect -398 -3636 -396 -3634
rect -390 -3636 -388 -3634
rect -374 -3636 -372 -3634
rect -358 -3636 -356 -3634
rect -350 -3636 -348 -3634
rect -340 -3636 -338 -3634
rect -214 -3636 -212 -3634
rect -204 -3636 -202 -3634
rect -188 -3636 -186 -3634
rect -178 -3636 -176 -3634
rect -162 -3636 -160 -3634
rect -152 -3636 -150 -3634
rect -144 -3636 -142 -3634
rect -134 -3636 -132 -3634
rect -118 -3636 -116 -3634
rect -110 -3636 -108 -3634
rect -100 -3636 -98 -3634
rect -84 -3636 -82 -3634
rect -74 -3636 -72 -3634
rect -66 -3636 -64 -3634
rect -56 -3636 -54 -3634
rect -40 -3636 -38 -3634
rect -32 -3636 -30 -3634
rect -16 -3636 -14 -3634
rect 0 -3636 2 -3634
rect 8 -3636 10 -3634
rect 18 -3636 20 -3634
rect 214 -3636 216 -3634
rect 224 -3636 226 -3634
rect 240 -3636 242 -3634
rect 250 -3636 252 -3634
rect 266 -3636 268 -3634
rect 276 -3636 278 -3634
rect 284 -3636 286 -3634
rect 294 -3636 296 -3634
rect 310 -3636 312 -3634
rect 318 -3636 320 -3634
rect 328 -3636 330 -3634
rect 344 -3636 346 -3634
rect 354 -3636 356 -3634
rect 362 -3636 364 -3634
rect 372 -3636 374 -3634
rect 388 -3636 390 -3634
rect 396 -3636 398 -3634
rect 412 -3636 414 -3634
rect 428 -3636 430 -3634
rect 436 -3636 438 -3634
rect 446 -3636 448 -3634
rect 570 -3636 572 -3634
rect 580 -3636 582 -3634
rect 596 -3636 598 -3634
rect 606 -3636 608 -3634
rect 622 -3636 624 -3634
rect 632 -3636 634 -3634
rect 640 -3636 642 -3634
rect 650 -3636 652 -3634
rect 666 -3636 668 -3634
rect 674 -3636 676 -3634
rect 684 -3636 686 -3634
rect 700 -3636 702 -3634
rect 710 -3636 712 -3634
rect 718 -3636 720 -3634
rect 728 -3636 730 -3634
rect 744 -3636 746 -3634
rect 752 -3636 754 -3634
rect 768 -3636 770 -3634
rect 784 -3636 786 -3634
rect 792 -3636 794 -3634
rect 802 -3636 804 -3634
rect 968 -3636 970 -3634
rect 978 -3636 980 -3634
rect 994 -3636 996 -3634
rect 1004 -3636 1006 -3634
rect 1020 -3636 1022 -3634
rect 1030 -3636 1032 -3634
rect 1038 -3636 1040 -3634
rect 1048 -3636 1050 -3634
rect 1064 -3636 1066 -3634
rect 1072 -3636 1074 -3634
rect 1082 -3636 1084 -3634
rect 1098 -3636 1100 -3634
rect 1108 -3636 1110 -3634
rect 1116 -3636 1118 -3634
rect 1126 -3636 1128 -3634
rect 1142 -3636 1144 -3634
rect 1150 -3636 1152 -3634
rect 1166 -3636 1168 -3634
rect 1182 -3636 1184 -3634
rect 1190 -3636 1192 -3634
rect 1200 -3636 1202 -3634
rect 1326 -3636 1328 -3634
rect 1336 -3636 1338 -3634
rect 1352 -3636 1354 -3634
rect 1362 -3636 1364 -3634
rect 1378 -3636 1380 -3634
rect 1388 -3636 1390 -3634
rect 1396 -3636 1398 -3634
rect 1406 -3636 1408 -3634
rect 1422 -3636 1424 -3634
rect 1430 -3636 1432 -3634
rect 1440 -3636 1442 -3634
rect 1456 -3636 1458 -3634
rect 1466 -3636 1468 -3634
rect 1474 -3636 1476 -3634
rect 1484 -3636 1486 -3634
rect 1500 -3636 1502 -3634
rect 1508 -3636 1510 -3634
rect 1524 -3636 1526 -3634
rect 1540 -3636 1542 -3634
rect 1548 -3636 1550 -3634
rect 1558 -3636 1560 -3634
rect -1259 -3684 -1257 -3682
rect -1249 -3684 -1247 -3682
rect -1233 -3684 -1231 -3682
rect -1225 -3684 -1223 -3682
rect -1209 -3684 -1207 -3682
rect -1201 -3684 -1199 -3682
rect -1191 -3684 -1189 -3682
rect -1183 -3684 -1181 -3682
rect -1167 -3684 -1165 -3682
rect -1159 -3684 -1157 -3682
rect -1149 -3684 -1147 -3682
rect -1141 -3684 -1139 -3682
rect -1125 -3684 -1123 -3682
rect -1117 -3684 -1115 -3682
rect -1107 -3684 -1105 -3682
rect -1099 -3684 -1097 -3682
rect -1083 -3684 -1081 -3682
rect -1075 -3684 -1073 -3682
rect -930 -3684 -928 -3682
rect -920 -3684 -918 -3682
rect -904 -3684 -902 -3682
rect -896 -3684 -894 -3682
rect -880 -3684 -878 -3682
rect -872 -3684 -870 -3682
rect -862 -3684 -860 -3682
rect -854 -3684 -852 -3682
rect -838 -3684 -836 -3682
rect -830 -3684 -828 -3682
rect -820 -3684 -818 -3682
rect -812 -3684 -810 -3682
rect -796 -3684 -794 -3682
rect -788 -3684 -786 -3682
rect -778 -3684 -776 -3682
rect -770 -3684 -768 -3682
rect -754 -3684 -752 -3682
rect -746 -3684 -744 -3682
rect -572 -3684 -570 -3682
rect -562 -3684 -560 -3682
rect -546 -3684 -544 -3682
rect -538 -3684 -536 -3682
rect -522 -3684 -520 -3682
rect -514 -3684 -512 -3682
rect -504 -3684 -502 -3682
rect -496 -3684 -494 -3682
rect -480 -3684 -478 -3682
rect -472 -3684 -470 -3682
rect -462 -3684 -460 -3682
rect -454 -3684 -452 -3682
rect -438 -3684 -436 -3682
rect -430 -3684 -428 -3682
rect -420 -3684 -418 -3682
rect -412 -3684 -410 -3682
rect -396 -3684 -394 -3682
rect -388 -3684 -386 -3682
rect -214 -3684 -212 -3682
rect -204 -3684 -202 -3682
rect -188 -3684 -186 -3682
rect -180 -3684 -178 -3682
rect -164 -3684 -162 -3682
rect -156 -3684 -154 -3682
rect -146 -3684 -144 -3682
rect -138 -3684 -136 -3682
rect -122 -3684 -120 -3682
rect -114 -3684 -112 -3682
rect -104 -3684 -102 -3682
rect -96 -3684 -94 -3682
rect -80 -3684 -78 -3682
rect -72 -3684 -70 -3682
rect -62 -3684 -60 -3682
rect -54 -3684 -52 -3682
rect -38 -3684 -36 -3682
rect -30 -3684 -28 -3682
rect -1259 -3760 -1257 -3692
rect -1249 -3760 -1247 -3692
rect -1233 -3760 -1231 -3692
rect -1225 -3760 -1223 -3692
rect -1209 -3760 -1207 -3692
rect -1201 -3760 -1199 -3692
rect -1191 -3760 -1189 -3692
rect -1183 -3760 -1181 -3692
rect -1167 -3760 -1165 -3692
rect -1159 -3725 -1157 -3692
rect -1149 -3725 -1147 -3692
rect -1159 -3727 -1147 -3725
rect -1159 -3760 -1157 -3727
rect -1149 -3760 -1147 -3727
rect -1141 -3760 -1139 -3692
rect -1125 -3760 -1123 -3692
rect -1117 -3760 -1115 -3692
rect -1107 -3760 -1105 -3692
rect -1099 -3760 -1097 -3692
rect -1083 -3760 -1081 -3692
rect -1075 -3760 -1073 -3692
rect -930 -3760 -928 -3692
rect -920 -3760 -918 -3692
rect -904 -3760 -902 -3692
rect -896 -3760 -894 -3692
rect -880 -3760 -878 -3692
rect -872 -3760 -870 -3692
rect -862 -3760 -860 -3692
rect -854 -3760 -852 -3692
rect -838 -3760 -836 -3692
rect -830 -3725 -828 -3692
rect -820 -3725 -818 -3692
rect -830 -3727 -818 -3725
rect -830 -3760 -828 -3727
rect -820 -3760 -818 -3727
rect -812 -3760 -810 -3692
rect -796 -3760 -794 -3692
rect -788 -3760 -786 -3692
rect -778 -3760 -776 -3692
rect -770 -3760 -768 -3692
rect -754 -3760 -752 -3692
rect -746 -3760 -744 -3692
rect -572 -3760 -570 -3692
rect -562 -3760 -560 -3692
rect -546 -3760 -544 -3692
rect -538 -3760 -536 -3692
rect -522 -3760 -520 -3692
rect -514 -3760 -512 -3692
rect -504 -3760 -502 -3692
rect -496 -3760 -494 -3692
rect -480 -3760 -478 -3692
rect -472 -3725 -470 -3692
rect -462 -3725 -460 -3692
rect -472 -3727 -460 -3725
rect -472 -3760 -470 -3727
rect -462 -3760 -460 -3727
rect -454 -3760 -452 -3692
rect -438 -3760 -436 -3692
rect -430 -3760 -428 -3692
rect -420 -3760 -418 -3692
rect -412 -3760 -410 -3692
rect -396 -3760 -394 -3692
rect -388 -3760 -386 -3692
rect -214 -3760 -212 -3692
rect -204 -3760 -202 -3692
rect -188 -3760 -186 -3692
rect -180 -3760 -178 -3692
rect -164 -3760 -162 -3692
rect -156 -3760 -154 -3692
rect -146 -3760 -144 -3692
rect -138 -3760 -136 -3692
rect -122 -3760 -120 -3692
rect -114 -3725 -112 -3692
rect -104 -3725 -102 -3692
rect -114 -3727 -102 -3725
rect -114 -3760 -112 -3727
rect -104 -3760 -102 -3727
rect -96 -3760 -94 -3692
rect -80 -3760 -78 -3692
rect -72 -3760 -70 -3692
rect -62 -3760 -60 -3692
rect -54 -3760 -52 -3692
rect -38 -3760 -36 -3692
rect -30 -3760 -28 -3692
rect -1259 -3766 -1257 -3764
rect -1249 -3766 -1247 -3764
rect -1233 -3766 -1231 -3764
rect -1225 -3766 -1223 -3764
rect -1209 -3766 -1207 -3764
rect -1201 -3766 -1199 -3764
rect -1191 -3766 -1189 -3764
rect -1183 -3766 -1181 -3764
rect -1167 -3766 -1165 -3764
rect -1159 -3766 -1157 -3764
rect -1149 -3766 -1147 -3764
rect -1141 -3766 -1139 -3764
rect -1125 -3766 -1123 -3764
rect -1117 -3766 -1115 -3764
rect -1107 -3766 -1105 -3764
rect -1099 -3766 -1097 -3764
rect -1083 -3766 -1081 -3764
rect -1075 -3766 -1073 -3764
rect -930 -3766 -928 -3764
rect -920 -3766 -918 -3764
rect -904 -3766 -902 -3764
rect -896 -3766 -894 -3764
rect -880 -3766 -878 -3764
rect -872 -3766 -870 -3764
rect -862 -3766 -860 -3764
rect -854 -3766 -852 -3764
rect -838 -3766 -836 -3764
rect -830 -3766 -828 -3764
rect -820 -3766 -818 -3764
rect -812 -3766 -810 -3764
rect -796 -3766 -794 -3764
rect -788 -3766 -786 -3764
rect -778 -3766 -776 -3764
rect -770 -3766 -768 -3764
rect -754 -3766 -752 -3764
rect -746 -3766 -744 -3764
rect -572 -3766 -570 -3764
rect -562 -3766 -560 -3764
rect -546 -3766 -544 -3764
rect -538 -3766 -536 -3764
rect -522 -3766 -520 -3764
rect -514 -3766 -512 -3764
rect -504 -3766 -502 -3764
rect -496 -3766 -494 -3764
rect -480 -3766 -478 -3764
rect -472 -3766 -470 -3764
rect -462 -3766 -460 -3764
rect -454 -3766 -452 -3764
rect -438 -3766 -436 -3764
rect -430 -3766 -428 -3764
rect -420 -3766 -418 -3764
rect -412 -3766 -410 -3764
rect -396 -3766 -394 -3764
rect -388 -3766 -386 -3764
rect -214 -3766 -212 -3764
rect -204 -3766 -202 -3764
rect -188 -3766 -186 -3764
rect -180 -3766 -178 -3764
rect -164 -3766 -162 -3764
rect -156 -3766 -154 -3764
rect -146 -3766 -144 -3764
rect -138 -3766 -136 -3764
rect -122 -3766 -120 -3764
rect -114 -3766 -112 -3764
rect -104 -3766 -102 -3764
rect -96 -3766 -94 -3764
rect -80 -3766 -78 -3764
rect -72 -3766 -70 -3764
rect -62 -3766 -60 -3764
rect -54 -3766 -52 -3764
rect -38 -3766 -36 -3764
rect -30 -3766 -28 -3764
rect 73 -3799 75 -3797
rect 73 -3863 75 -3831
rect 73 -3881 75 -3879
rect -1259 -3915 -1257 -3913
rect -1249 -3915 -1247 -3913
rect -1233 -3915 -1231 -3913
rect -1225 -3915 -1223 -3913
rect -1209 -3915 -1207 -3913
rect -1201 -3915 -1199 -3913
rect -1191 -3915 -1189 -3913
rect -1183 -3915 -1181 -3913
rect -1167 -3915 -1165 -3913
rect -1159 -3915 -1157 -3913
rect -1149 -3915 -1147 -3913
rect -1141 -3915 -1139 -3913
rect -1125 -3915 -1123 -3913
rect -1117 -3915 -1115 -3913
rect -1107 -3915 -1105 -3913
rect -1099 -3915 -1097 -3913
rect -1083 -3915 -1081 -3913
rect -1075 -3915 -1073 -3913
rect -930 -3915 -928 -3913
rect -920 -3915 -918 -3913
rect -904 -3915 -902 -3913
rect -896 -3915 -894 -3913
rect -880 -3915 -878 -3913
rect -872 -3915 -870 -3913
rect -862 -3915 -860 -3913
rect -854 -3915 -852 -3913
rect -838 -3915 -836 -3913
rect -830 -3915 -828 -3913
rect -820 -3915 -818 -3913
rect -812 -3915 -810 -3913
rect -796 -3915 -794 -3913
rect -788 -3915 -786 -3913
rect -778 -3915 -776 -3913
rect -770 -3915 -768 -3913
rect -754 -3915 -752 -3913
rect -746 -3915 -744 -3913
rect -572 -3915 -570 -3913
rect -562 -3915 -560 -3913
rect -546 -3915 -544 -3913
rect -538 -3915 -536 -3913
rect -522 -3915 -520 -3913
rect -514 -3915 -512 -3913
rect -504 -3915 -502 -3913
rect -496 -3915 -494 -3913
rect -480 -3915 -478 -3913
rect -472 -3915 -470 -3913
rect -462 -3915 -460 -3913
rect -454 -3915 -452 -3913
rect -438 -3915 -436 -3913
rect -430 -3915 -428 -3913
rect -420 -3915 -418 -3913
rect -412 -3915 -410 -3913
rect -396 -3915 -394 -3913
rect -388 -3915 -386 -3913
rect -214 -3915 -212 -3913
rect -204 -3915 -202 -3913
rect -188 -3915 -186 -3913
rect -180 -3915 -178 -3913
rect -164 -3915 -162 -3913
rect -156 -3915 -154 -3913
rect -146 -3915 -144 -3913
rect -138 -3915 -136 -3913
rect -122 -3915 -120 -3913
rect -114 -3915 -112 -3913
rect -104 -3915 -102 -3913
rect -96 -3915 -94 -3913
rect -80 -3915 -78 -3913
rect -72 -3915 -70 -3913
rect -62 -3915 -60 -3913
rect -54 -3915 -52 -3913
rect -38 -3915 -36 -3913
rect -30 -3915 -28 -3913
rect 214 -3915 216 -3913
rect 224 -3915 226 -3913
rect 240 -3915 242 -3913
rect 248 -3915 250 -3913
rect 264 -3915 266 -3913
rect 272 -3915 274 -3913
rect 282 -3915 284 -3913
rect 290 -3915 292 -3913
rect 306 -3915 308 -3913
rect 314 -3915 316 -3913
rect 324 -3915 326 -3913
rect 332 -3915 334 -3913
rect 348 -3915 350 -3913
rect 356 -3915 358 -3913
rect 366 -3915 368 -3913
rect 374 -3915 376 -3913
rect 390 -3915 392 -3913
rect 398 -3915 400 -3913
rect 570 -3915 572 -3913
rect 580 -3915 582 -3913
rect 596 -3915 598 -3913
rect 604 -3915 606 -3913
rect 620 -3915 622 -3913
rect 628 -3915 630 -3913
rect 638 -3915 640 -3913
rect 646 -3915 648 -3913
rect 662 -3915 664 -3913
rect 670 -3915 672 -3913
rect 680 -3915 682 -3913
rect 688 -3915 690 -3913
rect 704 -3915 706 -3913
rect 712 -3915 714 -3913
rect 722 -3915 724 -3913
rect 730 -3915 732 -3913
rect 746 -3915 748 -3913
rect 754 -3915 756 -3913
rect 968 -3915 970 -3913
rect 978 -3915 980 -3913
rect 994 -3915 996 -3913
rect 1002 -3915 1004 -3913
rect 1018 -3915 1020 -3913
rect 1026 -3915 1028 -3913
rect 1036 -3915 1038 -3913
rect 1044 -3915 1046 -3913
rect 1060 -3915 1062 -3913
rect 1068 -3915 1070 -3913
rect 1078 -3915 1080 -3913
rect 1086 -3915 1088 -3913
rect 1102 -3915 1104 -3913
rect 1110 -3915 1112 -3913
rect 1120 -3915 1122 -3913
rect 1128 -3915 1130 -3913
rect 1144 -3915 1146 -3913
rect 1152 -3915 1154 -3913
rect 1326 -3915 1328 -3913
rect 1336 -3915 1338 -3913
rect 1352 -3915 1354 -3913
rect 1360 -3915 1362 -3913
rect 1376 -3915 1378 -3913
rect 1384 -3915 1386 -3913
rect 1394 -3915 1396 -3913
rect 1402 -3915 1404 -3913
rect 1418 -3915 1420 -3913
rect 1426 -3915 1428 -3913
rect 1436 -3915 1438 -3913
rect 1444 -3915 1446 -3913
rect 1460 -3915 1462 -3913
rect 1468 -3915 1470 -3913
rect 1478 -3915 1480 -3913
rect 1486 -3915 1488 -3913
rect 1502 -3915 1504 -3913
rect 1510 -3915 1512 -3913
rect -1259 -3991 -1257 -3923
rect -1249 -3991 -1247 -3923
rect -1233 -3991 -1231 -3923
rect -1225 -3991 -1223 -3923
rect -1209 -3991 -1207 -3923
rect -1201 -3991 -1199 -3923
rect -1191 -3991 -1189 -3923
rect -1183 -3991 -1181 -3923
rect -1167 -3991 -1165 -3923
rect -1159 -3956 -1157 -3923
rect -1149 -3956 -1147 -3923
rect -1159 -3958 -1147 -3956
rect -1159 -3991 -1157 -3958
rect -1149 -3991 -1147 -3958
rect -1141 -3991 -1139 -3923
rect -1125 -3991 -1123 -3923
rect -1117 -3991 -1115 -3923
rect -1107 -3991 -1105 -3923
rect -1099 -3991 -1097 -3923
rect -1083 -3991 -1081 -3923
rect -1075 -3991 -1073 -3923
rect -930 -3991 -928 -3923
rect -920 -3991 -918 -3923
rect -904 -3991 -902 -3923
rect -896 -3991 -894 -3923
rect -880 -3991 -878 -3923
rect -872 -3991 -870 -3923
rect -862 -3991 -860 -3923
rect -854 -3991 -852 -3923
rect -838 -3991 -836 -3923
rect -830 -3956 -828 -3923
rect -820 -3956 -818 -3923
rect -830 -3958 -818 -3956
rect -830 -3991 -828 -3958
rect -820 -3991 -818 -3958
rect -812 -3991 -810 -3923
rect -796 -3991 -794 -3923
rect -788 -3991 -786 -3923
rect -778 -3991 -776 -3923
rect -770 -3991 -768 -3923
rect -754 -3991 -752 -3923
rect -746 -3991 -744 -3923
rect -572 -3991 -570 -3923
rect -562 -3991 -560 -3923
rect -546 -3991 -544 -3923
rect -538 -3991 -536 -3923
rect -522 -3991 -520 -3923
rect -514 -3991 -512 -3923
rect -504 -3991 -502 -3923
rect -496 -3991 -494 -3923
rect -480 -3991 -478 -3923
rect -472 -3956 -470 -3923
rect -462 -3956 -460 -3923
rect -472 -3958 -460 -3956
rect -472 -3991 -470 -3958
rect -462 -3991 -460 -3958
rect -454 -3991 -452 -3923
rect -438 -3991 -436 -3923
rect -430 -3991 -428 -3923
rect -420 -3991 -418 -3923
rect -412 -3991 -410 -3923
rect -396 -3991 -394 -3923
rect -388 -3991 -386 -3923
rect -214 -3991 -212 -3923
rect -204 -3991 -202 -3923
rect -188 -3991 -186 -3923
rect -180 -3991 -178 -3923
rect -164 -3991 -162 -3923
rect -156 -3991 -154 -3923
rect -146 -3991 -144 -3923
rect -138 -3991 -136 -3923
rect -122 -3991 -120 -3923
rect -114 -3956 -112 -3923
rect -104 -3956 -102 -3923
rect -114 -3958 -102 -3956
rect -114 -3991 -112 -3958
rect -104 -3991 -102 -3958
rect -96 -3991 -94 -3923
rect -80 -3991 -78 -3923
rect -72 -3991 -70 -3923
rect -62 -3991 -60 -3923
rect -54 -3991 -52 -3923
rect -38 -3991 -36 -3923
rect -30 -3991 -28 -3923
rect 214 -3991 216 -3923
rect 224 -3991 226 -3923
rect 240 -3991 242 -3923
rect 248 -3991 250 -3923
rect 264 -3991 266 -3923
rect 272 -3991 274 -3923
rect 282 -3991 284 -3923
rect 290 -3991 292 -3923
rect 306 -3991 308 -3923
rect 314 -3956 316 -3923
rect 324 -3956 326 -3923
rect 314 -3958 326 -3956
rect 314 -3991 316 -3958
rect 324 -3991 326 -3958
rect 332 -3991 334 -3923
rect 348 -3991 350 -3923
rect 356 -3991 358 -3923
rect 366 -3991 368 -3923
rect 374 -3991 376 -3923
rect 390 -3991 392 -3923
rect 398 -3991 400 -3923
rect 570 -3991 572 -3923
rect 580 -3991 582 -3923
rect 596 -3991 598 -3923
rect 604 -3991 606 -3923
rect 620 -3991 622 -3923
rect 628 -3991 630 -3923
rect 638 -3991 640 -3923
rect 646 -3991 648 -3923
rect 662 -3991 664 -3923
rect 670 -3956 672 -3923
rect 680 -3956 682 -3923
rect 670 -3958 682 -3956
rect 670 -3991 672 -3958
rect 680 -3991 682 -3958
rect 688 -3991 690 -3923
rect 704 -3991 706 -3923
rect 712 -3991 714 -3923
rect 722 -3991 724 -3923
rect 730 -3991 732 -3923
rect 746 -3991 748 -3923
rect 754 -3991 756 -3923
rect 968 -3991 970 -3923
rect 978 -3991 980 -3923
rect 994 -3991 996 -3923
rect 1002 -3991 1004 -3923
rect 1018 -3991 1020 -3923
rect 1026 -3991 1028 -3923
rect 1036 -3991 1038 -3923
rect 1044 -3991 1046 -3923
rect 1060 -3991 1062 -3923
rect 1068 -3956 1070 -3923
rect 1078 -3956 1080 -3923
rect 1068 -3958 1080 -3956
rect 1068 -3991 1070 -3958
rect 1078 -3991 1080 -3958
rect 1086 -3991 1088 -3923
rect 1102 -3991 1104 -3923
rect 1110 -3991 1112 -3923
rect 1120 -3991 1122 -3923
rect 1128 -3991 1130 -3923
rect 1144 -3991 1146 -3923
rect 1152 -3991 1154 -3923
rect 1326 -3991 1328 -3923
rect 1336 -3991 1338 -3923
rect 1352 -3991 1354 -3923
rect 1360 -3991 1362 -3923
rect 1376 -3991 1378 -3923
rect 1384 -3991 1386 -3923
rect 1394 -3991 1396 -3923
rect 1402 -3991 1404 -3923
rect 1418 -3991 1420 -3923
rect 1426 -3956 1428 -3923
rect 1436 -3956 1438 -3923
rect 1426 -3958 1438 -3956
rect 1426 -3991 1428 -3958
rect 1436 -3991 1438 -3958
rect 1444 -3991 1446 -3923
rect 1460 -3991 1462 -3923
rect 1468 -3991 1470 -3923
rect 1478 -3991 1480 -3923
rect 1486 -3991 1488 -3923
rect 1502 -3991 1504 -3923
rect 1510 -3991 1512 -3923
rect -1259 -3997 -1257 -3995
rect -1249 -3997 -1247 -3995
rect -1233 -3997 -1231 -3995
rect -1225 -3997 -1223 -3995
rect -1209 -3997 -1207 -3995
rect -1201 -3997 -1199 -3995
rect -1191 -3997 -1189 -3995
rect -1183 -3997 -1181 -3995
rect -1167 -3997 -1165 -3995
rect -1159 -3997 -1157 -3995
rect -1149 -3997 -1147 -3995
rect -1141 -3997 -1139 -3995
rect -1125 -3997 -1123 -3995
rect -1117 -3997 -1115 -3995
rect -1107 -3997 -1105 -3995
rect -1099 -3997 -1097 -3995
rect -1083 -3997 -1081 -3995
rect -1075 -3997 -1073 -3995
rect -930 -3997 -928 -3995
rect -920 -3997 -918 -3995
rect -904 -3997 -902 -3995
rect -896 -3997 -894 -3995
rect -880 -3997 -878 -3995
rect -872 -3997 -870 -3995
rect -862 -3997 -860 -3995
rect -854 -3997 -852 -3995
rect -838 -3997 -836 -3995
rect -830 -3997 -828 -3995
rect -820 -3997 -818 -3995
rect -812 -3997 -810 -3995
rect -796 -3997 -794 -3995
rect -788 -3997 -786 -3995
rect -778 -3997 -776 -3995
rect -770 -3997 -768 -3995
rect -754 -3997 -752 -3995
rect -746 -3997 -744 -3995
rect -572 -3997 -570 -3995
rect -562 -3997 -560 -3995
rect -546 -3997 -544 -3995
rect -538 -3997 -536 -3995
rect -522 -3997 -520 -3995
rect -514 -3997 -512 -3995
rect -504 -3997 -502 -3995
rect -496 -3997 -494 -3995
rect -480 -3997 -478 -3995
rect -472 -3997 -470 -3995
rect -462 -3997 -460 -3995
rect -454 -3997 -452 -3995
rect -438 -3997 -436 -3995
rect -430 -3997 -428 -3995
rect -420 -3997 -418 -3995
rect -412 -3997 -410 -3995
rect -396 -3997 -394 -3995
rect -388 -3997 -386 -3995
rect -214 -3997 -212 -3995
rect -204 -3997 -202 -3995
rect -188 -3997 -186 -3995
rect -180 -3997 -178 -3995
rect -164 -3997 -162 -3995
rect -156 -3997 -154 -3995
rect -146 -3997 -144 -3995
rect -138 -3997 -136 -3995
rect -122 -3997 -120 -3995
rect -114 -3997 -112 -3995
rect -104 -3997 -102 -3995
rect -96 -3997 -94 -3995
rect -80 -3997 -78 -3995
rect -72 -3997 -70 -3995
rect -62 -3997 -60 -3995
rect -54 -3997 -52 -3995
rect -38 -3997 -36 -3995
rect -30 -3997 -28 -3995
rect 214 -3997 216 -3995
rect 224 -3997 226 -3995
rect 240 -3997 242 -3995
rect 248 -3997 250 -3995
rect 264 -3997 266 -3995
rect 272 -3997 274 -3995
rect 282 -3997 284 -3995
rect 290 -3997 292 -3995
rect 306 -3997 308 -3995
rect 314 -3997 316 -3995
rect 324 -3997 326 -3995
rect 332 -3997 334 -3995
rect 348 -3997 350 -3995
rect 356 -3997 358 -3995
rect 366 -3997 368 -3995
rect 374 -3997 376 -3995
rect 390 -3997 392 -3995
rect 398 -3997 400 -3995
rect 570 -3997 572 -3995
rect 580 -3997 582 -3995
rect 596 -3997 598 -3995
rect 604 -3997 606 -3995
rect 620 -3997 622 -3995
rect 628 -3997 630 -3995
rect 638 -3997 640 -3995
rect 646 -3997 648 -3995
rect 662 -3997 664 -3995
rect 670 -3997 672 -3995
rect 680 -3997 682 -3995
rect 688 -3997 690 -3995
rect 704 -3997 706 -3995
rect 712 -3997 714 -3995
rect 722 -3997 724 -3995
rect 730 -3997 732 -3995
rect 746 -3997 748 -3995
rect 754 -3997 756 -3995
rect 968 -3997 970 -3995
rect 978 -3997 980 -3995
rect 994 -3997 996 -3995
rect 1002 -3997 1004 -3995
rect 1018 -3997 1020 -3995
rect 1026 -3997 1028 -3995
rect 1036 -3997 1038 -3995
rect 1044 -3997 1046 -3995
rect 1060 -3997 1062 -3995
rect 1068 -3997 1070 -3995
rect 1078 -3997 1080 -3995
rect 1086 -3997 1088 -3995
rect 1102 -3997 1104 -3995
rect 1110 -3997 1112 -3995
rect 1120 -3997 1122 -3995
rect 1128 -3997 1130 -3995
rect 1144 -3997 1146 -3995
rect 1152 -3997 1154 -3995
rect 1326 -3997 1328 -3995
rect 1336 -3997 1338 -3995
rect 1352 -3997 1354 -3995
rect 1360 -3997 1362 -3995
rect 1376 -3997 1378 -3995
rect 1384 -3997 1386 -3995
rect 1394 -3997 1396 -3995
rect 1402 -3997 1404 -3995
rect 1418 -3997 1420 -3995
rect 1426 -3997 1428 -3995
rect 1436 -3997 1438 -3995
rect 1444 -3997 1446 -3995
rect 1460 -3997 1462 -3995
rect 1468 -3997 1470 -3995
rect 1478 -3997 1480 -3995
rect 1486 -3997 1488 -3995
rect 1502 -3997 1504 -3995
rect 1510 -3997 1512 -3995
rect -1259 -4040 -1257 -4038
rect -1249 -4040 -1247 -4038
rect -1233 -4040 -1231 -4038
rect -1225 -4040 -1223 -4038
rect -1209 -4040 -1207 -4038
rect -1201 -4040 -1199 -4038
rect -1191 -4040 -1189 -4038
rect -1183 -4040 -1181 -4038
rect -1167 -4040 -1165 -4038
rect -1159 -4040 -1157 -4038
rect -1149 -4040 -1147 -4038
rect -1141 -4040 -1139 -4038
rect -1125 -4040 -1123 -4038
rect -1117 -4040 -1115 -4038
rect -1107 -4040 -1105 -4038
rect -1099 -4040 -1097 -4038
rect -1083 -4040 -1081 -4038
rect -1075 -4040 -1073 -4038
rect -930 -4040 -928 -4038
rect -920 -4040 -918 -4038
rect -904 -4040 -902 -4038
rect -896 -4040 -894 -4038
rect -880 -4040 -878 -4038
rect -872 -4040 -870 -4038
rect -862 -4040 -860 -4038
rect -854 -4040 -852 -4038
rect -838 -4040 -836 -4038
rect -830 -4040 -828 -4038
rect -820 -4040 -818 -4038
rect -812 -4040 -810 -4038
rect -796 -4040 -794 -4038
rect -788 -4040 -786 -4038
rect -778 -4040 -776 -4038
rect -770 -4040 -768 -4038
rect -754 -4040 -752 -4038
rect -746 -4040 -744 -4038
rect -572 -4040 -570 -4038
rect -562 -4040 -560 -4038
rect -546 -4040 -544 -4038
rect -538 -4040 -536 -4038
rect -522 -4040 -520 -4038
rect -514 -4040 -512 -4038
rect -504 -4040 -502 -4038
rect -496 -4040 -494 -4038
rect -480 -4040 -478 -4038
rect -472 -4040 -470 -4038
rect -462 -4040 -460 -4038
rect -454 -4040 -452 -4038
rect -438 -4040 -436 -4038
rect -430 -4040 -428 -4038
rect -420 -4040 -418 -4038
rect -412 -4040 -410 -4038
rect -396 -4040 -394 -4038
rect -388 -4040 -386 -4038
rect -214 -4040 -212 -4038
rect -204 -4040 -202 -4038
rect -188 -4040 -186 -4038
rect -180 -4040 -178 -4038
rect -164 -4040 -162 -4038
rect -156 -4040 -154 -4038
rect -146 -4040 -144 -4038
rect -138 -4040 -136 -4038
rect -122 -4040 -120 -4038
rect -114 -4040 -112 -4038
rect -104 -4040 -102 -4038
rect -96 -4040 -94 -4038
rect -80 -4040 -78 -4038
rect -72 -4040 -70 -4038
rect -62 -4040 -60 -4038
rect -54 -4040 -52 -4038
rect -38 -4040 -36 -4038
rect -30 -4040 -28 -4038
rect 214 -4040 216 -4038
rect 224 -4040 226 -4038
rect 240 -4040 242 -4038
rect 248 -4040 250 -4038
rect 264 -4040 266 -4038
rect 272 -4040 274 -4038
rect 282 -4040 284 -4038
rect 290 -4040 292 -4038
rect 306 -4040 308 -4038
rect 314 -4040 316 -4038
rect 324 -4040 326 -4038
rect 332 -4040 334 -4038
rect 348 -4040 350 -4038
rect 356 -4040 358 -4038
rect 366 -4040 368 -4038
rect 374 -4040 376 -4038
rect 390 -4040 392 -4038
rect 398 -4040 400 -4038
rect 570 -4040 572 -4038
rect 580 -4040 582 -4038
rect 596 -4040 598 -4038
rect 604 -4040 606 -4038
rect 620 -4040 622 -4038
rect 628 -4040 630 -4038
rect 638 -4040 640 -4038
rect 646 -4040 648 -4038
rect 662 -4040 664 -4038
rect 670 -4040 672 -4038
rect 680 -4040 682 -4038
rect 688 -4040 690 -4038
rect 704 -4040 706 -4038
rect 712 -4040 714 -4038
rect 722 -4040 724 -4038
rect 730 -4040 732 -4038
rect 746 -4040 748 -4038
rect 754 -4040 756 -4038
rect 968 -4040 970 -4038
rect 978 -4040 980 -4038
rect 994 -4040 996 -4038
rect 1002 -4040 1004 -4038
rect 1018 -4040 1020 -4038
rect 1026 -4040 1028 -4038
rect 1036 -4040 1038 -4038
rect 1044 -4040 1046 -4038
rect 1060 -4040 1062 -4038
rect 1068 -4040 1070 -4038
rect 1078 -4040 1080 -4038
rect 1086 -4040 1088 -4038
rect 1102 -4040 1104 -4038
rect 1110 -4040 1112 -4038
rect 1120 -4040 1122 -4038
rect 1128 -4040 1130 -4038
rect 1144 -4040 1146 -4038
rect 1152 -4040 1154 -4038
rect 1326 -4040 1328 -4038
rect 1336 -4040 1338 -4038
rect 1352 -4040 1354 -4038
rect 1360 -4040 1362 -4038
rect 1376 -4040 1378 -4038
rect 1384 -4040 1386 -4038
rect 1394 -4040 1396 -4038
rect 1402 -4040 1404 -4038
rect 1418 -4040 1420 -4038
rect 1426 -4040 1428 -4038
rect 1436 -4040 1438 -4038
rect 1444 -4040 1446 -4038
rect 1460 -4040 1462 -4038
rect 1468 -4040 1470 -4038
rect 1478 -4040 1480 -4038
rect 1486 -4040 1488 -4038
rect 1502 -4040 1504 -4038
rect 1510 -4040 1512 -4038
rect -1259 -4116 -1257 -4048
rect -1249 -4116 -1247 -4048
rect -1233 -4116 -1231 -4048
rect -1225 -4116 -1223 -4048
rect -1209 -4116 -1207 -4048
rect -1201 -4116 -1199 -4048
rect -1191 -4116 -1189 -4048
rect -1183 -4116 -1181 -4048
rect -1167 -4116 -1165 -4048
rect -1159 -4081 -1157 -4048
rect -1149 -4081 -1147 -4048
rect -1159 -4083 -1147 -4081
rect -1159 -4116 -1157 -4083
rect -1149 -4116 -1147 -4083
rect -1141 -4116 -1139 -4048
rect -1125 -4116 -1123 -4048
rect -1117 -4116 -1115 -4048
rect -1107 -4116 -1105 -4048
rect -1099 -4116 -1097 -4048
rect -1083 -4116 -1081 -4048
rect -1075 -4116 -1073 -4048
rect -930 -4116 -928 -4048
rect -920 -4116 -918 -4048
rect -904 -4116 -902 -4048
rect -896 -4116 -894 -4048
rect -880 -4116 -878 -4048
rect -872 -4116 -870 -4048
rect -862 -4116 -860 -4048
rect -854 -4116 -852 -4048
rect -838 -4116 -836 -4048
rect -830 -4081 -828 -4048
rect -820 -4081 -818 -4048
rect -830 -4083 -818 -4081
rect -830 -4116 -828 -4083
rect -820 -4116 -818 -4083
rect -812 -4116 -810 -4048
rect -796 -4116 -794 -4048
rect -788 -4116 -786 -4048
rect -778 -4116 -776 -4048
rect -770 -4116 -768 -4048
rect -754 -4116 -752 -4048
rect -746 -4116 -744 -4048
rect -572 -4116 -570 -4048
rect -562 -4116 -560 -4048
rect -546 -4116 -544 -4048
rect -538 -4116 -536 -4048
rect -522 -4116 -520 -4048
rect -514 -4116 -512 -4048
rect -504 -4116 -502 -4048
rect -496 -4116 -494 -4048
rect -480 -4116 -478 -4048
rect -472 -4081 -470 -4048
rect -462 -4081 -460 -4048
rect -472 -4083 -460 -4081
rect -472 -4116 -470 -4083
rect -462 -4116 -460 -4083
rect -454 -4116 -452 -4048
rect -438 -4116 -436 -4048
rect -430 -4116 -428 -4048
rect -420 -4116 -418 -4048
rect -412 -4116 -410 -4048
rect -396 -4116 -394 -4048
rect -388 -4116 -386 -4048
rect -214 -4116 -212 -4048
rect -204 -4116 -202 -4048
rect -188 -4116 -186 -4048
rect -180 -4116 -178 -4048
rect -164 -4116 -162 -4048
rect -156 -4116 -154 -4048
rect -146 -4116 -144 -4048
rect -138 -4116 -136 -4048
rect -122 -4116 -120 -4048
rect -114 -4081 -112 -4048
rect -104 -4081 -102 -4048
rect -114 -4083 -102 -4081
rect -114 -4116 -112 -4083
rect -104 -4116 -102 -4083
rect -96 -4116 -94 -4048
rect -80 -4116 -78 -4048
rect -72 -4116 -70 -4048
rect -62 -4116 -60 -4048
rect -54 -4116 -52 -4048
rect -38 -4116 -36 -4048
rect -30 -4116 -28 -4048
rect 214 -4116 216 -4048
rect 224 -4116 226 -4048
rect 240 -4116 242 -4048
rect 248 -4116 250 -4048
rect 264 -4116 266 -4048
rect 272 -4116 274 -4048
rect 282 -4116 284 -4048
rect 290 -4116 292 -4048
rect 306 -4116 308 -4048
rect 314 -4081 316 -4048
rect 324 -4081 326 -4048
rect 314 -4083 326 -4081
rect 314 -4116 316 -4083
rect 324 -4116 326 -4083
rect 332 -4116 334 -4048
rect 348 -4116 350 -4048
rect 356 -4116 358 -4048
rect 366 -4116 368 -4048
rect 374 -4116 376 -4048
rect 390 -4116 392 -4048
rect 398 -4116 400 -4048
rect 570 -4116 572 -4048
rect 580 -4116 582 -4048
rect 596 -4116 598 -4048
rect 604 -4116 606 -4048
rect 620 -4116 622 -4048
rect 628 -4116 630 -4048
rect 638 -4116 640 -4048
rect 646 -4116 648 -4048
rect 662 -4116 664 -4048
rect 670 -4081 672 -4048
rect 680 -4081 682 -4048
rect 670 -4083 682 -4081
rect 670 -4116 672 -4083
rect 680 -4116 682 -4083
rect 688 -4116 690 -4048
rect 704 -4116 706 -4048
rect 712 -4116 714 -4048
rect 722 -4116 724 -4048
rect 730 -4116 732 -4048
rect 746 -4116 748 -4048
rect 754 -4116 756 -4048
rect 968 -4116 970 -4048
rect 978 -4116 980 -4048
rect 994 -4116 996 -4048
rect 1002 -4116 1004 -4048
rect 1018 -4116 1020 -4048
rect 1026 -4116 1028 -4048
rect 1036 -4116 1038 -4048
rect 1044 -4116 1046 -4048
rect 1060 -4116 1062 -4048
rect 1068 -4081 1070 -4048
rect 1078 -4081 1080 -4048
rect 1068 -4083 1080 -4081
rect 1068 -4116 1070 -4083
rect 1078 -4116 1080 -4083
rect 1086 -4116 1088 -4048
rect 1102 -4116 1104 -4048
rect 1110 -4116 1112 -4048
rect 1120 -4116 1122 -4048
rect 1128 -4116 1130 -4048
rect 1144 -4116 1146 -4048
rect 1152 -4116 1154 -4048
rect 1326 -4116 1328 -4048
rect 1336 -4116 1338 -4048
rect 1352 -4116 1354 -4048
rect 1360 -4116 1362 -4048
rect 1376 -4116 1378 -4048
rect 1384 -4116 1386 -4048
rect 1394 -4116 1396 -4048
rect 1402 -4116 1404 -4048
rect 1418 -4116 1420 -4048
rect 1426 -4081 1428 -4048
rect 1436 -4081 1438 -4048
rect 1426 -4083 1438 -4081
rect 1426 -4116 1428 -4083
rect 1436 -4116 1438 -4083
rect 1444 -4116 1446 -4048
rect 1460 -4116 1462 -4048
rect 1468 -4116 1470 -4048
rect 1478 -4116 1480 -4048
rect 1486 -4116 1488 -4048
rect 1502 -4116 1504 -4048
rect 1510 -4116 1512 -4048
rect -1259 -4122 -1257 -4120
rect -1249 -4122 -1247 -4120
rect -1233 -4122 -1231 -4120
rect -1225 -4122 -1223 -4120
rect -1209 -4122 -1207 -4120
rect -1201 -4122 -1199 -4120
rect -1191 -4122 -1189 -4120
rect -1183 -4122 -1181 -4120
rect -1167 -4122 -1165 -4120
rect -1159 -4122 -1157 -4120
rect -1149 -4122 -1147 -4120
rect -1141 -4122 -1139 -4120
rect -1125 -4122 -1123 -4120
rect -1117 -4122 -1115 -4120
rect -1107 -4122 -1105 -4120
rect -1099 -4122 -1097 -4120
rect -1083 -4122 -1081 -4120
rect -1075 -4122 -1073 -4120
rect -930 -4122 -928 -4120
rect -920 -4122 -918 -4120
rect -904 -4122 -902 -4120
rect -896 -4122 -894 -4120
rect -880 -4122 -878 -4120
rect -872 -4122 -870 -4120
rect -862 -4122 -860 -4120
rect -854 -4122 -852 -4120
rect -838 -4122 -836 -4120
rect -830 -4122 -828 -4120
rect -820 -4122 -818 -4120
rect -812 -4122 -810 -4120
rect -796 -4122 -794 -4120
rect -788 -4122 -786 -4120
rect -778 -4122 -776 -4120
rect -770 -4122 -768 -4120
rect -754 -4122 -752 -4120
rect -746 -4122 -744 -4120
rect -572 -4122 -570 -4120
rect -562 -4122 -560 -4120
rect -546 -4122 -544 -4120
rect -538 -4122 -536 -4120
rect -522 -4122 -520 -4120
rect -514 -4122 -512 -4120
rect -504 -4122 -502 -4120
rect -496 -4122 -494 -4120
rect -480 -4122 -478 -4120
rect -472 -4122 -470 -4120
rect -462 -4122 -460 -4120
rect -454 -4122 -452 -4120
rect -438 -4122 -436 -4120
rect -430 -4122 -428 -4120
rect -420 -4122 -418 -4120
rect -412 -4122 -410 -4120
rect -396 -4122 -394 -4120
rect -388 -4122 -386 -4120
rect -214 -4122 -212 -4120
rect -204 -4122 -202 -4120
rect -188 -4122 -186 -4120
rect -180 -4122 -178 -4120
rect -164 -4122 -162 -4120
rect -156 -4122 -154 -4120
rect -146 -4122 -144 -4120
rect -138 -4122 -136 -4120
rect -122 -4122 -120 -4120
rect -114 -4122 -112 -4120
rect -104 -4122 -102 -4120
rect -96 -4122 -94 -4120
rect -80 -4122 -78 -4120
rect -72 -4122 -70 -4120
rect -62 -4122 -60 -4120
rect -54 -4122 -52 -4120
rect -38 -4122 -36 -4120
rect -30 -4122 -28 -4120
rect 214 -4122 216 -4120
rect 224 -4122 226 -4120
rect 240 -4122 242 -4120
rect 248 -4122 250 -4120
rect 264 -4122 266 -4120
rect 272 -4122 274 -4120
rect 282 -4122 284 -4120
rect 290 -4122 292 -4120
rect 306 -4122 308 -4120
rect 314 -4122 316 -4120
rect 324 -4122 326 -4120
rect 332 -4122 334 -4120
rect 348 -4122 350 -4120
rect 356 -4122 358 -4120
rect 366 -4122 368 -4120
rect 374 -4122 376 -4120
rect 390 -4122 392 -4120
rect 398 -4122 400 -4120
rect 570 -4122 572 -4120
rect 580 -4122 582 -4120
rect 596 -4122 598 -4120
rect 604 -4122 606 -4120
rect 620 -4122 622 -4120
rect 628 -4122 630 -4120
rect 638 -4122 640 -4120
rect 646 -4122 648 -4120
rect 662 -4122 664 -4120
rect 670 -4122 672 -4120
rect 680 -4122 682 -4120
rect 688 -4122 690 -4120
rect 704 -4122 706 -4120
rect 712 -4122 714 -4120
rect 722 -4122 724 -4120
rect 730 -4122 732 -4120
rect 746 -4122 748 -4120
rect 754 -4122 756 -4120
rect 968 -4122 970 -4120
rect 978 -4122 980 -4120
rect 994 -4122 996 -4120
rect 1002 -4122 1004 -4120
rect 1018 -4122 1020 -4120
rect 1026 -4122 1028 -4120
rect 1036 -4122 1038 -4120
rect 1044 -4122 1046 -4120
rect 1060 -4122 1062 -4120
rect 1068 -4122 1070 -4120
rect 1078 -4122 1080 -4120
rect 1086 -4122 1088 -4120
rect 1102 -4122 1104 -4120
rect 1110 -4122 1112 -4120
rect 1120 -4122 1122 -4120
rect 1128 -4122 1130 -4120
rect 1144 -4122 1146 -4120
rect 1152 -4122 1154 -4120
rect 1326 -4122 1328 -4120
rect 1336 -4122 1338 -4120
rect 1352 -4122 1354 -4120
rect 1360 -4122 1362 -4120
rect 1376 -4122 1378 -4120
rect 1384 -4122 1386 -4120
rect 1394 -4122 1396 -4120
rect 1402 -4122 1404 -4120
rect 1418 -4122 1420 -4120
rect 1426 -4122 1428 -4120
rect 1436 -4122 1438 -4120
rect 1444 -4122 1446 -4120
rect 1460 -4122 1462 -4120
rect 1468 -4122 1470 -4120
rect 1478 -4122 1480 -4120
rect 1486 -4122 1488 -4120
rect 1502 -4122 1504 -4120
rect 1510 -4122 1512 -4120
rect -1259 -4164 -1257 -4162
rect -1249 -4164 -1247 -4162
rect -1233 -4164 -1231 -4162
rect -1225 -4164 -1223 -4162
rect -1209 -4164 -1207 -4162
rect -1201 -4164 -1199 -4162
rect -1191 -4164 -1189 -4162
rect -1183 -4164 -1181 -4162
rect -1167 -4164 -1165 -4162
rect -1159 -4164 -1157 -4162
rect -1149 -4164 -1147 -4162
rect -1141 -4164 -1139 -4162
rect -1125 -4164 -1123 -4162
rect -1117 -4164 -1115 -4162
rect -1107 -4164 -1105 -4162
rect -1099 -4164 -1097 -4162
rect -1083 -4164 -1081 -4162
rect -1075 -4164 -1073 -4162
rect -1024 -4164 -1022 -4162
rect -930 -4164 -928 -4162
rect -920 -4164 -918 -4162
rect -904 -4164 -902 -4162
rect -896 -4164 -894 -4162
rect -880 -4164 -878 -4162
rect -872 -4164 -870 -4162
rect -862 -4164 -860 -4162
rect -854 -4164 -852 -4162
rect -838 -4164 -836 -4162
rect -830 -4164 -828 -4162
rect -820 -4164 -818 -4162
rect -812 -4164 -810 -4162
rect -796 -4164 -794 -4162
rect -788 -4164 -786 -4162
rect -778 -4164 -776 -4162
rect -770 -4164 -768 -4162
rect -754 -4164 -752 -4162
rect -746 -4164 -744 -4162
rect -572 -4164 -570 -4162
rect -562 -4164 -560 -4162
rect -546 -4164 -544 -4162
rect -538 -4164 -536 -4162
rect -522 -4164 -520 -4162
rect -514 -4164 -512 -4162
rect -504 -4164 -502 -4162
rect -496 -4164 -494 -4162
rect -480 -4164 -478 -4162
rect -472 -4164 -470 -4162
rect -462 -4164 -460 -4162
rect -454 -4164 -452 -4162
rect -438 -4164 -436 -4162
rect -430 -4164 -428 -4162
rect -420 -4164 -418 -4162
rect -412 -4164 -410 -4162
rect -396 -4164 -394 -4162
rect -388 -4164 -386 -4162
rect -327 -4164 -325 -4162
rect -214 -4164 -212 -4162
rect -204 -4164 -202 -4162
rect -188 -4164 -186 -4162
rect -180 -4164 -178 -4162
rect -164 -4164 -162 -4162
rect -156 -4164 -154 -4162
rect -146 -4164 -144 -4162
rect -138 -4164 -136 -4162
rect -122 -4164 -120 -4162
rect -114 -4164 -112 -4162
rect -104 -4164 -102 -4162
rect -96 -4164 -94 -4162
rect -80 -4164 -78 -4162
rect -72 -4164 -70 -4162
rect -62 -4164 -60 -4162
rect -54 -4164 -52 -4162
rect -38 -4164 -36 -4162
rect -30 -4164 -28 -4162
rect 461 -4164 463 -4162
rect 1206 -4164 1208 -4162
rect -1259 -4240 -1257 -4172
rect -1249 -4240 -1247 -4172
rect -1233 -4240 -1231 -4172
rect -1225 -4240 -1223 -4172
rect -1209 -4240 -1207 -4172
rect -1201 -4240 -1199 -4172
rect -1191 -4240 -1189 -4172
rect -1183 -4240 -1181 -4172
rect -1167 -4240 -1165 -4172
rect -1159 -4205 -1157 -4172
rect -1149 -4205 -1147 -4172
rect -1159 -4207 -1147 -4205
rect -1159 -4240 -1157 -4207
rect -1149 -4240 -1147 -4207
rect -1141 -4240 -1139 -4172
rect -1125 -4240 -1123 -4172
rect -1117 -4240 -1115 -4172
rect -1107 -4240 -1105 -4172
rect -1099 -4240 -1097 -4172
rect -1083 -4240 -1081 -4172
rect -1075 -4240 -1073 -4172
rect -1024 -4240 -1022 -4172
rect -930 -4240 -928 -4172
rect -920 -4240 -918 -4172
rect -904 -4240 -902 -4172
rect -896 -4240 -894 -4172
rect -880 -4240 -878 -4172
rect -872 -4240 -870 -4172
rect -862 -4240 -860 -4172
rect -854 -4240 -852 -4172
rect -838 -4240 -836 -4172
rect -830 -4205 -828 -4172
rect -820 -4205 -818 -4172
rect -830 -4207 -818 -4205
rect -830 -4240 -828 -4207
rect -820 -4240 -818 -4207
rect -812 -4240 -810 -4172
rect -796 -4240 -794 -4172
rect -788 -4240 -786 -4172
rect -778 -4240 -776 -4172
rect -770 -4240 -768 -4172
rect -754 -4240 -752 -4172
rect -746 -4240 -744 -4172
rect -572 -4240 -570 -4172
rect -562 -4240 -560 -4172
rect -546 -4240 -544 -4172
rect -538 -4240 -536 -4172
rect -522 -4240 -520 -4172
rect -514 -4240 -512 -4172
rect -504 -4240 -502 -4172
rect -496 -4240 -494 -4172
rect -480 -4240 -478 -4172
rect -472 -4205 -470 -4172
rect -462 -4205 -460 -4172
rect -472 -4207 -460 -4205
rect -472 -4240 -470 -4207
rect -462 -4240 -460 -4207
rect -454 -4240 -452 -4172
rect -438 -4240 -436 -4172
rect -430 -4240 -428 -4172
rect -420 -4240 -418 -4172
rect -412 -4240 -410 -4172
rect -396 -4240 -394 -4172
rect -388 -4240 -386 -4172
rect -327 -4240 -325 -4172
rect -214 -4240 -212 -4172
rect -204 -4240 -202 -4172
rect -188 -4240 -186 -4172
rect -180 -4240 -178 -4172
rect -164 -4240 -162 -4172
rect -156 -4240 -154 -4172
rect -146 -4240 -144 -4172
rect -138 -4240 -136 -4172
rect -122 -4240 -120 -4172
rect -114 -4205 -112 -4172
rect -104 -4205 -102 -4172
rect -114 -4207 -102 -4205
rect -114 -4240 -112 -4207
rect -104 -4240 -102 -4207
rect -96 -4240 -94 -4172
rect -80 -4240 -78 -4172
rect -72 -4240 -70 -4172
rect -62 -4240 -60 -4172
rect -54 -4240 -52 -4172
rect -38 -4240 -36 -4172
rect -30 -4240 -28 -4172
rect 461 -4240 463 -4172
rect 1206 -4240 1208 -4172
rect -1259 -4246 -1257 -4244
rect -1249 -4246 -1247 -4244
rect -1233 -4246 -1231 -4244
rect -1225 -4246 -1223 -4244
rect -1209 -4246 -1207 -4244
rect -1201 -4246 -1199 -4244
rect -1191 -4246 -1189 -4244
rect -1183 -4246 -1181 -4244
rect -1167 -4246 -1165 -4244
rect -1159 -4246 -1157 -4244
rect -1149 -4246 -1147 -4244
rect -1141 -4246 -1139 -4244
rect -1125 -4246 -1123 -4244
rect -1117 -4246 -1115 -4244
rect -1107 -4246 -1105 -4244
rect -1099 -4246 -1097 -4244
rect -1083 -4246 -1081 -4244
rect -1075 -4246 -1073 -4244
rect -1024 -4246 -1022 -4244
rect -930 -4246 -928 -4244
rect -920 -4246 -918 -4244
rect -904 -4246 -902 -4244
rect -896 -4246 -894 -4244
rect -880 -4246 -878 -4244
rect -872 -4246 -870 -4244
rect -862 -4246 -860 -4244
rect -854 -4246 -852 -4244
rect -838 -4246 -836 -4244
rect -830 -4246 -828 -4244
rect -820 -4246 -818 -4244
rect -812 -4246 -810 -4244
rect -796 -4246 -794 -4244
rect -788 -4246 -786 -4244
rect -778 -4246 -776 -4244
rect -770 -4246 -768 -4244
rect -754 -4246 -752 -4244
rect -746 -4246 -744 -4244
rect -572 -4246 -570 -4244
rect -562 -4246 -560 -4244
rect -546 -4246 -544 -4244
rect -538 -4246 -536 -4244
rect -522 -4246 -520 -4244
rect -514 -4246 -512 -4244
rect -504 -4246 -502 -4244
rect -496 -4246 -494 -4244
rect -480 -4246 -478 -4244
rect -472 -4246 -470 -4244
rect -462 -4246 -460 -4244
rect -454 -4246 -452 -4244
rect -438 -4246 -436 -4244
rect -430 -4246 -428 -4244
rect -420 -4246 -418 -4244
rect -412 -4246 -410 -4244
rect -396 -4246 -394 -4244
rect -388 -4246 -386 -4244
rect -327 -4246 -325 -4244
rect -214 -4246 -212 -4244
rect -204 -4246 -202 -4244
rect -188 -4246 -186 -4244
rect -180 -4246 -178 -4244
rect -164 -4246 -162 -4244
rect -156 -4246 -154 -4244
rect -146 -4246 -144 -4244
rect -138 -4246 -136 -4244
rect -122 -4246 -120 -4244
rect -114 -4246 -112 -4244
rect -104 -4246 -102 -4244
rect -96 -4246 -94 -4244
rect -80 -4246 -78 -4244
rect -72 -4246 -70 -4244
rect -62 -4246 -60 -4244
rect -54 -4246 -52 -4244
rect -38 -4246 -36 -4244
rect -30 -4246 -28 -4244
rect 461 -4246 463 -4244
rect 1206 -4246 1208 -4244
rect -1334 -4275 -1332 -4273
rect -1326 -4275 -1324 -4273
rect -1316 -4275 -1314 -4273
rect -1024 -4275 -1022 -4273
rect -930 -4275 -928 -4273
rect -922 -4275 -920 -4273
rect -912 -4275 -910 -4273
rect -668 -4275 -666 -4273
rect -572 -4275 -570 -4273
rect -564 -4275 -562 -4273
rect -554 -4275 -552 -4273
rect -327 -4275 -325 -4273
rect -214 -4275 -212 -4273
rect -206 -4275 -204 -4273
rect -196 -4275 -194 -4273
rect 214 -4275 216 -4273
rect 222 -4275 224 -4273
rect 232 -4275 234 -4273
rect 461 -4275 463 -4273
rect 570 -4275 572 -4273
rect 578 -4275 580 -4273
rect 588 -4275 590 -4273
rect 865 -4275 867 -4273
rect 968 -4275 970 -4273
rect 976 -4275 978 -4273
rect 986 -4275 988 -4273
rect 1206 -4275 1208 -4273
rect 1326 -4275 1328 -4273
rect 1334 -4275 1336 -4273
rect 1344 -4275 1346 -4273
rect -1334 -4351 -1332 -4283
rect -1326 -4307 -1324 -4283
rect -1326 -4351 -1324 -4311
rect -1316 -4351 -1314 -4283
rect -1024 -4351 -1022 -4283
rect -930 -4351 -928 -4283
rect -922 -4307 -920 -4283
rect -922 -4351 -920 -4311
rect -912 -4351 -910 -4283
rect -668 -4347 -666 -4291
rect -572 -4351 -570 -4283
rect -564 -4307 -562 -4283
rect -564 -4351 -562 -4311
rect -554 -4351 -552 -4283
rect -327 -4351 -325 -4283
rect -214 -4351 -212 -4283
rect -206 -4307 -204 -4283
rect -206 -4351 -204 -4311
rect -196 -4351 -194 -4283
rect 214 -4351 216 -4283
rect 222 -4307 224 -4283
rect 222 -4351 224 -4311
rect 232 -4351 234 -4283
rect 461 -4351 463 -4283
rect 570 -4351 572 -4283
rect 578 -4307 580 -4283
rect 578 -4351 580 -4311
rect 588 -4351 590 -4283
rect 865 -4347 867 -4291
rect 968 -4351 970 -4283
rect 976 -4307 978 -4283
rect 976 -4351 978 -4311
rect 986 -4351 988 -4283
rect 1206 -4351 1208 -4283
rect 1326 -4351 1328 -4283
rect 1334 -4307 1336 -4283
rect 1334 -4351 1336 -4311
rect 1344 -4351 1346 -4283
rect -1334 -4357 -1332 -4355
rect -1326 -4357 -1324 -4355
rect -1316 -4357 -1314 -4355
rect -1024 -4357 -1022 -4355
rect -930 -4357 -928 -4355
rect -922 -4357 -920 -4355
rect -912 -4357 -910 -4355
rect -668 -4357 -666 -4355
rect -572 -4357 -570 -4355
rect -564 -4357 -562 -4355
rect -554 -4357 -552 -4355
rect -327 -4357 -325 -4355
rect -214 -4357 -212 -4355
rect -206 -4357 -204 -4355
rect -196 -4357 -194 -4355
rect 214 -4357 216 -4355
rect 222 -4357 224 -4355
rect 232 -4357 234 -4355
rect 461 -4357 463 -4355
rect 570 -4357 572 -4355
rect 578 -4357 580 -4355
rect 588 -4357 590 -4355
rect 865 -4357 867 -4355
rect 968 -4357 970 -4355
rect 976 -4357 978 -4355
rect 986 -4357 988 -4355
rect 1206 -4357 1208 -4355
rect 1326 -4357 1328 -4355
rect 1334 -4357 1336 -4355
rect 1344 -4357 1346 -4355
rect -1259 -4394 -1257 -4392
rect -1249 -4394 -1247 -4392
rect -1233 -4394 -1231 -4392
rect -1223 -4394 -1221 -4392
rect -1215 -4394 -1213 -4392
rect -1205 -4394 -1203 -4392
rect -1189 -4394 -1187 -4392
rect -1181 -4394 -1179 -4392
rect -1171 -4394 -1169 -4392
rect -930 -4394 -928 -4392
rect -920 -4394 -918 -4392
rect -904 -4394 -902 -4392
rect -894 -4394 -892 -4392
rect -878 -4394 -876 -4392
rect -868 -4394 -866 -4392
rect -860 -4394 -858 -4392
rect -850 -4394 -848 -4392
rect -834 -4394 -832 -4392
rect -826 -4394 -824 -4392
rect -816 -4394 -814 -4392
rect -800 -4394 -798 -4392
rect -790 -4394 -788 -4392
rect -782 -4394 -780 -4392
rect -772 -4394 -770 -4392
rect -756 -4394 -754 -4392
rect -748 -4394 -746 -4392
rect -732 -4394 -730 -4392
rect -716 -4394 -714 -4392
rect -708 -4394 -706 -4392
rect -698 -4394 -696 -4392
rect -572 -4394 -570 -4392
rect -562 -4394 -560 -4392
rect -546 -4394 -544 -4392
rect -536 -4394 -534 -4392
rect -520 -4394 -518 -4392
rect -510 -4394 -508 -4392
rect -502 -4394 -500 -4392
rect -492 -4394 -490 -4392
rect -476 -4394 -474 -4392
rect -468 -4394 -466 -4392
rect -458 -4394 -456 -4392
rect -442 -4394 -440 -4392
rect -432 -4394 -430 -4392
rect -424 -4394 -422 -4392
rect -414 -4394 -412 -4392
rect -398 -4394 -396 -4392
rect -390 -4394 -388 -4392
rect -374 -4394 -372 -4392
rect -358 -4394 -356 -4392
rect -350 -4394 -348 -4392
rect -340 -4394 -338 -4392
rect -214 -4394 -212 -4392
rect -204 -4394 -202 -4392
rect -188 -4394 -186 -4392
rect -178 -4394 -176 -4392
rect -162 -4394 -160 -4392
rect -152 -4394 -150 -4392
rect -144 -4394 -142 -4392
rect -134 -4394 -132 -4392
rect -118 -4394 -116 -4392
rect -110 -4394 -108 -4392
rect -100 -4394 -98 -4392
rect -84 -4394 -82 -4392
rect -74 -4394 -72 -4392
rect -66 -4394 -64 -4392
rect -56 -4394 -54 -4392
rect -40 -4394 -38 -4392
rect -32 -4394 -30 -4392
rect -16 -4394 -14 -4392
rect 0 -4394 2 -4392
rect 8 -4394 10 -4392
rect 18 -4394 20 -4392
rect 214 -4394 216 -4392
rect 224 -4394 226 -4392
rect 240 -4394 242 -4392
rect 250 -4394 252 -4392
rect 266 -4394 268 -4392
rect 276 -4394 278 -4392
rect 284 -4394 286 -4392
rect 294 -4394 296 -4392
rect 310 -4394 312 -4392
rect 318 -4394 320 -4392
rect 328 -4394 330 -4392
rect 344 -4394 346 -4392
rect 354 -4394 356 -4392
rect 362 -4394 364 -4392
rect 372 -4394 374 -4392
rect 388 -4394 390 -4392
rect 396 -4394 398 -4392
rect 412 -4394 414 -4392
rect 428 -4394 430 -4392
rect 436 -4394 438 -4392
rect 446 -4394 448 -4392
rect 570 -4394 572 -4392
rect 580 -4394 582 -4392
rect 596 -4394 598 -4392
rect 606 -4394 608 -4392
rect 622 -4394 624 -4392
rect 632 -4394 634 -4392
rect 640 -4394 642 -4392
rect 650 -4394 652 -4392
rect 666 -4394 668 -4392
rect 674 -4394 676 -4392
rect 684 -4394 686 -4392
rect 700 -4394 702 -4392
rect 710 -4394 712 -4392
rect 718 -4394 720 -4392
rect 728 -4394 730 -4392
rect 744 -4394 746 -4392
rect 752 -4394 754 -4392
rect 768 -4394 770 -4392
rect 784 -4394 786 -4392
rect 792 -4394 794 -4392
rect 802 -4394 804 -4392
rect 968 -4394 970 -4392
rect 978 -4394 980 -4392
rect 994 -4394 996 -4392
rect 1004 -4394 1006 -4392
rect 1020 -4394 1022 -4392
rect 1030 -4394 1032 -4392
rect 1038 -4394 1040 -4392
rect 1048 -4394 1050 -4392
rect 1064 -4394 1066 -4392
rect 1072 -4394 1074 -4392
rect 1082 -4394 1084 -4392
rect 1098 -4394 1100 -4392
rect 1108 -4394 1110 -4392
rect 1116 -4394 1118 -4392
rect 1126 -4394 1128 -4392
rect 1142 -4394 1144 -4392
rect 1150 -4394 1152 -4392
rect 1166 -4394 1168 -4392
rect 1182 -4394 1184 -4392
rect 1190 -4394 1192 -4392
rect 1200 -4394 1202 -4392
rect 1326 -4394 1328 -4392
rect 1336 -4394 1338 -4392
rect 1352 -4394 1354 -4392
rect 1362 -4394 1364 -4392
rect 1378 -4394 1380 -4392
rect 1388 -4394 1390 -4392
rect 1396 -4394 1398 -4392
rect 1406 -4394 1408 -4392
rect 1422 -4394 1424 -4392
rect 1430 -4394 1432 -4392
rect 1440 -4394 1442 -4392
rect 1456 -4394 1458 -4392
rect 1466 -4394 1468 -4392
rect 1474 -4394 1476 -4392
rect 1484 -4394 1486 -4392
rect 1500 -4394 1502 -4392
rect 1508 -4394 1510 -4392
rect 1524 -4394 1526 -4392
rect 1540 -4394 1542 -4392
rect 1548 -4394 1550 -4392
rect 1558 -4394 1560 -4392
rect -1259 -4470 -1257 -4402
rect -1249 -4470 -1247 -4402
rect -1233 -4470 -1231 -4402
rect -1223 -4470 -1221 -4402
rect -1215 -4470 -1213 -4402
rect -1205 -4470 -1203 -4402
rect -1189 -4470 -1187 -4402
rect -1181 -4470 -1179 -4402
rect -1171 -4470 -1169 -4402
rect -930 -4470 -928 -4402
rect -920 -4470 -918 -4402
rect -904 -4470 -902 -4402
rect -894 -4470 -892 -4402
rect -878 -4470 -876 -4402
rect -868 -4470 -866 -4402
rect -860 -4470 -858 -4402
rect -850 -4470 -848 -4402
rect -834 -4470 -832 -4402
rect -826 -4470 -824 -4402
rect -816 -4470 -814 -4402
rect -800 -4470 -798 -4402
rect -790 -4470 -788 -4402
rect -782 -4470 -780 -4402
rect -772 -4470 -770 -4402
rect -756 -4470 -754 -4402
rect -748 -4470 -746 -4402
rect -732 -4470 -730 -4402
rect -716 -4470 -714 -4402
rect -708 -4470 -706 -4402
rect -698 -4470 -696 -4402
rect -572 -4470 -570 -4402
rect -562 -4470 -560 -4402
rect -546 -4470 -544 -4402
rect -536 -4470 -534 -4402
rect -520 -4470 -518 -4402
rect -510 -4470 -508 -4402
rect -502 -4470 -500 -4402
rect -492 -4470 -490 -4402
rect -476 -4470 -474 -4402
rect -468 -4470 -466 -4402
rect -458 -4470 -456 -4402
rect -442 -4470 -440 -4402
rect -432 -4470 -430 -4402
rect -424 -4470 -422 -4402
rect -414 -4470 -412 -4402
rect -398 -4470 -396 -4402
rect -390 -4470 -388 -4402
rect -374 -4470 -372 -4402
rect -358 -4470 -356 -4402
rect -350 -4470 -348 -4402
rect -340 -4470 -338 -4402
rect -214 -4470 -212 -4402
rect -204 -4470 -202 -4402
rect -188 -4470 -186 -4402
rect -178 -4470 -176 -4402
rect -162 -4470 -160 -4402
rect -152 -4470 -150 -4402
rect -144 -4470 -142 -4402
rect -134 -4470 -132 -4402
rect -118 -4470 -116 -4402
rect -110 -4470 -108 -4402
rect -100 -4470 -98 -4402
rect -84 -4470 -82 -4402
rect -74 -4470 -72 -4402
rect -66 -4470 -64 -4402
rect -56 -4470 -54 -4402
rect -40 -4470 -38 -4402
rect -32 -4470 -30 -4402
rect -16 -4470 -14 -4402
rect 0 -4470 2 -4402
rect 8 -4470 10 -4402
rect 18 -4470 20 -4402
rect 214 -4470 216 -4402
rect 224 -4470 226 -4402
rect 240 -4470 242 -4402
rect 250 -4470 252 -4402
rect 266 -4470 268 -4402
rect 276 -4470 278 -4402
rect 284 -4470 286 -4402
rect 294 -4470 296 -4402
rect 310 -4470 312 -4402
rect 318 -4470 320 -4402
rect 328 -4470 330 -4402
rect 344 -4470 346 -4402
rect 354 -4470 356 -4402
rect 362 -4470 364 -4402
rect 372 -4470 374 -4402
rect 388 -4470 390 -4402
rect 396 -4470 398 -4402
rect 412 -4470 414 -4402
rect 428 -4470 430 -4402
rect 436 -4470 438 -4402
rect 446 -4470 448 -4402
rect 570 -4470 572 -4402
rect 580 -4470 582 -4402
rect 596 -4470 598 -4402
rect 606 -4470 608 -4402
rect 622 -4470 624 -4402
rect 632 -4470 634 -4402
rect 640 -4470 642 -4402
rect 650 -4470 652 -4402
rect 666 -4470 668 -4402
rect 674 -4470 676 -4402
rect 684 -4470 686 -4402
rect 700 -4470 702 -4402
rect 710 -4470 712 -4402
rect 718 -4470 720 -4402
rect 728 -4470 730 -4402
rect 744 -4470 746 -4402
rect 752 -4470 754 -4402
rect 768 -4470 770 -4402
rect 784 -4470 786 -4402
rect 792 -4470 794 -4402
rect 802 -4470 804 -4402
rect 968 -4470 970 -4402
rect 978 -4470 980 -4402
rect 994 -4470 996 -4402
rect 1004 -4470 1006 -4402
rect 1020 -4470 1022 -4402
rect 1030 -4470 1032 -4402
rect 1038 -4470 1040 -4402
rect 1048 -4470 1050 -4402
rect 1064 -4470 1066 -4402
rect 1072 -4470 1074 -4402
rect 1082 -4470 1084 -4402
rect 1098 -4470 1100 -4402
rect 1108 -4470 1110 -4402
rect 1116 -4470 1118 -4402
rect 1126 -4470 1128 -4402
rect 1142 -4470 1144 -4402
rect 1150 -4470 1152 -4402
rect 1166 -4470 1168 -4402
rect 1182 -4470 1184 -4402
rect 1190 -4470 1192 -4402
rect 1200 -4470 1202 -4402
rect 1326 -4470 1328 -4402
rect 1336 -4470 1338 -4402
rect 1352 -4470 1354 -4402
rect 1362 -4470 1364 -4402
rect 1378 -4470 1380 -4402
rect 1388 -4470 1390 -4402
rect 1396 -4470 1398 -4402
rect 1406 -4470 1408 -4402
rect 1422 -4470 1424 -4402
rect 1430 -4470 1432 -4402
rect 1440 -4470 1442 -4402
rect 1456 -4470 1458 -4402
rect 1466 -4470 1468 -4402
rect 1474 -4470 1476 -4402
rect 1484 -4470 1486 -4402
rect 1500 -4470 1502 -4402
rect 1508 -4470 1510 -4402
rect 1524 -4470 1526 -4402
rect 1540 -4470 1542 -4402
rect 1548 -4470 1550 -4402
rect 1558 -4470 1560 -4402
rect -1259 -4476 -1257 -4474
rect -1249 -4476 -1247 -4474
rect -1233 -4476 -1231 -4474
rect -1223 -4476 -1221 -4474
rect -1215 -4476 -1213 -4474
rect -1205 -4476 -1203 -4474
rect -1189 -4476 -1187 -4474
rect -1181 -4476 -1179 -4474
rect -1171 -4476 -1169 -4474
rect -930 -4476 -928 -4474
rect -920 -4476 -918 -4474
rect -904 -4476 -902 -4474
rect -894 -4476 -892 -4474
rect -878 -4476 -876 -4474
rect -868 -4476 -866 -4474
rect -860 -4476 -858 -4474
rect -850 -4476 -848 -4474
rect -834 -4476 -832 -4474
rect -826 -4476 -824 -4474
rect -816 -4476 -814 -4474
rect -800 -4476 -798 -4474
rect -790 -4476 -788 -4474
rect -782 -4476 -780 -4474
rect -772 -4476 -770 -4474
rect -756 -4476 -754 -4474
rect -748 -4476 -746 -4474
rect -732 -4476 -730 -4474
rect -716 -4476 -714 -4474
rect -708 -4476 -706 -4474
rect -698 -4476 -696 -4474
rect -572 -4476 -570 -4474
rect -562 -4476 -560 -4474
rect -546 -4476 -544 -4474
rect -536 -4476 -534 -4474
rect -520 -4476 -518 -4474
rect -510 -4476 -508 -4474
rect -502 -4476 -500 -4474
rect -492 -4476 -490 -4474
rect -476 -4476 -474 -4474
rect -468 -4476 -466 -4474
rect -458 -4476 -456 -4474
rect -442 -4476 -440 -4474
rect -432 -4476 -430 -4474
rect -424 -4476 -422 -4474
rect -414 -4476 -412 -4474
rect -398 -4476 -396 -4474
rect -390 -4476 -388 -4474
rect -374 -4476 -372 -4474
rect -358 -4476 -356 -4474
rect -350 -4476 -348 -4474
rect -340 -4476 -338 -4474
rect -214 -4476 -212 -4474
rect -204 -4476 -202 -4474
rect -188 -4476 -186 -4474
rect -178 -4476 -176 -4474
rect -162 -4476 -160 -4474
rect -152 -4476 -150 -4474
rect -144 -4476 -142 -4474
rect -134 -4476 -132 -4474
rect -118 -4476 -116 -4474
rect -110 -4476 -108 -4474
rect -100 -4476 -98 -4474
rect -84 -4476 -82 -4474
rect -74 -4476 -72 -4474
rect -66 -4476 -64 -4474
rect -56 -4476 -54 -4474
rect -40 -4476 -38 -4474
rect -32 -4476 -30 -4474
rect -16 -4476 -14 -4474
rect 0 -4476 2 -4474
rect 8 -4476 10 -4474
rect 18 -4476 20 -4474
rect 214 -4476 216 -4474
rect 224 -4476 226 -4474
rect 240 -4476 242 -4474
rect 250 -4476 252 -4474
rect 266 -4476 268 -4474
rect 276 -4476 278 -4474
rect 284 -4476 286 -4474
rect 294 -4476 296 -4474
rect 310 -4476 312 -4474
rect 318 -4476 320 -4474
rect 328 -4476 330 -4474
rect 344 -4476 346 -4474
rect 354 -4476 356 -4474
rect 362 -4476 364 -4474
rect 372 -4476 374 -4474
rect 388 -4476 390 -4474
rect 396 -4476 398 -4474
rect 412 -4476 414 -4474
rect 428 -4476 430 -4474
rect 436 -4476 438 -4474
rect 446 -4476 448 -4474
rect 570 -4476 572 -4474
rect 580 -4476 582 -4474
rect 596 -4476 598 -4474
rect 606 -4476 608 -4474
rect 622 -4476 624 -4474
rect 632 -4476 634 -4474
rect 640 -4476 642 -4474
rect 650 -4476 652 -4474
rect 666 -4476 668 -4474
rect 674 -4476 676 -4474
rect 684 -4476 686 -4474
rect 700 -4476 702 -4474
rect 710 -4476 712 -4474
rect 718 -4476 720 -4474
rect 728 -4476 730 -4474
rect 744 -4476 746 -4474
rect 752 -4476 754 -4474
rect 768 -4476 770 -4474
rect 784 -4476 786 -4474
rect 792 -4476 794 -4474
rect 802 -4476 804 -4474
rect 968 -4476 970 -4474
rect 978 -4476 980 -4474
rect 994 -4476 996 -4474
rect 1004 -4476 1006 -4474
rect 1020 -4476 1022 -4474
rect 1030 -4476 1032 -4474
rect 1038 -4476 1040 -4474
rect 1048 -4476 1050 -4474
rect 1064 -4476 1066 -4474
rect 1072 -4476 1074 -4474
rect 1082 -4476 1084 -4474
rect 1098 -4476 1100 -4474
rect 1108 -4476 1110 -4474
rect 1116 -4476 1118 -4474
rect 1126 -4476 1128 -4474
rect 1142 -4476 1144 -4474
rect 1150 -4476 1152 -4474
rect 1166 -4476 1168 -4474
rect 1182 -4476 1184 -4474
rect 1190 -4476 1192 -4474
rect 1200 -4476 1202 -4474
rect 1326 -4476 1328 -4474
rect 1336 -4476 1338 -4474
rect 1352 -4476 1354 -4474
rect 1362 -4476 1364 -4474
rect 1378 -4476 1380 -4474
rect 1388 -4476 1390 -4474
rect 1396 -4476 1398 -4474
rect 1406 -4476 1408 -4474
rect 1422 -4476 1424 -4474
rect 1430 -4476 1432 -4474
rect 1440 -4476 1442 -4474
rect 1456 -4476 1458 -4474
rect 1466 -4476 1468 -4474
rect 1474 -4476 1476 -4474
rect 1484 -4476 1486 -4474
rect 1500 -4476 1502 -4474
rect 1508 -4476 1510 -4474
rect 1524 -4476 1526 -4474
rect 1540 -4476 1542 -4474
rect 1548 -4476 1550 -4474
rect 1558 -4476 1560 -4474
rect -1259 -4517 -1257 -4515
rect -1249 -4517 -1247 -4515
rect -1233 -4517 -1231 -4515
rect -1225 -4517 -1223 -4515
rect -1209 -4517 -1207 -4515
rect -1201 -4517 -1199 -4515
rect -1191 -4517 -1189 -4515
rect -1183 -4517 -1181 -4515
rect -1167 -4517 -1165 -4515
rect -1159 -4517 -1157 -4515
rect -1149 -4517 -1147 -4515
rect -1141 -4517 -1139 -4515
rect -1125 -4517 -1123 -4515
rect -1117 -4517 -1115 -4515
rect -1107 -4517 -1105 -4515
rect -1099 -4517 -1097 -4515
rect -1083 -4517 -1081 -4515
rect -1075 -4517 -1073 -4515
rect -930 -4517 -928 -4515
rect -920 -4517 -918 -4515
rect -904 -4517 -902 -4515
rect -896 -4517 -894 -4515
rect -880 -4517 -878 -4515
rect -872 -4517 -870 -4515
rect -862 -4517 -860 -4515
rect -854 -4517 -852 -4515
rect -838 -4517 -836 -4515
rect -830 -4517 -828 -4515
rect -820 -4517 -818 -4515
rect -812 -4517 -810 -4515
rect -796 -4517 -794 -4515
rect -788 -4517 -786 -4515
rect -778 -4517 -776 -4515
rect -770 -4517 -768 -4515
rect -754 -4517 -752 -4515
rect -746 -4517 -744 -4515
rect -572 -4517 -570 -4515
rect -562 -4517 -560 -4515
rect -546 -4517 -544 -4515
rect -538 -4517 -536 -4515
rect -522 -4517 -520 -4515
rect -514 -4517 -512 -4515
rect -504 -4517 -502 -4515
rect -496 -4517 -494 -4515
rect -480 -4517 -478 -4515
rect -472 -4517 -470 -4515
rect -462 -4517 -460 -4515
rect -454 -4517 -452 -4515
rect -438 -4517 -436 -4515
rect -430 -4517 -428 -4515
rect -420 -4517 -418 -4515
rect -412 -4517 -410 -4515
rect -396 -4517 -394 -4515
rect -388 -4517 -386 -4515
rect -1259 -4593 -1257 -4525
rect -1249 -4593 -1247 -4525
rect -1233 -4593 -1231 -4525
rect -1225 -4593 -1223 -4525
rect -1209 -4593 -1207 -4525
rect -1201 -4593 -1199 -4525
rect -1191 -4593 -1189 -4525
rect -1183 -4593 -1181 -4525
rect -1167 -4593 -1165 -4525
rect -1159 -4558 -1157 -4525
rect -1149 -4558 -1147 -4525
rect -1159 -4560 -1147 -4558
rect -1159 -4593 -1157 -4560
rect -1149 -4593 -1147 -4560
rect -1141 -4593 -1139 -4525
rect -1125 -4593 -1123 -4525
rect -1117 -4593 -1115 -4525
rect -1107 -4593 -1105 -4525
rect -1099 -4593 -1097 -4525
rect -1083 -4593 -1081 -4525
rect -1075 -4593 -1073 -4525
rect -930 -4593 -928 -4525
rect -920 -4593 -918 -4525
rect -904 -4593 -902 -4525
rect -896 -4593 -894 -4525
rect -880 -4593 -878 -4525
rect -872 -4593 -870 -4525
rect -862 -4593 -860 -4525
rect -854 -4593 -852 -4525
rect -838 -4593 -836 -4525
rect -830 -4558 -828 -4525
rect -820 -4558 -818 -4525
rect -830 -4560 -818 -4558
rect -830 -4593 -828 -4560
rect -820 -4593 -818 -4560
rect -812 -4593 -810 -4525
rect -796 -4593 -794 -4525
rect -788 -4593 -786 -4525
rect -778 -4593 -776 -4525
rect -770 -4593 -768 -4525
rect -754 -4593 -752 -4525
rect -746 -4593 -744 -4525
rect -572 -4593 -570 -4525
rect -562 -4593 -560 -4525
rect -546 -4593 -544 -4525
rect -538 -4593 -536 -4525
rect -522 -4593 -520 -4525
rect -514 -4593 -512 -4525
rect -504 -4593 -502 -4525
rect -496 -4593 -494 -4525
rect -480 -4593 -478 -4525
rect -472 -4558 -470 -4525
rect -462 -4558 -460 -4525
rect -472 -4560 -460 -4558
rect -472 -4593 -470 -4560
rect -462 -4593 -460 -4560
rect -454 -4593 -452 -4525
rect -438 -4593 -436 -4525
rect -430 -4593 -428 -4525
rect -420 -4593 -418 -4525
rect -412 -4593 -410 -4525
rect -396 -4593 -394 -4525
rect -388 -4593 -386 -4525
rect -1259 -4599 -1257 -4597
rect -1249 -4599 -1247 -4597
rect -1233 -4599 -1231 -4597
rect -1225 -4599 -1223 -4597
rect -1209 -4599 -1207 -4597
rect -1201 -4599 -1199 -4597
rect -1191 -4599 -1189 -4597
rect -1183 -4599 -1181 -4597
rect -1167 -4599 -1165 -4597
rect -1159 -4599 -1157 -4597
rect -1149 -4599 -1147 -4597
rect -1141 -4599 -1139 -4597
rect -1125 -4599 -1123 -4597
rect -1117 -4599 -1115 -4597
rect -1107 -4599 -1105 -4597
rect -1099 -4599 -1097 -4597
rect -1083 -4599 -1081 -4597
rect -1075 -4599 -1073 -4597
rect -930 -4599 -928 -4597
rect -920 -4599 -918 -4597
rect -904 -4599 -902 -4597
rect -896 -4599 -894 -4597
rect -880 -4599 -878 -4597
rect -872 -4599 -870 -4597
rect -862 -4599 -860 -4597
rect -854 -4599 -852 -4597
rect -838 -4599 -836 -4597
rect -830 -4599 -828 -4597
rect -820 -4599 -818 -4597
rect -812 -4599 -810 -4597
rect -796 -4599 -794 -4597
rect -788 -4599 -786 -4597
rect -778 -4599 -776 -4597
rect -770 -4599 -768 -4597
rect -754 -4599 -752 -4597
rect -746 -4599 -744 -4597
rect -572 -4599 -570 -4597
rect -562 -4599 -560 -4597
rect -546 -4599 -544 -4597
rect -538 -4599 -536 -4597
rect -522 -4599 -520 -4597
rect -514 -4599 -512 -4597
rect -504 -4599 -502 -4597
rect -496 -4599 -494 -4597
rect -480 -4599 -478 -4597
rect -472 -4599 -470 -4597
rect -462 -4599 -460 -4597
rect -454 -4599 -452 -4597
rect -438 -4599 -436 -4597
rect -430 -4599 -428 -4597
rect -420 -4599 -418 -4597
rect -412 -4599 -410 -4597
rect -396 -4599 -394 -4597
rect -388 -4599 -386 -4597
rect -1259 -4638 -1257 -4636
rect -1249 -4638 -1247 -4636
rect -1233 -4638 -1231 -4636
rect -1225 -4638 -1223 -4636
rect -1209 -4638 -1207 -4636
rect -1201 -4638 -1199 -4636
rect -1191 -4638 -1189 -4636
rect -1183 -4638 -1181 -4636
rect -1167 -4638 -1165 -4636
rect -1159 -4638 -1157 -4636
rect -1149 -4638 -1147 -4636
rect -1141 -4638 -1139 -4636
rect -1125 -4638 -1123 -4636
rect -1117 -4638 -1115 -4636
rect -1107 -4638 -1105 -4636
rect -1099 -4638 -1097 -4636
rect -1083 -4638 -1081 -4636
rect -1075 -4638 -1073 -4636
rect -930 -4638 -928 -4636
rect -920 -4638 -918 -4636
rect -904 -4638 -902 -4636
rect -896 -4638 -894 -4636
rect -880 -4638 -878 -4636
rect -872 -4638 -870 -4636
rect -862 -4638 -860 -4636
rect -854 -4638 -852 -4636
rect -838 -4638 -836 -4636
rect -830 -4638 -828 -4636
rect -820 -4638 -818 -4636
rect -812 -4638 -810 -4636
rect -796 -4638 -794 -4636
rect -788 -4638 -786 -4636
rect -778 -4638 -776 -4636
rect -770 -4638 -768 -4636
rect -754 -4638 -752 -4636
rect -746 -4638 -744 -4636
rect -572 -4638 -570 -4636
rect -562 -4638 -560 -4636
rect -546 -4638 -544 -4636
rect -538 -4638 -536 -4636
rect -522 -4638 -520 -4636
rect -514 -4638 -512 -4636
rect -504 -4638 -502 -4636
rect -496 -4638 -494 -4636
rect -480 -4638 -478 -4636
rect -472 -4638 -470 -4636
rect -462 -4638 -460 -4636
rect -454 -4638 -452 -4636
rect -438 -4638 -436 -4636
rect -430 -4638 -428 -4636
rect -420 -4638 -418 -4636
rect -412 -4638 -410 -4636
rect -396 -4638 -394 -4636
rect -388 -4638 -386 -4636
rect -214 -4638 -212 -4636
rect -204 -4638 -202 -4636
rect -188 -4638 -186 -4636
rect -180 -4638 -178 -4636
rect -164 -4638 -162 -4636
rect -156 -4638 -154 -4636
rect -146 -4638 -144 -4636
rect -138 -4638 -136 -4636
rect -122 -4638 -120 -4636
rect -114 -4638 -112 -4636
rect -104 -4638 -102 -4636
rect -96 -4638 -94 -4636
rect -80 -4638 -78 -4636
rect -72 -4638 -70 -4636
rect -62 -4638 -60 -4636
rect -54 -4638 -52 -4636
rect -38 -4638 -36 -4636
rect -30 -4638 -28 -4636
rect 214 -4638 216 -4636
rect 224 -4638 226 -4636
rect 240 -4638 242 -4636
rect 248 -4638 250 -4636
rect 264 -4638 266 -4636
rect 272 -4638 274 -4636
rect 282 -4638 284 -4636
rect 290 -4638 292 -4636
rect 306 -4638 308 -4636
rect 314 -4638 316 -4636
rect 324 -4638 326 -4636
rect 332 -4638 334 -4636
rect 348 -4638 350 -4636
rect 356 -4638 358 -4636
rect 366 -4638 368 -4636
rect 374 -4638 376 -4636
rect 390 -4638 392 -4636
rect 398 -4638 400 -4636
rect 570 -4638 572 -4636
rect 580 -4638 582 -4636
rect 596 -4638 598 -4636
rect 604 -4638 606 -4636
rect 620 -4638 622 -4636
rect 628 -4638 630 -4636
rect 638 -4638 640 -4636
rect 646 -4638 648 -4636
rect 662 -4638 664 -4636
rect 670 -4638 672 -4636
rect 680 -4638 682 -4636
rect 688 -4638 690 -4636
rect 704 -4638 706 -4636
rect 712 -4638 714 -4636
rect 722 -4638 724 -4636
rect 730 -4638 732 -4636
rect 746 -4638 748 -4636
rect 754 -4638 756 -4636
rect 968 -4638 970 -4636
rect 978 -4638 980 -4636
rect 994 -4638 996 -4636
rect 1002 -4638 1004 -4636
rect 1018 -4638 1020 -4636
rect 1026 -4638 1028 -4636
rect 1036 -4638 1038 -4636
rect 1044 -4638 1046 -4636
rect 1060 -4638 1062 -4636
rect 1068 -4638 1070 -4636
rect 1078 -4638 1080 -4636
rect 1086 -4638 1088 -4636
rect 1102 -4638 1104 -4636
rect 1110 -4638 1112 -4636
rect 1120 -4638 1122 -4636
rect 1128 -4638 1130 -4636
rect 1144 -4638 1146 -4636
rect 1152 -4638 1154 -4636
rect 1326 -4638 1328 -4636
rect 1336 -4638 1338 -4636
rect 1352 -4638 1354 -4636
rect 1360 -4638 1362 -4636
rect 1376 -4638 1378 -4636
rect 1384 -4638 1386 -4636
rect 1394 -4638 1396 -4636
rect 1402 -4638 1404 -4636
rect 1418 -4638 1420 -4636
rect 1426 -4638 1428 -4636
rect 1436 -4638 1438 -4636
rect 1444 -4638 1446 -4636
rect 1460 -4638 1462 -4636
rect 1468 -4638 1470 -4636
rect 1478 -4638 1480 -4636
rect 1486 -4638 1488 -4636
rect 1502 -4638 1504 -4636
rect 1510 -4638 1512 -4636
rect -1259 -4714 -1257 -4646
rect -1249 -4714 -1247 -4646
rect -1233 -4714 -1231 -4646
rect -1225 -4714 -1223 -4646
rect -1209 -4714 -1207 -4646
rect -1201 -4714 -1199 -4646
rect -1191 -4714 -1189 -4646
rect -1183 -4714 -1181 -4646
rect -1167 -4714 -1165 -4646
rect -1159 -4679 -1157 -4646
rect -1149 -4679 -1147 -4646
rect -1159 -4681 -1147 -4679
rect -1159 -4714 -1157 -4681
rect -1149 -4714 -1147 -4681
rect -1141 -4714 -1139 -4646
rect -1125 -4714 -1123 -4646
rect -1117 -4714 -1115 -4646
rect -1107 -4714 -1105 -4646
rect -1099 -4714 -1097 -4646
rect -1083 -4714 -1081 -4646
rect -1075 -4714 -1073 -4646
rect -930 -4714 -928 -4646
rect -920 -4714 -918 -4646
rect -904 -4714 -902 -4646
rect -896 -4714 -894 -4646
rect -880 -4714 -878 -4646
rect -872 -4714 -870 -4646
rect -862 -4714 -860 -4646
rect -854 -4714 -852 -4646
rect -838 -4714 -836 -4646
rect -830 -4679 -828 -4646
rect -820 -4679 -818 -4646
rect -830 -4681 -818 -4679
rect -830 -4714 -828 -4681
rect -820 -4714 -818 -4681
rect -812 -4714 -810 -4646
rect -796 -4714 -794 -4646
rect -788 -4714 -786 -4646
rect -778 -4714 -776 -4646
rect -770 -4714 -768 -4646
rect -754 -4714 -752 -4646
rect -746 -4714 -744 -4646
rect -572 -4714 -570 -4646
rect -562 -4714 -560 -4646
rect -546 -4714 -544 -4646
rect -538 -4714 -536 -4646
rect -522 -4714 -520 -4646
rect -514 -4714 -512 -4646
rect -504 -4714 -502 -4646
rect -496 -4714 -494 -4646
rect -480 -4714 -478 -4646
rect -472 -4679 -470 -4646
rect -462 -4679 -460 -4646
rect -472 -4681 -460 -4679
rect -472 -4714 -470 -4681
rect -462 -4714 -460 -4681
rect -454 -4714 -452 -4646
rect -438 -4714 -436 -4646
rect -430 -4714 -428 -4646
rect -420 -4714 -418 -4646
rect -412 -4714 -410 -4646
rect -396 -4714 -394 -4646
rect -388 -4714 -386 -4646
rect -214 -4714 -212 -4646
rect -204 -4714 -202 -4646
rect -188 -4714 -186 -4646
rect -180 -4714 -178 -4646
rect -164 -4714 -162 -4646
rect -156 -4714 -154 -4646
rect -146 -4714 -144 -4646
rect -138 -4714 -136 -4646
rect -122 -4714 -120 -4646
rect -114 -4679 -112 -4646
rect -104 -4679 -102 -4646
rect -114 -4681 -102 -4679
rect -114 -4714 -112 -4681
rect -104 -4714 -102 -4681
rect -96 -4714 -94 -4646
rect -80 -4714 -78 -4646
rect -72 -4714 -70 -4646
rect -62 -4714 -60 -4646
rect -54 -4714 -52 -4646
rect -38 -4714 -36 -4646
rect -30 -4714 -28 -4646
rect 214 -4714 216 -4646
rect 224 -4714 226 -4646
rect 240 -4714 242 -4646
rect 248 -4714 250 -4646
rect 264 -4714 266 -4646
rect 272 -4714 274 -4646
rect 282 -4714 284 -4646
rect 290 -4714 292 -4646
rect 306 -4714 308 -4646
rect 314 -4679 316 -4646
rect 324 -4679 326 -4646
rect 314 -4681 326 -4679
rect 314 -4714 316 -4681
rect 324 -4714 326 -4681
rect 332 -4714 334 -4646
rect 348 -4714 350 -4646
rect 356 -4714 358 -4646
rect 366 -4714 368 -4646
rect 374 -4714 376 -4646
rect 390 -4714 392 -4646
rect 398 -4714 400 -4646
rect 570 -4714 572 -4646
rect 580 -4714 582 -4646
rect 596 -4714 598 -4646
rect 604 -4714 606 -4646
rect 620 -4714 622 -4646
rect 628 -4714 630 -4646
rect 638 -4714 640 -4646
rect 646 -4714 648 -4646
rect 662 -4714 664 -4646
rect 670 -4679 672 -4646
rect 680 -4679 682 -4646
rect 670 -4681 682 -4679
rect 670 -4714 672 -4681
rect 680 -4714 682 -4681
rect 688 -4714 690 -4646
rect 704 -4714 706 -4646
rect 712 -4714 714 -4646
rect 722 -4714 724 -4646
rect 730 -4714 732 -4646
rect 746 -4714 748 -4646
rect 754 -4714 756 -4646
rect 968 -4714 970 -4646
rect 978 -4714 980 -4646
rect 994 -4714 996 -4646
rect 1002 -4714 1004 -4646
rect 1018 -4714 1020 -4646
rect 1026 -4714 1028 -4646
rect 1036 -4714 1038 -4646
rect 1044 -4714 1046 -4646
rect 1060 -4714 1062 -4646
rect 1068 -4679 1070 -4646
rect 1078 -4679 1080 -4646
rect 1068 -4681 1080 -4679
rect 1068 -4714 1070 -4681
rect 1078 -4714 1080 -4681
rect 1086 -4714 1088 -4646
rect 1102 -4714 1104 -4646
rect 1110 -4714 1112 -4646
rect 1120 -4714 1122 -4646
rect 1128 -4714 1130 -4646
rect 1144 -4714 1146 -4646
rect 1152 -4714 1154 -4646
rect 1326 -4714 1328 -4646
rect 1336 -4714 1338 -4646
rect 1352 -4714 1354 -4646
rect 1360 -4714 1362 -4646
rect 1376 -4714 1378 -4646
rect 1384 -4714 1386 -4646
rect 1394 -4714 1396 -4646
rect 1402 -4714 1404 -4646
rect 1418 -4714 1420 -4646
rect 1426 -4679 1428 -4646
rect 1436 -4679 1438 -4646
rect 1426 -4681 1438 -4679
rect 1426 -4714 1428 -4681
rect 1436 -4714 1438 -4681
rect 1444 -4714 1446 -4646
rect 1460 -4714 1462 -4646
rect 1468 -4714 1470 -4646
rect 1478 -4714 1480 -4646
rect 1486 -4714 1488 -4646
rect 1502 -4714 1504 -4646
rect 1510 -4714 1512 -4646
rect -1259 -4720 -1257 -4718
rect -1249 -4720 -1247 -4718
rect -1233 -4720 -1231 -4718
rect -1225 -4720 -1223 -4718
rect -1209 -4720 -1207 -4718
rect -1201 -4720 -1199 -4718
rect -1191 -4720 -1189 -4718
rect -1183 -4720 -1181 -4718
rect -1167 -4720 -1165 -4718
rect -1159 -4720 -1157 -4718
rect -1149 -4720 -1147 -4718
rect -1141 -4720 -1139 -4718
rect -1125 -4720 -1123 -4718
rect -1117 -4720 -1115 -4718
rect -1107 -4720 -1105 -4718
rect -1099 -4720 -1097 -4718
rect -1083 -4720 -1081 -4718
rect -1075 -4720 -1073 -4718
rect -930 -4720 -928 -4718
rect -920 -4720 -918 -4718
rect -904 -4720 -902 -4718
rect -896 -4720 -894 -4718
rect -880 -4720 -878 -4718
rect -872 -4720 -870 -4718
rect -862 -4720 -860 -4718
rect -854 -4720 -852 -4718
rect -838 -4720 -836 -4718
rect -830 -4720 -828 -4718
rect -820 -4720 -818 -4718
rect -812 -4720 -810 -4718
rect -796 -4720 -794 -4718
rect -788 -4720 -786 -4718
rect -778 -4720 -776 -4718
rect -770 -4720 -768 -4718
rect -754 -4720 -752 -4718
rect -746 -4720 -744 -4718
rect -572 -4720 -570 -4718
rect -562 -4720 -560 -4718
rect -546 -4720 -544 -4718
rect -538 -4720 -536 -4718
rect -522 -4720 -520 -4718
rect -514 -4720 -512 -4718
rect -504 -4720 -502 -4718
rect -496 -4720 -494 -4718
rect -480 -4720 -478 -4718
rect -472 -4720 -470 -4718
rect -462 -4720 -460 -4718
rect -454 -4720 -452 -4718
rect -438 -4720 -436 -4718
rect -430 -4720 -428 -4718
rect -420 -4720 -418 -4718
rect -412 -4720 -410 -4718
rect -396 -4720 -394 -4718
rect -388 -4720 -386 -4718
rect -214 -4720 -212 -4718
rect -204 -4720 -202 -4718
rect -188 -4720 -186 -4718
rect -180 -4720 -178 -4718
rect -164 -4720 -162 -4718
rect -156 -4720 -154 -4718
rect -146 -4720 -144 -4718
rect -138 -4720 -136 -4718
rect -122 -4720 -120 -4718
rect -114 -4720 -112 -4718
rect -104 -4720 -102 -4718
rect -96 -4720 -94 -4718
rect -80 -4720 -78 -4718
rect -72 -4720 -70 -4718
rect -62 -4720 -60 -4718
rect -54 -4720 -52 -4718
rect -38 -4720 -36 -4718
rect -30 -4720 -28 -4718
rect 214 -4720 216 -4718
rect 224 -4720 226 -4718
rect 240 -4720 242 -4718
rect 248 -4720 250 -4718
rect 264 -4720 266 -4718
rect 272 -4720 274 -4718
rect 282 -4720 284 -4718
rect 290 -4720 292 -4718
rect 306 -4720 308 -4718
rect 314 -4720 316 -4718
rect 324 -4720 326 -4718
rect 332 -4720 334 -4718
rect 348 -4720 350 -4718
rect 356 -4720 358 -4718
rect 366 -4720 368 -4718
rect 374 -4720 376 -4718
rect 390 -4720 392 -4718
rect 398 -4720 400 -4718
rect 570 -4720 572 -4718
rect 580 -4720 582 -4718
rect 596 -4720 598 -4718
rect 604 -4720 606 -4718
rect 620 -4720 622 -4718
rect 628 -4720 630 -4718
rect 638 -4720 640 -4718
rect 646 -4720 648 -4718
rect 662 -4720 664 -4718
rect 670 -4720 672 -4718
rect 680 -4720 682 -4718
rect 688 -4720 690 -4718
rect 704 -4720 706 -4718
rect 712 -4720 714 -4718
rect 722 -4720 724 -4718
rect 730 -4720 732 -4718
rect 746 -4720 748 -4718
rect 754 -4720 756 -4718
rect 968 -4720 970 -4718
rect 978 -4720 980 -4718
rect 994 -4720 996 -4718
rect 1002 -4720 1004 -4718
rect 1018 -4720 1020 -4718
rect 1026 -4720 1028 -4718
rect 1036 -4720 1038 -4718
rect 1044 -4720 1046 -4718
rect 1060 -4720 1062 -4718
rect 1068 -4720 1070 -4718
rect 1078 -4720 1080 -4718
rect 1086 -4720 1088 -4718
rect 1102 -4720 1104 -4718
rect 1110 -4720 1112 -4718
rect 1120 -4720 1122 -4718
rect 1128 -4720 1130 -4718
rect 1144 -4720 1146 -4718
rect 1152 -4720 1154 -4718
rect 1326 -4720 1328 -4718
rect 1336 -4720 1338 -4718
rect 1352 -4720 1354 -4718
rect 1360 -4720 1362 -4718
rect 1376 -4720 1378 -4718
rect 1384 -4720 1386 -4718
rect 1394 -4720 1396 -4718
rect 1402 -4720 1404 -4718
rect 1418 -4720 1420 -4718
rect 1426 -4720 1428 -4718
rect 1436 -4720 1438 -4718
rect 1444 -4720 1446 -4718
rect 1460 -4720 1462 -4718
rect 1468 -4720 1470 -4718
rect 1478 -4720 1480 -4718
rect 1486 -4720 1488 -4718
rect 1502 -4720 1504 -4718
rect 1510 -4720 1512 -4718
rect -1259 -4759 -1257 -4757
rect -1249 -4759 -1247 -4757
rect -1233 -4759 -1231 -4757
rect -1225 -4759 -1223 -4757
rect -1209 -4759 -1207 -4757
rect -1201 -4759 -1199 -4757
rect -1191 -4759 -1189 -4757
rect -1183 -4759 -1181 -4757
rect -1167 -4759 -1165 -4757
rect -1159 -4759 -1157 -4757
rect -1149 -4759 -1147 -4757
rect -1141 -4759 -1139 -4757
rect -1125 -4759 -1123 -4757
rect -1117 -4759 -1115 -4757
rect -1107 -4759 -1105 -4757
rect -1099 -4759 -1097 -4757
rect -1083 -4759 -1081 -4757
rect -1075 -4759 -1073 -4757
rect -930 -4759 -928 -4757
rect -920 -4759 -918 -4757
rect -904 -4759 -902 -4757
rect -896 -4759 -894 -4757
rect -880 -4759 -878 -4757
rect -872 -4759 -870 -4757
rect -862 -4759 -860 -4757
rect -854 -4759 -852 -4757
rect -838 -4759 -836 -4757
rect -830 -4759 -828 -4757
rect -820 -4759 -818 -4757
rect -812 -4759 -810 -4757
rect -796 -4759 -794 -4757
rect -788 -4759 -786 -4757
rect -778 -4759 -776 -4757
rect -770 -4759 -768 -4757
rect -754 -4759 -752 -4757
rect -746 -4759 -744 -4757
rect -572 -4759 -570 -4757
rect -562 -4759 -560 -4757
rect -546 -4759 -544 -4757
rect -538 -4759 -536 -4757
rect -522 -4759 -520 -4757
rect -514 -4759 -512 -4757
rect -504 -4759 -502 -4757
rect -496 -4759 -494 -4757
rect -480 -4759 -478 -4757
rect -472 -4759 -470 -4757
rect -462 -4759 -460 -4757
rect -454 -4759 -452 -4757
rect -438 -4759 -436 -4757
rect -430 -4759 -428 -4757
rect -420 -4759 -418 -4757
rect -412 -4759 -410 -4757
rect -396 -4759 -394 -4757
rect -388 -4759 -386 -4757
rect -214 -4759 -212 -4757
rect -204 -4759 -202 -4757
rect -188 -4759 -186 -4757
rect -180 -4759 -178 -4757
rect -164 -4759 -162 -4757
rect -156 -4759 -154 -4757
rect -146 -4759 -144 -4757
rect -138 -4759 -136 -4757
rect -122 -4759 -120 -4757
rect -114 -4759 -112 -4757
rect -104 -4759 -102 -4757
rect -96 -4759 -94 -4757
rect -80 -4759 -78 -4757
rect -72 -4759 -70 -4757
rect -62 -4759 -60 -4757
rect -54 -4759 -52 -4757
rect -38 -4759 -36 -4757
rect -30 -4759 -28 -4757
rect 95 -4759 97 -4757
rect 214 -4759 216 -4757
rect 224 -4759 226 -4757
rect 240 -4759 242 -4757
rect 248 -4759 250 -4757
rect 264 -4759 266 -4757
rect 272 -4759 274 -4757
rect 282 -4759 284 -4757
rect 290 -4759 292 -4757
rect 306 -4759 308 -4757
rect 314 -4759 316 -4757
rect 324 -4759 326 -4757
rect 332 -4759 334 -4757
rect 348 -4759 350 -4757
rect 356 -4759 358 -4757
rect 366 -4759 368 -4757
rect 374 -4759 376 -4757
rect 390 -4759 392 -4757
rect 398 -4759 400 -4757
rect 570 -4759 572 -4757
rect 580 -4759 582 -4757
rect 596 -4759 598 -4757
rect 604 -4759 606 -4757
rect 620 -4759 622 -4757
rect 628 -4759 630 -4757
rect 638 -4759 640 -4757
rect 646 -4759 648 -4757
rect 662 -4759 664 -4757
rect 670 -4759 672 -4757
rect 680 -4759 682 -4757
rect 688 -4759 690 -4757
rect 704 -4759 706 -4757
rect 712 -4759 714 -4757
rect 722 -4759 724 -4757
rect 730 -4759 732 -4757
rect 746 -4759 748 -4757
rect 754 -4759 756 -4757
rect 968 -4759 970 -4757
rect 978 -4759 980 -4757
rect 994 -4759 996 -4757
rect 1002 -4759 1004 -4757
rect 1018 -4759 1020 -4757
rect 1026 -4759 1028 -4757
rect 1036 -4759 1038 -4757
rect 1044 -4759 1046 -4757
rect 1060 -4759 1062 -4757
rect 1068 -4759 1070 -4757
rect 1078 -4759 1080 -4757
rect 1086 -4759 1088 -4757
rect 1102 -4759 1104 -4757
rect 1110 -4759 1112 -4757
rect 1120 -4759 1122 -4757
rect 1128 -4759 1130 -4757
rect 1144 -4759 1146 -4757
rect 1152 -4759 1154 -4757
rect 1326 -4759 1328 -4757
rect 1336 -4759 1338 -4757
rect 1352 -4759 1354 -4757
rect 1360 -4759 1362 -4757
rect 1376 -4759 1378 -4757
rect 1384 -4759 1386 -4757
rect 1394 -4759 1396 -4757
rect 1402 -4759 1404 -4757
rect 1418 -4759 1420 -4757
rect 1426 -4759 1428 -4757
rect 1436 -4759 1438 -4757
rect 1444 -4759 1446 -4757
rect 1460 -4759 1462 -4757
rect 1468 -4759 1470 -4757
rect 1478 -4759 1480 -4757
rect 1486 -4759 1488 -4757
rect 1502 -4759 1504 -4757
rect 1510 -4759 1512 -4757
rect -1259 -4835 -1257 -4767
rect -1249 -4835 -1247 -4767
rect -1233 -4835 -1231 -4767
rect -1225 -4835 -1223 -4767
rect -1209 -4835 -1207 -4767
rect -1201 -4835 -1199 -4767
rect -1191 -4835 -1189 -4767
rect -1183 -4835 -1181 -4767
rect -1167 -4835 -1165 -4767
rect -1159 -4800 -1157 -4767
rect -1149 -4800 -1147 -4767
rect -1159 -4802 -1147 -4800
rect -1159 -4835 -1157 -4802
rect -1149 -4835 -1147 -4802
rect -1141 -4835 -1139 -4767
rect -1125 -4835 -1123 -4767
rect -1117 -4835 -1115 -4767
rect -1107 -4835 -1105 -4767
rect -1099 -4835 -1097 -4767
rect -1083 -4835 -1081 -4767
rect -1075 -4835 -1073 -4767
rect -930 -4835 -928 -4767
rect -920 -4835 -918 -4767
rect -904 -4835 -902 -4767
rect -896 -4835 -894 -4767
rect -880 -4835 -878 -4767
rect -872 -4835 -870 -4767
rect -862 -4835 -860 -4767
rect -854 -4835 -852 -4767
rect -838 -4835 -836 -4767
rect -830 -4800 -828 -4767
rect -820 -4800 -818 -4767
rect -830 -4802 -818 -4800
rect -830 -4835 -828 -4802
rect -820 -4835 -818 -4802
rect -812 -4835 -810 -4767
rect -796 -4835 -794 -4767
rect -788 -4835 -786 -4767
rect -778 -4835 -776 -4767
rect -770 -4835 -768 -4767
rect -754 -4835 -752 -4767
rect -746 -4835 -744 -4767
rect -572 -4835 -570 -4767
rect -562 -4835 -560 -4767
rect -546 -4835 -544 -4767
rect -538 -4835 -536 -4767
rect -522 -4835 -520 -4767
rect -514 -4835 -512 -4767
rect -504 -4835 -502 -4767
rect -496 -4835 -494 -4767
rect -480 -4835 -478 -4767
rect -472 -4800 -470 -4767
rect -462 -4800 -460 -4767
rect -472 -4802 -460 -4800
rect -472 -4835 -470 -4802
rect -462 -4835 -460 -4802
rect -454 -4835 -452 -4767
rect -438 -4835 -436 -4767
rect -430 -4835 -428 -4767
rect -420 -4835 -418 -4767
rect -412 -4835 -410 -4767
rect -396 -4835 -394 -4767
rect -388 -4835 -386 -4767
rect -214 -4835 -212 -4767
rect -204 -4835 -202 -4767
rect -188 -4835 -186 -4767
rect -180 -4835 -178 -4767
rect -164 -4835 -162 -4767
rect -156 -4835 -154 -4767
rect -146 -4835 -144 -4767
rect -138 -4835 -136 -4767
rect -122 -4835 -120 -4767
rect -114 -4800 -112 -4767
rect -104 -4800 -102 -4767
rect -114 -4802 -102 -4800
rect -114 -4835 -112 -4802
rect -104 -4835 -102 -4802
rect -96 -4835 -94 -4767
rect -80 -4835 -78 -4767
rect -72 -4835 -70 -4767
rect -62 -4835 -60 -4767
rect -54 -4835 -52 -4767
rect -38 -4835 -36 -4767
rect -30 -4835 -28 -4767
rect 95 -4823 97 -4791
rect 214 -4835 216 -4767
rect 224 -4835 226 -4767
rect 240 -4835 242 -4767
rect 248 -4835 250 -4767
rect 264 -4835 266 -4767
rect 272 -4835 274 -4767
rect 282 -4835 284 -4767
rect 290 -4835 292 -4767
rect 306 -4835 308 -4767
rect 314 -4800 316 -4767
rect 324 -4800 326 -4767
rect 314 -4802 326 -4800
rect 314 -4835 316 -4802
rect 324 -4835 326 -4802
rect 332 -4835 334 -4767
rect 348 -4835 350 -4767
rect 356 -4835 358 -4767
rect 366 -4835 368 -4767
rect 374 -4835 376 -4767
rect 390 -4835 392 -4767
rect 398 -4835 400 -4767
rect 570 -4835 572 -4767
rect 580 -4835 582 -4767
rect 596 -4835 598 -4767
rect 604 -4835 606 -4767
rect 620 -4835 622 -4767
rect 628 -4835 630 -4767
rect 638 -4835 640 -4767
rect 646 -4835 648 -4767
rect 662 -4835 664 -4767
rect 670 -4800 672 -4767
rect 680 -4800 682 -4767
rect 670 -4802 682 -4800
rect 670 -4835 672 -4802
rect 680 -4835 682 -4802
rect 688 -4835 690 -4767
rect 704 -4835 706 -4767
rect 712 -4835 714 -4767
rect 722 -4835 724 -4767
rect 730 -4835 732 -4767
rect 746 -4835 748 -4767
rect 754 -4835 756 -4767
rect 968 -4835 970 -4767
rect 978 -4835 980 -4767
rect 994 -4835 996 -4767
rect 1002 -4835 1004 -4767
rect 1018 -4835 1020 -4767
rect 1026 -4835 1028 -4767
rect 1036 -4835 1038 -4767
rect 1044 -4835 1046 -4767
rect 1060 -4835 1062 -4767
rect 1068 -4800 1070 -4767
rect 1078 -4800 1080 -4767
rect 1068 -4802 1080 -4800
rect 1068 -4835 1070 -4802
rect 1078 -4835 1080 -4802
rect 1086 -4835 1088 -4767
rect 1102 -4835 1104 -4767
rect 1110 -4835 1112 -4767
rect 1120 -4835 1122 -4767
rect 1128 -4835 1130 -4767
rect 1144 -4835 1146 -4767
rect 1152 -4835 1154 -4767
rect 1326 -4835 1328 -4767
rect 1336 -4835 1338 -4767
rect 1352 -4835 1354 -4767
rect 1360 -4835 1362 -4767
rect 1376 -4835 1378 -4767
rect 1384 -4835 1386 -4767
rect 1394 -4835 1396 -4767
rect 1402 -4835 1404 -4767
rect 1418 -4835 1420 -4767
rect 1426 -4800 1428 -4767
rect 1436 -4800 1438 -4767
rect 1426 -4802 1438 -4800
rect 1426 -4835 1428 -4802
rect 1436 -4835 1438 -4802
rect 1444 -4835 1446 -4767
rect 1460 -4835 1462 -4767
rect 1468 -4835 1470 -4767
rect 1478 -4835 1480 -4767
rect 1486 -4835 1488 -4767
rect 1502 -4835 1504 -4767
rect 1510 -4835 1512 -4767
rect -1259 -4841 -1257 -4839
rect -1249 -4841 -1247 -4839
rect -1233 -4841 -1231 -4839
rect -1225 -4841 -1223 -4839
rect -1209 -4841 -1207 -4839
rect -1201 -4841 -1199 -4839
rect -1191 -4841 -1189 -4839
rect -1183 -4841 -1181 -4839
rect -1167 -4841 -1165 -4839
rect -1159 -4841 -1157 -4839
rect -1149 -4841 -1147 -4839
rect -1141 -4841 -1139 -4839
rect -1125 -4841 -1123 -4839
rect -1117 -4841 -1115 -4839
rect -1107 -4841 -1105 -4839
rect -1099 -4841 -1097 -4839
rect -1083 -4841 -1081 -4839
rect -1075 -4841 -1073 -4839
rect -930 -4841 -928 -4839
rect -920 -4841 -918 -4839
rect -904 -4841 -902 -4839
rect -896 -4841 -894 -4839
rect -880 -4841 -878 -4839
rect -872 -4841 -870 -4839
rect -862 -4841 -860 -4839
rect -854 -4841 -852 -4839
rect -838 -4841 -836 -4839
rect -830 -4841 -828 -4839
rect -820 -4841 -818 -4839
rect -812 -4841 -810 -4839
rect -796 -4841 -794 -4839
rect -788 -4841 -786 -4839
rect -778 -4841 -776 -4839
rect -770 -4841 -768 -4839
rect -754 -4841 -752 -4839
rect -746 -4841 -744 -4839
rect -572 -4841 -570 -4839
rect -562 -4841 -560 -4839
rect -546 -4841 -544 -4839
rect -538 -4841 -536 -4839
rect -522 -4841 -520 -4839
rect -514 -4841 -512 -4839
rect -504 -4841 -502 -4839
rect -496 -4841 -494 -4839
rect -480 -4841 -478 -4839
rect -472 -4841 -470 -4839
rect -462 -4841 -460 -4839
rect -454 -4841 -452 -4839
rect -438 -4841 -436 -4839
rect -430 -4841 -428 -4839
rect -420 -4841 -418 -4839
rect -412 -4841 -410 -4839
rect -396 -4841 -394 -4839
rect -388 -4841 -386 -4839
rect -214 -4841 -212 -4839
rect -204 -4841 -202 -4839
rect -188 -4841 -186 -4839
rect -180 -4841 -178 -4839
rect -164 -4841 -162 -4839
rect -156 -4841 -154 -4839
rect -146 -4841 -144 -4839
rect -138 -4841 -136 -4839
rect -122 -4841 -120 -4839
rect -114 -4841 -112 -4839
rect -104 -4841 -102 -4839
rect -96 -4841 -94 -4839
rect -80 -4841 -78 -4839
rect -72 -4841 -70 -4839
rect -62 -4841 -60 -4839
rect -54 -4841 -52 -4839
rect -38 -4841 -36 -4839
rect -30 -4841 -28 -4839
rect 95 -4841 97 -4839
rect 214 -4841 216 -4839
rect 224 -4841 226 -4839
rect 240 -4841 242 -4839
rect 248 -4841 250 -4839
rect 264 -4841 266 -4839
rect 272 -4841 274 -4839
rect 282 -4841 284 -4839
rect 290 -4841 292 -4839
rect 306 -4841 308 -4839
rect 314 -4841 316 -4839
rect 324 -4841 326 -4839
rect 332 -4841 334 -4839
rect 348 -4841 350 -4839
rect 356 -4841 358 -4839
rect 366 -4841 368 -4839
rect 374 -4841 376 -4839
rect 390 -4841 392 -4839
rect 398 -4841 400 -4839
rect 570 -4841 572 -4839
rect 580 -4841 582 -4839
rect 596 -4841 598 -4839
rect 604 -4841 606 -4839
rect 620 -4841 622 -4839
rect 628 -4841 630 -4839
rect 638 -4841 640 -4839
rect 646 -4841 648 -4839
rect 662 -4841 664 -4839
rect 670 -4841 672 -4839
rect 680 -4841 682 -4839
rect 688 -4841 690 -4839
rect 704 -4841 706 -4839
rect 712 -4841 714 -4839
rect 722 -4841 724 -4839
rect 730 -4841 732 -4839
rect 746 -4841 748 -4839
rect 754 -4841 756 -4839
rect 968 -4841 970 -4839
rect 978 -4841 980 -4839
rect 994 -4841 996 -4839
rect 1002 -4841 1004 -4839
rect 1018 -4841 1020 -4839
rect 1026 -4841 1028 -4839
rect 1036 -4841 1038 -4839
rect 1044 -4841 1046 -4839
rect 1060 -4841 1062 -4839
rect 1068 -4841 1070 -4839
rect 1078 -4841 1080 -4839
rect 1086 -4841 1088 -4839
rect 1102 -4841 1104 -4839
rect 1110 -4841 1112 -4839
rect 1120 -4841 1122 -4839
rect 1128 -4841 1130 -4839
rect 1144 -4841 1146 -4839
rect 1152 -4841 1154 -4839
rect 1326 -4841 1328 -4839
rect 1336 -4841 1338 -4839
rect 1352 -4841 1354 -4839
rect 1360 -4841 1362 -4839
rect 1376 -4841 1378 -4839
rect 1384 -4841 1386 -4839
rect 1394 -4841 1396 -4839
rect 1402 -4841 1404 -4839
rect 1418 -4841 1420 -4839
rect 1426 -4841 1428 -4839
rect 1436 -4841 1438 -4839
rect 1444 -4841 1446 -4839
rect 1460 -4841 1462 -4839
rect 1468 -4841 1470 -4839
rect 1478 -4841 1480 -4839
rect 1486 -4841 1488 -4839
rect 1502 -4841 1504 -4839
rect 1510 -4841 1512 -4839
rect -1259 -4877 -1257 -4875
rect -1249 -4877 -1247 -4875
rect -1233 -4877 -1231 -4875
rect -1225 -4877 -1223 -4875
rect -1209 -4877 -1207 -4875
rect -1201 -4877 -1199 -4875
rect -1191 -4877 -1189 -4875
rect -1183 -4877 -1181 -4875
rect -1167 -4877 -1165 -4875
rect -1159 -4877 -1157 -4875
rect -1149 -4877 -1147 -4875
rect -1141 -4877 -1139 -4875
rect -1125 -4877 -1123 -4875
rect -1117 -4877 -1115 -4875
rect -1107 -4877 -1105 -4875
rect -1099 -4877 -1097 -4875
rect -1083 -4877 -1081 -4875
rect -1075 -4877 -1073 -4875
rect -930 -4877 -928 -4875
rect -920 -4877 -918 -4875
rect -904 -4877 -902 -4875
rect -896 -4877 -894 -4875
rect -880 -4877 -878 -4875
rect -872 -4877 -870 -4875
rect -862 -4877 -860 -4875
rect -854 -4877 -852 -4875
rect -838 -4877 -836 -4875
rect -830 -4877 -828 -4875
rect -820 -4877 -818 -4875
rect -812 -4877 -810 -4875
rect -796 -4877 -794 -4875
rect -788 -4877 -786 -4875
rect -778 -4877 -776 -4875
rect -770 -4877 -768 -4875
rect -754 -4877 -752 -4875
rect -746 -4877 -744 -4875
rect -572 -4877 -570 -4875
rect -562 -4877 -560 -4875
rect -546 -4877 -544 -4875
rect -538 -4877 -536 -4875
rect -522 -4877 -520 -4875
rect -514 -4877 -512 -4875
rect -504 -4877 -502 -4875
rect -496 -4877 -494 -4875
rect -480 -4877 -478 -4875
rect -472 -4877 -470 -4875
rect -462 -4877 -460 -4875
rect -454 -4877 -452 -4875
rect -438 -4877 -436 -4875
rect -430 -4877 -428 -4875
rect -420 -4877 -418 -4875
rect -412 -4877 -410 -4875
rect -396 -4877 -394 -4875
rect -388 -4877 -386 -4875
rect -214 -4877 -212 -4875
rect -204 -4877 -202 -4875
rect -188 -4877 -186 -4875
rect -180 -4877 -178 -4875
rect -164 -4877 -162 -4875
rect -156 -4877 -154 -4875
rect -146 -4877 -144 -4875
rect -138 -4877 -136 -4875
rect -122 -4877 -120 -4875
rect -114 -4877 -112 -4875
rect -104 -4877 -102 -4875
rect -96 -4877 -94 -4875
rect -80 -4877 -78 -4875
rect -72 -4877 -70 -4875
rect -62 -4877 -60 -4875
rect -54 -4877 -52 -4875
rect -38 -4877 -36 -4875
rect -30 -4877 -28 -4875
rect 214 -4877 216 -4875
rect 224 -4877 226 -4875
rect 240 -4877 242 -4875
rect 248 -4877 250 -4875
rect 264 -4877 266 -4875
rect 272 -4877 274 -4875
rect 282 -4877 284 -4875
rect 290 -4877 292 -4875
rect 306 -4877 308 -4875
rect 314 -4877 316 -4875
rect 324 -4877 326 -4875
rect 332 -4877 334 -4875
rect 348 -4877 350 -4875
rect 356 -4877 358 -4875
rect 366 -4877 368 -4875
rect 374 -4877 376 -4875
rect 390 -4877 392 -4875
rect 398 -4877 400 -4875
rect -1259 -4953 -1257 -4885
rect -1249 -4953 -1247 -4885
rect -1233 -4953 -1231 -4885
rect -1225 -4953 -1223 -4885
rect -1209 -4953 -1207 -4885
rect -1201 -4953 -1199 -4885
rect -1191 -4953 -1189 -4885
rect -1183 -4953 -1181 -4885
rect -1167 -4953 -1165 -4885
rect -1159 -4918 -1157 -4885
rect -1149 -4918 -1147 -4885
rect -1159 -4920 -1147 -4918
rect -1159 -4953 -1157 -4920
rect -1149 -4953 -1147 -4920
rect -1141 -4953 -1139 -4885
rect -1125 -4953 -1123 -4885
rect -1117 -4953 -1115 -4885
rect -1107 -4953 -1105 -4885
rect -1099 -4953 -1097 -4885
rect -1083 -4953 -1081 -4885
rect -1075 -4953 -1073 -4885
rect -930 -4953 -928 -4885
rect -920 -4953 -918 -4885
rect -904 -4953 -902 -4885
rect -896 -4953 -894 -4885
rect -880 -4953 -878 -4885
rect -872 -4953 -870 -4885
rect -862 -4953 -860 -4885
rect -854 -4953 -852 -4885
rect -838 -4953 -836 -4885
rect -830 -4918 -828 -4885
rect -820 -4918 -818 -4885
rect -830 -4920 -818 -4918
rect -830 -4953 -828 -4920
rect -820 -4953 -818 -4920
rect -812 -4953 -810 -4885
rect -796 -4953 -794 -4885
rect -788 -4953 -786 -4885
rect -778 -4953 -776 -4885
rect -770 -4953 -768 -4885
rect -754 -4953 -752 -4885
rect -746 -4953 -744 -4885
rect -572 -4953 -570 -4885
rect -562 -4953 -560 -4885
rect -546 -4953 -544 -4885
rect -538 -4953 -536 -4885
rect -522 -4953 -520 -4885
rect -514 -4953 -512 -4885
rect -504 -4953 -502 -4885
rect -496 -4953 -494 -4885
rect -480 -4953 -478 -4885
rect -472 -4918 -470 -4885
rect -462 -4918 -460 -4885
rect -472 -4920 -460 -4918
rect -472 -4953 -470 -4920
rect -462 -4953 -460 -4920
rect -454 -4953 -452 -4885
rect -438 -4953 -436 -4885
rect -430 -4953 -428 -4885
rect -420 -4953 -418 -4885
rect -412 -4953 -410 -4885
rect -396 -4953 -394 -4885
rect -388 -4953 -386 -4885
rect -214 -4953 -212 -4885
rect -204 -4953 -202 -4885
rect -188 -4953 -186 -4885
rect -180 -4953 -178 -4885
rect -164 -4953 -162 -4885
rect -156 -4953 -154 -4885
rect -146 -4953 -144 -4885
rect -138 -4953 -136 -4885
rect -122 -4953 -120 -4885
rect -114 -4918 -112 -4885
rect -104 -4918 -102 -4885
rect -114 -4920 -102 -4918
rect -114 -4953 -112 -4920
rect -104 -4953 -102 -4920
rect -96 -4953 -94 -4885
rect -80 -4953 -78 -4885
rect -72 -4953 -70 -4885
rect -62 -4953 -60 -4885
rect -54 -4953 -52 -4885
rect -38 -4953 -36 -4885
rect -30 -4953 -28 -4885
rect 214 -4953 216 -4885
rect 224 -4953 226 -4885
rect 240 -4953 242 -4885
rect 248 -4953 250 -4885
rect 264 -4953 266 -4885
rect 272 -4953 274 -4885
rect 282 -4953 284 -4885
rect 290 -4953 292 -4885
rect 306 -4953 308 -4885
rect 314 -4918 316 -4885
rect 324 -4918 326 -4885
rect 314 -4920 326 -4918
rect 314 -4953 316 -4920
rect 324 -4953 326 -4920
rect 332 -4953 334 -4885
rect 348 -4953 350 -4885
rect 356 -4953 358 -4885
rect 366 -4953 368 -4885
rect 374 -4953 376 -4885
rect 390 -4953 392 -4885
rect 398 -4953 400 -4885
rect -1259 -4959 -1257 -4957
rect -1249 -4959 -1247 -4957
rect -1233 -4959 -1231 -4957
rect -1225 -4959 -1223 -4957
rect -1209 -4959 -1207 -4957
rect -1201 -4959 -1199 -4957
rect -1191 -4959 -1189 -4957
rect -1183 -4959 -1181 -4957
rect -1167 -4959 -1165 -4957
rect -1159 -4959 -1157 -4957
rect -1149 -4959 -1147 -4957
rect -1141 -4959 -1139 -4957
rect -1125 -4959 -1123 -4957
rect -1117 -4959 -1115 -4957
rect -1107 -4959 -1105 -4957
rect -1099 -4959 -1097 -4957
rect -1083 -4959 -1081 -4957
rect -1075 -4959 -1073 -4957
rect -930 -4959 -928 -4957
rect -920 -4959 -918 -4957
rect -904 -4959 -902 -4957
rect -896 -4959 -894 -4957
rect -880 -4959 -878 -4957
rect -872 -4959 -870 -4957
rect -862 -4959 -860 -4957
rect -854 -4959 -852 -4957
rect -838 -4959 -836 -4957
rect -830 -4959 -828 -4957
rect -820 -4959 -818 -4957
rect -812 -4959 -810 -4957
rect -796 -4959 -794 -4957
rect -788 -4959 -786 -4957
rect -778 -4959 -776 -4957
rect -770 -4959 -768 -4957
rect -754 -4959 -752 -4957
rect -746 -4959 -744 -4957
rect -572 -4959 -570 -4957
rect -562 -4959 -560 -4957
rect -546 -4959 -544 -4957
rect -538 -4959 -536 -4957
rect -522 -4959 -520 -4957
rect -514 -4959 -512 -4957
rect -504 -4959 -502 -4957
rect -496 -4959 -494 -4957
rect -480 -4959 -478 -4957
rect -472 -4959 -470 -4957
rect -462 -4959 -460 -4957
rect -454 -4959 -452 -4957
rect -438 -4959 -436 -4957
rect -430 -4959 -428 -4957
rect -420 -4959 -418 -4957
rect -412 -4959 -410 -4957
rect -396 -4959 -394 -4957
rect -388 -4959 -386 -4957
rect -214 -4959 -212 -4957
rect -204 -4959 -202 -4957
rect -188 -4959 -186 -4957
rect -180 -4959 -178 -4957
rect -164 -4959 -162 -4957
rect -156 -4959 -154 -4957
rect -146 -4959 -144 -4957
rect -138 -4959 -136 -4957
rect -122 -4959 -120 -4957
rect -114 -4959 -112 -4957
rect -104 -4959 -102 -4957
rect -96 -4959 -94 -4957
rect -80 -4959 -78 -4957
rect -72 -4959 -70 -4957
rect -62 -4959 -60 -4957
rect -54 -4959 -52 -4957
rect -38 -4959 -36 -4957
rect -30 -4959 -28 -4957
rect 214 -4959 216 -4957
rect 224 -4959 226 -4957
rect 240 -4959 242 -4957
rect 248 -4959 250 -4957
rect 264 -4959 266 -4957
rect 272 -4959 274 -4957
rect 282 -4959 284 -4957
rect 290 -4959 292 -4957
rect 306 -4959 308 -4957
rect 314 -4959 316 -4957
rect 324 -4959 326 -4957
rect 332 -4959 334 -4957
rect 348 -4959 350 -4957
rect 356 -4959 358 -4957
rect 366 -4959 368 -4957
rect 374 -4959 376 -4957
rect 390 -4959 392 -4957
rect 398 -4959 400 -4957
rect -1334 -4994 -1332 -4992
rect -1326 -4994 -1324 -4992
rect -1316 -4994 -1314 -4992
rect -930 -4994 -928 -4992
rect -922 -4994 -920 -4992
rect -912 -4994 -910 -4992
rect -572 -4994 -570 -4992
rect -564 -4994 -562 -4992
rect -554 -4994 -552 -4992
rect -214 -4994 -212 -4992
rect -206 -4994 -204 -4992
rect -196 -4994 -194 -4992
rect 214 -4994 216 -4992
rect 222 -4994 224 -4992
rect 232 -4994 234 -4992
rect 570 -4994 572 -4992
rect 578 -4994 580 -4992
rect 588 -4994 590 -4992
rect 968 -4994 970 -4992
rect 976 -4994 978 -4992
rect 986 -4994 988 -4992
rect 1326 -4994 1328 -4992
rect 1334 -4994 1336 -4992
rect 1344 -4994 1346 -4992
rect -1334 -5070 -1332 -5002
rect -1326 -5026 -1324 -5002
rect -1326 -5070 -1324 -5030
rect -1316 -5070 -1314 -5002
rect -930 -5070 -928 -5002
rect -922 -5026 -920 -5002
rect -922 -5070 -920 -5030
rect -912 -5070 -910 -5002
rect -572 -5070 -570 -5002
rect -564 -5026 -562 -5002
rect -564 -5070 -562 -5030
rect -554 -5070 -552 -5002
rect -214 -5070 -212 -5002
rect -206 -5026 -204 -5002
rect -206 -5070 -204 -5030
rect -196 -5070 -194 -5002
rect 214 -5070 216 -5002
rect 222 -5026 224 -5002
rect 222 -5070 224 -5030
rect 232 -5070 234 -5002
rect 570 -5070 572 -5002
rect 578 -5026 580 -5002
rect 578 -5070 580 -5030
rect 588 -5070 590 -5002
rect 968 -5070 970 -5002
rect 976 -5026 978 -5002
rect 976 -5070 978 -5030
rect 986 -5070 988 -5002
rect 1326 -5070 1328 -5002
rect 1334 -5026 1336 -5002
rect 1334 -5070 1336 -5030
rect 1344 -5070 1346 -5002
rect -1334 -5076 -1332 -5074
rect -1326 -5076 -1324 -5074
rect -1316 -5076 -1314 -5074
rect -930 -5076 -928 -5074
rect -922 -5076 -920 -5074
rect -912 -5076 -910 -5074
rect -572 -5076 -570 -5074
rect -564 -5076 -562 -5074
rect -554 -5076 -552 -5074
rect -214 -5076 -212 -5074
rect -206 -5076 -204 -5074
rect -196 -5076 -194 -5074
rect 214 -5076 216 -5074
rect 222 -5076 224 -5074
rect 232 -5076 234 -5074
rect 570 -5076 572 -5074
rect 578 -5076 580 -5074
rect 588 -5076 590 -5074
rect 968 -5076 970 -5074
rect 976 -5076 978 -5074
rect 986 -5076 988 -5074
rect 1326 -5076 1328 -5074
rect 1334 -5076 1336 -5074
rect 1344 -5076 1346 -5074
rect -1259 -5113 -1257 -5111
rect -1249 -5113 -1247 -5111
rect -1233 -5113 -1231 -5111
rect -1223 -5113 -1221 -5111
rect -1215 -5113 -1213 -5111
rect -1205 -5113 -1203 -5111
rect -1189 -5113 -1187 -5111
rect -1181 -5113 -1179 -5111
rect -1171 -5113 -1169 -5111
rect -930 -5113 -928 -5111
rect -920 -5113 -918 -5111
rect -904 -5113 -902 -5111
rect -894 -5113 -892 -5111
rect -878 -5113 -876 -5111
rect -868 -5113 -866 -5111
rect -860 -5113 -858 -5111
rect -850 -5113 -848 -5111
rect -834 -5113 -832 -5111
rect -826 -5113 -824 -5111
rect -816 -5113 -814 -5111
rect -800 -5113 -798 -5111
rect -790 -5113 -788 -5111
rect -782 -5113 -780 -5111
rect -772 -5113 -770 -5111
rect -756 -5113 -754 -5111
rect -748 -5113 -746 -5111
rect -732 -5113 -730 -5111
rect -716 -5113 -714 -5111
rect -708 -5113 -706 -5111
rect -698 -5113 -696 -5111
rect -572 -5113 -570 -5111
rect -562 -5113 -560 -5111
rect -546 -5113 -544 -5111
rect -536 -5113 -534 -5111
rect -520 -5113 -518 -5111
rect -510 -5113 -508 -5111
rect -502 -5113 -500 -5111
rect -492 -5113 -490 -5111
rect -476 -5113 -474 -5111
rect -468 -5113 -466 -5111
rect -458 -5113 -456 -5111
rect -442 -5113 -440 -5111
rect -432 -5113 -430 -5111
rect -424 -5113 -422 -5111
rect -414 -5113 -412 -5111
rect -398 -5113 -396 -5111
rect -390 -5113 -388 -5111
rect -374 -5113 -372 -5111
rect -358 -5113 -356 -5111
rect -350 -5113 -348 -5111
rect -340 -5113 -338 -5111
rect -214 -5113 -212 -5111
rect -204 -5113 -202 -5111
rect -188 -5113 -186 -5111
rect -178 -5113 -176 -5111
rect -162 -5113 -160 -5111
rect -152 -5113 -150 -5111
rect -144 -5113 -142 -5111
rect -134 -5113 -132 -5111
rect -118 -5113 -116 -5111
rect -110 -5113 -108 -5111
rect -100 -5113 -98 -5111
rect -84 -5113 -82 -5111
rect -74 -5113 -72 -5111
rect -66 -5113 -64 -5111
rect -56 -5113 -54 -5111
rect -40 -5113 -38 -5111
rect -32 -5113 -30 -5111
rect -16 -5113 -14 -5111
rect 0 -5113 2 -5111
rect 8 -5113 10 -5111
rect 18 -5113 20 -5111
rect 214 -5113 216 -5111
rect 224 -5113 226 -5111
rect 240 -5113 242 -5111
rect 250 -5113 252 -5111
rect 266 -5113 268 -5111
rect 276 -5113 278 -5111
rect 284 -5113 286 -5111
rect 294 -5113 296 -5111
rect 310 -5113 312 -5111
rect 318 -5113 320 -5111
rect 328 -5113 330 -5111
rect 344 -5113 346 -5111
rect 354 -5113 356 -5111
rect 362 -5113 364 -5111
rect 372 -5113 374 -5111
rect 388 -5113 390 -5111
rect 396 -5113 398 -5111
rect 412 -5113 414 -5111
rect 428 -5113 430 -5111
rect 436 -5113 438 -5111
rect 446 -5113 448 -5111
rect 570 -5113 572 -5111
rect 580 -5113 582 -5111
rect 596 -5113 598 -5111
rect 606 -5113 608 -5111
rect 622 -5113 624 -5111
rect 632 -5113 634 -5111
rect 640 -5113 642 -5111
rect 650 -5113 652 -5111
rect 666 -5113 668 -5111
rect 674 -5113 676 -5111
rect 684 -5113 686 -5111
rect 700 -5113 702 -5111
rect 710 -5113 712 -5111
rect 718 -5113 720 -5111
rect 728 -5113 730 -5111
rect 744 -5113 746 -5111
rect 752 -5113 754 -5111
rect 768 -5113 770 -5111
rect 784 -5113 786 -5111
rect 792 -5113 794 -5111
rect 802 -5113 804 -5111
rect 968 -5113 970 -5111
rect 978 -5113 980 -5111
rect 994 -5113 996 -5111
rect 1004 -5113 1006 -5111
rect 1020 -5113 1022 -5111
rect 1030 -5113 1032 -5111
rect 1038 -5113 1040 -5111
rect 1048 -5113 1050 -5111
rect 1064 -5113 1066 -5111
rect 1072 -5113 1074 -5111
rect 1082 -5113 1084 -5111
rect 1098 -5113 1100 -5111
rect 1108 -5113 1110 -5111
rect 1116 -5113 1118 -5111
rect 1126 -5113 1128 -5111
rect 1142 -5113 1144 -5111
rect 1150 -5113 1152 -5111
rect 1166 -5113 1168 -5111
rect 1182 -5113 1184 -5111
rect 1190 -5113 1192 -5111
rect 1200 -5113 1202 -5111
rect 1326 -5113 1328 -5111
rect 1336 -5113 1338 -5111
rect 1352 -5113 1354 -5111
rect 1362 -5113 1364 -5111
rect 1378 -5113 1380 -5111
rect 1388 -5113 1390 -5111
rect 1396 -5113 1398 -5111
rect 1406 -5113 1408 -5111
rect 1422 -5113 1424 -5111
rect 1430 -5113 1432 -5111
rect 1440 -5113 1442 -5111
rect 1456 -5113 1458 -5111
rect 1466 -5113 1468 -5111
rect 1474 -5113 1476 -5111
rect 1484 -5113 1486 -5111
rect 1500 -5113 1502 -5111
rect 1508 -5113 1510 -5111
rect 1524 -5113 1526 -5111
rect 1540 -5113 1542 -5111
rect 1548 -5113 1550 -5111
rect 1558 -5113 1560 -5111
rect -1259 -5189 -1257 -5121
rect -1249 -5189 -1247 -5121
rect -1233 -5189 -1231 -5121
rect -1223 -5189 -1221 -5121
rect -1215 -5189 -1213 -5121
rect -1205 -5189 -1203 -5121
rect -1189 -5189 -1187 -5121
rect -1181 -5189 -1179 -5121
rect -1171 -5189 -1169 -5121
rect -930 -5189 -928 -5121
rect -920 -5189 -918 -5121
rect -904 -5189 -902 -5121
rect -894 -5189 -892 -5121
rect -878 -5189 -876 -5121
rect -868 -5189 -866 -5121
rect -860 -5189 -858 -5121
rect -850 -5189 -848 -5121
rect -834 -5189 -832 -5121
rect -826 -5189 -824 -5121
rect -816 -5189 -814 -5121
rect -800 -5189 -798 -5121
rect -790 -5189 -788 -5121
rect -782 -5189 -780 -5121
rect -772 -5189 -770 -5121
rect -756 -5189 -754 -5121
rect -748 -5189 -746 -5121
rect -732 -5189 -730 -5121
rect -716 -5189 -714 -5121
rect -708 -5189 -706 -5121
rect -698 -5189 -696 -5121
rect -572 -5189 -570 -5121
rect -562 -5189 -560 -5121
rect -546 -5189 -544 -5121
rect -536 -5189 -534 -5121
rect -520 -5189 -518 -5121
rect -510 -5189 -508 -5121
rect -502 -5189 -500 -5121
rect -492 -5189 -490 -5121
rect -476 -5189 -474 -5121
rect -468 -5189 -466 -5121
rect -458 -5189 -456 -5121
rect -442 -5189 -440 -5121
rect -432 -5189 -430 -5121
rect -424 -5189 -422 -5121
rect -414 -5189 -412 -5121
rect -398 -5189 -396 -5121
rect -390 -5189 -388 -5121
rect -374 -5189 -372 -5121
rect -358 -5189 -356 -5121
rect -350 -5189 -348 -5121
rect -340 -5189 -338 -5121
rect -214 -5189 -212 -5121
rect -204 -5189 -202 -5121
rect -188 -5189 -186 -5121
rect -178 -5189 -176 -5121
rect -162 -5189 -160 -5121
rect -152 -5189 -150 -5121
rect -144 -5189 -142 -5121
rect -134 -5189 -132 -5121
rect -118 -5189 -116 -5121
rect -110 -5189 -108 -5121
rect -100 -5189 -98 -5121
rect -84 -5189 -82 -5121
rect -74 -5189 -72 -5121
rect -66 -5189 -64 -5121
rect -56 -5189 -54 -5121
rect -40 -5189 -38 -5121
rect -32 -5189 -30 -5121
rect -16 -5189 -14 -5121
rect 0 -5189 2 -5121
rect 8 -5189 10 -5121
rect 18 -5189 20 -5121
rect 214 -5189 216 -5121
rect 224 -5189 226 -5121
rect 240 -5189 242 -5121
rect 250 -5189 252 -5121
rect 266 -5189 268 -5121
rect 276 -5189 278 -5121
rect 284 -5189 286 -5121
rect 294 -5189 296 -5121
rect 310 -5189 312 -5121
rect 318 -5189 320 -5121
rect 328 -5189 330 -5121
rect 344 -5189 346 -5121
rect 354 -5189 356 -5121
rect 362 -5189 364 -5121
rect 372 -5189 374 -5121
rect 388 -5189 390 -5121
rect 396 -5189 398 -5121
rect 412 -5189 414 -5121
rect 428 -5189 430 -5121
rect 436 -5189 438 -5121
rect 446 -5189 448 -5121
rect 570 -5189 572 -5121
rect 580 -5189 582 -5121
rect 596 -5189 598 -5121
rect 606 -5189 608 -5121
rect 622 -5189 624 -5121
rect 632 -5189 634 -5121
rect 640 -5189 642 -5121
rect 650 -5189 652 -5121
rect 666 -5189 668 -5121
rect 674 -5189 676 -5121
rect 684 -5189 686 -5121
rect 700 -5189 702 -5121
rect 710 -5189 712 -5121
rect 718 -5189 720 -5121
rect 728 -5189 730 -5121
rect 744 -5189 746 -5121
rect 752 -5189 754 -5121
rect 768 -5189 770 -5121
rect 784 -5189 786 -5121
rect 792 -5189 794 -5121
rect 802 -5189 804 -5121
rect 968 -5189 970 -5121
rect 978 -5189 980 -5121
rect 994 -5189 996 -5121
rect 1004 -5189 1006 -5121
rect 1020 -5189 1022 -5121
rect 1030 -5189 1032 -5121
rect 1038 -5189 1040 -5121
rect 1048 -5189 1050 -5121
rect 1064 -5189 1066 -5121
rect 1072 -5189 1074 -5121
rect 1082 -5189 1084 -5121
rect 1098 -5189 1100 -5121
rect 1108 -5189 1110 -5121
rect 1116 -5189 1118 -5121
rect 1126 -5189 1128 -5121
rect 1142 -5189 1144 -5121
rect 1150 -5189 1152 -5121
rect 1166 -5189 1168 -5121
rect 1182 -5189 1184 -5121
rect 1190 -5189 1192 -5121
rect 1200 -5189 1202 -5121
rect 1326 -5189 1328 -5121
rect 1336 -5189 1338 -5121
rect 1352 -5189 1354 -5121
rect 1362 -5189 1364 -5121
rect 1378 -5189 1380 -5121
rect 1388 -5189 1390 -5121
rect 1396 -5189 1398 -5121
rect 1406 -5189 1408 -5121
rect 1422 -5189 1424 -5121
rect 1430 -5189 1432 -5121
rect 1440 -5189 1442 -5121
rect 1456 -5189 1458 -5121
rect 1466 -5189 1468 -5121
rect 1474 -5189 1476 -5121
rect 1484 -5189 1486 -5121
rect 1500 -5189 1502 -5121
rect 1508 -5189 1510 -5121
rect 1524 -5189 1526 -5121
rect 1540 -5189 1542 -5121
rect 1548 -5189 1550 -5121
rect 1558 -5189 1560 -5121
rect -1259 -5195 -1257 -5193
rect -1249 -5195 -1247 -5193
rect -1233 -5195 -1231 -5193
rect -1223 -5195 -1221 -5193
rect -1215 -5195 -1213 -5193
rect -1205 -5195 -1203 -5193
rect -1189 -5195 -1187 -5193
rect -1181 -5195 -1179 -5193
rect -1171 -5195 -1169 -5193
rect -930 -5195 -928 -5193
rect -920 -5195 -918 -5193
rect -904 -5195 -902 -5193
rect -894 -5195 -892 -5193
rect -878 -5195 -876 -5193
rect -868 -5195 -866 -5193
rect -860 -5195 -858 -5193
rect -850 -5195 -848 -5193
rect -834 -5195 -832 -5193
rect -826 -5195 -824 -5193
rect -816 -5195 -814 -5193
rect -800 -5195 -798 -5193
rect -790 -5195 -788 -5193
rect -782 -5195 -780 -5193
rect -772 -5195 -770 -5193
rect -756 -5195 -754 -5193
rect -748 -5195 -746 -5193
rect -732 -5195 -730 -5193
rect -716 -5195 -714 -5193
rect -708 -5195 -706 -5193
rect -698 -5195 -696 -5193
rect -572 -5195 -570 -5193
rect -562 -5195 -560 -5193
rect -546 -5195 -544 -5193
rect -536 -5195 -534 -5193
rect -520 -5195 -518 -5193
rect -510 -5195 -508 -5193
rect -502 -5195 -500 -5193
rect -492 -5195 -490 -5193
rect -476 -5195 -474 -5193
rect -468 -5195 -466 -5193
rect -458 -5195 -456 -5193
rect -442 -5195 -440 -5193
rect -432 -5195 -430 -5193
rect -424 -5195 -422 -5193
rect -414 -5195 -412 -5193
rect -398 -5195 -396 -5193
rect -390 -5195 -388 -5193
rect -374 -5195 -372 -5193
rect -358 -5195 -356 -5193
rect -350 -5195 -348 -5193
rect -340 -5195 -338 -5193
rect -214 -5195 -212 -5193
rect -204 -5195 -202 -5193
rect -188 -5195 -186 -5193
rect -178 -5195 -176 -5193
rect -162 -5195 -160 -5193
rect -152 -5195 -150 -5193
rect -144 -5195 -142 -5193
rect -134 -5195 -132 -5193
rect -118 -5195 -116 -5193
rect -110 -5195 -108 -5193
rect -100 -5195 -98 -5193
rect -84 -5195 -82 -5193
rect -74 -5195 -72 -5193
rect -66 -5195 -64 -5193
rect -56 -5195 -54 -5193
rect -40 -5195 -38 -5193
rect -32 -5195 -30 -5193
rect -16 -5195 -14 -5193
rect 0 -5195 2 -5193
rect 8 -5195 10 -5193
rect 18 -5195 20 -5193
rect 214 -5195 216 -5193
rect 224 -5195 226 -5193
rect 240 -5195 242 -5193
rect 250 -5195 252 -5193
rect 266 -5195 268 -5193
rect 276 -5195 278 -5193
rect 284 -5195 286 -5193
rect 294 -5195 296 -5193
rect 310 -5195 312 -5193
rect 318 -5195 320 -5193
rect 328 -5195 330 -5193
rect 344 -5195 346 -5193
rect 354 -5195 356 -5193
rect 362 -5195 364 -5193
rect 372 -5195 374 -5193
rect 388 -5195 390 -5193
rect 396 -5195 398 -5193
rect 412 -5195 414 -5193
rect 428 -5195 430 -5193
rect 436 -5195 438 -5193
rect 446 -5195 448 -5193
rect 570 -5195 572 -5193
rect 580 -5195 582 -5193
rect 596 -5195 598 -5193
rect 606 -5195 608 -5193
rect 622 -5195 624 -5193
rect 632 -5195 634 -5193
rect 640 -5195 642 -5193
rect 650 -5195 652 -5193
rect 666 -5195 668 -5193
rect 674 -5195 676 -5193
rect 684 -5195 686 -5193
rect 700 -5195 702 -5193
rect 710 -5195 712 -5193
rect 718 -5195 720 -5193
rect 728 -5195 730 -5193
rect 744 -5195 746 -5193
rect 752 -5195 754 -5193
rect 768 -5195 770 -5193
rect 784 -5195 786 -5193
rect 792 -5195 794 -5193
rect 802 -5195 804 -5193
rect 968 -5195 970 -5193
rect 978 -5195 980 -5193
rect 994 -5195 996 -5193
rect 1004 -5195 1006 -5193
rect 1020 -5195 1022 -5193
rect 1030 -5195 1032 -5193
rect 1038 -5195 1040 -5193
rect 1048 -5195 1050 -5193
rect 1064 -5195 1066 -5193
rect 1072 -5195 1074 -5193
rect 1082 -5195 1084 -5193
rect 1098 -5195 1100 -5193
rect 1108 -5195 1110 -5193
rect 1116 -5195 1118 -5193
rect 1126 -5195 1128 -5193
rect 1142 -5195 1144 -5193
rect 1150 -5195 1152 -5193
rect 1166 -5195 1168 -5193
rect 1182 -5195 1184 -5193
rect 1190 -5195 1192 -5193
rect 1200 -5195 1202 -5193
rect 1326 -5195 1328 -5193
rect 1336 -5195 1338 -5193
rect 1352 -5195 1354 -5193
rect 1362 -5195 1364 -5193
rect 1378 -5195 1380 -5193
rect 1388 -5195 1390 -5193
rect 1396 -5195 1398 -5193
rect 1406 -5195 1408 -5193
rect 1422 -5195 1424 -5193
rect 1430 -5195 1432 -5193
rect 1440 -5195 1442 -5193
rect 1456 -5195 1458 -5193
rect 1466 -5195 1468 -5193
rect 1474 -5195 1476 -5193
rect 1484 -5195 1486 -5193
rect 1500 -5195 1502 -5193
rect 1508 -5195 1510 -5193
rect 1524 -5195 1526 -5193
rect 1540 -5195 1542 -5193
rect 1548 -5195 1550 -5193
rect 1558 -5195 1560 -5193
rect -1259 -5232 -1257 -5230
rect -1249 -5232 -1247 -5230
rect -1233 -5232 -1231 -5230
rect -1225 -5232 -1223 -5230
rect -1209 -5232 -1207 -5230
rect -1201 -5232 -1199 -5230
rect -1191 -5232 -1189 -5230
rect -1183 -5232 -1181 -5230
rect -1167 -5232 -1165 -5230
rect -1159 -5232 -1157 -5230
rect -1149 -5232 -1147 -5230
rect -1141 -5232 -1139 -5230
rect -1125 -5232 -1123 -5230
rect -1117 -5232 -1115 -5230
rect -1107 -5232 -1105 -5230
rect -1099 -5232 -1097 -5230
rect -1083 -5232 -1081 -5230
rect -1075 -5232 -1073 -5230
rect -930 -5232 -928 -5230
rect -920 -5232 -918 -5230
rect -904 -5232 -902 -5230
rect -896 -5232 -894 -5230
rect -880 -5232 -878 -5230
rect -872 -5232 -870 -5230
rect -862 -5232 -860 -5230
rect -854 -5232 -852 -5230
rect -838 -5232 -836 -5230
rect -830 -5232 -828 -5230
rect -820 -5232 -818 -5230
rect -812 -5232 -810 -5230
rect -796 -5232 -794 -5230
rect -788 -5232 -786 -5230
rect -778 -5232 -776 -5230
rect -770 -5232 -768 -5230
rect -754 -5232 -752 -5230
rect -746 -5232 -744 -5230
rect -1259 -5308 -1257 -5240
rect -1249 -5308 -1247 -5240
rect -1233 -5308 -1231 -5240
rect -1225 -5308 -1223 -5240
rect -1209 -5308 -1207 -5240
rect -1201 -5308 -1199 -5240
rect -1191 -5308 -1189 -5240
rect -1183 -5308 -1181 -5240
rect -1167 -5308 -1165 -5240
rect -1159 -5273 -1157 -5240
rect -1149 -5273 -1147 -5240
rect -1159 -5275 -1147 -5273
rect -1159 -5308 -1157 -5275
rect -1149 -5308 -1147 -5275
rect -1141 -5308 -1139 -5240
rect -1125 -5308 -1123 -5240
rect -1117 -5308 -1115 -5240
rect -1107 -5308 -1105 -5240
rect -1099 -5308 -1097 -5240
rect -1083 -5308 -1081 -5240
rect -1075 -5308 -1073 -5240
rect -930 -5308 -928 -5240
rect -920 -5308 -918 -5240
rect -904 -5308 -902 -5240
rect -896 -5308 -894 -5240
rect -880 -5308 -878 -5240
rect -872 -5308 -870 -5240
rect -862 -5308 -860 -5240
rect -854 -5308 -852 -5240
rect -838 -5308 -836 -5240
rect -830 -5273 -828 -5240
rect -820 -5273 -818 -5240
rect -830 -5275 -818 -5273
rect -830 -5308 -828 -5275
rect -820 -5308 -818 -5275
rect -812 -5308 -810 -5240
rect -796 -5308 -794 -5240
rect -788 -5308 -786 -5240
rect -778 -5308 -776 -5240
rect -770 -5308 -768 -5240
rect -754 -5308 -752 -5240
rect -746 -5308 -744 -5240
rect -1259 -5314 -1257 -5312
rect -1249 -5314 -1247 -5312
rect -1233 -5314 -1231 -5312
rect -1225 -5314 -1223 -5312
rect -1209 -5314 -1207 -5312
rect -1201 -5314 -1199 -5312
rect -1191 -5314 -1189 -5312
rect -1183 -5314 -1181 -5312
rect -1167 -5314 -1165 -5312
rect -1159 -5314 -1157 -5312
rect -1149 -5314 -1147 -5312
rect -1141 -5314 -1139 -5312
rect -1125 -5314 -1123 -5312
rect -1117 -5314 -1115 -5312
rect -1107 -5314 -1105 -5312
rect -1099 -5314 -1097 -5312
rect -1083 -5314 -1081 -5312
rect -1075 -5314 -1073 -5312
rect -930 -5314 -928 -5312
rect -920 -5314 -918 -5312
rect -904 -5314 -902 -5312
rect -896 -5314 -894 -5312
rect -880 -5314 -878 -5312
rect -872 -5314 -870 -5312
rect -862 -5314 -860 -5312
rect -854 -5314 -852 -5312
rect -838 -5314 -836 -5312
rect -830 -5314 -828 -5312
rect -820 -5314 -818 -5312
rect -812 -5314 -810 -5312
rect -796 -5314 -794 -5312
rect -788 -5314 -786 -5312
rect -778 -5314 -776 -5312
rect -770 -5314 -768 -5312
rect -754 -5314 -752 -5312
rect -746 -5314 -744 -5312
rect -1259 -5353 -1257 -5351
rect -1249 -5353 -1247 -5351
rect -1233 -5353 -1231 -5351
rect -1225 -5353 -1223 -5351
rect -1209 -5353 -1207 -5351
rect -1201 -5353 -1199 -5351
rect -1191 -5353 -1189 -5351
rect -1183 -5353 -1181 -5351
rect -1167 -5353 -1165 -5351
rect -1159 -5353 -1157 -5351
rect -1149 -5353 -1147 -5351
rect -1141 -5353 -1139 -5351
rect -1125 -5353 -1123 -5351
rect -1117 -5353 -1115 -5351
rect -1107 -5353 -1105 -5351
rect -1099 -5353 -1097 -5351
rect -1083 -5353 -1081 -5351
rect -1075 -5353 -1073 -5351
rect -1021 -5353 -1019 -5351
rect -930 -5353 -928 -5351
rect -920 -5353 -918 -5351
rect -904 -5353 -902 -5351
rect -896 -5353 -894 -5351
rect -880 -5353 -878 -5351
rect -872 -5353 -870 -5351
rect -862 -5353 -860 -5351
rect -854 -5353 -852 -5351
rect -838 -5353 -836 -5351
rect -830 -5353 -828 -5351
rect -820 -5353 -818 -5351
rect -812 -5353 -810 -5351
rect -796 -5353 -794 -5351
rect -788 -5353 -786 -5351
rect -778 -5353 -776 -5351
rect -770 -5353 -768 -5351
rect -754 -5353 -752 -5351
rect -746 -5353 -744 -5351
rect -668 -5353 -666 -5351
rect -572 -5353 -570 -5351
rect -562 -5353 -560 -5351
rect -546 -5353 -544 -5351
rect -538 -5353 -536 -5351
rect -522 -5353 -520 -5351
rect -514 -5353 -512 -5351
rect -504 -5353 -502 -5351
rect -496 -5353 -494 -5351
rect -480 -5353 -478 -5351
rect -472 -5353 -470 -5351
rect -462 -5353 -460 -5351
rect -454 -5353 -452 -5351
rect -438 -5353 -436 -5351
rect -430 -5353 -428 -5351
rect -420 -5353 -418 -5351
rect -412 -5353 -410 -5351
rect -396 -5353 -394 -5351
rect -388 -5353 -386 -5351
rect -322 -5353 -320 -5351
rect -214 -5353 -212 -5351
rect -204 -5353 -202 -5351
rect -188 -5353 -186 -5351
rect -180 -5353 -178 -5351
rect -164 -5353 -162 -5351
rect -156 -5353 -154 -5351
rect -146 -5353 -144 -5351
rect -138 -5353 -136 -5351
rect -122 -5353 -120 -5351
rect -114 -5353 -112 -5351
rect -104 -5353 -102 -5351
rect -96 -5353 -94 -5351
rect -80 -5353 -78 -5351
rect -72 -5353 -70 -5351
rect -62 -5353 -60 -5351
rect -54 -5353 -52 -5351
rect -38 -5353 -36 -5351
rect -30 -5353 -28 -5351
rect 214 -5353 216 -5351
rect 224 -5353 226 -5351
rect 240 -5353 242 -5351
rect 248 -5353 250 -5351
rect 264 -5353 266 -5351
rect 272 -5353 274 -5351
rect 282 -5353 284 -5351
rect 290 -5353 292 -5351
rect 306 -5353 308 -5351
rect 314 -5353 316 -5351
rect 324 -5353 326 -5351
rect 332 -5353 334 -5351
rect 348 -5353 350 -5351
rect 356 -5353 358 -5351
rect 366 -5353 368 -5351
rect 374 -5353 376 -5351
rect 390 -5353 392 -5351
rect 398 -5353 400 -5351
rect 471 -5353 473 -5351
rect 570 -5353 572 -5351
rect 580 -5353 582 -5351
rect 596 -5353 598 -5351
rect 604 -5353 606 -5351
rect 620 -5353 622 -5351
rect 628 -5353 630 -5351
rect 638 -5353 640 -5351
rect 646 -5353 648 -5351
rect 662 -5353 664 -5351
rect 670 -5353 672 -5351
rect 680 -5353 682 -5351
rect 688 -5353 690 -5351
rect 704 -5353 706 -5351
rect 712 -5353 714 -5351
rect 722 -5353 724 -5351
rect 730 -5353 732 -5351
rect 746 -5353 748 -5351
rect 754 -5353 756 -5351
rect 872 -5353 874 -5351
rect 968 -5353 970 -5351
rect 978 -5353 980 -5351
rect 994 -5353 996 -5351
rect 1002 -5353 1004 -5351
rect 1018 -5353 1020 -5351
rect 1026 -5353 1028 -5351
rect 1036 -5353 1038 -5351
rect 1044 -5353 1046 -5351
rect 1060 -5353 1062 -5351
rect 1068 -5353 1070 -5351
rect 1078 -5353 1080 -5351
rect 1086 -5353 1088 -5351
rect 1102 -5353 1104 -5351
rect 1110 -5353 1112 -5351
rect 1120 -5353 1122 -5351
rect 1128 -5353 1130 -5351
rect 1144 -5353 1146 -5351
rect 1152 -5353 1154 -5351
rect 1215 -5353 1217 -5351
rect 1326 -5353 1328 -5351
rect 1336 -5353 1338 -5351
rect 1352 -5353 1354 -5351
rect 1360 -5353 1362 -5351
rect 1376 -5353 1378 -5351
rect 1384 -5353 1386 -5351
rect 1394 -5353 1396 -5351
rect 1402 -5353 1404 -5351
rect 1418 -5353 1420 -5351
rect 1426 -5353 1428 -5351
rect 1436 -5353 1438 -5351
rect 1444 -5353 1446 -5351
rect 1460 -5353 1462 -5351
rect 1468 -5353 1470 -5351
rect 1478 -5353 1480 -5351
rect 1486 -5353 1488 -5351
rect 1502 -5353 1504 -5351
rect 1510 -5353 1512 -5351
rect -1259 -5429 -1257 -5361
rect -1249 -5429 -1247 -5361
rect -1233 -5429 -1231 -5361
rect -1225 -5429 -1223 -5361
rect -1209 -5429 -1207 -5361
rect -1201 -5429 -1199 -5361
rect -1191 -5429 -1189 -5361
rect -1183 -5429 -1181 -5361
rect -1167 -5429 -1165 -5361
rect -1159 -5394 -1157 -5361
rect -1149 -5394 -1147 -5361
rect -1159 -5396 -1147 -5394
rect -1159 -5429 -1157 -5396
rect -1149 -5429 -1147 -5396
rect -1141 -5429 -1139 -5361
rect -1125 -5429 -1123 -5361
rect -1117 -5429 -1115 -5361
rect -1107 -5429 -1105 -5361
rect -1099 -5429 -1097 -5361
rect -1083 -5429 -1081 -5361
rect -1075 -5429 -1073 -5361
rect -1021 -5429 -1019 -5361
rect -930 -5429 -928 -5361
rect -920 -5429 -918 -5361
rect -904 -5429 -902 -5361
rect -896 -5429 -894 -5361
rect -880 -5429 -878 -5361
rect -872 -5429 -870 -5361
rect -862 -5429 -860 -5361
rect -854 -5429 -852 -5361
rect -838 -5429 -836 -5361
rect -830 -5394 -828 -5361
rect -820 -5394 -818 -5361
rect -830 -5396 -818 -5394
rect -830 -5429 -828 -5396
rect -820 -5429 -818 -5396
rect -812 -5429 -810 -5361
rect -796 -5429 -794 -5361
rect -788 -5429 -786 -5361
rect -778 -5429 -776 -5361
rect -770 -5429 -768 -5361
rect -754 -5429 -752 -5361
rect -746 -5429 -744 -5361
rect -668 -5425 -666 -5369
rect -572 -5429 -570 -5361
rect -562 -5429 -560 -5361
rect -546 -5429 -544 -5361
rect -538 -5429 -536 -5361
rect -522 -5429 -520 -5361
rect -514 -5429 -512 -5361
rect -504 -5429 -502 -5361
rect -496 -5429 -494 -5361
rect -480 -5429 -478 -5361
rect -472 -5394 -470 -5361
rect -462 -5394 -460 -5361
rect -472 -5396 -460 -5394
rect -472 -5429 -470 -5396
rect -462 -5429 -460 -5396
rect -454 -5429 -452 -5361
rect -438 -5429 -436 -5361
rect -430 -5429 -428 -5361
rect -420 -5429 -418 -5361
rect -412 -5429 -410 -5361
rect -396 -5429 -394 -5361
rect -388 -5429 -386 -5361
rect -322 -5429 -320 -5361
rect -214 -5429 -212 -5361
rect -204 -5429 -202 -5361
rect -188 -5429 -186 -5361
rect -180 -5429 -178 -5361
rect -164 -5429 -162 -5361
rect -156 -5429 -154 -5361
rect -146 -5429 -144 -5361
rect -138 -5429 -136 -5361
rect -122 -5429 -120 -5361
rect -114 -5394 -112 -5361
rect -104 -5394 -102 -5361
rect -114 -5396 -102 -5394
rect -114 -5429 -112 -5396
rect -104 -5429 -102 -5396
rect -96 -5429 -94 -5361
rect -80 -5429 -78 -5361
rect -72 -5429 -70 -5361
rect -62 -5429 -60 -5361
rect -54 -5429 -52 -5361
rect -38 -5429 -36 -5361
rect -30 -5429 -28 -5361
rect 214 -5429 216 -5361
rect 224 -5429 226 -5361
rect 240 -5429 242 -5361
rect 248 -5429 250 -5361
rect 264 -5429 266 -5361
rect 272 -5429 274 -5361
rect 282 -5429 284 -5361
rect 290 -5429 292 -5361
rect 306 -5429 308 -5361
rect 314 -5394 316 -5361
rect 324 -5394 326 -5361
rect 314 -5396 326 -5394
rect 314 -5429 316 -5396
rect 324 -5429 326 -5396
rect 332 -5429 334 -5361
rect 348 -5429 350 -5361
rect 356 -5429 358 -5361
rect 366 -5429 368 -5361
rect 374 -5429 376 -5361
rect 390 -5429 392 -5361
rect 398 -5429 400 -5361
rect 471 -5429 473 -5361
rect 570 -5429 572 -5361
rect 580 -5429 582 -5361
rect 596 -5429 598 -5361
rect 604 -5429 606 -5361
rect 620 -5429 622 -5361
rect 628 -5429 630 -5361
rect 638 -5429 640 -5361
rect 646 -5429 648 -5361
rect 662 -5429 664 -5361
rect 670 -5394 672 -5361
rect 680 -5394 682 -5361
rect 670 -5396 682 -5394
rect 670 -5429 672 -5396
rect 680 -5429 682 -5396
rect 688 -5429 690 -5361
rect 704 -5429 706 -5361
rect 712 -5429 714 -5361
rect 722 -5429 724 -5361
rect 730 -5429 732 -5361
rect 746 -5429 748 -5361
rect 754 -5429 756 -5361
rect 872 -5425 874 -5369
rect 968 -5429 970 -5361
rect 978 -5429 980 -5361
rect 994 -5429 996 -5361
rect 1002 -5429 1004 -5361
rect 1018 -5429 1020 -5361
rect 1026 -5429 1028 -5361
rect 1036 -5429 1038 -5361
rect 1044 -5429 1046 -5361
rect 1060 -5429 1062 -5361
rect 1068 -5394 1070 -5361
rect 1078 -5394 1080 -5361
rect 1068 -5396 1080 -5394
rect 1068 -5429 1070 -5396
rect 1078 -5429 1080 -5396
rect 1086 -5429 1088 -5361
rect 1102 -5429 1104 -5361
rect 1110 -5429 1112 -5361
rect 1120 -5429 1122 -5361
rect 1128 -5429 1130 -5361
rect 1144 -5429 1146 -5361
rect 1152 -5429 1154 -5361
rect 1215 -5429 1217 -5361
rect 1326 -5429 1328 -5361
rect 1336 -5429 1338 -5361
rect 1352 -5429 1354 -5361
rect 1360 -5429 1362 -5361
rect 1376 -5429 1378 -5361
rect 1384 -5429 1386 -5361
rect 1394 -5429 1396 -5361
rect 1402 -5429 1404 -5361
rect 1418 -5429 1420 -5361
rect 1426 -5394 1428 -5361
rect 1436 -5394 1438 -5361
rect 1426 -5396 1438 -5394
rect 1426 -5429 1428 -5396
rect 1436 -5429 1438 -5396
rect 1444 -5429 1446 -5361
rect 1460 -5429 1462 -5361
rect 1468 -5429 1470 -5361
rect 1478 -5429 1480 -5361
rect 1486 -5429 1488 -5361
rect 1502 -5429 1504 -5361
rect 1510 -5429 1512 -5361
rect -1259 -5435 -1257 -5433
rect -1249 -5435 -1247 -5433
rect -1233 -5435 -1231 -5433
rect -1225 -5435 -1223 -5433
rect -1209 -5435 -1207 -5433
rect -1201 -5435 -1199 -5433
rect -1191 -5435 -1189 -5433
rect -1183 -5435 -1181 -5433
rect -1167 -5435 -1165 -5433
rect -1159 -5435 -1157 -5433
rect -1149 -5435 -1147 -5433
rect -1141 -5435 -1139 -5433
rect -1125 -5435 -1123 -5433
rect -1117 -5435 -1115 -5433
rect -1107 -5435 -1105 -5433
rect -1099 -5435 -1097 -5433
rect -1083 -5435 -1081 -5433
rect -1075 -5435 -1073 -5433
rect -1021 -5435 -1019 -5433
rect -930 -5435 -928 -5433
rect -920 -5435 -918 -5433
rect -904 -5435 -902 -5433
rect -896 -5435 -894 -5433
rect -880 -5435 -878 -5433
rect -872 -5435 -870 -5433
rect -862 -5435 -860 -5433
rect -854 -5435 -852 -5433
rect -838 -5435 -836 -5433
rect -830 -5435 -828 -5433
rect -820 -5435 -818 -5433
rect -812 -5435 -810 -5433
rect -796 -5435 -794 -5433
rect -788 -5435 -786 -5433
rect -778 -5435 -776 -5433
rect -770 -5435 -768 -5433
rect -754 -5435 -752 -5433
rect -746 -5435 -744 -5433
rect -668 -5435 -666 -5433
rect -572 -5435 -570 -5433
rect -562 -5435 -560 -5433
rect -546 -5435 -544 -5433
rect -538 -5435 -536 -5433
rect -522 -5435 -520 -5433
rect -514 -5435 -512 -5433
rect -504 -5435 -502 -5433
rect -496 -5435 -494 -5433
rect -480 -5435 -478 -5433
rect -472 -5435 -470 -5433
rect -462 -5435 -460 -5433
rect -454 -5435 -452 -5433
rect -438 -5435 -436 -5433
rect -430 -5435 -428 -5433
rect -420 -5435 -418 -5433
rect -412 -5435 -410 -5433
rect -396 -5435 -394 -5433
rect -388 -5435 -386 -5433
rect -322 -5435 -320 -5433
rect -214 -5435 -212 -5433
rect -204 -5435 -202 -5433
rect -188 -5435 -186 -5433
rect -180 -5435 -178 -5433
rect -164 -5435 -162 -5433
rect -156 -5435 -154 -5433
rect -146 -5435 -144 -5433
rect -138 -5435 -136 -5433
rect -122 -5435 -120 -5433
rect -114 -5435 -112 -5433
rect -104 -5435 -102 -5433
rect -96 -5435 -94 -5433
rect -80 -5435 -78 -5433
rect -72 -5435 -70 -5433
rect -62 -5435 -60 -5433
rect -54 -5435 -52 -5433
rect -38 -5435 -36 -5433
rect -30 -5435 -28 -5433
rect 214 -5435 216 -5433
rect 224 -5435 226 -5433
rect 240 -5435 242 -5433
rect 248 -5435 250 -5433
rect 264 -5435 266 -5433
rect 272 -5435 274 -5433
rect 282 -5435 284 -5433
rect 290 -5435 292 -5433
rect 306 -5435 308 -5433
rect 314 -5435 316 -5433
rect 324 -5435 326 -5433
rect 332 -5435 334 -5433
rect 348 -5435 350 -5433
rect 356 -5435 358 -5433
rect 366 -5435 368 -5433
rect 374 -5435 376 -5433
rect 390 -5435 392 -5433
rect 398 -5435 400 -5433
rect 471 -5435 473 -5433
rect 570 -5435 572 -5433
rect 580 -5435 582 -5433
rect 596 -5435 598 -5433
rect 604 -5435 606 -5433
rect 620 -5435 622 -5433
rect 628 -5435 630 -5433
rect 638 -5435 640 -5433
rect 646 -5435 648 -5433
rect 662 -5435 664 -5433
rect 670 -5435 672 -5433
rect 680 -5435 682 -5433
rect 688 -5435 690 -5433
rect 704 -5435 706 -5433
rect 712 -5435 714 -5433
rect 722 -5435 724 -5433
rect 730 -5435 732 -5433
rect 746 -5435 748 -5433
rect 754 -5435 756 -5433
rect 872 -5435 874 -5433
rect 968 -5435 970 -5433
rect 978 -5435 980 -5433
rect 994 -5435 996 -5433
rect 1002 -5435 1004 -5433
rect 1018 -5435 1020 -5433
rect 1026 -5435 1028 -5433
rect 1036 -5435 1038 -5433
rect 1044 -5435 1046 -5433
rect 1060 -5435 1062 -5433
rect 1068 -5435 1070 -5433
rect 1078 -5435 1080 -5433
rect 1086 -5435 1088 -5433
rect 1102 -5435 1104 -5433
rect 1110 -5435 1112 -5433
rect 1120 -5435 1122 -5433
rect 1128 -5435 1130 -5433
rect 1144 -5435 1146 -5433
rect 1152 -5435 1154 -5433
rect 1215 -5435 1217 -5433
rect 1326 -5435 1328 -5433
rect 1336 -5435 1338 -5433
rect 1352 -5435 1354 -5433
rect 1360 -5435 1362 -5433
rect 1376 -5435 1378 -5433
rect 1384 -5435 1386 -5433
rect 1394 -5435 1396 -5433
rect 1402 -5435 1404 -5433
rect 1418 -5435 1420 -5433
rect 1426 -5435 1428 -5433
rect 1436 -5435 1438 -5433
rect 1444 -5435 1446 -5433
rect 1460 -5435 1462 -5433
rect 1468 -5435 1470 -5433
rect 1478 -5435 1480 -5433
rect 1486 -5435 1488 -5433
rect 1502 -5435 1504 -5433
rect 1510 -5435 1512 -5433
rect -1259 -5473 -1257 -5471
rect -1249 -5473 -1247 -5471
rect -1233 -5473 -1231 -5471
rect -1225 -5473 -1223 -5471
rect -1209 -5473 -1207 -5471
rect -1201 -5473 -1199 -5471
rect -1191 -5473 -1189 -5471
rect -1183 -5473 -1181 -5471
rect -1167 -5473 -1165 -5471
rect -1159 -5473 -1157 -5471
rect -1149 -5473 -1147 -5471
rect -1141 -5473 -1139 -5471
rect -1125 -5473 -1123 -5471
rect -1117 -5473 -1115 -5471
rect -1107 -5473 -1105 -5471
rect -1099 -5473 -1097 -5471
rect -1083 -5473 -1081 -5471
rect -1075 -5473 -1073 -5471
rect -1021 -5473 -1019 -5471
rect -930 -5473 -928 -5471
rect -920 -5473 -918 -5471
rect -904 -5473 -902 -5471
rect -896 -5473 -894 -5471
rect -880 -5473 -878 -5471
rect -872 -5473 -870 -5471
rect -862 -5473 -860 -5471
rect -854 -5473 -852 -5471
rect -838 -5473 -836 -5471
rect -830 -5473 -828 -5471
rect -820 -5473 -818 -5471
rect -812 -5473 -810 -5471
rect -796 -5473 -794 -5471
rect -788 -5473 -786 -5471
rect -778 -5473 -776 -5471
rect -770 -5473 -768 -5471
rect -754 -5473 -752 -5471
rect -746 -5473 -744 -5471
rect -572 -5473 -570 -5471
rect -562 -5473 -560 -5471
rect -546 -5473 -544 -5471
rect -538 -5473 -536 -5471
rect -522 -5473 -520 -5471
rect -514 -5473 -512 -5471
rect -504 -5473 -502 -5471
rect -496 -5473 -494 -5471
rect -480 -5473 -478 -5471
rect -472 -5473 -470 -5471
rect -462 -5473 -460 -5471
rect -454 -5473 -452 -5471
rect -438 -5473 -436 -5471
rect -430 -5473 -428 -5471
rect -420 -5473 -418 -5471
rect -412 -5473 -410 -5471
rect -396 -5473 -394 -5471
rect -388 -5473 -386 -5471
rect -322 -5473 -320 -5471
rect -214 -5473 -212 -5471
rect -204 -5473 -202 -5471
rect -188 -5473 -186 -5471
rect -180 -5473 -178 -5471
rect -164 -5473 -162 -5471
rect -156 -5473 -154 -5471
rect -146 -5473 -144 -5471
rect -138 -5473 -136 -5471
rect -122 -5473 -120 -5471
rect -114 -5473 -112 -5471
rect -104 -5473 -102 -5471
rect -96 -5473 -94 -5471
rect -80 -5473 -78 -5471
rect -72 -5473 -70 -5471
rect -62 -5473 -60 -5471
rect -54 -5473 -52 -5471
rect -38 -5473 -36 -5471
rect -30 -5473 -28 -5471
rect 214 -5473 216 -5471
rect 224 -5473 226 -5471
rect 240 -5473 242 -5471
rect 248 -5473 250 -5471
rect 264 -5473 266 -5471
rect 272 -5473 274 -5471
rect 282 -5473 284 -5471
rect 290 -5473 292 -5471
rect 306 -5473 308 -5471
rect 314 -5473 316 -5471
rect 324 -5473 326 -5471
rect 332 -5473 334 -5471
rect 348 -5473 350 -5471
rect 356 -5473 358 -5471
rect 366 -5473 368 -5471
rect 374 -5473 376 -5471
rect 390 -5473 392 -5471
rect 398 -5473 400 -5471
rect 471 -5473 473 -5471
rect 570 -5473 572 -5471
rect 580 -5473 582 -5471
rect 596 -5473 598 -5471
rect 604 -5473 606 -5471
rect 620 -5473 622 -5471
rect 628 -5473 630 -5471
rect 638 -5473 640 -5471
rect 646 -5473 648 -5471
rect 662 -5473 664 -5471
rect 670 -5473 672 -5471
rect 680 -5473 682 -5471
rect 688 -5473 690 -5471
rect 704 -5473 706 -5471
rect 712 -5473 714 -5471
rect 722 -5473 724 -5471
rect 730 -5473 732 -5471
rect 746 -5473 748 -5471
rect 754 -5473 756 -5471
rect 968 -5473 970 -5471
rect 978 -5473 980 -5471
rect 994 -5473 996 -5471
rect 1002 -5473 1004 -5471
rect 1018 -5473 1020 -5471
rect 1026 -5473 1028 -5471
rect 1036 -5473 1038 -5471
rect 1044 -5473 1046 -5471
rect 1060 -5473 1062 -5471
rect 1068 -5473 1070 -5471
rect 1078 -5473 1080 -5471
rect 1086 -5473 1088 -5471
rect 1102 -5473 1104 -5471
rect 1110 -5473 1112 -5471
rect 1120 -5473 1122 -5471
rect 1128 -5473 1130 -5471
rect 1144 -5473 1146 -5471
rect 1152 -5473 1154 -5471
rect 1215 -5473 1217 -5471
rect 1326 -5473 1328 -5471
rect 1336 -5473 1338 -5471
rect 1352 -5473 1354 -5471
rect 1360 -5473 1362 -5471
rect 1376 -5473 1378 -5471
rect 1384 -5473 1386 -5471
rect 1394 -5473 1396 -5471
rect 1402 -5473 1404 -5471
rect 1418 -5473 1420 -5471
rect 1426 -5473 1428 -5471
rect 1436 -5473 1438 -5471
rect 1444 -5473 1446 -5471
rect 1460 -5473 1462 -5471
rect 1468 -5473 1470 -5471
rect 1478 -5473 1480 -5471
rect 1486 -5473 1488 -5471
rect 1502 -5473 1504 -5471
rect 1510 -5473 1512 -5471
rect -1259 -5549 -1257 -5481
rect -1249 -5549 -1247 -5481
rect -1233 -5549 -1231 -5481
rect -1225 -5549 -1223 -5481
rect -1209 -5549 -1207 -5481
rect -1201 -5549 -1199 -5481
rect -1191 -5549 -1189 -5481
rect -1183 -5549 -1181 -5481
rect -1167 -5549 -1165 -5481
rect -1159 -5514 -1157 -5481
rect -1149 -5514 -1147 -5481
rect -1159 -5516 -1147 -5514
rect -1159 -5549 -1157 -5516
rect -1149 -5549 -1147 -5516
rect -1141 -5549 -1139 -5481
rect -1125 -5549 -1123 -5481
rect -1117 -5549 -1115 -5481
rect -1107 -5549 -1105 -5481
rect -1099 -5549 -1097 -5481
rect -1083 -5549 -1081 -5481
rect -1075 -5549 -1073 -5481
rect -1021 -5549 -1019 -5481
rect -930 -5549 -928 -5481
rect -920 -5549 -918 -5481
rect -904 -5549 -902 -5481
rect -896 -5549 -894 -5481
rect -880 -5549 -878 -5481
rect -872 -5549 -870 -5481
rect -862 -5549 -860 -5481
rect -854 -5549 -852 -5481
rect -838 -5549 -836 -5481
rect -830 -5514 -828 -5481
rect -820 -5514 -818 -5481
rect -830 -5516 -818 -5514
rect -830 -5549 -828 -5516
rect -820 -5549 -818 -5516
rect -812 -5549 -810 -5481
rect -796 -5549 -794 -5481
rect -788 -5549 -786 -5481
rect -778 -5549 -776 -5481
rect -770 -5549 -768 -5481
rect -754 -5549 -752 -5481
rect -746 -5549 -744 -5481
rect -572 -5549 -570 -5481
rect -562 -5549 -560 -5481
rect -546 -5549 -544 -5481
rect -538 -5549 -536 -5481
rect -522 -5549 -520 -5481
rect -514 -5549 -512 -5481
rect -504 -5549 -502 -5481
rect -496 -5549 -494 -5481
rect -480 -5549 -478 -5481
rect -472 -5514 -470 -5481
rect -462 -5514 -460 -5481
rect -472 -5516 -460 -5514
rect -472 -5549 -470 -5516
rect -462 -5549 -460 -5516
rect -454 -5549 -452 -5481
rect -438 -5549 -436 -5481
rect -430 -5549 -428 -5481
rect -420 -5549 -418 -5481
rect -412 -5549 -410 -5481
rect -396 -5549 -394 -5481
rect -388 -5549 -386 -5481
rect -322 -5549 -320 -5481
rect -214 -5549 -212 -5481
rect -204 -5549 -202 -5481
rect -188 -5549 -186 -5481
rect -180 -5549 -178 -5481
rect -164 -5549 -162 -5481
rect -156 -5549 -154 -5481
rect -146 -5549 -144 -5481
rect -138 -5549 -136 -5481
rect -122 -5549 -120 -5481
rect -114 -5514 -112 -5481
rect -104 -5514 -102 -5481
rect -114 -5516 -102 -5514
rect -114 -5549 -112 -5516
rect -104 -5549 -102 -5516
rect -96 -5549 -94 -5481
rect -80 -5549 -78 -5481
rect -72 -5549 -70 -5481
rect -62 -5549 -60 -5481
rect -54 -5549 -52 -5481
rect -38 -5549 -36 -5481
rect -30 -5549 -28 -5481
rect 214 -5549 216 -5481
rect 224 -5549 226 -5481
rect 240 -5549 242 -5481
rect 248 -5549 250 -5481
rect 264 -5549 266 -5481
rect 272 -5549 274 -5481
rect 282 -5549 284 -5481
rect 290 -5549 292 -5481
rect 306 -5549 308 -5481
rect 314 -5514 316 -5481
rect 324 -5514 326 -5481
rect 314 -5516 326 -5514
rect 314 -5549 316 -5516
rect 324 -5549 326 -5516
rect 332 -5549 334 -5481
rect 348 -5549 350 -5481
rect 356 -5549 358 -5481
rect 366 -5549 368 -5481
rect 374 -5549 376 -5481
rect 390 -5549 392 -5481
rect 398 -5549 400 -5481
rect 471 -5549 473 -5481
rect 570 -5549 572 -5481
rect 580 -5549 582 -5481
rect 596 -5549 598 -5481
rect 604 -5549 606 -5481
rect 620 -5549 622 -5481
rect 628 -5549 630 -5481
rect 638 -5549 640 -5481
rect 646 -5549 648 -5481
rect 662 -5549 664 -5481
rect 670 -5514 672 -5481
rect 680 -5514 682 -5481
rect 670 -5516 682 -5514
rect 670 -5549 672 -5516
rect 680 -5549 682 -5516
rect 688 -5549 690 -5481
rect 704 -5549 706 -5481
rect 712 -5549 714 -5481
rect 722 -5549 724 -5481
rect 730 -5549 732 -5481
rect 746 -5549 748 -5481
rect 754 -5549 756 -5481
rect 968 -5549 970 -5481
rect 978 -5549 980 -5481
rect 994 -5549 996 -5481
rect 1002 -5549 1004 -5481
rect 1018 -5549 1020 -5481
rect 1026 -5549 1028 -5481
rect 1036 -5549 1038 -5481
rect 1044 -5549 1046 -5481
rect 1060 -5549 1062 -5481
rect 1068 -5514 1070 -5481
rect 1078 -5514 1080 -5481
rect 1068 -5516 1080 -5514
rect 1068 -5549 1070 -5516
rect 1078 -5549 1080 -5516
rect 1086 -5549 1088 -5481
rect 1102 -5549 1104 -5481
rect 1110 -5549 1112 -5481
rect 1120 -5549 1122 -5481
rect 1128 -5549 1130 -5481
rect 1144 -5549 1146 -5481
rect 1152 -5549 1154 -5481
rect 1215 -5549 1217 -5481
rect 1326 -5549 1328 -5481
rect 1336 -5549 1338 -5481
rect 1352 -5549 1354 -5481
rect 1360 -5549 1362 -5481
rect 1376 -5549 1378 -5481
rect 1384 -5549 1386 -5481
rect 1394 -5549 1396 -5481
rect 1402 -5549 1404 -5481
rect 1418 -5549 1420 -5481
rect 1426 -5514 1428 -5481
rect 1436 -5514 1438 -5481
rect 1426 -5516 1438 -5514
rect 1426 -5549 1428 -5516
rect 1436 -5549 1438 -5516
rect 1444 -5549 1446 -5481
rect 1460 -5549 1462 -5481
rect 1468 -5549 1470 -5481
rect 1478 -5549 1480 -5481
rect 1486 -5549 1488 -5481
rect 1502 -5549 1504 -5481
rect 1510 -5549 1512 -5481
rect -1259 -5555 -1257 -5553
rect -1249 -5555 -1247 -5553
rect -1233 -5555 -1231 -5553
rect -1225 -5555 -1223 -5553
rect -1209 -5555 -1207 -5553
rect -1201 -5555 -1199 -5553
rect -1191 -5555 -1189 -5553
rect -1183 -5555 -1181 -5553
rect -1167 -5555 -1165 -5553
rect -1159 -5555 -1157 -5553
rect -1149 -5555 -1147 -5553
rect -1141 -5555 -1139 -5553
rect -1125 -5555 -1123 -5553
rect -1117 -5555 -1115 -5553
rect -1107 -5555 -1105 -5553
rect -1099 -5555 -1097 -5553
rect -1083 -5555 -1081 -5553
rect -1075 -5555 -1073 -5553
rect -1021 -5555 -1019 -5553
rect -930 -5555 -928 -5553
rect -920 -5555 -918 -5553
rect -904 -5555 -902 -5553
rect -896 -5555 -894 -5553
rect -880 -5555 -878 -5553
rect -872 -5555 -870 -5553
rect -862 -5555 -860 -5553
rect -854 -5555 -852 -5553
rect -838 -5555 -836 -5553
rect -830 -5555 -828 -5553
rect -820 -5555 -818 -5553
rect -812 -5555 -810 -5553
rect -796 -5555 -794 -5553
rect -788 -5555 -786 -5553
rect -778 -5555 -776 -5553
rect -770 -5555 -768 -5553
rect -754 -5555 -752 -5553
rect -746 -5555 -744 -5553
rect -572 -5555 -570 -5553
rect -562 -5555 -560 -5553
rect -546 -5555 -544 -5553
rect -538 -5555 -536 -5553
rect -522 -5555 -520 -5553
rect -514 -5555 -512 -5553
rect -504 -5555 -502 -5553
rect -496 -5555 -494 -5553
rect -480 -5555 -478 -5553
rect -472 -5555 -470 -5553
rect -462 -5555 -460 -5553
rect -454 -5555 -452 -5553
rect -438 -5555 -436 -5553
rect -430 -5555 -428 -5553
rect -420 -5555 -418 -5553
rect -412 -5555 -410 -5553
rect -396 -5555 -394 -5553
rect -388 -5555 -386 -5553
rect -322 -5555 -320 -5553
rect -214 -5555 -212 -5553
rect -204 -5555 -202 -5553
rect -188 -5555 -186 -5553
rect -180 -5555 -178 -5553
rect -164 -5555 -162 -5553
rect -156 -5555 -154 -5553
rect -146 -5555 -144 -5553
rect -138 -5555 -136 -5553
rect -122 -5555 -120 -5553
rect -114 -5555 -112 -5553
rect -104 -5555 -102 -5553
rect -96 -5555 -94 -5553
rect -80 -5555 -78 -5553
rect -72 -5555 -70 -5553
rect -62 -5555 -60 -5553
rect -54 -5555 -52 -5553
rect -38 -5555 -36 -5553
rect -30 -5555 -28 -5553
rect 214 -5555 216 -5553
rect 224 -5555 226 -5553
rect 240 -5555 242 -5553
rect 248 -5555 250 -5553
rect 264 -5555 266 -5553
rect 272 -5555 274 -5553
rect 282 -5555 284 -5553
rect 290 -5555 292 -5553
rect 306 -5555 308 -5553
rect 314 -5555 316 -5553
rect 324 -5555 326 -5553
rect 332 -5555 334 -5553
rect 348 -5555 350 -5553
rect 356 -5555 358 -5553
rect 366 -5555 368 -5553
rect 374 -5555 376 -5553
rect 390 -5555 392 -5553
rect 398 -5555 400 -5553
rect 471 -5555 473 -5553
rect 570 -5555 572 -5553
rect 580 -5555 582 -5553
rect 596 -5555 598 -5553
rect 604 -5555 606 -5553
rect 620 -5555 622 -5553
rect 628 -5555 630 -5553
rect 638 -5555 640 -5553
rect 646 -5555 648 -5553
rect 662 -5555 664 -5553
rect 670 -5555 672 -5553
rect 680 -5555 682 -5553
rect 688 -5555 690 -5553
rect 704 -5555 706 -5553
rect 712 -5555 714 -5553
rect 722 -5555 724 -5553
rect 730 -5555 732 -5553
rect 746 -5555 748 -5553
rect 754 -5555 756 -5553
rect 968 -5555 970 -5553
rect 978 -5555 980 -5553
rect 994 -5555 996 -5553
rect 1002 -5555 1004 -5553
rect 1018 -5555 1020 -5553
rect 1026 -5555 1028 -5553
rect 1036 -5555 1038 -5553
rect 1044 -5555 1046 -5553
rect 1060 -5555 1062 -5553
rect 1068 -5555 1070 -5553
rect 1078 -5555 1080 -5553
rect 1086 -5555 1088 -5553
rect 1102 -5555 1104 -5553
rect 1110 -5555 1112 -5553
rect 1120 -5555 1122 -5553
rect 1128 -5555 1130 -5553
rect 1144 -5555 1146 -5553
rect 1152 -5555 1154 -5553
rect 1215 -5555 1217 -5553
rect 1326 -5555 1328 -5553
rect 1336 -5555 1338 -5553
rect 1352 -5555 1354 -5553
rect 1360 -5555 1362 -5553
rect 1376 -5555 1378 -5553
rect 1384 -5555 1386 -5553
rect 1394 -5555 1396 -5553
rect 1402 -5555 1404 -5553
rect 1418 -5555 1420 -5553
rect 1426 -5555 1428 -5553
rect 1436 -5555 1438 -5553
rect 1444 -5555 1446 -5553
rect 1460 -5555 1462 -5553
rect 1468 -5555 1470 -5553
rect 1478 -5555 1480 -5553
rect 1486 -5555 1488 -5553
rect 1502 -5555 1504 -5553
rect 1510 -5555 1512 -5553
rect -1259 -5590 -1257 -5588
rect -1249 -5590 -1247 -5588
rect -1233 -5590 -1231 -5588
rect -1225 -5590 -1223 -5588
rect -1209 -5590 -1207 -5588
rect -1201 -5590 -1199 -5588
rect -1191 -5590 -1189 -5588
rect -1183 -5590 -1181 -5588
rect -1167 -5590 -1165 -5588
rect -1159 -5590 -1157 -5588
rect -1149 -5590 -1147 -5588
rect -1141 -5590 -1139 -5588
rect -1125 -5590 -1123 -5588
rect -1117 -5590 -1115 -5588
rect -1107 -5590 -1105 -5588
rect -1099 -5590 -1097 -5588
rect -1083 -5590 -1081 -5588
rect -1075 -5590 -1073 -5588
rect -930 -5590 -928 -5588
rect -920 -5590 -918 -5588
rect -904 -5590 -902 -5588
rect -896 -5590 -894 -5588
rect -880 -5590 -878 -5588
rect -872 -5590 -870 -5588
rect -862 -5590 -860 -5588
rect -854 -5590 -852 -5588
rect -838 -5590 -836 -5588
rect -830 -5590 -828 -5588
rect -820 -5590 -818 -5588
rect -812 -5590 -810 -5588
rect -796 -5590 -794 -5588
rect -788 -5590 -786 -5588
rect -778 -5590 -776 -5588
rect -770 -5590 -768 -5588
rect -754 -5590 -752 -5588
rect -746 -5590 -744 -5588
rect -572 -5590 -570 -5588
rect -562 -5590 -560 -5588
rect -546 -5590 -544 -5588
rect -538 -5590 -536 -5588
rect -522 -5590 -520 -5588
rect -514 -5590 -512 -5588
rect -504 -5590 -502 -5588
rect -496 -5590 -494 -5588
rect -480 -5590 -478 -5588
rect -472 -5590 -470 -5588
rect -462 -5590 -460 -5588
rect -454 -5590 -452 -5588
rect -438 -5590 -436 -5588
rect -430 -5590 -428 -5588
rect -420 -5590 -418 -5588
rect -412 -5590 -410 -5588
rect -396 -5590 -394 -5588
rect -388 -5590 -386 -5588
rect -214 -5590 -212 -5588
rect -204 -5590 -202 -5588
rect -188 -5590 -186 -5588
rect -180 -5590 -178 -5588
rect -164 -5590 -162 -5588
rect -156 -5590 -154 -5588
rect -146 -5590 -144 -5588
rect -138 -5590 -136 -5588
rect -122 -5590 -120 -5588
rect -114 -5590 -112 -5588
rect -104 -5590 -102 -5588
rect -96 -5590 -94 -5588
rect -80 -5590 -78 -5588
rect -72 -5590 -70 -5588
rect -62 -5590 -60 -5588
rect -54 -5590 -52 -5588
rect -38 -5590 -36 -5588
rect -30 -5590 -28 -5588
rect 214 -5590 216 -5588
rect 224 -5590 226 -5588
rect 240 -5590 242 -5588
rect 248 -5590 250 -5588
rect 264 -5590 266 -5588
rect 272 -5590 274 -5588
rect 282 -5590 284 -5588
rect 290 -5590 292 -5588
rect 306 -5590 308 -5588
rect 314 -5590 316 -5588
rect 324 -5590 326 -5588
rect 332 -5590 334 -5588
rect 348 -5590 350 -5588
rect 356 -5590 358 -5588
rect 366 -5590 368 -5588
rect 374 -5590 376 -5588
rect 390 -5590 392 -5588
rect 398 -5590 400 -5588
rect 570 -5590 572 -5588
rect 580 -5590 582 -5588
rect 596 -5590 598 -5588
rect 604 -5590 606 -5588
rect 620 -5590 622 -5588
rect 628 -5590 630 -5588
rect 638 -5590 640 -5588
rect 646 -5590 648 -5588
rect 662 -5590 664 -5588
rect 670 -5590 672 -5588
rect 680 -5590 682 -5588
rect 688 -5590 690 -5588
rect 704 -5590 706 -5588
rect 712 -5590 714 -5588
rect 722 -5590 724 -5588
rect 730 -5590 732 -5588
rect 746 -5590 748 -5588
rect 754 -5590 756 -5588
rect -1259 -5666 -1257 -5598
rect -1249 -5666 -1247 -5598
rect -1233 -5666 -1231 -5598
rect -1225 -5666 -1223 -5598
rect -1209 -5666 -1207 -5598
rect -1201 -5666 -1199 -5598
rect -1191 -5666 -1189 -5598
rect -1183 -5666 -1181 -5598
rect -1167 -5666 -1165 -5598
rect -1159 -5631 -1157 -5598
rect -1149 -5631 -1147 -5598
rect -1159 -5633 -1147 -5631
rect -1159 -5666 -1157 -5633
rect -1149 -5666 -1147 -5633
rect -1141 -5666 -1139 -5598
rect -1125 -5666 -1123 -5598
rect -1117 -5666 -1115 -5598
rect -1107 -5666 -1105 -5598
rect -1099 -5666 -1097 -5598
rect -1083 -5666 -1081 -5598
rect -1075 -5666 -1073 -5598
rect -930 -5666 -928 -5598
rect -920 -5666 -918 -5598
rect -904 -5666 -902 -5598
rect -896 -5666 -894 -5598
rect -880 -5666 -878 -5598
rect -872 -5666 -870 -5598
rect -862 -5666 -860 -5598
rect -854 -5666 -852 -5598
rect -838 -5666 -836 -5598
rect -830 -5631 -828 -5598
rect -820 -5631 -818 -5598
rect -830 -5633 -818 -5631
rect -830 -5666 -828 -5633
rect -820 -5666 -818 -5633
rect -812 -5666 -810 -5598
rect -796 -5666 -794 -5598
rect -788 -5666 -786 -5598
rect -778 -5666 -776 -5598
rect -770 -5666 -768 -5598
rect -754 -5666 -752 -5598
rect -746 -5666 -744 -5598
rect -572 -5666 -570 -5598
rect -562 -5666 -560 -5598
rect -546 -5666 -544 -5598
rect -538 -5666 -536 -5598
rect -522 -5666 -520 -5598
rect -514 -5666 -512 -5598
rect -504 -5666 -502 -5598
rect -496 -5666 -494 -5598
rect -480 -5666 -478 -5598
rect -472 -5631 -470 -5598
rect -462 -5631 -460 -5598
rect -472 -5633 -460 -5631
rect -472 -5666 -470 -5633
rect -462 -5666 -460 -5633
rect -454 -5666 -452 -5598
rect -438 -5666 -436 -5598
rect -430 -5666 -428 -5598
rect -420 -5666 -418 -5598
rect -412 -5666 -410 -5598
rect -396 -5666 -394 -5598
rect -388 -5666 -386 -5598
rect -214 -5666 -212 -5598
rect -204 -5666 -202 -5598
rect -188 -5666 -186 -5598
rect -180 -5666 -178 -5598
rect -164 -5666 -162 -5598
rect -156 -5666 -154 -5598
rect -146 -5666 -144 -5598
rect -138 -5666 -136 -5598
rect -122 -5666 -120 -5598
rect -114 -5631 -112 -5598
rect -104 -5631 -102 -5598
rect -114 -5633 -102 -5631
rect -114 -5666 -112 -5633
rect -104 -5666 -102 -5633
rect -96 -5666 -94 -5598
rect -80 -5666 -78 -5598
rect -72 -5666 -70 -5598
rect -62 -5666 -60 -5598
rect -54 -5666 -52 -5598
rect -38 -5666 -36 -5598
rect -30 -5666 -28 -5598
rect 214 -5666 216 -5598
rect 224 -5666 226 -5598
rect 240 -5666 242 -5598
rect 248 -5666 250 -5598
rect 264 -5666 266 -5598
rect 272 -5666 274 -5598
rect 282 -5666 284 -5598
rect 290 -5666 292 -5598
rect 306 -5666 308 -5598
rect 314 -5631 316 -5598
rect 324 -5631 326 -5598
rect 314 -5633 326 -5631
rect 314 -5666 316 -5633
rect 324 -5666 326 -5633
rect 332 -5666 334 -5598
rect 348 -5666 350 -5598
rect 356 -5666 358 -5598
rect 366 -5666 368 -5598
rect 374 -5666 376 -5598
rect 390 -5666 392 -5598
rect 398 -5666 400 -5598
rect 570 -5666 572 -5598
rect 580 -5666 582 -5598
rect 596 -5666 598 -5598
rect 604 -5666 606 -5598
rect 620 -5666 622 -5598
rect 628 -5666 630 -5598
rect 638 -5666 640 -5598
rect 646 -5666 648 -5598
rect 662 -5666 664 -5598
rect 670 -5631 672 -5598
rect 680 -5631 682 -5598
rect 670 -5633 682 -5631
rect 670 -5666 672 -5633
rect 680 -5666 682 -5633
rect 688 -5666 690 -5598
rect 704 -5666 706 -5598
rect 712 -5666 714 -5598
rect 722 -5666 724 -5598
rect 730 -5666 732 -5598
rect 746 -5666 748 -5598
rect 754 -5666 756 -5598
rect -1259 -5672 -1257 -5670
rect -1249 -5672 -1247 -5670
rect -1233 -5672 -1231 -5670
rect -1225 -5672 -1223 -5670
rect -1209 -5672 -1207 -5670
rect -1201 -5672 -1199 -5670
rect -1191 -5672 -1189 -5670
rect -1183 -5672 -1181 -5670
rect -1167 -5672 -1165 -5670
rect -1159 -5672 -1157 -5670
rect -1149 -5672 -1147 -5670
rect -1141 -5672 -1139 -5670
rect -1125 -5672 -1123 -5670
rect -1117 -5672 -1115 -5670
rect -1107 -5672 -1105 -5670
rect -1099 -5672 -1097 -5670
rect -1083 -5672 -1081 -5670
rect -1075 -5672 -1073 -5670
rect -930 -5672 -928 -5670
rect -920 -5672 -918 -5670
rect -904 -5672 -902 -5670
rect -896 -5672 -894 -5670
rect -880 -5672 -878 -5670
rect -872 -5672 -870 -5670
rect -862 -5672 -860 -5670
rect -854 -5672 -852 -5670
rect -838 -5672 -836 -5670
rect -830 -5672 -828 -5670
rect -820 -5672 -818 -5670
rect -812 -5672 -810 -5670
rect -796 -5672 -794 -5670
rect -788 -5672 -786 -5670
rect -778 -5672 -776 -5670
rect -770 -5672 -768 -5670
rect -754 -5672 -752 -5670
rect -746 -5672 -744 -5670
rect -572 -5672 -570 -5670
rect -562 -5672 -560 -5670
rect -546 -5672 -544 -5670
rect -538 -5672 -536 -5670
rect -522 -5672 -520 -5670
rect -514 -5672 -512 -5670
rect -504 -5672 -502 -5670
rect -496 -5672 -494 -5670
rect -480 -5672 -478 -5670
rect -472 -5672 -470 -5670
rect -462 -5672 -460 -5670
rect -454 -5672 -452 -5670
rect -438 -5672 -436 -5670
rect -430 -5672 -428 -5670
rect -420 -5672 -418 -5670
rect -412 -5672 -410 -5670
rect -396 -5672 -394 -5670
rect -388 -5672 -386 -5670
rect -214 -5672 -212 -5670
rect -204 -5672 -202 -5670
rect -188 -5672 -186 -5670
rect -180 -5672 -178 -5670
rect -164 -5672 -162 -5670
rect -156 -5672 -154 -5670
rect -146 -5672 -144 -5670
rect -138 -5672 -136 -5670
rect -122 -5672 -120 -5670
rect -114 -5672 -112 -5670
rect -104 -5672 -102 -5670
rect -96 -5672 -94 -5670
rect -80 -5672 -78 -5670
rect -72 -5672 -70 -5670
rect -62 -5672 -60 -5670
rect -54 -5672 -52 -5670
rect -38 -5672 -36 -5670
rect -30 -5672 -28 -5670
rect 214 -5672 216 -5670
rect 224 -5672 226 -5670
rect 240 -5672 242 -5670
rect 248 -5672 250 -5670
rect 264 -5672 266 -5670
rect 272 -5672 274 -5670
rect 282 -5672 284 -5670
rect 290 -5672 292 -5670
rect 306 -5672 308 -5670
rect 314 -5672 316 -5670
rect 324 -5672 326 -5670
rect 332 -5672 334 -5670
rect 348 -5672 350 -5670
rect 356 -5672 358 -5670
rect 366 -5672 368 -5670
rect 374 -5672 376 -5670
rect 390 -5672 392 -5670
rect 398 -5672 400 -5670
rect 570 -5672 572 -5670
rect 580 -5672 582 -5670
rect 596 -5672 598 -5670
rect 604 -5672 606 -5670
rect 620 -5672 622 -5670
rect 628 -5672 630 -5670
rect 638 -5672 640 -5670
rect 646 -5672 648 -5670
rect 662 -5672 664 -5670
rect 670 -5672 672 -5670
rect 680 -5672 682 -5670
rect 688 -5672 690 -5670
rect 704 -5672 706 -5670
rect 712 -5672 714 -5670
rect 722 -5672 724 -5670
rect 730 -5672 732 -5670
rect 746 -5672 748 -5670
rect 754 -5672 756 -5670
rect -1334 -5707 -1332 -5705
rect -1326 -5707 -1324 -5705
rect -1316 -5707 -1314 -5705
rect -930 -5707 -928 -5705
rect -922 -5707 -920 -5705
rect -912 -5707 -910 -5705
rect -572 -5707 -570 -5705
rect -564 -5707 -562 -5705
rect -554 -5707 -552 -5705
rect -214 -5707 -212 -5705
rect -206 -5707 -204 -5705
rect -196 -5707 -194 -5705
rect 214 -5707 216 -5705
rect 222 -5707 224 -5705
rect 232 -5707 234 -5705
rect 570 -5707 572 -5705
rect 578 -5707 580 -5705
rect 588 -5707 590 -5705
rect 968 -5707 970 -5705
rect 976 -5707 978 -5705
rect 986 -5707 988 -5705
rect 1326 -5707 1328 -5705
rect 1334 -5707 1336 -5705
rect 1344 -5707 1346 -5705
rect -1334 -5783 -1332 -5715
rect -1326 -5739 -1324 -5715
rect -1326 -5783 -1324 -5743
rect -1316 -5783 -1314 -5715
rect -930 -5783 -928 -5715
rect -922 -5739 -920 -5715
rect -922 -5783 -920 -5743
rect -912 -5783 -910 -5715
rect -572 -5783 -570 -5715
rect -564 -5739 -562 -5715
rect -564 -5783 -562 -5743
rect -554 -5783 -552 -5715
rect -214 -5783 -212 -5715
rect -206 -5739 -204 -5715
rect -206 -5783 -204 -5743
rect -196 -5783 -194 -5715
rect 214 -5783 216 -5715
rect 222 -5739 224 -5715
rect 222 -5783 224 -5743
rect 232 -5783 234 -5715
rect 570 -5783 572 -5715
rect 578 -5739 580 -5715
rect 578 -5783 580 -5743
rect 588 -5783 590 -5715
rect 968 -5783 970 -5715
rect 976 -5739 978 -5715
rect 976 -5783 978 -5743
rect 986 -5783 988 -5715
rect 1326 -5783 1328 -5715
rect 1334 -5739 1336 -5715
rect 1334 -5783 1336 -5743
rect 1344 -5783 1346 -5715
rect -1334 -5789 -1332 -5787
rect -1326 -5789 -1324 -5787
rect -1316 -5789 -1314 -5787
rect -930 -5789 -928 -5787
rect -922 -5789 -920 -5787
rect -912 -5789 -910 -5787
rect -572 -5789 -570 -5787
rect -564 -5789 -562 -5787
rect -554 -5789 -552 -5787
rect -214 -5789 -212 -5787
rect -206 -5789 -204 -5787
rect -196 -5789 -194 -5787
rect 214 -5789 216 -5787
rect 222 -5789 224 -5787
rect 232 -5789 234 -5787
rect 570 -5789 572 -5787
rect 578 -5789 580 -5787
rect 588 -5789 590 -5787
rect 968 -5789 970 -5787
rect 976 -5789 978 -5787
rect 986 -5789 988 -5787
rect 1326 -5789 1328 -5787
rect 1334 -5789 1336 -5787
rect 1344 -5789 1346 -5787
rect -1259 -5826 -1257 -5824
rect -1249 -5826 -1247 -5824
rect -1233 -5826 -1231 -5824
rect -1223 -5826 -1221 -5824
rect -1215 -5826 -1213 -5824
rect -1205 -5826 -1203 -5824
rect -1189 -5826 -1187 -5824
rect -1181 -5826 -1179 -5824
rect -1171 -5826 -1169 -5824
rect -930 -5826 -928 -5824
rect -920 -5826 -918 -5824
rect -904 -5826 -902 -5824
rect -894 -5826 -892 -5824
rect -878 -5826 -876 -5824
rect -868 -5826 -866 -5824
rect -860 -5826 -858 -5824
rect -850 -5826 -848 -5824
rect -834 -5826 -832 -5824
rect -826 -5826 -824 -5824
rect -816 -5826 -814 -5824
rect -800 -5826 -798 -5824
rect -790 -5826 -788 -5824
rect -782 -5826 -780 -5824
rect -772 -5826 -770 -5824
rect -756 -5826 -754 -5824
rect -748 -5826 -746 -5824
rect -732 -5826 -730 -5824
rect -716 -5826 -714 -5824
rect -708 -5826 -706 -5824
rect -698 -5826 -696 -5824
rect -572 -5826 -570 -5824
rect -562 -5826 -560 -5824
rect -546 -5826 -544 -5824
rect -536 -5826 -534 -5824
rect -520 -5826 -518 -5824
rect -510 -5826 -508 -5824
rect -502 -5826 -500 -5824
rect -492 -5826 -490 -5824
rect -476 -5826 -474 -5824
rect -468 -5826 -466 -5824
rect -458 -5826 -456 -5824
rect -442 -5826 -440 -5824
rect -432 -5826 -430 -5824
rect -424 -5826 -422 -5824
rect -414 -5826 -412 -5824
rect -398 -5826 -396 -5824
rect -390 -5826 -388 -5824
rect -374 -5826 -372 -5824
rect -358 -5826 -356 -5824
rect -350 -5826 -348 -5824
rect -340 -5826 -338 -5824
rect -214 -5826 -212 -5824
rect -204 -5826 -202 -5824
rect -188 -5826 -186 -5824
rect -178 -5826 -176 -5824
rect -162 -5826 -160 -5824
rect -152 -5826 -150 -5824
rect -144 -5826 -142 -5824
rect -134 -5826 -132 -5824
rect -118 -5826 -116 -5824
rect -110 -5826 -108 -5824
rect -100 -5826 -98 -5824
rect -84 -5826 -82 -5824
rect -74 -5826 -72 -5824
rect -66 -5826 -64 -5824
rect -56 -5826 -54 -5824
rect -40 -5826 -38 -5824
rect -32 -5826 -30 -5824
rect -16 -5826 -14 -5824
rect 0 -5826 2 -5824
rect 8 -5826 10 -5824
rect 18 -5826 20 -5824
rect 214 -5826 216 -5824
rect 224 -5826 226 -5824
rect 240 -5826 242 -5824
rect 250 -5826 252 -5824
rect 266 -5826 268 -5824
rect 276 -5826 278 -5824
rect 284 -5826 286 -5824
rect 294 -5826 296 -5824
rect 310 -5826 312 -5824
rect 318 -5826 320 -5824
rect 328 -5826 330 -5824
rect 344 -5826 346 -5824
rect 354 -5826 356 -5824
rect 362 -5826 364 -5824
rect 372 -5826 374 -5824
rect 388 -5826 390 -5824
rect 396 -5826 398 -5824
rect 412 -5826 414 -5824
rect 428 -5826 430 -5824
rect 436 -5826 438 -5824
rect 446 -5826 448 -5824
rect 570 -5826 572 -5824
rect 580 -5826 582 -5824
rect 596 -5826 598 -5824
rect 606 -5826 608 -5824
rect 622 -5826 624 -5824
rect 632 -5826 634 -5824
rect 640 -5826 642 -5824
rect 650 -5826 652 -5824
rect 666 -5826 668 -5824
rect 674 -5826 676 -5824
rect 684 -5826 686 -5824
rect 700 -5826 702 -5824
rect 710 -5826 712 -5824
rect 718 -5826 720 -5824
rect 728 -5826 730 -5824
rect 744 -5826 746 -5824
rect 752 -5826 754 -5824
rect 768 -5826 770 -5824
rect 784 -5826 786 -5824
rect 792 -5826 794 -5824
rect 802 -5826 804 -5824
rect 968 -5826 970 -5824
rect 978 -5826 980 -5824
rect 994 -5826 996 -5824
rect 1004 -5826 1006 -5824
rect 1020 -5826 1022 -5824
rect 1030 -5826 1032 -5824
rect 1038 -5826 1040 -5824
rect 1048 -5826 1050 -5824
rect 1064 -5826 1066 -5824
rect 1072 -5826 1074 -5824
rect 1082 -5826 1084 -5824
rect 1098 -5826 1100 -5824
rect 1108 -5826 1110 -5824
rect 1116 -5826 1118 -5824
rect 1126 -5826 1128 -5824
rect 1142 -5826 1144 -5824
rect 1150 -5826 1152 -5824
rect 1166 -5826 1168 -5824
rect 1182 -5826 1184 -5824
rect 1190 -5826 1192 -5824
rect 1200 -5826 1202 -5824
rect 1326 -5826 1328 -5824
rect 1336 -5826 1338 -5824
rect 1352 -5826 1354 -5824
rect 1362 -5826 1364 -5824
rect 1378 -5826 1380 -5824
rect 1388 -5826 1390 -5824
rect 1396 -5826 1398 -5824
rect 1406 -5826 1408 -5824
rect 1422 -5826 1424 -5824
rect 1430 -5826 1432 -5824
rect 1440 -5826 1442 -5824
rect 1456 -5826 1458 -5824
rect 1466 -5826 1468 -5824
rect 1474 -5826 1476 -5824
rect 1484 -5826 1486 -5824
rect 1500 -5826 1502 -5824
rect 1508 -5826 1510 -5824
rect 1524 -5826 1526 -5824
rect 1540 -5826 1542 -5824
rect 1548 -5826 1550 -5824
rect 1558 -5826 1560 -5824
rect -1259 -5902 -1257 -5834
rect -1249 -5902 -1247 -5834
rect -1233 -5902 -1231 -5834
rect -1223 -5902 -1221 -5834
rect -1215 -5902 -1213 -5834
rect -1205 -5902 -1203 -5834
rect -1189 -5902 -1187 -5834
rect -1181 -5902 -1179 -5834
rect -1171 -5902 -1169 -5834
rect -930 -5902 -928 -5834
rect -920 -5902 -918 -5834
rect -904 -5902 -902 -5834
rect -894 -5902 -892 -5834
rect -878 -5902 -876 -5834
rect -868 -5902 -866 -5834
rect -860 -5902 -858 -5834
rect -850 -5902 -848 -5834
rect -834 -5902 -832 -5834
rect -826 -5902 -824 -5834
rect -816 -5902 -814 -5834
rect -800 -5902 -798 -5834
rect -790 -5902 -788 -5834
rect -782 -5902 -780 -5834
rect -772 -5902 -770 -5834
rect -756 -5902 -754 -5834
rect -748 -5902 -746 -5834
rect -732 -5902 -730 -5834
rect -716 -5902 -714 -5834
rect -708 -5902 -706 -5834
rect -698 -5902 -696 -5834
rect -572 -5902 -570 -5834
rect -562 -5902 -560 -5834
rect -546 -5902 -544 -5834
rect -536 -5902 -534 -5834
rect -520 -5902 -518 -5834
rect -510 -5902 -508 -5834
rect -502 -5902 -500 -5834
rect -492 -5902 -490 -5834
rect -476 -5902 -474 -5834
rect -468 -5902 -466 -5834
rect -458 -5902 -456 -5834
rect -442 -5902 -440 -5834
rect -432 -5902 -430 -5834
rect -424 -5902 -422 -5834
rect -414 -5902 -412 -5834
rect -398 -5902 -396 -5834
rect -390 -5902 -388 -5834
rect -374 -5902 -372 -5834
rect -358 -5902 -356 -5834
rect -350 -5902 -348 -5834
rect -340 -5902 -338 -5834
rect -214 -5902 -212 -5834
rect -204 -5902 -202 -5834
rect -188 -5902 -186 -5834
rect -178 -5902 -176 -5834
rect -162 -5902 -160 -5834
rect -152 -5902 -150 -5834
rect -144 -5902 -142 -5834
rect -134 -5902 -132 -5834
rect -118 -5902 -116 -5834
rect -110 -5902 -108 -5834
rect -100 -5902 -98 -5834
rect -84 -5902 -82 -5834
rect -74 -5902 -72 -5834
rect -66 -5902 -64 -5834
rect -56 -5902 -54 -5834
rect -40 -5902 -38 -5834
rect -32 -5902 -30 -5834
rect -16 -5902 -14 -5834
rect 0 -5902 2 -5834
rect 8 -5902 10 -5834
rect 18 -5902 20 -5834
rect 214 -5902 216 -5834
rect 224 -5902 226 -5834
rect 240 -5902 242 -5834
rect 250 -5902 252 -5834
rect 266 -5902 268 -5834
rect 276 -5902 278 -5834
rect 284 -5902 286 -5834
rect 294 -5902 296 -5834
rect 310 -5902 312 -5834
rect 318 -5902 320 -5834
rect 328 -5902 330 -5834
rect 344 -5902 346 -5834
rect 354 -5902 356 -5834
rect 362 -5902 364 -5834
rect 372 -5902 374 -5834
rect 388 -5902 390 -5834
rect 396 -5902 398 -5834
rect 412 -5902 414 -5834
rect 428 -5902 430 -5834
rect 436 -5902 438 -5834
rect 446 -5902 448 -5834
rect 570 -5902 572 -5834
rect 580 -5902 582 -5834
rect 596 -5902 598 -5834
rect 606 -5902 608 -5834
rect 622 -5902 624 -5834
rect 632 -5902 634 -5834
rect 640 -5902 642 -5834
rect 650 -5902 652 -5834
rect 666 -5902 668 -5834
rect 674 -5902 676 -5834
rect 684 -5902 686 -5834
rect 700 -5902 702 -5834
rect 710 -5902 712 -5834
rect 718 -5902 720 -5834
rect 728 -5902 730 -5834
rect 744 -5902 746 -5834
rect 752 -5902 754 -5834
rect 768 -5902 770 -5834
rect 784 -5902 786 -5834
rect 792 -5902 794 -5834
rect 802 -5902 804 -5834
rect 968 -5902 970 -5834
rect 978 -5902 980 -5834
rect 994 -5902 996 -5834
rect 1004 -5902 1006 -5834
rect 1020 -5902 1022 -5834
rect 1030 -5902 1032 -5834
rect 1038 -5902 1040 -5834
rect 1048 -5902 1050 -5834
rect 1064 -5902 1066 -5834
rect 1072 -5902 1074 -5834
rect 1082 -5902 1084 -5834
rect 1098 -5902 1100 -5834
rect 1108 -5902 1110 -5834
rect 1116 -5902 1118 -5834
rect 1126 -5902 1128 -5834
rect 1142 -5902 1144 -5834
rect 1150 -5902 1152 -5834
rect 1166 -5902 1168 -5834
rect 1182 -5902 1184 -5834
rect 1190 -5902 1192 -5834
rect 1200 -5902 1202 -5834
rect 1326 -5902 1328 -5834
rect 1336 -5902 1338 -5834
rect 1352 -5902 1354 -5834
rect 1362 -5902 1364 -5834
rect 1378 -5902 1380 -5834
rect 1388 -5902 1390 -5834
rect 1396 -5902 1398 -5834
rect 1406 -5902 1408 -5834
rect 1422 -5902 1424 -5834
rect 1430 -5902 1432 -5834
rect 1440 -5902 1442 -5834
rect 1456 -5902 1458 -5834
rect 1466 -5902 1468 -5834
rect 1474 -5902 1476 -5834
rect 1484 -5902 1486 -5834
rect 1500 -5902 1502 -5834
rect 1508 -5902 1510 -5834
rect 1524 -5902 1526 -5834
rect 1540 -5902 1542 -5834
rect 1548 -5902 1550 -5834
rect 1558 -5902 1560 -5834
rect -1259 -5908 -1257 -5906
rect -1249 -5908 -1247 -5906
rect -1233 -5908 -1231 -5906
rect -1223 -5908 -1221 -5906
rect -1215 -5908 -1213 -5906
rect -1205 -5908 -1203 -5906
rect -1189 -5908 -1187 -5906
rect -1181 -5908 -1179 -5906
rect -1171 -5908 -1169 -5906
rect -930 -5908 -928 -5906
rect -920 -5908 -918 -5906
rect -904 -5908 -902 -5906
rect -894 -5908 -892 -5906
rect -878 -5908 -876 -5906
rect -868 -5908 -866 -5906
rect -860 -5908 -858 -5906
rect -850 -5908 -848 -5906
rect -834 -5908 -832 -5906
rect -826 -5908 -824 -5906
rect -816 -5908 -814 -5906
rect -800 -5908 -798 -5906
rect -790 -5908 -788 -5906
rect -782 -5908 -780 -5906
rect -772 -5908 -770 -5906
rect -756 -5908 -754 -5906
rect -748 -5908 -746 -5906
rect -732 -5908 -730 -5906
rect -716 -5908 -714 -5906
rect -708 -5908 -706 -5906
rect -698 -5908 -696 -5906
rect -572 -5908 -570 -5906
rect -562 -5908 -560 -5906
rect -546 -5908 -544 -5906
rect -536 -5908 -534 -5906
rect -520 -5908 -518 -5906
rect -510 -5908 -508 -5906
rect -502 -5908 -500 -5906
rect -492 -5908 -490 -5906
rect -476 -5908 -474 -5906
rect -468 -5908 -466 -5906
rect -458 -5908 -456 -5906
rect -442 -5908 -440 -5906
rect -432 -5908 -430 -5906
rect -424 -5908 -422 -5906
rect -414 -5908 -412 -5906
rect -398 -5908 -396 -5906
rect -390 -5908 -388 -5906
rect -374 -5908 -372 -5906
rect -358 -5908 -356 -5906
rect -350 -5908 -348 -5906
rect -340 -5908 -338 -5906
rect -214 -5908 -212 -5906
rect -204 -5908 -202 -5906
rect -188 -5908 -186 -5906
rect -178 -5908 -176 -5906
rect -162 -5908 -160 -5906
rect -152 -5908 -150 -5906
rect -144 -5908 -142 -5906
rect -134 -5908 -132 -5906
rect -118 -5908 -116 -5906
rect -110 -5908 -108 -5906
rect -100 -5908 -98 -5906
rect -84 -5908 -82 -5906
rect -74 -5908 -72 -5906
rect -66 -5908 -64 -5906
rect -56 -5908 -54 -5906
rect -40 -5908 -38 -5906
rect -32 -5908 -30 -5906
rect -16 -5908 -14 -5906
rect 0 -5908 2 -5906
rect 8 -5908 10 -5906
rect 18 -5908 20 -5906
rect 214 -5908 216 -5906
rect 224 -5908 226 -5906
rect 240 -5908 242 -5906
rect 250 -5908 252 -5906
rect 266 -5908 268 -5906
rect 276 -5908 278 -5906
rect 284 -5908 286 -5906
rect 294 -5908 296 -5906
rect 310 -5908 312 -5906
rect 318 -5908 320 -5906
rect 328 -5908 330 -5906
rect 344 -5908 346 -5906
rect 354 -5908 356 -5906
rect 362 -5908 364 -5906
rect 372 -5908 374 -5906
rect 388 -5908 390 -5906
rect 396 -5908 398 -5906
rect 412 -5908 414 -5906
rect 428 -5908 430 -5906
rect 436 -5908 438 -5906
rect 446 -5908 448 -5906
rect 570 -5908 572 -5906
rect 580 -5908 582 -5906
rect 596 -5908 598 -5906
rect 606 -5908 608 -5906
rect 622 -5908 624 -5906
rect 632 -5908 634 -5906
rect 640 -5908 642 -5906
rect 650 -5908 652 -5906
rect 666 -5908 668 -5906
rect 674 -5908 676 -5906
rect 684 -5908 686 -5906
rect 700 -5908 702 -5906
rect 710 -5908 712 -5906
rect 718 -5908 720 -5906
rect 728 -5908 730 -5906
rect 744 -5908 746 -5906
rect 752 -5908 754 -5906
rect 768 -5908 770 -5906
rect 784 -5908 786 -5906
rect 792 -5908 794 -5906
rect 802 -5908 804 -5906
rect 968 -5908 970 -5906
rect 978 -5908 980 -5906
rect 994 -5908 996 -5906
rect 1004 -5908 1006 -5906
rect 1020 -5908 1022 -5906
rect 1030 -5908 1032 -5906
rect 1038 -5908 1040 -5906
rect 1048 -5908 1050 -5906
rect 1064 -5908 1066 -5906
rect 1072 -5908 1074 -5906
rect 1082 -5908 1084 -5906
rect 1098 -5908 1100 -5906
rect 1108 -5908 1110 -5906
rect 1116 -5908 1118 -5906
rect 1126 -5908 1128 -5906
rect 1142 -5908 1144 -5906
rect 1150 -5908 1152 -5906
rect 1166 -5908 1168 -5906
rect 1182 -5908 1184 -5906
rect 1190 -5908 1192 -5906
rect 1200 -5908 1202 -5906
rect 1326 -5908 1328 -5906
rect 1336 -5908 1338 -5906
rect 1352 -5908 1354 -5906
rect 1362 -5908 1364 -5906
rect 1378 -5908 1380 -5906
rect 1388 -5908 1390 -5906
rect 1396 -5908 1398 -5906
rect 1406 -5908 1408 -5906
rect 1422 -5908 1424 -5906
rect 1430 -5908 1432 -5906
rect 1440 -5908 1442 -5906
rect 1456 -5908 1458 -5906
rect 1466 -5908 1468 -5906
rect 1474 -5908 1476 -5906
rect 1484 -5908 1486 -5906
rect 1500 -5908 1502 -5906
rect 1508 -5908 1510 -5906
rect 1524 -5908 1526 -5906
rect 1540 -5908 1542 -5906
rect 1548 -5908 1550 -5906
rect 1558 -5908 1560 -5906
rect -1259 -5949 -1257 -5947
rect -1249 -5949 -1247 -5947
rect -1233 -5949 -1231 -5947
rect -1225 -5949 -1223 -5947
rect -1209 -5949 -1207 -5947
rect -1201 -5949 -1199 -5947
rect -1191 -5949 -1189 -5947
rect -1183 -5949 -1181 -5947
rect -1167 -5949 -1165 -5947
rect -1159 -5949 -1157 -5947
rect -1149 -5949 -1147 -5947
rect -1141 -5949 -1139 -5947
rect -1125 -5949 -1123 -5947
rect -1117 -5949 -1115 -5947
rect -1107 -5949 -1105 -5947
rect -1099 -5949 -1097 -5947
rect -1083 -5949 -1081 -5947
rect -1075 -5949 -1073 -5947
rect -930 -5949 -928 -5947
rect -920 -5949 -918 -5947
rect -904 -5949 -902 -5947
rect -896 -5949 -894 -5947
rect -880 -5949 -878 -5947
rect -872 -5949 -870 -5947
rect -862 -5949 -860 -5947
rect -854 -5949 -852 -5947
rect -838 -5949 -836 -5947
rect -830 -5949 -828 -5947
rect -820 -5949 -818 -5947
rect -812 -5949 -810 -5947
rect -796 -5949 -794 -5947
rect -788 -5949 -786 -5947
rect -778 -5949 -776 -5947
rect -770 -5949 -768 -5947
rect -754 -5949 -752 -5947
rect -746 -5949 -744 -5947
rect -572 -5949 -570 -5947
rect -562 -5949 -560 -5947
rect -546 -5949 -544 -5947
rect -538 -5949 -536 -5947
rect -522 -5949 -520 -5947
rect -514 -5949 -512 -5947
rect -504 -5949 -502 -5947
rect -496 -5949 -494 -5947
rect -480 -5949 -478 -5947
rect -472 -5949 -470 -5947
rect -462 -5949 -460 -5947
rect -454 -5949 -452 -5947
rect -438 -5949 -436 -5947
rect -430 -5949 -428 -5947
rect -420 -5949 -418 -5947
rect -412 -5949 -410 -5947
rect -396 -5949 -394 -5947
rect -388 -5949 -386 -5947
rect -214 -5949 -212 -5947
rect -204 -5949 -202 -5947
rect -188 -5949 -186 -5947
rect -180 -5949 -178 -5947
rect -164 -5949 -162 -5947
rect -156 -5949 -154 -5947
rect -146 -5949 -144 -5947
rect -138 -5949 -136 -5947
rect -122 -5949 -120 -5947
rect -114 -5949 -112 -5947
rect -104 -5949 -102 -5947
rect -96 -5949 -94 -5947
rect -80 -5949 -78 -5947
rect -72 -5949 -70 -5947
rect -62 -5949 -60 -5947
rect -54 -5949 -52 -5947
rect -38 -5949 -36 -5947
rect -30 -5949 -28 -5947
rect 214 -5949 216 -5947
rect 224 -5949 226 -5947
rect 240 -5949 242 -5947
rect 248 -5949 250 -5947
rect 264 -5949 266 -5947
rect 272 -5949 274 -5947
rect 282 -5949 284 -5947
rect 290 -5949 292 -5947
rect 306 -5949 308 -5947
rect 314 -5949 316 -5947
rect 324 -5949 326 -5947
rect 332 -5949 334 -5947
rect 348 -5949 350 -5947
rect 356 -5949 358 -5947
rect 366 -5949 368 -5947
rect 374 -5949 376 -5947
rect 390 -5949 392 -5947
rect 398 -5949 400 -5947
rect 570 -5949 572 -5947
rect 580 -5949 582 -5947
rect 596 -5949 598 -5947
rect 604 -5949 606 -5947
rect 620 -5949 622 -5947
rect 628 -5949 630 -5947
rect 638 -5949 640 -5947
rect 646 -5949 648 -5947
rect 662 -5949 664 -5947
rect 670 -5949 672 -5947
rect 680 -5949 682 -5947
rect 688 -5949 690 -5947
rect 704 -5949 706 -5947
rect 712 -5949 714 -5947
rect 722 -5949 724 -5947
rect 730 -5949 732 -5947
rect 746 -5949 748 -5947
rect 754 -5949 756 -5947
rect 968 -5949 970 -5947
rect 978 -5949 980 -5947
rect 994 -5949 996 -5947
rect 1002 -5949 1004 -5947
rect 1018 -5949 1020 -5947
rect 1026 -5949 1028 -5947
rect 1036 -5949 1038 -5947
rect 1044 -5949 1046 -5947
rect 1060 -5949 1062 -5947
rect 1068 -5949 1070 -5947
rect 1078 -5949 1080 -5947
rect 1086 -5949 1088 -5947
rect 1102 -5949 1104 -5947
rect 1110 -5949 1112 -5947
rect 1120 -5949 1122 -5947
rect 1128 -5949 1130 -5947
rect 1144 -5949 1146 -5947
rect 1152 -5949 1154 -5947
rect 1326 -5949 1328 -5947
rect 1336 -5949 1338 -5947
rect 1352 -5949 1354 -5947
rect 1360 -5949 1362 -5947
rect 1376 -5949 1378 -5947
rect 1384 -5949 1386 -5947
rect 1394 -5949 1396 -5947
rect 1402 -5949 1404 -5947
rect 1418 -5949 1420 -5947
rect 1426 -5949 1428 -5947
rect 1436 -5949 1438 -5947
rect 1444 -5949 1446 -5947
rect 1460 -5949 1462 -5947
rect 1468 -5949 1470 -5947
rect 1478 -5949 1480 -5947
rect 1486 -5949 1488 -5947
rect 1502 -5949 1504 -5947
rect 1510 -5949 1512 -5947
rect -1259 -6025 -1257 -5957
rect -1249 -6025 -1247 -5957
rect -1233 -6025 -1231 -5957
rect -1225 -6025 -1223 -5957
rect -1209 -6025 -1207 -5957
rect -1201 -6025 -1199 -5957
rect -1191 -6025 -1189 -5957
rect -1183 -6025 -1181 -5957
rect -1167 -6025 -1165 -5957
rect -1159 -5990 -1157 -5957
rect -1149 -5990 -1147 -5957
rect -1159 -5992 -1147 -5990
rect -1159 -6025 -1157 -5992
rect -1149 -6025 -1147 -5992
rect -1141 -6025 -1139 -5957
rect -1125 -6025 -1123 -5957
rect -1117 -6025 -1115 -5957
rect -1107 -6025 -1105 -5957
rect -1099 -6025 -1097 -5957
rect -1083 -6025 -1081 -5957
rect -1075 -6025 -1073 -5957
rect -930 -6025 -928 -5957
rect -920 -6025 -918 -5957
rect -904 -6025 -902 -5957
rect -896 -6025 -894 -5957
rect -880 -6025 -878 -5957
rect -872 -6025 -870 -5957
rect -862 -6025 -860 -5957
rect -854 -6025 -852 -5957
rect -838 -6025 -836 -5957
rect -830 -5990 -828 -5957
rect -820 -5990 -818 -5957
rect -830 -5992 -818 -5990
rect -830 -6025 -828 -5992
rect -820 -6025 -818 -5992
rect -812 -6025 -810 -5957
rect -796 -6025 -794 -5957
rect -788 -6025 -786 -5957
rect -778 -6025 -776 -5957
rect -770 -6025 -768 -5957
rect -754 -6025 -752 -5957
rect -746 -6025 -744 -5957
rect -572 -6025 -570 -5957
rect -562 -6025 -560 -5957
rect -546 -6025 -544 -5957
rect -538 -6025 -536 -5957
rect -522 -6025 -520 -5957
rect -514 -6025 -512 -5957
rect -504 -6025 -502 -5957
rect -496 -6025 -494 -5957
rect -480 -6025 -478 -5957
rect -472 -5990 -470 -5957
rect -462 -5990 -460 -5957
rect -472 -5992 -460 -5990
rect -472 -6025 -470 -5992
rect -462 -6025 -460 -5992
rect -454 -6025 -452 -5957
rect -438 -6025 -436 -5957
rect -430 -6025 -428 -5957
rect -420 -6025 -418 -5957
rect -412 -6025 -410 -5957
rect -396 -6025 -394 -5957
rect -388 -6025 -386 -5957
rect -214 -6025 -212 -5957
rect -204 -6025 -202 -5957
rect -188 -6025 -186 -5957
rect -180 -6025 -178 -5957
rect -164 -6025 -162 -5957
rect -156 -6025 -154 -5957
rect -146 -6025 -144 -5957
rect -138 -6025 -136 -5957
rect -122 -6025 -120 -5957
rect -114 -5990 -112 -5957
rect -104 -5990 -102 -5957
rect -114 -5992 -102 -5990
rect -114 -6025 -112 -5992
rect -104 -6025 -102 -5992
rect -96 -6025 -94 -5957
rect -80 -6025 -78 -5957
rect -72 -6025 -70 -5957
rect -62 -6025 -60 -5957
rect -54 -6025 -52 -5957
rect -38 -6025 -36 -5957
rect -30 -6025 -28 -5957
rect 214 -6025 216 -5957
rect 224 -6025 226 -5957
rect 240 -6025 242 -5957
rect 248 -6025 250 -5957
rect 264 -6025 266 -5957
rect 272 -6025 274 -5957
rect 282 -6025 284 -5957
rect 290 -6025 292 -5957
rect 306 -6025 308 -5957
rect 314 -5990 316 -5957
rect 324 -5990 326 -5957
rect 314 -5992 326 -5990
rect 314 -6025 316 -5992
rect 324 -6025 326 -5992
rect 332 -6025 334 -5957
rect 348 -6025 350 -5957
rect 356 -6025 358 -5957
rect 366 -6025 368 -5957
rect 374 -6025 376 -5957
rect 390 -6025 392 -5957
rect 398 -6025 400 -5957
rect 570 -6025 572 -5957
rect 580 -6025 582 -5957
rect 596 -6025 598 -5957
rect 604 -6025 606 -5957
rect 620 -6025 622 -5957
rect 628 -6025 630 -5957
rect 638 -6025 640 -5957
rect 646 -6025 648 -5957
rect 662 -6025 664 -5957
rect 670 -5990 672 -5957
rect 680 -5990 682 -5957
rect 670 -5992 682 -5990
rect 670 -6025 672 -5992
rect 680 -6025 682 -5992
rect 688 -6025 690 -5957
rect 704 -6025 706 -5957
rect 712 -6025 714 -5957
rect 722 -6025 724 -5957
rect 730 -6025 732 -5957
rect 746 -6025 748 -5957
rect 754 -6025 756 -5957
rect 968 -6025 970 -5957
rect 978 -6025 980 -5957
rect 994 -6025 996 -5957
rect 1002 -6025 1004 -5957
rect 1018 -6025 1020 -5957
rect 1026 -6025 1028 -5957
rect 1036 -6025 1038 -5957
rect 1044 -6025 1046 -5957
rect 1060 -6025 1062 -5957
rect 1068 -5990 1070 -5957
rect 1078 -5990 1080 -5957
rect 1068 -5992 1080 -5990
rect 1068 -6025 1070 -5992
rect 1078 -6025 1080 -5992
rect 1086 -6025 1088 -5957
rect 1102 -6025 1104 -5957
rect 1110 -6025 1112 -5957
rect 1120 -6025 1122 -5957
rect 1128 -6025 1130 -5957
rect 1144 -6025 1146 -5957
rect 1152 -6025 1154 -5957
rect 1326 -6025 1328 -5957
rect 1336 -6025 1338 -5957
rect 1352 -6025 1354 -5957
rect 1360 -6025 1362 -5957
rect 1376 -6025 1378 -5957
rect 1384 -6025 1386 -5957
rect 1394 -6025 1396 -5957
rect 1402 -6025 1404 -5957
rect 1418 -6025 1420 -5957
rect 1426 -5990 1428 -5957
rect 1436 -5990 1438 -5957
rect 1426 -5992 1438 -5990
rect 1426 -6025 1428 -5992
rect 1436 -6025 1438 -5992
rect 1444 -6025 1446 -5957
rect 1460 -6025 1462 -5957
rect 1468 -6025 1470 -5957
rect 1478 -6025 1480 -5957
rect 1486 -6025 1488 -5957
rect 1502 -6025 1504 -5957
rect 1510 -6025 1512 -5957
rect -1259 -6031 -1257 -6029
rect -1249 -6031 -1247 -6029
rect -1233 -6031 -1231 -6029
rect -1225 -6031 -1223 -6029
rect -1209 -6031 -1207 -6029
rect -1201 -6031 -1199 -6029
rect -1191 -6031 -1189 -6029
rect -1183 -6031 -1181 -6029
rect -1167 -6031 -1165 -6029
rect -1159 -6031 -1157 -6029
rect -1149 -6031 -1147 -6029
rect -1141 -6031 -1139 -6029
rect -1125 -6031 -1123 -6029
rect -1117 -6031 -1115 -6029
rect -1107 -6031 -1105 -6029
rect -1099 -6031 -1097 -6029
rect -1083 -6031 -1081 -6029
rect -1075 -6031 -1073 -6029
rect -930 -6031 -928 -6029
rect -920 -6031 -918 -6029
rect -904 -6031 -902 -6029
rect -896 -6031 -894 -6029
rect -880 -6031 -878 -6029
rect -872 -6031 -870 -6029
rect -862 -6031 -860 -6029
rect -854 -6031 -852 -6029
rect -838 -6031 -836 -6029
rect -830 -6031 -828 -6029
rect -820 -6031 -818 -6029
rect -812 -6031 -810 -6029
rect -796 -6031 -794 -6029
rect -788 -6031 -786 -6029
rect -778 -6031 -776 -6029
rect -770 -6031 -768 -6029
rect -754 -6031 -752 -6029
rect -746 -6031 -744 -6029
rect -572 -6031 -570 -6029
rect -562 -6031 -560 -6029
rect -546 -6031 -544 -6029
rect -538 -6031 -536 -6029
rect -522 -6031 -520 -6029
rect -514 -6031 -512 -6029
rect -504 -6031 -502 -6029
rect -496 -6031 -494 -6029
rect -480 -6031 -478 -6029
rect -472 -6031 -470 -6029
rect -462 -6031 -460 -6029
rect -454 -6031 -452 -6029
rect -438 -6031 -436 -6029
rect -430 -6031 -428 -6029
rect -420 -6031 -418 -6029
rect -412 -6031 -410 -6029
rect -396 -6031 -394 -6029
rect -388 -6031 -386 -6029
rect -214 -6031 -212 -6029
rect -204 -6031 -202 -6029
rect -188 -6031 -186 -6029
rect -180 -6031 -178 -6029
rect -164 -6031 -162 -6029
rect -156 -6031 -154 -6029
rect -146 -6031 -144 -6029
rect -138 -6031 -136 -6029
rect -122 -6031 -120 -6029
rect -114 -6031 -112 -6029
rect -104 -6031 -102 -6029
rect -96 -6031 -94 -6029
rect -80 -6031 -78 -6029
rect -72 -6031 -70 -6029
rect -62 -6031 -60 -6029
rect -54 -6031 -52 -6029
rect -38 -6031 -36 -6029
rect -30 -6031 -28 -6029
rect 214 -6031 216 -6029
rect 224 -6031 226 -6029
rect 240 -6031 242 -6029
rect 248 -6031 250 -6029
rect 264 -6031 266 -6029
rect 272 -6031 274 -6029
rect 282 -6031 284 -6029
rect 290 -6031 292 -6029
rect 306 -6031 308 -6029
rect 314 -6031 316 -6029
rect 324 -6031 326 -6029
rect 332 -6031 334 -6029
rect 348 -6031 350 -6029
rect 356 -6031 358 -6029
rect 366 -6031 368 -6029
rect 374 -6031 376 -6029
rect 390 -6031 392 -6029
rect 398 -6031 400 -6029
rect 570 -6031 572 -6029
rect 580 -6031 582 -6029
rect 596 -6031 598 -6029
rect 604 -6031 606 -6029
rect 620 -6031 622 -6029
rect 628 -6031 630 -6029
rect 638 -6031 640 -6029
rect 646 -6031 648 -6029
rect 662 -6031 664 -6029
rect 670 -6031 672 -6029
rect 680 -6031 682 -6029
rect 688 -6031 690 -6029
rect 704 -6031 706 -6029
rect 712 -6031 714 -6029
rect 722 -6031 724 -6029
rect 730 -6031 732 -6029
rect 746 -6031 748 -6029
rect 754 -6031 756 -6029
rect 968 -6031 970 -6029
rect 978 -6031 980 -6029
rect 994 -6031 996 -6029
rect 1002 -6031 1004 -6029
rect 1018 -6031 1020 -6029
rect 1026 -6031 1028 -6029
rect 1036 -6031 1038 -6029
rect 1044 -6031 1046 -6029
rect 1060 -6031 1062 -6029
rect 1068 -6031 1070 -6029
rect 1078 -6031 1080 -6029
rect 1086 -6031 1088 -6029
rect 1102 -6031 1104 -6029
rect 1110 -6031 1112 -6029
rect 1120 -6031 1122 -6029
rect 1128 -6031 1130 -6029
rect 1144 -6031 1146 -6029
rect 1152 -6031 1154 -6029
rect 1326 -6031 1328 -6029
rect 1336 -6031 1338 -6029
rect 1352 -6031 1354 -6029
rect 1360 -6031 1362 -6029
rect 1376 -6031 1378 -6029
rect 1384 -6031 1386 -6029
rect 1394 -6031 1396 -6029
rect 1402 -6031 1404 -6029
rect 1418 -6031 1420 -6029
rect 1426 -6031 1428 -6029
rect 1436 -6031 1438 -6029
rect 1444 -6031 1446 -6029
rect 1460 -6031 1462 -6029
rect 1468 -6031 1470 -6029
rect 1478 -6031 1480 -6029
rect 1486 -6031 1488 -6029
rect 1502 -6031 1504 -6029
rect 1510 -6031 1512 -6029
rect 1326 -6067 1328 -6065
rect 1336 -6067 1338 -6065
rect 1352 -6067 1354 -6065
rect 1360 -6067 1362 -6065
rect 1376 -6067 1378 -6065
rect 1384 -6067 1386 -6065
rect 1394 -6067 1396 -6065
rect 1402 -6067 1404 -6065
rect 1418 -6067 1420 -6065
rect 1426 -6067 1428 -6065
rect 1436 -6067 1438 -6065
rect 1444 -6067 1446 -6065
rect 1460 -6067 1462 -6065
rect 1468 -6067 1470 -6065
rect 1478 -6067 1480 -6065
rect 1486 -6067 1488 -6065
rect 1502 -6067 1504 -6065
rect 1510 -6067 1512 -6065
rect 1326 -6143 1328 -6075
rect 1336 -6143 1338 -6075
rect 1352 -6143 1354 -6075
rect 1360 -6143 1362 -6075
rect 1376 -6143 1378 -6075
rect 1384 -6143 1386 -6075
rect 1394 -6143 1396 -6075
rect 1402 -6143 1404 -6075
rect 1418 -6143 1420 -6075
rect 1426 -6108 1428 -6075
rect 1436 -6108 1438 -6075
rect 1426 -6110 1438 -6108
rect 1426 -6143 1428 -6110
rect 1436 -6143 1438 -6110
rect 1444 -6143 1446 -6075
rect 1460 -6143 1462 -6075
rect 1468 -6143 1470 -6075
rect 1478 -6143 1480 -6075
rect 1486 -6143 1488 -6075
rect 1502 -6143 1504 -6075
rect 1510 -6143 1512 -6075
rect 1326 -6149 1328 -6147
rect 1336 -6149 1338 -6147
rect 1352 -6149 1354 -6147
rect 1360 -6149 1362 -6147
rect 1376 -6149 1378 -6147
rect 1384 -6149 1386 -6147
rect 1394 -6149 1396 -6147
rect 1402 -6149 1404 -6147
rect 1418 -6149 1420 -6147
rect 1426 -6149 1428 -6147
rect 1436 -6149 1438 -6147
rect 1444 -6149 1446 -6147
rect 1460 -6149 1462 -6147
rect 1468 -6149 1470 -6147
rect 1478 -6149 1480 -6147
rect 1486 -6149 1488 -6147
rect 1502 -6149 1504 -6147
rect 1510 -6149 1512 -6147
<< ndiffusion >>
rect -1333 -1118 -1332 -1114
rect -1330 -1118 -1324 -1114
rect -1322 -1118 -1320 -1114
rect -1316 -1118 -1314 -1114
rect -1312 -1118 -1311 -1114
rect -932 -1118 -931 -1114
rect -929 -1118 -923 -1114
rect -921 -1118 -919 -1114
rect -915 -1118 -913 -1114
rect -911 -1118 -910 -1114
rect -573 -1118 -572 -1114
rect -570 -1118 -564 -1114
rect -562 -1118 -560 -1114
rect -556 -1118 -554 -1114
rect -552 -1118 -551 -1114
rect -215 -1118 -214 -1114
rect -212 -1118 -206 -1114
rect -204 -1118 -202 -1114
rect -198 -1118 -196 -1114
rect -194 -1118 -193 -1114
rect 213 -1118 214 -1114
rect 216 -1118 222 -1114
rect 224 -1118 226 -1114
rect 230 -1118 232 -1114
rect 234 -1118 235 -1114
rect 569 -1118 570 -1114
rect 572 -1118 578 -1114
rect 580 -1118 582 -1114
rect 586 -1118 588 -1114
rect 590 -1118 591 -1114
rect 967 -1118 968 -1114
rect 970 -1118 976 -1114
rect 978 -1118 980 -1114
rect 984 -1118 986 -1114
rect 988 -1118 989 -1114
rect 1325 -1118 1326 -1114
rect 1328 -1118 1334 -1114
rect 1336 -1118 1338 -1114
rect 1342 -1118 1344 -1114
rect 1346 -1118 1347 -1114
rect -1256 -1232 -1255 -1228
rect -1253 -1232 -1251 -1228
rect -1247 -1232 -1245 -1228
rect -1243 -1232 -1242 -1228
rect -1230 -1232 -1229 -1228
rect -1227 -1232 -1221 -1228
rect -1219 -1232 -1218 -1228
rect -1206 -1232 -1205 -1228
rect -1203 -1232 -1197 -1228
rect -1195 -1232 -1193 -1228
rect -1189 -1232 -1187 -1228
rect -1185 -1232 -1179 -1228
rect -1177 -1232 -1176 -1228
rect -1164 -1232 -1163 -1228
rect -1161 -1232 -1155 -1228
rect -1153 -1232 -1151 -1228
rect -1147 -1232 -1145 -1228
rect -1143 -1232 -1137 -1228
rect -1135 -1232 -1134 -1228
rect -1122 -1232 -1121 -1228
rect -1119 -1232 -1113 -1228
rect -1111 -1232 -1109 -1228
rect -1105 -1232 -1103 -1228
rect -1101 -1232 -1095 -1228
rect -1093 -1232 -1092 -1228
rect -1080 -1232 -1079 -1228
rect -1077 -1232 -1071 -1228
rect -1069 -1232 -1068 -1228
rect -931 -1232 -930 -1228
rect -928 -1232 -926 -1228
rect -922 -1232 -920 -1228
rect -918 -1232 -917 -1228
rect -905 -1232 -904 -1228
rect -902 -1232 -896 -1228
rect -894 -1232 -893 -1228
rect -881 -1232 -880 -1228
rect -878 -1232 -872 -1228
rect -870 -1232 -868 -1228
rect -864 -1232 -862 -1228
rect -860 -1232 -854 -1228
rect -852 -1232 -851 -1228
rect -839 -1232 -838 -1228
rect -836 -1232 -830 -1228
rect -828 -1232 -826 -1228
rect -822 -1232 -820 -1228
rect -818 -1232 -812 -1228
rect -810 -1232 -809 -1228
rect -797 -1232 -796 -1228
rect -794 -1232 -788 -1228
rect -786 -1232 -784 -1228
rect -780 -1232 -778 -1228
rect -776 -1232 -770 -1228
rect -768 -1232 -767 -1228
rect -755 -1232 -754 -1228
rect -752 -1232 -746 -1228
rect -744 -1232 -743 -1228
rect -573 -1232 -572 -1228
rect -570 -1232 -568 -1228
rect -564 -1232 -562 -1228
rect -560 -1232 -559 -1228
rect -547 -1232 -546 -1228
rect -544 -1232 -538 -1228
rect -536 -1232 -535 -1228
rect -523 -1232 -522 -1228
rect -520 -1232 -514 -1228
rect -512 -1232 -510 -1228
rect -506 -1232 -504 -1228
rect -502 -1232 -496 -1228
rect -494 -1232 -493 -1228
rect -481 -1232 -480 -1228
rect -478 -1232 -472 -1228
rect -470 -1232 -468 -1228
rect -464 -1232 -462 -1228
rect -460 -1232 -454 -1228
rect -452 -1232 -451 -1228
rect -439 -1232 -438 -1228
rect -436 -1232 -430 -1228
rect -428 -1232 -426 -1228
rect -422 -1232 -420 -1228
rect -418 -1232 -412 -1228
rect -410 -1232 -409 -1228
rect -397 -1232 -396 -1228
rect -394 -1232 -388 -1228
rect -386 -1232 -385 -1228
rect -215 -1232 -214 -1228
rect -212 -1232 -210 -1228
rect -206 -1232 -204 -1228
rect -202 -1232 -201 -1228
rect -189 -1232 -188 -1228
rect -186 -1232 -180 -1228
rect -178 -1232 -177 -1228
rect -165 -1232 -164 -1228
rect -162 -1232 -156 -1228
rect -154 -1232 -152 -1228
rect -148 -1232 -146 -1228
rect -144 -1232 -138 -1228
rect -136 -1232 -135 -1228
rect -123 -1232 -122 -1228
rect -120 -1232 -114 -1228
rect -112 -1232 -110 -1228
rect -106 -1232 -104 -1228
rect -102 -1232 -96 -1228
rect -94 -1232 -93 -1228
rect -81 -1232 -80 -1228
rect -78 -1232 -72 -1228
rect -70 -1232 -68 -1228
rect -64 -1232 -62 -1228
rect -60 -1232 -54 -1228
rect -52 -1232 -51 -1228
rect -39 -1232 -38 -1228
rect -36 -1232 -30 -1228
rect -28 -1232 -27 -1228
rect 213 -1232 214 -1228
rect 216 -1232 218 -1228
rect 222 -1232 224 -1228
rect 226 -1232 227 -1228
rect 239 -1232 240 -1228
rect 242 -1232 248 -1228
rect 250 -1232 251 -1228
rect 263 -1232 264 -1228
rect 266 -1232 272 -1228
rect 274 -1232 276 -1228
rect 280 -1232 282 -1228
rect 284 -1232 290 -1228
rect 292 -1232 293 -1228
rect 305 -1232 306 -1228
rect 308 -1232 314 -1228
rect 316 -1232 318 -1228
rect 322 -1232 324 -1228
rect 326 -1232 332 -1228
rect 334 -1232 335 -1228
rect 347 -1232 348 -1228
rect 350 -1232 356 -1228
rect 358 -1232 360 -1228
rect 364 -1232 366 -1228
rect 368 -1232 374 -1228
rect 376 -1232 377 -1228
rect 389 -1232 390 -1228
rect 392 -1232 398 -1228
rect 400 -1232 401 -1228
rect 569 -1232 570 -1228
rect 572 -1232 574 -1228
rect 578 -1232 580 -1228
rect 582 -1232 583 -1228
rect 595 -1232 596 -1228
rect 598 -1232 604 -1228
rect 606 -1232 607 -1228
rect 619 -1232 620 -1228
rect 622 -1232 628 -1228
rect 630 -1232 632 -1228
rect 636 -1232 638 -1228
rect 640 -1232 646 -1228
rect 648 -1232 649 -1228
rect 661 -1232 662 -1228
rect 664 -1232 670 -1228
rect 672 -1232 674 -1228
rect 678 -1232 680 -1228
rect 682 -1232 688 -1228
rect 690 -1232 691 -1228
rect 703 -1232 704 -1228
rect 706 -1232 712 -1228
rect 714 -1232 716 -1228
rect 720 -1232 722 -1228
rect 724 -1232 730 -1228
rect 732 -1232 733 -1228
rect 745 -1232 746 -1228
rect 748 -1232 754 -1228
rect 756 -1232 757 -1228
rect 967 -1232 968 -1228
rect 970 -1232 972 -1228
rect 976 -1232 978 -1228
rect 980 -1232 981 -1228
rect 993 -1232 994 -1228
rect 996 -1232 1002 -1228
rect 1004 -1232 1005 -1228
rect 1017 -1232 1018 -1228
rect 1020 -1232 1026 -1228
rect 1028 -1232 1030 -1228
rect 1034 -1232 1036 -1228
rect 1038 -1232 1044 -1228
rect 1046 -1232 1047 -1228
rect 1059 -1232 1060 -1228
rect 1062 -1232 1068 -1228
rect 1070 -1232 1072 -1228
rect 1076 -1232 1078 -1228
rect 1080 -1232 1086 -1228
rect 1088 -1232 1089 -1228
rect 1101 -1232 1102 -1228
rect 1104 -1232 1110 -1228
rect 1112 -1232 1114 -1228
rect 1118 -1232 1120 -1228
rect 1122 -1232 1128 -1228
rect 1130 -1232 1131 -1228
rect 1143 -1232 1144 -1228
rect 1146 -1232 1152 -1228
rect 1154 -1232 1155 -1228
rect -1335 -1348 -1334 -1344
rect -1332 -1348 -1326 -1344
rect -1324 -1348 -1322 -1344
rect -1318 -1348 -1316 -1344
rect -1314 -1348 -1313 -1344
rect -931 -1348 -930 -1344
rect -928 -1348 -922 -1344
rect -920 -1348 -918 -1344
rect -914 -1348 -912 -1344
rect -910 -1348 -909 -1344
rect -573 -1348 -572 -1344
rect -570 -1348 -564 -1344
rect -562 -1348 -560 -1344
rect -556 -1348 -554 -1344
rect -552 -1348 -551 -1344
rect -215 -1348 -214 -1344
rect -212 -1348 -206 -1344
rect -204 -1348 -202 -1344
rect -198 -1348 -196 -1344
rect -194 -1348 -193 -1344
rect 213 -1348 214 -1344
rect 216 -1348 222 -1344
rect 224 -1348 226 -1344
rect 230 -1348 232 -1344
rect 234 -1348 235 -1344
rect 569 -1348 570 -1344
rect 572 -1348 578 -1344
rect 580 -1348 582 -1344
rect 586 -1348 588 -1344
rect 590 -1348 591 -1344
rect 967 -1348 968 -1344
rect 970 -1348 976 -1344
rect 978 -1348 980 -1344
rect 984 -1348 986 -1344
rect 988 -1348 989 -1344
rect 1325 -1348 1326 -1344
rect 1328 -1348 1334 -1344
rect 1336 -1348 1338 -1344
rect 1342 -1348 1344 -1344
rect 1346 -1348 1347 -1344
rect -1256 -1462 -1255 -1458
rect -1253 -1462 -1251 -1458
rect -1247 -1462 -1245 -1458
rect -1243 -1462 -1242 -1458
rect -1230 -1462 -1229 -1458
rect -1227 -1462 -1225 -1458
rect -1221 -1462 -1219 -1458
rect -1217 -1462 -1211 -1458
rect -1209 -1462 -1207 -1458
rect -1203 -1462 -1201 -1458
rect -1199 -1462 -1198 -1458
rect -1186 -1462 -1185 -1458
rect -1183 -1462 -1177 -1458
rect -1175 -1462 -1173 -1458
rect -1169 -1462 -1167 -1458
rect -1165 -1462 -1164 -1458
rect -931 -1462 -930 -1458
rect -928 -1462 -926 -1458
rect -922 -1462 -920 -1458
rect -918 -1462 -917 -1458
rect -905 -1462 -904 -1458
rect -902 -1462 -900 -1458
rect -896 -1462 -894 -1458
rect -892 -1462 -891 -1458
rect -879 -1462 -878 -1458
rect -876 -1462 -875 -1458
rect -871 -1462 -868 -1458
rect -866 -1462 -860 -1458
rect -858 -1462 -857 -1458
rect -853 -1462 -850 -1458
rect -848 -1462 -847 -1458
rect -835 -1462 -834 -1458
rect -832 -1462 -826 -1458
rect -824 -1462 -822 -1458
rect -818 -1462 -816 -1458
rect -814 -1462 -813 -1458
rect -801 -1462 -800 -1458
rect -798 -1462 -796 -1458
rect -792 -1462 -790 -1458
rect -788 -1462 -782 -1458
rect -780 -1462 -778 -1458
rect -774 -1462 -772 -1458
rect -770 -1462 -769 -1458
rect -757 -1462 -756 -1458
rect -754 -1462 -748 -1458
rect -746 -1462 -745 -1458
rect -733 -1462 -732 -1458
rect -730 -1462 -725 -1458
rect -721 -1462 -716 -1458
rect -714 -1462 -713 -1458
rect -709 -1462 -708 -1458
rect -706 -1462 -704 -1458
rect -700 -1462 -698 -1458
rect -696 -1462 -695 -1458
rect -573 -1462 -572 -1458
rect -570 -1462 -568 -1458
rect -564 -1462 -562 -1458
rect -560 -1462 -559 -1458
rect -547 -1462 -546 -1458
rect -544 -1462 -542 -1458
rect -538 -1462 -536 -1458
rect -534 -1462 -533 -1458
rect -521 -1462 -520 -1458
rect -518 -1462 -517 -1458
rect -513 -1462 -510 -1458
rect -508 -1462 -502 -1458
rect -500 -1462 -499 -1458
rect -495 -1462 -492 -1458
rect -490 -1462 -489 -1458
rect -477 -1462 -476 -1458
rect -474 -1462 -468 -1458
rect -466 -1462 -464 -1458
rect -460 -1462 -458 -1458
rect -456 -1462 -455 -1458
rect -443 -1462 -442 -1458
rect -440 -1462 -438 -1458
rect -434 -1462 -432 -1458
rect -430 -1462 -424 -1458
rect -422 -1462 -420 -1458
rect -416 -1462 -414 -1458
rect -412 -1462 -411 -1458
rect -399 -1462 -398 -1458
rect -396 -1462 -390 -1458
rect -388 -1462 -387 -1458
rect -375 -1462 -374 -1458
rect -372 -1462 -367 -1458
rect -363 -1462 -358 -1458
rect -356 -1462 -355 -1458
rect -351 -1462 -350 -1458
rect -348 -1462 -346 -1458
rect -342 -1462 -340 -1458
rect -338 -1462 -337 -1458
rect -215 -1462 -214 -1458
rect -212 -1462 -210 -1458
rect -206 -1462 -204 -1458
rect -202 -1462 -201 -1458
rect -189 -1462 -188 -1458
rect -186 -1462 -184 -1458
rect -180 -1462 -178 -1458
rect -176 -1462 -175 -1458
rect -163 -1462 -162 -1458
rect -160 -1462 -159 -1458
rect -155 -1462 -152 -1458
rect -150 -1462 -144 -1458
rect -142 -1462 -141 -1458
rect -137 -1462 -134 -1458
rect -132 -1462 -131 -1458
rect -119 -1462 -118 -1458
rect -116 -1462 -110 -1458
rect -108 -1462 -106 -1458
rect -102 -1462 -100 -1458
rect -98 -1462 -97 -1458
rect -85 -1462 -84 -1458
rect -82 -1462 -80 -1458
rect -76 -1462 -74 -1458
rect -72 -1462 -66 -1458
rect -64 -1462 -62 -1458
rect -58 -1462 -56 -1458
rect -54 -1462 -53 -1458
rect -41 -1462 -40 -1458
rect -38 -1462 -32 -1458
rect -30 -1462 -29 -1458
rect -17 -1462 -16 -1458
rect -14 -1462 -9 -1458
rect -5 -1462 0 -1458
rect 2 -1462 3 -1458
rect 7 -1462 8 -1458
rect 10 -1462 12 -1458
rect 16 -1462 18 -1458
rect 20 -1462 21 -1458
rect 213 -1462 214 -1458
rect 216 -1462 218 -1458
rect 222 -1462 224 -1458
rect 226 -1462 227 -1458
rect 239 -1462 240 -1458
rect 242 -1462 244 -1458
rect 248 -1462 250 -1458
rect 252 -1462 253 -1458
rect 265 -1462 266 -1458
rect 268 -1462 269 -1458
rect 273 -1462 276 -1458
rect 278 -1462 284 -1458
rect 286 -1462 287 -1458
rect 291 -1462 294 -1458
rect 296 -1462 297 -1458
rect 309 -1462 310 -1458
rect 312 -1462 318 -1458
rect 320 -1462 322 -1458
rect 326 -1462 328 -1458
rect 330 -1462 331 -1458
rect 343 -1462 344 -1458
rect 346 -1462 348 -1458
rect 352 -1462 354 -1458
rect 356 -1462 362 -1458
rect 364 -1462 366 -1458
rect 370 -1462 372 -1458
rect 374 -1462 375 -1458
rect 387 -1462 388 -1458
rect 390 -1462 396 -1458
rect 398 -1462 399 -1458
rect 411 -1462 412 -1458
rect 414 -1462 419 -1458
rect 423 -1462 428 -1458
rect 430 -1462 431 -1458
rect 435 -1462 436 -1458
rect 438 -1462 440 -1458
rect 444 -1462 446 -1458
rect 448 -1462 449 -1458
rect 569 -1462 570 -1458
rect 572 -1462 574 -1458
rect 578 -1462 580 -1458
rect 582 -1462 583 -1458
rect 595 -1462 596 -1458
rect 598 -1462 600 -1458
rect 604 -1462 606 -1458
rect 608 -1462 609 -1458
rect 621 -1462 622 -1458
rect 624 -1462 625 -1458
rect 629 -1462 632 -1458
rect 634 -1462 640 -1458
rect 642 -1462 643 -1458
rect 647 -1462 650 -1458
rect 652 -1462 653 -1458
rect 665 -1462 666 -1458
rect 668 -1462 674 -1458
rect 676 -1462 678 -1458
rect 682 -1462 684 -1458
rect 686 -1462 687 -1458
rect 699 -1462 700 -1458
rect 702 -1462 704 -1458
rect 708 -1462 710 -1458
rect 712 -1462 718 -1458
rect 720 -1462 722 -1458
rect 726 -1462 728 -1458
rect 730 -1462 731 -1458
rect 743 -1462 744 -1458
rect 746 -1462 752 -1458
rect 754 -1462 755 -1458
rect 767 -1462 768 -1458
rect 770 -1462 775 -1458
rect 779 -1462 784 -1458
rect 786 -1462 787 -1458
rect 791 -1462 792 -1458
rect 794 -1462 796 -1458
rect 800 -1462 802 -1458
rect 804 -1462 805 -1458
rect 967 -1462 968 -1458
rect 970 -1462 972 -1458
rect 976 -1462 978 -1458
rect 980 -1462 981 -1458
rect 993 -1462 994 -1458
rect 996 -1462 998 -1458
rect 1002 -1462 1004 -1458
rect 1006 -1462 1007 -1458
rect 1019 -1462 1020 -1458
rect 1022 -1462 1023 -1458
rect 1027 -1462 1030 -1458
rect 1032 -1462 1038 -1458
rect 1040 -1462 1041 -1458
rect 1045 -1462 1048 -1458
rect 1050 -1462 1051 -1458
rect 1063 -1462 1064 -1458
rect 1066 -1462 1072 -1458
rect 1074 -1462 1076 -1458
rect 1080 -1462 1082 -1458
rect 1084 -1462 1085 -1458
rect 1097 -1462 1098 -1458
rect 1100 -1462 1102 -1458
rect 1106 -1462 1108 -1458
rect 1110 -1462 1116 -1458
rect 1118 -1462 1120 -1458
rect 1124 -1462 1126 -1458
rect 1128 -1462 1129 -1458
rect 1141 -1462 1142 -1458
rect 1144 -1462 1150 -1458
rect 1152 -1462 1153 -1458
rect 1165 -1462 1166 -1458
rect 1168 -1462 1173 -1458
rect 1177 -1462 1182 -1458
rect 1184 -1462 1185 -1458
rect 1189 -1462 1190 -1458
rect 1192 -1462 1194 -1458
rect 1198 -1462 1200 -1458
rect 1202 -1462 1203 -1458
rect 1325 -1462 1326 -1458
rect 1328 -1462 1330 -1458
rect 1334 -1462 1336 -1458
rect 1338 -1462 1339 -1458
rect 1351 -1462 1352 -1458
rect 1354 -1462 1356 -1458
rect 1360 -1462 1362 -1458
rect 1364 -1462 1370 -1458
rect 1372 -1462 1374 -1458
rect 1378 -1462 1380 -1458
rect 1382 -1462 1383 -1458
rect 1395 -1462 1396 -1458
rect 1398 -1462 1404 -1458
rect 1406 -1462 1408 -1458
rect 1412 -1462 1414 -1458
rect 1416 -1462 1417 -1458
rect -1256 -1585 -1255 -1581
rect -1253 -1585 -1251 -1581
rect -1247 -1585 -1245 -1581
rect -1243 -1585 -1242 -1581
rect -1230 -1585 -1229 -1581
rect -1227 -1585 -1221 -1581
rect -1219 -1585 -1218 -1581
rect -1206 -1585 -1205 -1581
rect -1203 -1585 -1197 -1581
rect -1195 -1585 -1193 -1581
rect -1189 -1585 -1187 -1581
rect -1185 -1585 -1179 -1581
rect -1177 -1585 -1176 -1581
rect -1164 -1585 -1163 -1581
rect -1161 -1585 -1155 -1581
rect -1153 -1585 -1151 -1581
rect -1147 -1585 -1145 -1581
rect -1143 -1585 -1137 -1581
rect -1135 -1585 -1134 -1581
rect -1122 -1585 -1121 -1581
rect -1119 -1585 -1113 -1581
rect -1111 -1585 -1109 -1581
rect -1105 -1585 -1103 -1581
rect -1101 -1585 -1095 -1581
rect -1093 -1585 -1092 -1581
rect -1080 -1585 -1079 -1581
rect -1077 -1585 -1071 -1581
rect -1069 -1585 -1068 -1581
rect -931 -1585 -930 -1581
rect -928 -1585 -926 -1581
rect -922 -1585 -920 -1581
rect -918 -1585 -917 -1581
rect -905 -1585 -904 -1581
rect -902 -1585 -896 -1581
rect -894 -1585 -893 -1581
rect -881 -1585 -880 -1581
rect -878 -1585 -872 -1581
rect -870 -1585 -868 -1581
rect -864 -1585 -862 -1581
rect -860 -1585 -854 -1581
rect -852 -1585 -851 -1581
rect -839 -1585 -838 -1581
rect -836 -1585 -830 -1581
rect -828 -1585 -826 -1581
rect -822 -1585 -820 -1581
rect -818 -1585 -812 -1581
rect -810 -1585 -809 -1581
rect -797 -1585 -796 -1581
rect -794 -1585 -788 -1581
rect -786 -1585 -784 -1581
rect -780 -1585 -778 -1581
rect -776 -1585 -770 -1581
rect -768 -1585 -767 -1581
rect -755 -1585 -754 -1581
rect -752 -1585 -746 -1581
rect -744 -1585 -743 -1581
rect -573 -1585 -572 -1581
rect -570 -1585 -568 -1581
rect -564 -1585 -562 -1581
rect -560 -1585 -559 -1581
rect -547 -1585 -546 -1581
rect -544 -1585 -538 -1581
rect -536 -1585 -535 -1581
rect -523 -1585 -522 -1581
rect -520 -1585 -514 -1581
rect -512 -1585 -510 -1581
rect -506 -1585 -504 -1581
rect -502 -1585 -496 -1581
rect -494 -1585 -493 -1581
rect -481 -1585 -480 -1581
rect -478 -1585 -472 -1581
rect -470 -1585 -468 -1581
rect -464 -1585 -462 -1581
rect -460 -1585 -454 -1581
rect -452 -1585 -451 -1581
rect -439 -1585 -438 -1581
rect -436 -1585 -430 -1581
rect -428 -1585 -426 -1581
rect -422 -1585 -420 -1581
rect -418 -1585 -412 -1581
rect -410 -1585 -409 -1581
rect -397 -1585 -396 -1581
rect -394 -1585 -388 -1581
rect -386 -1585 -385 -1581
rect -215 -1585 -214 -1581
rect -212 -1585 -210 -1581
rect -206 -1585 -204 -1581
rect -202 -1585 -201 -1581
rect -189 -1585 -188 -1581
rect -186 -1585 -180 -1581
rect -178 -1585 -177 -1581
rect -165 -1585 -164 -1581
rect -162 -1585 -156 -1581
rect -154 -1585 -152 -1581
rect -148 -1585 -146 -1581
rect -144 -1585 -138 -1581
rect -136 -1585 -135 -1581
rect -123 -1585 -122 -1581
rect -120 -1585 -114 -1581
rect -112 -1585 -110 -1581
rect -106 -1585 -104 -1581
rect -102 -1585 -96 -1581
rect -94 -1585 -93 -1581
rect -81 -1585 -80 -1581
rect -78 -1585 -72 -1581
rect -70 -1585 -68 -1581
rect -64 -1585 -62 -1581
rect -60 -1585 -54 -1581
rect -52 -1585 -51 -1581
rect -39 -1585 -38 -1581
rect -36 -1585 -30 -1581
rect -28 -1585 -27 -1581
rect 213 -1585 214 -1581
rect 216 -1585 218 -1581
rect 222 -1585 224 -1581
rect 226 -1585 227 -1581
rect 239 -1585 240 -1581
rect 242 -1585 248 -1581
rect 250 -1585 251 -1581
rect 263 -1585 264 -1581
rect 266 -1585 272 -1581
rect 274 -1585 276 -1581
rect 280 -1585 282 -1581
rect 284 -1585 290 -1581
rect 292 -1585 293 -1581
rect 305 -1585 306 -1581
rect 308 -1585 314 -1581
rect 316 -1585 318 -1581
rect 322 -1585 324 -1581
rect 326 -1585 332 -1581
rect 334 -1585 335 -1581
rect 347 -1585 348 -1581
rect 350 -1585 356 -1581
rect 358 -1585 360 -1581
rect 364 -1585 366 -1581
rect 368 -1585 374 -1581
rect 376 -1585 377 -1581
rect 389 -1585 390 -1581
rect 392 -1585 398 -1581
rect 400 -1585 401 -1581
rect 569 -1585 570 -1581
rect 572 -1585 574 -1581
rect 578 -1585 580 -1581
rect 582 -1585 583 -1581
rect 595 -1585 596 -1581
rect 598 -1585 604 -1581
rect 606 -1585 607 -1581
rect 619 -1585 620 -1581
rect 622 -1585 628 -1581
rect 630 -1585 632 -1581
rect 636 -1585 638 -1581
rect 640 -1585 646 -1581
rect 648 -1585 649 -1581
rect 661 -1585 662 -1581
rect 664 -1585 670 -1581
rect 672 -1585 674 -1581
rect 678 -1585 680 -1581
rect 682 -1585 688 -1581
rect 690 -1585 691 -1581
rect 703 -1585 704 -1581
rect 706 -1585 712 -1581
rect 714 -1585 716 -1581
rect 720 -1585 722 -1581
rect 724 -1585 730 -1581
rect 732 -1585 733 -1581
rect 745 -1585 746 -1581
rect 748 -1585 754 -1581
rect 756 -1585 757 -1581
rect 967 -1585 968 -1581
rect 970 -1585 972 -1581
rect 976 -1585 978 -1581
rect 980 -1585 981 -1581
rect 993 -1585 994 -1581
rect 996 -1585 1002 -1581
rect 1004 -1585 1005 -1581
rect 1017 -1585 1018 -1581
rect 1020 -1585 1026 -1581
rect 1028 -1585 1030 -1581
rect 1034 -1585 1036 -1581
rect 1038 -1585 1044 -1581
rect 1046 -1585 1047 -1581
rect 1059 -1585 1060 -1581
rect 1062 -1585 1068 -1581
rect 1070 -1585 1072 -1581
rect 1076 -1585 1078 -1581
rect 1080 -1585 1086 -1581
rect 1088 -1585 1089 -1581
rect 1101 -1585 1102 -1581
rect 1104 -1585 1110 -1581
rect 1112 -1585 1114 -1581
rect 1118 -1585 1120 -1581
rect 1122 -1585 1128 -1581
rect 1130 -1585 1131 -1581
rect 1143 -1585 1144 -1581
rect 1146 -1585 1152 -1581
rect 1154 -1585 1155 -1581
rect -1256 -1706 -1255 -1702
rect -1253 -1706 -1251 -1702
rect -1247 -1706 -1245 -1702
rect -1243 -1706 -1242 -1702
rect -1230 -1706 -1229 -1702
rect -1227 -1706 -1221 -1702
rect -1219 -1706 -1218 -1702
rect -1206 -1706 -1205 -1702
rect -1203 -1706 -1197 -1702
rect -1195 -1706 -1193 -1702
rect -1189 -1706 -1187 -1702
rect -1185 -1706 -1179 -1702
rect -1177 -1706 -1176 -1702
rect -1164 -1706 -1163 -1702
rect -1161 -1706 -1155 -1702
rect -1153 -1706 -1151 -1702
rect -1147 -1706 -1145 -1702
rect -1143 -1706 -1137 -1702
rect -1135 -1706 -1134 -1702
rect -1122 -1706 -1121 -1702
rect -1119 -1706 -1113 -1702
rect -1111 -1706 -1109 -1702
rect -1105 -1706 -1103 -1702
rect -1101 -1706 -1095 -1702
rect -1093 -1706 -1092 -1702
rect -1080 -1706 -1079 -1702
rect -1077 -1706 -1071 -1702
rect -1069 -1706 -1068 -1702
rect -931 -1706 -930 -1702
rect -928 -1706 -926 -1702
rect -922 -1706 -920 -1702
rect -918 -1706 -917 -1702
rect -905 -1706 -904 -1702
rect -902 -1706 -896 -1702
rect -894 -1706 -893 -1702
rect -881 -1706 -880 -1702
rect -878 -1706 -872 -1702
rect -870 -1706 -868 -1702
rect -864 -1706 -862 -1702
rect -860 -1706 -854 -1702
rect -852 -1706 -851 -1702
rect -839 -1706 -838 -1702
rect -836 -1706 -830 -1702
rect -828 -1706 -826 -1702
rect -822 -1706 -820 -1702
rect -818 -1706 -812 -1702
rect -810 -1706 -809 -1702
rect -797 -1706 -796 -1702
rect -794 -1706 -788 -1702
rect -786 -1706 -784 -1702
rect -780 -1706 -778 -1702
rect -776 -1706 -770 -1702
rect -768 -1706 -767 -1702
rect -755 -1706 -754 -1702
rect -752 -1706 -746 -1702
rect -744 -1706 -743 -1702
rect -573 -1706 -572 -1702
rect -570 -1706 -568 -1702
rect -564 -1706 -562 -1702
rect -560 -1706 -559 -1702
rect -547 -1706 -546 -1702
rect -544 -1706 -538 -1702
rect -536 -1706 -535 -1702
rect -523 -1706 -522 -1702
rect -520 -1706 -514 -1702
rect -512 -1706 -510 -1702
rect -506 -1706 -504 -1702
rect -502 -1706 -496 -1702
rect -494 -1706 -493 -1702
rect -481 -1706 -480 -1702
rect -478 -1706 -472 -1702
rect -470 -1706 -468 -1702
rect -464 -1706 -462 -1702
rect -460 -1706 -454 -1702
rect -452 -1706 -451 -1702
rect -439 -1706 -438 -1702
rect -436 -1706 -430 -1702
rect -428 -1706 -426 -1702
rect -422 -1706 -420 -1702
rect -418 -1706 -412 -1702
rect -410 -1706 -409 -1702
rect -397 -1706 -396 -1702
rect -394 -1706 -388 -1702
rect -386 -1706 -385 -1702
rect -215 -1706 -214 -1702
rect -212 -1706 -210 -1702
rect -206 -1706 -204 -1702
rect -202 -1706 -201 -1702
rect -189 -1706 -188 -1702
rect -186 -1706 -180 -1702
rect -178 -1706 -177 -1702
rect -165 -1706 -164 -1702
rect -162 -1706 -156 -1702
rect -154 -1706 -152 -1702
rect -148 -1706 -146 -1702
rect -144 -1706 -138 -1702
rect -136 -1706 -135 -1702
rect -123 -1706 -122 -1702
rect -120 -1706 -114 -1702
rect -112 -1706 -110 -1702
rect -106 -1706 -104 -1702
rect -102 -1706 -96 -1702
rect -94 -1706 -93 -1702
rect -81 -1706 -80 -1702
rect -78 -1706 -72 -1702
rect -70 -1706 -68 -1702
rect -64 -1706 -62 -1702
rect -60 -1706 -54 -1702
rect -52 -1706 -51 -1702
rect -39 -1706 -38 -1702
rect -36 -1706 -30 -1702
rect -28 -1706 -27 -1702
rect 213 -1706 214 -1702
rect 216 -1706 218 -1702
rect 222 -1706 224 -1702
rect 226 -1706 227 -1702
rect 239 -1706 240 -1702
rect 242 -1706 248 -1702
rect 250 -1706 251 -1702
rect 263 -1706 264 -1702
rect 266 -1706 272 -1702
rect 274 -1706 276 -1702
rect 280 -1706 282 -1702
rect 284 -1706 290 -1702
rect 292 -1706 293 -1702
rect 305 -1706 306 -1702
rect 308 -1706 314 -1702
rect 316 -1706 318 -1702
rect 322 -1706 324 -1702
rect 326 -1706 332 -1702
rect 334 -1706 335 -1702
rect 347 -1706 348 -1702
rect 350 -1706 356 -1702
rect 358 -1706 360 -1702
rect 364 -1706 366 -1702
rect 368 -1706 374 -1702
rect 376 -1706 377 -1702
rect 389 -1706 390 -1702
rect 392 -1706 398 -1702
rect 400 -1706 401 -1702
rect 569 -1706 570 -1702
rect 572 -1706 574 -1702
rect 578 -1706 580 -1702
rect 582 -1706 583 -1702
rect 595 -1706 596 -1702
rect 598 -1706 604 -1702
rect 606 -1706 607 -1702
rect 619 -1706 620 -1702
rect 622 -1706 628 -1702
rect 630 -1706 632 -1702
rect 636 -1706 638 -1702
rect 640 -1706 646 -1702
rect 648 -1706 649 -1702
rect 661 -1706 662 -1702
rect 664 -1706 670 -1702
rect 672 -1706 674 -1702
rect 678 -1706 680 -1702
rect 682 -1706 688 -1702
rect 690 -1706 691 -1702
rect 703 -1706 704 -1702
rect 706 -1706 712 -1702
rect 714 -1706 716 -1702
rect 720 -1706 722 -1702
rect 724 -1706 730 -1702
rect 732 -1706 733 -1702
rect 745 -1706 746 -1702
rect 748 -1706 754 -1702
rect 756 -1706 757 -1702
rect 967 -1706 968 -1702
rect 970 -1706 972 -1702
rect 976 -1706 978 -1702
rect 980 -1706 981 -1702
rect 993 -1706 994 -1702
rect 996 -1706 1002 -1702
rect 1004 -1706 1005 -1702
rect 1017 -1706 1018 -1702
rect 1020 -1706 1026 -1702
rect 1028 -1706 1030 -1702
rect 1034 -1706 1036 -1702
rect 1038 -1706 1044 -1702
rect 1046 -1706 1047 -1702
rect 1059 -1706 1060 -1702
rect 1062 -1706 1068 -1702
rect 1070 -1706 1072 -1702
rect 1076 -1706 1078 -1702
rect 1080 -1706 1086 -1702
rect 1088 -1706 1089 -1702
rect 1101 -1706 1102 -1702
rect 1104 -1706 1110 -1702
rect 1112 -1706 1114 -1702
rect 1118 -1706 1120 -1702
rect 1122 -1706 1128 -1702
rect 1130 -1706 1131 -1702
rect 1143 -1706 1144 -1702
rect 1146 -1706 1152 -1702
rect 1154 -1706 1155 -1702
rect 1325 -1706 1326 -1702
rect 1328 -1706 1330 -1702
rect 1334 -1706 1336 -1702
rect 1338 -1706 1339 -1702
rect 1351 -1706 1352 -1702
rect 1354 -1706 1360 -1702
rect 1362 -1706 1363 -1702
rect 1375 -1706 1376 -1702
rect 1378 -1706 1384 -1702
rect 1386 -1706 1388 -1702
rect 1392 -1706 1394 -1702
rect 1396 -1706 1402 -1702
rect 1404 -1706 1405 -1702
rect 1417 -1706 1418 -1702
rect 1420 -1706 1426 -1702
rect 1428 -1706 1430 -1702
rect 1434 -1706 1436 -1702
rect 1438 -1706 1444 -1702
rect 1446 -1706 1447 -1702
rect 1459 -1706 1460 -1702
rect 1462 -1706 1468 -1702
rect 1470 -1706 1472 -1702
rect 1476 -1706 1478 -1702
rect 1480 -1706 1486 -1702
rect 1488 -1706 1489 -1702
rect 1501 -1706 1502 -1702
rect 1504 -1706 1510 -1702
rect 1512 -1706 1513 -1702
rect -1256 -1827 -1255 -1823
rect -1253 -1827 -1251 -1823
rect -1247 -1827 -1245 -1823
rect -1243 -1827 -1242 -1823
rect -1230 -1827 -1229 -1823
rect -1227 -1827 -1221 -1823
rect -1219 -1827 -1218 -1823
rect -1206 -1827 -1205 -1823
rect -1203 -1827 -1197 -1823
rect -1195 -1827 -1193 -1823
rect -1189 -1827 -1187 -1823
rect -1185 -1827 -1179 -1823
rect -1177 -1827 -1176 -1823
rect -1164 -1827 -1163 -1823
rect -1161 -1827 -1155 -1823
rect -1153 -1827 -1151 -1823
rect -1147 -1827 -1145 -1823
rect -1143 -1827 -1137 -1823
rect -1135 -1827 -1134 -1823
rect -1122 -1827 -1121 -1823
rect -1119 -1827 -1113 -1823
rect -1111 -1827 -1109 -1823
rect -1105 -1827 -1103 -1823
rect -1101 -1827 -1095 -1823
rect -1093 -1827 -1092 -1823
rect -1080 -1827 -1079 -1823
rect -1077 -1827 -1071 -1823
rect -1069 -1827 -1068 -1823
rect -1025 -1827 -1024 -1823
rect -1022 -1827 -1021 -1823
rect -931 -1827 -930 -1823
rect -928 -1827 -926 -1823
rect -922 -1827 -920 -1823
rect -918 -1827 -917 -1823
rect -905 -1827 -904 -1823
rect -902 -1827 -896 -1823
rect -894 -1827 -893 -1823
rect -881 -1827 -880 -1823
rect -878 -1827 -872 -1823
rect -870 -1827 -868 -1823
rect -864 -1827 -862 -1823
rect -860 -1827 -854 -1823
rect -852 -1827 -851 -1823
rect -839 -1827 -838 -1823
rect -836 -1827 -830 -1823
rect -828 -1827 -826 -1823
rect -822 -1827 -820 -1823
rect -818 -1827 -812 -1823
rect -810 -1827 -809 -1823
rect -797 -1827 -796 -1823
rect -794 -1827 -788 -1823
rect -786 -1827 -784 -1823
rect -780 -1827 -778 -1823
rect -776 -1827 -770 -1823
rect -768 -1827 -767 -1823
rect -755 -1827 -754 -1823
rect -752 -1827 -746 -1823
rect -744 -1827 -743 -1823
rect -573 -1827 -572 -1823
rect -570 -1827 -568 -1823
rect -564 -1827 -562 -1823
rect -560 -1827 -559 -1823
rect -547 -1827 -546 -1823
rect -544 -1827 -538 -1823
rect -536 -1827 -535 -1823
rect -523 -1827 -522 -1823
rect -520 -1827 -514 -1823
rect -512 -1827 -510 -1823
rect -506 -1827 -504 -1823
rect -502 -1827 -496 -1823
rect -494 -1827 -493 -1823
rect -481 -1827 -480 -1823
rect -478 -1827 -472 -1823
rect -470 -1827 -468 -1823
rect -464 -1827 -462 -1823
rect -460 -1827 -454 -1823
rect -452 -1827 -451 -1823
rect -439 -1827 -438 -1823
rect -436 -1827 -430 -1823
rect -428 -1827 -426 -1823
rect -422 -1827 -420 -1823
rect -418 -1827 -412 -1823
rect -410 -1827 -409 -1823
rect -397 -1827 -396 -1823
rect -394 -1827 -388 -1823
rect -386 -1827 -385 -1823
rect -328 -1827 -327 -1823
rect -325 -1827 -324 -1823
rect -215 -1827 -214 -1823
rect -212 -1827 -210 -1823
rect -206 -1827 -204 -1823
rect -202 -1827 -201 -1823
rect -189 -1827 -188 -1823
rect -186 -1827 -180 -1823
rect -178 -1827 -177 -1823
rect -165 -1827 -164 -1823
rect -162 -1827 -156 -1823
rect -154 -1827 -152 -1823
rect -148 -1827 -146 -1823
rect -144 -1827 -138 -1823
rect -136 -1827 -135 -1823
rect -123 -1827 -122 -1823
rect -120 -1827 -114 -1823
rect -112 -1827 -110 -1823
rect -106 -1827 -104 -1823
rect -102 -1827 -96 -1823
rect -94 -1827 -93 -1823
rect -81 -1827 -80 -1823
rect -78 -1827 -72 -1823
rect -70 -1827 -68 -1823
rect -64 -1827 -62 -1823
rect -60 -1827 -54 -1823
rect -52 -1827 -51 -1823
rect -39 -1827 -38 -1823
rect -36 -1827 -30 -1823
rect -28 -1827 -27 -1823
rect 213 -1827 214 -1823
rect 216 -1827 218 -1823
rect 222 -1827 224 -1823
rect 226 -1827 227 -1823
rect 239 -1827 240 -1823
rect 242 -1827 248 -1823
rect 250 -1827 251 -1823
rect 263 -1827 264 -1823
rect 266 -1827 272 -1823
rect 274 -1827 276 -1823
rect 280 -1827 282 -1823
rect 284 -1827 290 -1823
rect 292 -1827 293 -1823
rect 305 -1827 306 -1823
rect 308 -1827 314 -1823
rect 316 -1827 318 -1823
rect 322 -1827 324 -1823
rect 326 -1827 332 -1823
rect 334 -1827 335 -1823
rect 347 -1827 348 -1823
rect 350 -1827 356 -1823
rect 358 -1827 360 -1823
rect 364 -1827 366 -1823
rect 368 -1827 374 -1823
rect 376 -1827 377 -1823
rect 389 -1827 390 -1823
rect 392 -1827 398 -1823
rect 400 -1827 401 -1823
rect 468 -1827 469 -1823
rect 471 -1827 472 -1823
rect 569 -1827 570 -1823
rect 572 -1827 574 -1823
rect 578 -1827 580 -1823
rect 582 -1827 583 -1823
rect 595 -1827 596 -1823
rect 598 -1827 604 -1823
rect 606 -1827 607 -1823
rect 619 -1827 620 -1823
rect 622 -1827 628 -1823
rect 630 -1827 632 -1823
rect 636 -1827 638 -1823
rect 640 -1827 646 -1823
rect 648 -1827 649 -1823
rect 661 -1827 662 -1823
rect 664 -1827 670 -1823
rect 672 -1827 674 -1823
rect 678 -1827 680 -1823
rect 682 -1827 688 -1823
rect 690 -1827 691 -1823
rect 703 -1827 704 -1823
rect 706 -1827 712 -1823
rect 714 -1827 716 -1823
rect 720 -1827 722 -1823
rect 724 -1827 730 -1823
rect 732 -1827 733 -1823
rect 745 -1827 746 -1823
rect 748 -1827 754 -1823
rect 756 -1827 757 -1823
rect 967 -1827 968 -1823
rect 970 -1827 972 -1823
rect 976 -1827 978 -1823
rect 980 -1827 981 -1823
rect 993 -1827 994 -1823
rect 996 -1827 1002 -1823
rect 1004 -1827 1005 -1823
rect 1017 -1827 1018 -1823
rect 1020 -1827 1026 -1823
rect 1028 -1827 1030 -1823
rect 1034 -1827 1036 -1823
rect 1038 -1827 1044 -1823
rect 1046 -1827 1047 -1823
rect 1059 -1827 1060 -1823
rect 1062 -1827 1068 -1823
rect 1070 -1827 1072 -1823
rect 1076 -1827 1078 -1823
rect 1080 -1827 1086 -1823
rect 1088 -1827 1089 -1823
rect 1101 -1827 1102 -1823
rect 1104 -1827 1110 -1823
rect 1112 -1827 1114 -1823
rect 1118 -1827 1120 -1823
rect 1122 -1827 1128 -1823
rect 1130 -1827 1131 -1823
rect 1143 -1827 1144 -1823
rect 1146 -1827 1152 -1823
rect 1154 -1827 1155 -1823
rect 1207 -1827 1208 -1823
rect 1210 -1827 1211 -1823
rect 1325 -1827 1326 -1823
rect 1328 -1827 1330 -1823
rect 1334 -1827 1336 -1823
rect 1338 -1827 1339 -1823
rect 1351 -1827 1352 -1823
rect 1354 -1827 1360 -1823
rect 1362 -1827 1363 -1823
rect 1375 -1827 1376 -1823
rect 1378 -1827 1384 -1823
rect 1386 -1827 1388 -1823
rect 1392 -1827 1394 -1823
rect 1396 -1827 1402 -1823
rect 1404 -1827 1405 -1823
rect 1417 -1827 1418 -1823
rect 1420 -1827 1426 -1823
rect 1428 -1827 1430 -1823
rect 1434 -1827 1436 -1823
rect 1438 -1827 1444 -1823
rect 1446 -1827 1447 -1823
rect 1459 -1827 1460 -1823
rect 1462 -1827 1468 -1823
rect 1470 -1827 1472 -1823
rect 1476 -1827 1478 -1823
rect 1480 -1827 1486 -1823
rect 1488 -1827 1489 -1823
rect 1501 -1827 1502 -1823
rect 1504 -1827 1510 -1823
rect 1512 -1827 1513 -1823
rect -1256 -1942 -1255 -1938
rect -1253 -1942 -1251 -1938
rect -1247 -1942 -1245 -1938
rect -1243 -1942 -1242 -1938
rect -1230 -1942 -1229 -1938
rect -1227 -1942 -1221 -1938
rect -1219 -1942 -1218 -1938
rect -1206 -1942 -1205 -1938
rect -1203 -1942 -1197 -1938
rect -1195 -1942 -1193 -1938
rect -1189 -1942 -1187 -1938
rect -1185 -1942 -1179 -1938
rect -1177 -1942 -1176 -1938
rect -1164 -1942 -1163 -1938
rect -1161 -1942 -1155 -1938
rect -1153 -1942 -1151 -1938
rect -1147 -1942 -1145 -1938
rect -1143 -1942 -1137 -1938
rect -1135 -1942 -1134 -1938
rect -1122 -1942 -1121 -1938
rect -1119 -1942 -1113 -1938
rect -1111 -1942 -1109 -1938
rect -1105 -1942 -1103 -1938
rect -1101 -1942 -1095 -1938
rect -1093 -1942 -1092 -1938
rect -1080 -1942 -1079 -1938
rect -1077 -1942 -1071 -1938
rect -1069 -1942 -1068 -1938
rect -1025 -1942 -1024 -1938
rect -1022 -1942 -1021 -1938
rect -669 -1942 -668 -1934
rect -666 -1942 -665 -1934
rect -328 -1942 -327 -1938
rect -325 -1942 -324 -1938
rect 468 -1942 469 -1938
rect 471 -1942 472 -1938
rect 845 -1942 846 -1934
rect 848 -1942 849 -1934
rect 1207 -1942 1208 -1938
rect 1210 -1942 1211 -1938
rect -1335 -2054 -1334 -2050
rect -1332 -2054 -1326 -2050
rect -1324 -2054 -1322 -2050
rect -1318 -2054 -1316 -2050
rect -1314 -2054 -1313 -2050
rect -931 -2054 -930 -2050
rect -928 -2054 -922 -2050
rect -920 -2054 -918 -2050
rect -914 -2054 -912 -2050
rect -910 -2054 -909 -2050
rect -573 -2054 -572 -2050
rect -570 -2054 -564 -2050
rect -562 -2054 -560 -2050
rect -556 -2054 -554 -2050
rect -552 -2054 -551 -2050
rect -215 -2054 -214 -2050
rect -212 -2054 -206 -2050
rect -204 -2054 -202 -2050
rect -198 -2054 -196 -2050
rect -194 -2054 -193 -2050
rect 213 -2054 214 -2050
rect 216 -2054 222 -2050
rect 224 -2054 226 -2050
rect 230 -2054 232 -2050
rect 234 -2054 235 -2050
rect 569 -2054 570 -2050
rect 572 -2054 578 -2050
rect 580 -2054 582 -2050
rect 586 -2054 588 -2050
rect 590 -2054 591 -2050
rect 967 -2054 968 -2050
rect 970 -2054 976 -2050
rect 978 -2054 980 -2050
rect 984 -2054 986 -2050
rect 988 -2054 989 -2050
rect 1325 -2054 1326 -2050
rect 1328 -2054 1334 -2050
rect 1336 -2054 1338 -2050
rect 1342 -2054 1344 -2050
rect 1346 -2054 1347 -2050
rect -1256 -2173 -1255 -2169
rect -1253 -2173 -1251 -2169
rect -1247 -2173 -1245 -2169
rect -1243 -2173 -1242 -2169
rect -1230 -2173 -1229 -2169
rect -1227 -2173 -1225 -2169
rect -1221 -2173 -1219 -2169
rect -1217 -2173 -1211 -2169
rect -1209 -2173 -1207 -2169
rect -1203 -2173 -1201 -2169
rect -1199 -2173 -1198 -2169
rect -1186 -2173 -1185 -2169
rect -1183 -2173 -1177 -2169
rect -1175 -2173 -1173 -2169
rect -1169 -2173 -1167 -2169
rect -1165 -2173 -1164 -2169
rect -931 -2173 -930 -2169
rect -928 -2173 -926 -2169
rect -922 -2173 -920 -2169
rect -918 -2173 -917 -2169
rect -905 -2173 -904 -2169
rect -902 -2173 -900 -2169
rect -896 -2173 -894 -2169
rect -892 -2173 -891 -2169
rect -879 -2173 -878 -2169
rect -876 -2173 -875 -2169
rect -871 -2173 -868 -2169
rect -866 -2173 -860 -2169
rect -858 -2173 -857 -2169
rect -853 -2173 -850 -2169
rect -848 -2173 -847 -2169
rect -835 -2173 -834 -2169
rect -832 -2173 -826 -2169
rect -824 -2173 -822 -2169
rect -818 -2173 -816 -2169
rect -814 -2173 -813 -2169
rect -801 -2173 -800 -2169
rect -798 -2173 -796 -2169
rect -792 -2173 -790 -2169
rect -788 -2173 -782 -2169
rect -780 -2173 -778 -2169
rect -774 -2173 -772 -2169
rect -770 -2173 -769 -2169
rect -757 -2173 -756 -2169
rect -754 -2173 -748 -2169
rect -746 -2173 -745 -2169
rect -733 -2173 -732 -2169
rect -730 -2173 -725 -2169
rect -721 -2173 -716 -2169
rect -714 -2173 -713 -2169
rect -709 -2173 -708 -2169
rect -706 -2173 -704 -2169
rect -700 -2173 -698 -2169
rect -696 -2173 -695 -2169
rect -573 -2173 -572 -2169
rect -570 -2173 -568 -2169
rect -564 -2173 -562 -2169
rect -560 -2173 -559 -2169
rect -547 -2173 -546 -2169
rect -544 -2173 -542 -2169
rect -538 -2173 -536 -2169
rect -534 -2173 -533 -2169
rect -521 -2173 -520 -2169
rect -518 -2173 -517 -2169
rect -513 -2173 -510 -2169
rect -508 -2173 -502 -2169
rect -500 -2173 -499 -2169
rect -495 -2173 -492 -2169
rect -490 -2173 -489 -2169
rect -477 -2173 -476 -2169
rect -474 -2173 -468 -2169
rect -466 -2173 -464 -2169
rect -460 -2173 -458 -2169
rect -456 -2173 -455 -2169
rect -443 -2173 -442 -2169
rect -440 -2173 -438 -2169
rect -434 -2173 -432 -2169
rect -430 -2173 -424 -2169
rect -422 -2173 -420 -2169
rect -416 -2173 -414 -2169
rect -412 -2173 -411 -2169
rect -399 -2173 -398 -2169
rect -396 -2173 -390 -2169
rect -388 -2173 -387 -2169
rect -375 -2173 -374 -2169
rect -372 -2173 -367 -2169
rect -363 -2173 -358 -2169
rect -356 -2173 -355 -2169
rect -351 -2173 -350 -2169
rect -348 -2173 -346 -2169
rect -342 -2173 -340 -2169
rect -338 -2173 -337 -2169
rect -215 -2173 -214 -2169
rect -212 -2173 -210 -2169
rect -206 -2173 -204 -2169
rect -202 -2173 -201 -2169
rect -189 -2173 -188 -2169
rect -186 -2173 -184 -2169
rect -180 -2173 -178 -2169
rect -176 -2173 -175 -2169
rect -163 -2173 -162 -2169
rect -160 -2173 -159 -2169
rect -155 -2173 -152 -2169
rect -150 -2173 -144 -2169
rect -142 -2173 -141 -2169
rect -137 -2173 -134 -2169
rect -132 -2173 -131 -2169
rect -119 -2173 -118 -2169
rect -116 -2173 -110 -2169
rect -108 -2173 -106 -2169
rect -102 -2173 -100 -2169
rect -98 -2173 -97 -2169
rect -85 -2173 -84 -2169
rect -82 -2173 -80 -2169
rect -76 -2173 -74 -2169
rect -72 -2173 -66 -2169
rect -64 -2173 -62 -2169
rect -58 -2173 -56 -2169
rect -54 -2173 -53 -2169
rect -41 -2173 -40 -2169
rect -38 -2173 -32 -2169
rect -30 -2173 -29 -2169
rect -17 -2173 -16 -2169
rect -14 -2173 -9 -2169
rect -5 -2173 0 -2169
rect 2 -2173 3 -2169
rect 7 -2173 8 -2169
rect 10 -2173 12 -2169
rect 16 -2173 18 -2169
rect 20 -2173 21 -2169
rect 213 -2173 214 -2169
rect 216 -2173 218 -2169
rect 222 -2173 224 -2169
rect 226 -2173 227 -2169
rect 239 -2173 240 -2169
rect 242 -2173 244 -2169
rect 248 -2173 250 -2169
rect 252 -2173 253 -2169
rect 265 -2173 266 -2169
rect 268 -2173 269 -2169
rect 273 -2173 276 -2169
rect 278 -2173 284 -2169
rect 286 -2173 287 -2169
rect 291 -2173 294 -2169
rect 296 -2173 297 -2169
rect 309 -2173 310 -2169
rect 312 -2173 318 -2169
rect 320 -2173 322 -2169
rect 326 -2173 328 -2169
rect 330 -2173 331 -2169
rect 343 -2173 344 -2169
rect 346 -2173 348 -2169
rect 352 -2173 354 -2169
rect 356 -2173 362 -2169
rect 364 -2173 366 -2169
rect 370 -2173 372 -2169
rect 374 -2173 375 -2169
rect 387 -2173 388 -2169
rect 390 -2173 396 -2169
rect 398 -2173 399 -2169
rect 411 -2173 412 -2169
rect 414 -2173 419 -2169
rect 423 -2173 428 -2169
rect 430 -2173 431 -2169
rect 435 -2173 436 -2169
rect 438 -2173 440 -2169
rect 444 -2173 446 -2169
rect 448 -2173 449 -2169
rect 569 -2173 570 -2169
rect 572 -2173 574 -2169
rect 578 -2173 580 -2169
rect 582 -2173 583 -2169
rect 595 -2173 596 -2169
rect 598 -2173 600 -2169
rect 604 -2173 606 -2169
rect 608 -2173 609 -2169
rect 621 -2173 622 -2169
rect 624 -2173 625 -2169
rect 629 -2173 632 -2169
rect 634 -2173 640 -2169
rect 642 -2173 643 -2169
rect 647 -2173 650 -2169
rect 652 -2173 653 -2169
rect 665 -2173 666 -2169
rect 668 -2173 674 -2169
rect 676 -2173 678 -2169
rect 682 -2173 684 -2169
rect 686 -2173 687 -2169
rect 699 -2173 700 -2169
rect 702 -2173 704 -2169
rect 708 -2173 710 -2169
rect 712 -2173 718 -2169
rect 720 -2173 722 -2169
rect 726 -2173 728 -2169
rect 730 -2173 731 -2169
rect 743 -2173 744 -2169
rect 746 -2173 752 -2169
rect 754 -2173 755 -2169
rect 767 -2173 768 -2169
rect 770 -2173 775 -2169
rect 779 -2173 784 -2169
rect 786 -2173 787 -2169
rect 791 -2173 792 -2169
rect 794 -2173 796 -2169
rect 800 -2173 802 -2169
rect 804 -2173 805 -2169
rect 967 -2173 968 -2169
rect 970 -2173 972 -2169
rect 976 -2173 978 -2169
rect 980 -2173 981 -2169
rect 993 -2173 994 -2169
rect 996 -2173 998 -2169
rect 1002 -2173 1004 -2169
rect 1006 -2173 1007 -2169
rect 1019 -2173 1020 -2169
rect 1022 -2173 1023 -2169
rect 1027 -2173 1030 -2169
rect 1032 -2173 1038 -2169
rect 1040 -2173 1041 -2169
rect 1045 -2173 1048 -2169
rect 1050 -2173 1051 -2169
rect 1063 -2173 1064 -2169
rect 1066 -2173 1072 -2169
rect 1074 -2173 1076 -2169
rect 1080 -2173 1082 -2169
rect 1084 -2173 1085 -2169
rect 1097 -2173 1098 -2169
rect 1100 -2173 1102 -2169
rect 1106 -2173 1108 -2169
rect 1110 -2173 1116 -2169
rect 1118 -2173 1120 -2169
rect 1124 -2173 1126 -2169
rect 1128 -2173 1129 -2169
rect 1141 -2173 1142 -2169
rect 1144 -2173 1150 -2169
rect 1152 -2173 1153 -2169
rect 1165 -2173 1166 -2169
rect 1168 -2173 1173 -2169
rect 1177 -2173 1182 -2169
rect 1184 -2173 1185 -2169
rect 1189 -2173 1190 -2169
rect 1192 -2173 1194 -2169
rect 1198 -2173 1200 -2169
rect 1202 -2173 1203 -2169
rect 1325 -2173 1326 -2169
rect 1328 -2173 1330 -2169
rect 1334 -2173 1336 -2169
rect 1338 -2173 1339 -2169
rect 1351 -2173 1352 -2169
rect 1354 -2173 1356 -2169
rect 1360 -2173 1362 -2169
rect 1364 -2173 1365 -2169
rect 1377 -2173 1378 -2169
rect 1380 -2173 1381 -2169
rect 1385 -2173 1388 -2169
rect 1390 -2173 1396 -2169
rect 1398 -2173 1399 -2169
rect 1403 -2173 1406 -2169
rect 1408 -2173 1409 -2169
rect 1421 -2173 1422 -2169
rect 1424 -2173 1430 -2169
rect 1432 -2173 1434 -2169
rect 1438 -2173 1440 -2169
rect 1442 -2173 1443 -2169
rect 1455 -2173 1456 -2169
rect 1458 -2173 1460 -2169
rect 1464 -2173 1466 -2169
rect 1468 -2173 1474 -2169
rect 1476 -2173 1478 -2169
rect 1482 -2173 1484 -2169
rect 1486 -2173 1487 -2169
rect 1499 -2173 1500 -2169
rect 1502 -2173 1508 -2169
rect 1510 -2173 1511 -2169
rect 1523 -2173 1524 -2169
rect 1526 -2173 1531 -2169
rect 1535 -2173 1540 -2169
rect 1542 -2173 1543 -2169
rect 1547 -2173 1548 -2169
rect 1550 -2173 1552 -2169
rect 1556 -2173 1558 -2169
rect 1560 -2173 1561 -2169
rect -1260 -2317 -1259 -2313
rect -1257 -2317 -1255 -2313
rect -1251 -2317 -1249 -2313
rect -1247 -2317 -1246 -2313
rect -1234 -2317 -1233 -2313
rect -1231 -2317 -1225 -2313
rect -1223 -2317 -1222 -2313
rect -1210 -2317 -1209 -2313
rect -1207 -2317 -1201 -2313
rect -1199 -2317 -1197 -2313
rect -1193 -2317 -1191 -2313
rect -1189 -2317 -1183 -2313
rect -1181 -2317 -1180 -2313
rect -1168 -2317 -1167 -2313
rect -1165 -2317 -1159 -2313
rect -1157 -2317 -1155 -2313
rect -1151 -2317 -1149 -2313
rect -1147 -2317 -1141 -2313
rect -1139 -2317 -1138 -2313
rect -1126 -2317 -1125 -2313
rect -1123 -2317 -1117 -2313
rect -1115 -2317 -1113 -2313
rect -1109 -2317 -1107 -2313
rect -1105 -2317 -1099 -2313
rect -1097 -2317 -1096 -2313
rect -1084 -2317 -1083 -2313
rect -1081 -2317 -1075 -2313
rect -1073 -2317 -1072 -2313
rect -931 -2317 -930 -2313
rect -928 -2317 -926 -2313
rect -922 -2317 -920 -2313
rect -918 -2317 -917 -2313
rect -905 -2317 -904 -2313
rect -902 -2317 -896 -2313
rect -894 -2317 -893 -2313
rect -881 -2317 -880 -2313
rect -878 -2317 -872 -2313
rect -870 -2317 -868 -2313
rect -864 -2317 -862 -2313
rect -860 -2317 -854 -2313
rect -852 -2317 -851 -2313
rect -839 -2317 -838 -2313
rect -836 -2317 -830 -2313
rect -828 -2317 -826 -2313
rect -822 -2317 -820 -2313
rect -818 -2317 -812 -2313
rect -810 -2317 -809 -2313
rect -797 -2317 -796 -2313
rect -794 -2317 -788 -2313
rect -786 -2317 -784 -2313
rect -780 -2317 -778 -2313
rect -776 -2317 -770 -2313
rect -768 -2317 -767 -2313
rect -755 -2317 -754 -2313
rect -752 -2317 -746 -2313
rect -744 -2317 -743 -2313
rect -573 -2317 -572 -2313
rect -570 -2317 -568 -2313
rect -564 -2317 -562 -2313
rect -560 -2317 -559 -2313
rect -547 -2317 -546 -2313
rect -544 -2317 -538 -2313
rect -536 -2317 -535 -2313
rect -523 -2317 -522 -2313
rect -520 -2317 -514 -2313
rect -512 -2317 -510 -2313
rect -506 -2317 -504 -2313
rect -502 -2317 -496 -2313
rect -494 -2317 -493 -2313
rect -481 -2317 -480 -2313
rect -478 -2317 -472 -2313
rect -470 -2317 -468 -2313
rect -464 -2317 -462 -2313
rect -460 -2317 -454 -2313
rect -452 -2317 -451 -2313
rect -439 -2317 -438 -2313
rect -436 -2317 -430 -2313
rect -428 -2317 -426 -2313
rect -422 -2317 -420 -2313
rect -418 -2317 -412 -2313
rect -410 -2317 -409 -2313
rect -397 -2317 -396 -2313
rect -394 -2317 -388 -2313
rect -386 -2317 -385 -2313
rect -215 -2317 -214 -2313
rect -212 -2317 -210 -2313
rect -206 -2317 -204 -2313
rect -202 -2317 -201 -2313
rect -189 -2317 -188 -2313
rect -186 -2317 -180 -2313
rect -178 -2317 -177 -2313
rect -165 -2317 -164 -2313
rect -162 -2317 -156 -2313
rect -154 -2317 -152 -2313
rect -148 -2317 -146 -2313
rect -144 -2317 -138 -2313
rect -136 -2317 -135 -2313
rect -123 -2317 -122 -2313
rect -120 -2317 -114 -2313
rect -112 -2317 -110 -2313
rect -106 -2317 -104 -2313
rect -102 -2317 -96 -2313
rect -94 -2317 -93 -2313
rect -81 -2317 -80 -2313
rect -78 -2317 -72 -2313
rect -70 -2317 -68 -2313
rect -64 -2317 -62 -2313
rect -60 -2317 -54 -2313
rect -52 -2317 -51 -2313
rect -39 -2317 -38 -2313
rect -36 -2317 -30 -2313
rect -28 -2317 -27 -2313
rect 213 -2317 214 -2313
rect 216 -2317 218 -2313
rect 222 -2317 224 -2313
rect 226 -2317 227 -2313
rect 239 -2317 240 -2313
rect 242 -2317 248 -2313
rect 250 -2317 251 -2313
rect 263 -2317 264 -2313
rect 266 -2317 272 -2313
rect 274 -2317 276 -2313
rect 280 -2317 282 -2313
rect 284 -2317 290 -2313
rect 292 -2317 293 -2313
rect 305 -2317 306 -2313
rect 308 -2317 314 -2313
rect 316 -2317 318 -2313
rect 322 -2317 324 -2313
rect 326 -2317 332 -2313
rect 334 -2317 335 -2313
rect 347 -2317 348 -2313
rect 350 -2317 356 -2313
rect 358 -2317 360 -2313
rect 364 -2317 366 -2313
rect 368 -2317 374 -2313
rect 376 -2317 377 -2313
rect 389 -2317 390 -2313
rect 392 -2317 398 -2313
rect 400 -2317 401 -2313
rect 569 -2317 570 -2313
rect 572 -2317 574 -2313
rect 578 -2317 580 -2313
rect 582 -2317 583 -2313
rect 595 -2317 596 -2313
rect 598 -2317 604 -2313
rect 606 -2317 607 -2313
rect 619 -2317 620 -2313
rect 622 -2317 628 -2313
rect 630 -2317 632 -2313
rect 636 -2317 638 -2313
rect 640 -2317 646 -2313
rect 648 -2317 649 -2313
rect 661 -2317 662 -2313
rect 664 -2317 670 -2313
rect 672 -2317 674 -2313
rect 678 -2317 680 -2313
rect 682 -2317 688 -2313
rect 690 -2317 691 -2313
rect 703 -2317 704 -2313
rect 706 -2317 712 -2313
rect 714 -2317 716 -2313
rect 720 -2317 722 -2313
rect 724 -2317 730 -2313
rect 732 -2317 733 -2313
rect 745 -2317 746 -2313
rect 748 -2317 754 -2313
rect 756 -2317 757 -2313
rect -1260 -2448 -1259 -2444
rect -1257 -2448 -1255 -2444
rect -1251 -2448 -1249 -2444
rect -1247 -2448 -1246 -2444
rect -1234 -2448 -1233 -2444
rect -1231 -2448 -1225 -2444
rect -1223 -2448 -1222 -2444
rect -1210 -2448 -1209 -2444
rect -1207 -2448 -1201 -2444
rect -1199 -2448 -1197 -2444
rect -1193 -2448 -1191 -2444
rect -1189 -2448 -1183 -2444
rect -1181 -2448 -1180 -2444
rect -1168 -2448 -1167 -2444
rect -1165 -2448 -1159 -2444
rect -1157 -2448 -1155 -2444
rect -1151 -2448 -1149 -2444
rect -1147 -2448 -1141 -2444
rect -1139 -2448 -1138 -2444
rect -1126 -2448 -1125 -2444
rect -1123 -2448 -1117 -2444
rect -1115 -2448 -1113 -2444
rect -1109 -2448 -1107 -2444
rect -1105 -2448 -1099 -2444
rect -1097 -2448 -1096 -2444
rect -1084 -2448 -1083 -2444
rect -1081 -2448 -1075 -2444
rect -1073 -2448 -1072 -2444
rect -931 -2448 -930 -2444
rect -928 -2448 -926 -2444
rect -922 -2448 -920 -2444
rect -918 -2448 -917 -2444
rect -905 -2448 -904 -2444
rect -902 -2448 -896 -2444
rect -894 -2448 -893 -2444
rect -881 -2448 -880 -2444
rect -878 -2448 -872 -2444
rect -870 -2448 -868 -2444
rect -864 -2448 -862 -2444
rect -860 -2448 -854 -2444
rect -852 -2448 -851 -2444
rect -839 -2448 -838 -2444
rect -836 -2448 -830 -2444
rect -828 -2448 -826 -2444
rect -822 -2448 -820 -2444
rect -818 -2448 -812 -2444
rect -810 -2448 -809 -2444
rect -797 -2448 -796 -2444
rect -794 -2448 -788 -2444
rect -786 -2448 -784 -2444
rect -780 -2448 -778 -2444
rect -776 -2448 -770 -2444
rect -768 -2448 -767 -2444
rect -755 -2448 -754 -2444
rect -752 -2448 -746 -2444
rect -744 -2448 -743 -2444
rect -573 -2448 -572 -2444
rect -570 -2448 -568 -2444
rect -564 -2448 -562 -2444
rect -560 -2448 -559 -2444
rect -547 -2448 -546 -2444
rect -544 -2448 -538 -2444
rect -536 -2448 -535 -2444
rect -523 -2448 -522 -2444
rect -520 -2448 -514 -2444
rect -512 -2448 -510 -2444
rect -506 -2448 -504 -2444
rect -502 -2448 -496 -2444
rect -494 -2448 -493 -2444
rect -481 -2448 -480 -2444
rect -478 -2448 -472 -2444
rect -470 -2448 -468 -2444
rect -464 -2448 -462 -2444
rect -460 -2448 -454 -2444
rect -452 -2448 -451 -2444
rect -439 -2448 -438 -2444
rect -436 -2448 -430 -2444
rect -428 -2448 -426 -2444
rect -422 -2448 -420 -2444
rect -418 -2448 -412 -2444
rect -410 -2448 -409 -2444
rect -397 -2448 -396 -2444
rect -394 -2448 -388 -2444
rect -386 -2448 -385 -2444
rect -215 -2448 -214 -2444
rect -212 -2448 -210 -2444
rect -206 -2448 -204 -2444
rect -202 -2448 -201 -2444
rect -189 -2448 -188 -2444
rect -186 -2448 -180 -2444
rect -178 -2448 -177 -2444
rect -165 -2448 -164 -2444
rect -162 -2448 -156 -2444
rect -154 -2448 -152 -2444
rect -148 -2448 -146 -2444
rect -144 -2448 -138 -2444
rect -136 -2448 -135 -2444
rect -123 -2448 -122 -2444
rect -120 -2448 -114 -2444
rect -112 -2448 -110 -2444
rect -106 -2448 -104 -2444
rect -102 -2448 -96 -2444
rect -94 -2448 -93 -2444
rect -81 -2448 -80 -2444
rect -78 -2448 -72 -2444
rect -70 -2448 -68 -2444
rect -64 -2448 -62 -2444
rect -60 -2448 -54 -2444
rect -52 -2448 -51 -2444
rect -39 -2448 -38 -2444
rect -36 -2448 -30 -2444
rect -28 -2448 -27 -2444
rect 213 -2448 214 -2444
rect 216 -2448 218 -2444
rect 222 -2448 224 -2444
rect 226 -2448 227 -2444
rect 239 -2448 240 -2444
rect 242 -2448 248 -2444
rect 250 -2448 251 -2444
rect 263 -2448 264 -2444
rect 266 -2448 272 -2444
rect 274 -2448 276 -2444
rect 280 -2448 282 -2444
rect 284 -2448 290 -2444
rect 292 -2448 293 -2444
rect 305 -2448 306 -2444
rect 308 -2448 314 -2444
rect 316 -2448 318 -2444
rect 322 -2448 324 -2444
rect 326 -2448 332 -2444
rect 334 -2448 335 -2444
rect 347 -2448 348 -2444
rect 350 -2448 356 -2444
rect 358 -2448 360 -2444
rect 364 -2448 366 -2444
rect 368 -2448 374 -2444
rect 376 -2448 377 -2444
rect 389 -2448 390 -2444
rect 392 -2448 398 -2444
rect 400 -2448 401 -2444
rect 569 -2448 570 -2444
rect 572 -2448 574 -2444
rect 578 -2448 580 -2444
rect 582 -2448 583 -2444
rect 595 -2448 596 -2444
rect 598 -2448 604 -2444
rect 606 -2448 607 -2444
rect 619 -2448 620 -2444
rect 622 -2448 628 -2444
rect 630 -2448 632 -2444
rect 636 -2448 638 -2444
rect 640 -2448 646 -2444
rect 648 -2448 649 -2444
rect 661 -2448 662 -2444
rect 664 -2448 670 -2444
rect 672 -2448 674 -2444
rect 678 -2448 680 -2444
rect 682 -2448 688 -2444
rect 690 -2448 691 -2444
rect 703 -2448 704 -2444
rect 706 -2448 712 -2444
rect 714 -2448 716 -2444
rect 720 -2448 722 -2444
rect 724 -2448 730 -2444
rect 732 -2448 733 -2444
rect 745 -2448 746 -2444
rect 748 -2448 754 -2444
rect 756 -2448 757 -2444
rect 967 -2448 968 -2444
rect 970 -2448 972 -2444
rect 976 -2448 978 -2444
rect 980 -2448 981 -2444
rect 993 -2448 994 -2444
rect 996 -2448 1002 -2444
rect 1004 -2448 1005 -2444
rect 1017 -2448 1018 -2444
rect 1020 -2448 1026 -2444
rect 1028 -2448 1030 -2444
rect 1034 -2448 1036 -2444
rect 1038 -2448 1044 -2444
rect 1046 -2448 1047 -2444
rect 1059 -2448 1060 -2444
rect 1062 -2448 1068 -2444
rect 1070 -2448 1072 -2444
rect 1076 -2448 1078 -2444
rect 1080 -2448 1086 -2444
rect 1088 -2448 1089 -2444
rect 1101 -2448 1102 -2444
rect 1104 -2448 1110 -2444
rect 1112 -2448 1114 -2444
rect 1118 -2448 1120 -2444
rect 1122 -2448 1128 -2444
rect 1130 -2448 1131 -2444
rect 1143 -2448 1144 -2444
rect 1146 -2448 1152 -2444
rect 1154 -2448 1155 -2444
rect 1325 -2448 1326 -2444
rect 1328 -2448 1330 -2444
rect 1334 -2448 1336 -2444
rect 1338 -2448 1339 -2444
rect 1351 -2448 1352 -2444
rect 1354 -2448 1360 -2444
rect 1362 -2448 1363 -2444
rect 1375 -2448 1376 -2444
rect 1378 -2448 1384 -2444
rect 1386 -2448 1388 -2444
rect 1392 -2448 1394 -2444
rect 1396 -2448 1402 -2444
rect 1404 -2448 1405 -2444
rect 1417 -2448 1418 -2444
rect 1420 -2448 1426 -2444
rect 1428 -2448 1430 -2444
rect 1434 -2448 1436 -2444
rect 1438 -2448 1444 -2444
rect 1446 -2448 1447 -2444
rect 1459 -2448 1460 -2444
rect 1462 -2448 1468 -2444
rect 1470 -2448 1472 -2444
rect 1476 -2448 1478 -2444
rect 1480 -2448 1486 -2444
rect 1488 -2448 1489 -2444
rect 1501 -2448 1502 -2444
rect 1504 -2448 1510 -2444
rect 1512 -2448 1513 -2444
rect -1260 -2579 -1259 -2575
rect -1257 -2579 -1255 -2575
rect -1251 -2579 -1249 -2575
rect -1247 -2579 -1246 -2575
rect -1234 -2579 -1233 -2575
rect -1231 -2579 -1225 -2575
rect -1223 -2579 -1222 -2575
rect -1210 -2579 -1209 -2575
rect -1207 -2579 -1201 -2575
rect -1199 -2579 -1197 -2575
rect -1193 -2579 -1191 -2575
rect -1189 -2579 -1183 -2575
rect -1181 -2579 -1180 -2575
rect -1168 -2579 -1167 -2575
rect -1165 -2579 -1159 -2575
rect -1157 -2579 -1155 -2575
rect -1151 -2579 -1149 -2575
rect -1147 -2579 -1141 -2575
rect -1139 -2579 -1138 -2575
rect -1126 -2579 -1125 -2575
rect -1123 -2579 -1117 -2575
rect -1115 -2579 -1113 -2575
rect -1109 -2579 -1107 -2575
rect -1105 -2579 -1099 -2575
rect -1097 -2579 -1096 -2575
rect -1084 -2579 -1083 -2575
rect -1081 -2579 -1075 -2575
rect -1073 -2579 -1072 -2575
rect -931 -2579 -930 -2575
rect -928 -2579 -926 -2575
rect -922 -2579 -920 -2575
rect -918 -2579 -917 -2575
rect -905 -2579 -904 -2575
rect -902 -2579 -896 -2575
rect -894 -2579 -893 -2575
rect -881 -2579 -880 -2575
rect -878 -2579 -872 -2575
rect -870 -2579 -868 -2575
rect -864 -2579 -862 -2575
rect -860 -2579 -854 -2575
rect -852 -2579 -851 -2575
rect -839 -2579 -838 -2575
rect -836 -2579 -830 -2575
rect -828 -2579 -826 -2575
rect -822 -2579 -820 -2575
rect -818 -2579 -812 -2575
rect -810 -2579 -809 -2575
rect -797 -2579 -796 -2575
rect -794 -2579 -788 -2575
rect -786 -2579 -784 -2575
rect -780 -2579 -778 -2575
rect -776 -2579 -770 -2575
rect -768 -2579 -767 -2575
rect -755 -2579 -754 -2575
rect -752 -2579 -746 -2575
rect -744 -2579 -743 -2575
rect -573 -2579 -572 -2575
rect -570 -2579 -568 -2575
rect -564 -2579 -562 -2575
rect -560 -2579 -559 -2575
rect -547 -2579 -546 -2575
rect -544 -2579 -538 -2575
rect -536 -2579 -535 -2575
rect -523 -2579 -522 -2575
rect -520 -2579 -514 -2575
rect -512 -2579 -510 -2575
rect -506 -2579 -504 -2575
rect -502 -2579 -496 -2575
rect -494 -2579 -493 -2575
rect -481 -2579 -480 -2575
rect -478 -2579 -472 -2575
rect -470 -2579 -468 -2575
rect -464 -2579 -462 -2575
rect -460 -2579 -454 -2575
rect -452 -2579 -451 -2575
rect -439 -2579 -438 -2575
rect -436 -2579 -430 -2575
rect -428 -2579 -426 -2575
rect -422 -2579 -420 -2575
rect -418 -2579 -412 -2575
rect -410 -2579 -409 -2575
rect -397 -2579 -396 -2575
rect -394 -2579 -388 -2575
rect -386 -2579 -385 -2575
rect -215 -2579 -214 -2575
rect -212 -2579 -210 -2575
rect -206 -2579 -204 -2575
rect -202 -2579 -201 -2575
rect -189 -2579 -188 -2575
rect -186 -2579 -180 -2575
rect -178 -2579 -177 -2575
rect -165 -2579 -164 -2575
rect -162 -2579 -156 -2575
rect -154 -2579 -152 -2575
rect -148 -2579 -146 -2575
rect -144 -2579 -138 -2575
rect -136 -2579 -135 -2575
rect -123 -2579 -122 -2575
rect -120 -2579 -114 -2575
rect -112 -2579 -110 -2575
rect -106 -2579 -104 -2575
rect -102 -2579 -96 -2575
rect -94 -2579 -93 -2575
rect -81 -2579 -80 -2575
rect -78 -2579 -72 -2575
rect -70 -2579 -68 -2575
rect -64 -2579 -62 -2575
rect -60 -2579 -54 -2575
rect -52 -2579 -51 -2575
rect -39 -2579 -38 -2575
rect -36 -2579 -30 -2575
rect -28 -2579 -27 -2575
rect 94 -2579 95 -2563
rect 97 -2579 98 -2563
rect 213 -2579 214 -2575
rect 216 -2579 218 -2575
rect 222 -2579 224 -2575
rect 226 -2579 227 -2575
rect 239 -2579 240 -2575
rect 242 -2579 248 -2575
rect 250 -2579 251 -2575
rect 263 -2579 264 -2575
rect 266 -2579 272 -2575
rect 274 -2579 276 -2575
rect 280 -2579 282 -2575
rect 284 -2579 290 -2575
rect 292 -2579 293 -2575
rect 305 -2579 306 -2575
rect 308 -2579 314 -2575
rect 316 -2579 318 -2575
rect 322 -2579 324 -2575
rect 326 -2579 332 -2575
rect 334 -2579 335 -2575
rect 347 -2579 348 -2575
rect 350 -2579 356 -2575
rect 358 -2579 360 -2575
rect 364 -2579 366 -2575
rect 368 -2579 374 -2575
rect 376 -2579 377 -2575
rect 389 -2579 390 -2575
rect 392 -2579 398 -2575
rect 400 -2579 401 -2575
rect 569 -2579 570 -2575
rect 572 -2579 574 -2575
rect 578 -2579 580 -2575
rect 582 -2579 583 -2575
rect 595 -2579 596 -2575
rect 598 -2579 604 -2575
rect 606 -2579 607 -2575
rect 619 -2579 620 -2575
rect 622 -2579 628 -2575
rect 630 -2579 632 -2575
rect 636 -2579 638 -2575
rect 640 -2579 646 -2575
rect 648 -2579 649 -2575
rect 661 -2579 662 -2575
rect 664 -2579 670 -2575
rect 672 -2579 674 -2575
rect 678 -2579 680 -2575
rect 682 -2579 688 -2575
rect 690 -2579 691 -2575
rect 703 -2579 704 -2575
rect 706 -2579 712 -2575
rect 714 -2579 716 -2575
rect 720 -2579 722 -2575
rect 724 -2579 730 -2575
rect 732 -2579 733 -2575
rect 745 -2579 746 -2575
rect 748 -2579 754 -2575
rect 756 -2579 757 -2575
rect 967 -2579 968 -2575
rect 970 -2579 972 -2575
rect 976 -2579 978 -2575
rect 980 -2579 981 -2575
rect 993 -2579 994 -2575
rect 996 -2579 1002 -2575
rect 1004 -2579 1005 -2575
rect 1017 -2579 1018 -2575
rect 1020 -2579 1026 -2575
rect 1028 -2579 1030 -2575
rect 1034 -2579 1036 -2575
rect 1038 -2579 1044 -2575
rect 1046 -2579 1047 -2575
rect 1059 -2579 1060 -2575
rect 1062 -2579 1068 -2575
rect 1070 -2579 1072 -2575
rect 1076 -2579 1078 -2575
rect 1080 -2579 1086 -2575
rect 1088 -2579 1089 -2575
rect 1101 -2579 1102 -2575
rect 1104 -2579 1110 -2575
rect 1112 -2579 1114 -2575
rect 1118 -2579 1120 -2575
rect 1122 -2579 1128 -2575
rect 1130 -2579 1131 -2575
rect 1143 -2579 1144 -2575
rect 1146 -2579 1152 -2575
rect 1154 -2579 1155 -2575
rect 1325 -2579 1326 -2575
rect 1328 -2579 1330 -2575
rect 1334 -2579 1336 -2575
rect 1338 -2579 1339 -2575
rect 1351 -2579 1352 -2575
rect 1354 -2579 1360 -2575
rect 1362 -2579 1363 -2575
rect 1375 -2579 1376 -2575
rect 1378 -2579 1384 -2575
rect 1386 -2579 1388 -2575
rect 1392 -2579 1394 -2575
rect 1396 -2579 1402 -2575
rect 1404 -2579 1405 -2575
rect 1417 -2579 1418 -2575
rect 1420 -2579 1426 -2575
rect 1428 -2579 1430 -2575
rect 1434 -2579 1436 -2575
rect 1438 -2579 1444 -2575
rect 1446 -2579 1447 -2575
rect 1459 -2579 1460 -2575
rect 1462 -2579 1468 -2575
rect 1470 -2579 1472 -2575
rect 1476 -2579 1478 -2575
rect 1480 -2579 1486 -2575
rect 1488 -2579 1489 -2575
rect 1501 -2579 1502 -2575
rect 1504 -2579 1510 -2575
rect 1512 -2579 1513 -2575
rect -1260 -2691 -1259 -2687
rect -1257 -2691 -1255 -2687
rect -1251 -2691 -1249 -2687
rect -1247 -2691 -1246 -2687
rect -1234 -2691 -1233 -2687
rect -1231 -2691 -1225 -2687
rect -1223 -2691 -1222 -2687
rect -1210 -2691 -1209 -2687
rect -1207 -2691 -1201 -2687
rect -1199 -2691 -1197 -2687
rect -1193 -2691 -1191 -2687
rect -1189 -2691 -1183 -2687
rect -1181 -2691 -1180 -2687
rect -1168 -2691 -1167 -2687
rect -1165 -2691 -1159 -2687
rect -1157 -2691 -1155 -2687
rect -1151 -2691 -1149 -2687
rect -1147 -2691 -1141 -2687
rect -1139 -2691 -1138 -2687
rect -1126 -2691 -1125 -2687
rect -1123 -2691 -1117 -2687
rect -1115 -2691 -1113 -2687
rect -1109 -2691 -1107 -2687
rect -1105 -2691 -1099 -2687
rect -1097 -2691 -1096 -2687
rect -1084 -2691 -1083 -2687
rect -1081 -2691 -1075 -2687
rect -1073 -2691 -1072 -2687
rect -931 -2691 -930 -2687
rect -928 -2691 -926 -2687
rect -922 -2691 -920 -2687
rect -918 -2691 -917 -2687
rect -905 -2691 -904 -2687
rect -902 -2691 -896 -2687
rect -894 -2691 -893 -2687
rect -881 -2691 -880 -2687
rect -878 -2691 -872 -2687
rect -870 -2691 -868 -2687
rect -864 -2691 -862 -2687
rect -860 -2691 -854 -2687
rect -852 -2691 -851 -2687
rect -839 -2691 -838 -2687
rect -836 -2691 -830 -2687
rect -828 -2691 -826 -2687
rect -822 -2691 -820 -2687
rect -818 -2691 -812 -2687
rect -810 -2691 -809 -2687
rect -797 -2691 -796 -2687
rect -794 -2691 -788 -2687
rect -786 -2691 -784 -2687
rect -780 -2691 -778 -2687
rect -776 -2691 -770 -2687
rect -768 -2691 -767 -2687
rect -755 -2691 -754 -2687
rect -752 -2691 -746 -2687
rect -744 -2691 -743 -2687
rect -1335 -2804 -1334 -2800
rect -1332 -2804 -1326 -2800
rect -1324 -2804 -1322 -2800
rect -1318 -2804 -1316 -2800
rect -1314 -2804 -1313 -2800
rect -931 -2804 -930 -2800
rect -928 -2804 -922 -2800
rect -920 -2804 -918 -2800
rect -914 -2804 -912 -2800
rect -910 -2804 -909 -2800
rect -573 -2804 -572 -2800
rect -570 -2804 -564 -2800
rect -562 -2804 -560 -2800
rect -556 -2804 -554 -2800
rect -552 -2804 -551 -2800
rect -215 -2804 -214 -2800
rect -212 -2804 -206 -2800
rect -204 -2804 -202 -2800
rect -198 -2804 -196 -2800
rect -194 -2804 -193 -2800
rect 213 -2804 214 -2800
rect 216 -2804 222 -2800
rect 224 -2804 226 -2800
rect 230 -2804 232 -2800
rect 234 -2804 235 -2800
rect 569 -2804 570 -2800
rect 572 -2804 578 -2800
rect 580 -2804 582 -2800
rect 586 -2804 588 -2800
rect 590 -2804 591 -2800
rect 967 -2804 968 -2800
rect 970 -2804 976 -2800
rect 978 -2804 980 -2800
rect 984 -2804 986 -2800
rect 988 -2804 989 -2800
rect 1325 -2804 1326 -2800
rect 1328 -2804 1334 -2800
rect 1336 -2804 1338 -2800
rect 1342 -2804 1344 -2800
rect 1346 -2804 1347 -2800
rect -1260 -2923 -1259 -2919
rect -1257 -2923 -1255 -2919
rect -1251 -2923 -1249 -2919
rect -1247 -2923 -1246 -2919
rect -1234 -2923 -1233 -2919
rect -1231 -2923 -1229 -2919
rect -1225 -2923 -1223 -2919
rect -1221 -2923 -1215 -2919
rect -1213 -2923 -1211 -2919
rect -1207 -2923 -1205 -2919
rect -1203 -2923 -1202 -2919
rect -1190 -2923 -1189 -2919
rect -1187 -2923 -1181 -2919
rect -1179 -2923 -1177 -2919
rect -1173 -2923 -1171 -2919
rect -1169 -2923 -1168 -2919
rect -931 -2923 -930 -2919
rect -928 -2923 -926 -2919
rect -922 -2923 -920 -2919
rect -918 -2923 -917 -2919
rect -905 -2923 -904 -2919
rect -902 -2923 -900 -2919
rect -896 -2923 -894 -2919
rect -892 -2923 -891 -2919
rect -879 -2923 -878 -2919
rect -876 -2923 -875 -2919
rect -871 -2923 -868 -2919
rect -866 -2923 -860 -2919
rect -858 -2923 -857 -2919
rect -853 -2923 -850 -2919
rect -848 -2923 -847 -2919
rect -835 -2923 -834 -2919
rect -832 -2923 -826 -2919
rect -824 -2923 -822 -2919
rect -818 -2923 -816 -2919
rect -814 -2923 -813 -2919
rect -801 -2923 -800 -2919
rect -798 -2923 -796 -2919
rect -792 -2923 -790 -2919
rect -788 -2923 -782 -2919
rect -780 -2923 -778 -2919
rect -774 -2923 -772 -2919
rect -770 -2923 -769 -2919
rect -757 -2923 -756 -2919
rect -754 -2923 -748 -2919
rect -746 -2923 -745 -2919
rect -733 -2923 -732 -2919
rect -730 -2923 -725 -2919
rect -721 -2923 -716 -2919
rect -714 -2923 -713 -2919
rect -709 -2923 -708 -2919
rect -706 -2923 -704 -2919
rect -700 -2923 -698 -2919
rect -696 -2923 -695 -2919
rect -573 -2923 -572 -2919
rect -570 -2923 -568 -2919
rect -564 -2923 -562 -2919
rect -560 -2923 -559 -2919
rect -547 -2923 -546 -2919
rect -544 -2923 -542 -2919
rect -538 -2923 -536 -2919
rect -534 -2923 -533 -2919
rect -521 -2923 -520 -2919
rect -518 -2923 -517 -2919
rect -513 -2923 -510 -2919
rect -508 -2923 -502 -2919
rect -500 -2923 -499 -2919
rect -495 -2923 -492 -2919
rect -490 -2923 -489 -2919
rect -477 -2923 -476 -2919
rect -474 -2923 -468 -2919
rect -466 -2923 -464 -2919
rect -460 -2923 -458 -2919
rect -456 -2923 -455 -2919
rect -443 -2923 -442 -2919
rect -440 -2923 -438 -2919
rect -434 -2923 -432 -2919
rect -430 -2923 -424 -2919
rect -422 -2923 -420 -2919
rect -416 -2923 -414 -2919
rect -412 -2923 -411 -2919
rect -399 -2923 -398 -2919
rect -396 -2923 -390 -2919
rect -388 -2923 -387 -2919
rect -375 -2923 -374 -2919
rect -372 -2923 -367 -2919
rect -363 -2923 -358 -2919
rect -356 -2923 -355 -2919
rect -351 -2923 -350 -2919
rect -348 -2923 -346 -2919
rect -342 -2923 -340 -2919
rect -338 -2923 -337 -2919
rect -215 -2923 -214 -2919
rect -212 -2923 -210 -2919
rect -206 -2923 -204 -2919
rect -202 -2923 -201 -2919
rect -189 -2923 -188 -2919
rect -186 -2923 -184 -2919
rect -180 -2923 -178 -2919
rect -176 -2923 -175 -2919
rect -163 -2923 -162 -2919
rect -160 -2923 -159 -2919
rect -155 -2923 -152 -2919
rect -150 -2923 -144 -2919
rect -142 -2923 -141 -2919
rect -137 -2923 -134 -2919
rect -132 -2923 -131 -2919
rect -119 -2923 -118 -2919
rect -116 -2923 -110 -2919
rect -108 -2923 -106 -2919
rect -102 -2923 -100 -2919
rect -98 -2923 -97 -2919
rect -85 -2923 -84 -2919
rect -82 -2923 -80 -2919
rect -76 -2923 -74 -2919
rect -72 -2923 -66 -2919
rect -64 -2923 -62 -2919
rect -58 -2923 -56 -2919
rect -54 -2923 -53 -2919
rect -41 -2923 -40 -2919
rect -38 -2923 -32 -2919
rect -30 -2923 -29 -2919
rect -17 -2923 -16 -2919
rect -14 -2923 -9 -2919
rect -5 -2923 0 -2919
rect 2 -2923 3 -2919
rect 7 -2923 8 -2919
rect 10 -2923 12 -2919
rect 16 -2923 18 -2919
rect 20 -2923 21 -2919
rect 213 -2923 214 -2919
rect 216 -2923 218 -2919
rect 222 -2923 224 -2919
rect 226 -2923 227 -2919
rect 239 -2923 240 -2919
rect 242 -2923 244 -2919
rect 248 -2923 250 -2919
rect 252 -2923 253 -2919
rect 265 -2923 266 -2919
rect 268 -2923 269 -2919
rect 273 -2923 276 -2919
rect 278 -2923 284 -2919
rect 286 -2923 287 -2919
rect 291 -2923 294 -2919
rect 296 -2923 297 -2919
rect 309 -2923 310 -2919
rect 312 -2923 318 -2919
rect 320 -2923 322 -2919
rect 326 -2923 328 -2919
rect 330 -2923 331 -2919
rect 343 -2923 344 -2919
rect 346 -2923 348 -2919
rect 352 -2923 354 -2919
rect 356 -2923 362 -2919
rect 364 -2923 366 -2919
rect 370 -2923 372 -2919
rect 374 -2923 375 -2919
rect 387 -2923 388 -2919
rect 390 -2923 396 -2919
rect 398 -2923 399 -2919
rect 411 -2923 412 -2919
rect 414 -2923 419 -2919
rect 423 -2923 428 -2919
rect 430 -2923 431 -2919
rect 435 -2923 436 -2919
rect 438 -2923 440 -2919
rect 444 -2923 446 -2919
rect 448 -2923 449 -2919
rect 569 -2923 570 -2919
rect 572 -2923 574 -2919
rect 578 -2923 580 -2919
rect 582 -2923 583 -2919
rect 595 -2923 596 -2919
rect 598 -2923 600 -2919
rect 604 -2923 606 -2919
rect 608 -2923 609 -2919
rect 621 -2923 622 -2919
rect 624 -2923 625 -2919
rect 629 -2923 632 -2919
rect 634 -2923 640 -2919
rect 642 -2923 643 -2919
rect 647 -2923 650 -2919
rect 652 -2923 653 -2919
rect 665 -2923 666 -2919
rect 668 -2923 674 -2919
rect 676 -2923 678 -2919
rect 682 -2923 684 -2919
rect 686 -2923 687 -2919
rect 699 -2923 700 -2919
rect 702 -2923 704 -2919
rect 708 -2923 710 -2919
rect 712 -2923 718 -2919
rect 720 -2923 722 -2919
rect 726 -2923 728 -2919
rect 730 -2923 731 -2919
rect 743 -2923 744 -2919
rect 746 -2923 752 -2919
rect 754 -2923 755 -2919
rect 767 -2923 768 -2919
rect 770 -2923 775 -2919
rect 779 -2923 784 -2919
rect 786 -2923 787 -2919
rect 791 -2923 792 -2919
rect 794 -2923 796 -2919
rect 800 -2923 802 -2919
rect 804 -2923 805 -2919
rect 967 -2923 968 -2919
rect 970 -2923 972 -2919
rect 976 -2923 978 -2919
rect 980 -2923 981 -2919
rect 993 -2923 994 -2919
rect 996 -2923 998 -2919
rect 1002 -2923 1004 -2919
rect 1006 -2923 1007 -2919
rect 1019 -2923 1020 -2919
rect 1022 -2923 1023 -2919
rect 1027 -2923 1030 -2919
rect 1032 -2923 1038 -2919
rect 1040 -2923 1041 -2919
rect 1045 -2923 1048 -2919
rect 1050 -2923 1051 -2919
rect 1063 -2923 1064 -2919
rect 1066 -2923 1072 -2919
rect 1074 -2923 1076 -2919
rect 1080 -2923 1082 -2919
rect 1084 -2923 1085 -2919
rect 1097 -2923 1098 -2919
rect 1100 -2923 1102 -2919
rect 1106 -2923 1108 -2919
rect 1110 -2923 1116 -2919
rect 1118 -2923 1120 -2919
rect 1124 -2923 1126 -2919
rect 1128 -2923 1129 -2919
rect 1141 -2923 1142 -2919
rect 1144 -2923 1150 -2919
rect 1152 -2923 1153 -2919
rect 1165 -2923 1166 -2919
rect 1168 -2923 1173 -2919
rect 1177 -2923 1182 -2919
rect 1184 -2923 1185 -2919
rect 1189 -2923 1190 -2919
rect 1192 -2923 1194 -2919
rect 1198 -2923 1200 -2919
rect 1202 -2923 1203 -2919
rect 1325 -2923 1326 -2919
rect 1328 -2923 1330 -2919
rect 1334 -2923 1336 -2919
rect 1338 -2923 1339 -2919
rect 1351 -2923 1352 -2919
rect 1354 -2923 1356 -2919
rect 1360 -2923 1362 -2919
rect 1364 -2923 1365 -2919
rect 1377 -2923 1378 -2919
rect 1380 -2923 1381 -2919
rect 1385 -2923 1388 -2919
rect 1390 -2923 1396 -2919
rect 1398 -2923 1399 -2919
rect 1403 -2923 1406 -2919
rect 1408 -2923 1409 -2919
rect 1421 -2923 1422 -2919
rect 1424 -2923 1430 -2919
rect 1432 -2923 1434 -2919
rect 1438 -2923 1440 -2919
rect 1442 -2923 1443 -2919
rect 1455 -2923 1456 -2919
rect 1458 -2923 1460 -2919
rect 1464 -2923 1466 -2919
rect 1468 -2923 1474 -2919
rect 1476 -2923 1478 -2919
rect 1482 -2923 1484 -2919
rect 1486 -2923 1487 -2919
rect 1499 -2923 1500 -2919
rect 1502 -2923 1508 -2919
rect 1510 -2923 1511 -2919
rect 1523 -2923 1524 -2919
rect 1526 -2923 1531 -2919
rect 1535 -2923 1540 -2919
rect 1542 -2923 1543 -2919
rect 1547 -2923 1548 -2919
rect 1550 -2923 1552 -2919
rect 1556 -2923 1558 -2919
rect 1560 -2923 1561 -2919
rect -1260 -3042 -1259 -3038
rect -1257 -3042 -1255 -3038
rect -1251 -3042 -1249 -3038
rect -1247 -3042 -1246 -3038
rect -1234 -3042 -1233 -3038
rect -1231 -3042 -1225 -3038
rect -1223 -3042 -1222 -3038
rect -1210 -3042 -1209 -3038
rect -1207 -3042 -1201 -3038
rect -1199 -3042 -1197 -3038
rect -1193 -3042 -1191 -3038
rect -1189 -3042 -1183 -3038
rect -1181 -3042 -1180 -3038
rect -1168 -3042 -1167 -3038
rect -1165 -3042 -1159 -3038
rect -1157 -3042 -1155 -3038
rect -1151 -3042 -1149 -3038
rect -1147 -3042 -1141 -3038
rect -1139 -3042 -1138 -3038
rect -1126 -3042 -1125 -3038
rect -1123 -3042 -1117 -3038
rect -1115 -3042 -1113 -3038
rect -1109 -3042 -1107 -3038
rect -1105 -3042 -1099 -3038
rect -1097 -3042 -1096 -3038
rect -1084 -3042 -1083 -3038
rect -1081 -3042 -1075 -3038
rect -1073 -3042 -1072 -3038
rect -1022 -3042 -1021 -3038
rect -1019 -3042 -1018 -3038
rect -931 -3042 -930 -3038
rect -928 -3042 -926 -3038
rect -922 -3042 -920 -3038
rect -918 -3042 -917 -3038
rect -905 -3042 -904 -3038
rect -902 -3042 -896 -3038
rect -894 -3042 -893 -3038
rect -881 -3042 -880 -3038
rect -878 -3042 -872 -3038
rect -870 -3042 -868 -3038
rect -864 -3042 -862 -3038
rect -860 -3042 -854 -3038
rect -852 -3042 -851 -3038
rect -839 -3042 -838 -3038
rect -836 -3042 -830 -3038
rect -828 -3042 -826 -3038
rect -822 -3042 -820 -3038
rect -818 -3042 -812 -3038
rect -810 -3042 -809 -3038
rect -797 -3042 -796 -3038
rect -794 -3042 -788 -3038
rect -786 -3042 -784 -3038
rect -780 -3042 -778 -3038
rect -776 -3042 -770 -3038
rect -768 -3042 -767 -3038
rect -755 -3042 -754 -3038
rect -752 -3042 -746 -3038
rect -744 -3042 -743 -3038
rect -668 -3042 -667 -3034
rect -665 -3042 -664 -3034
rect -573 -3042 -572 -3038
rect -570 -3042 -568 -3038
rect -564 -3042 -562 -3038
rect -560 -3042 -559 -3038
rect -547 -3042 -546 -3038
rect -544 -3042 -538 -3038
rect -536 -3042 -535 -3038
rect -523 -3042 -522 -3038
rect -520 -3042 -514 -3038
rect -512 -3042 -510 -3038
rect -506 -3042 -504 -3038
rect -502 -3042 -496 -3038
rect -494 -3042 -493 -3038
rect -481 -3042 -480 -3038
rect -478 -3042 -472 -3038
rect -470 -3042 -468 -3038
rect -464 -3042 -462 -3038
rect -460 -3042 -454 -3038
rect -452 -3042 -451 -3038
rect -439 -3042 -438 -3038
rect -436 -3042 -430 -3038
rect -428 -3042 -426 -3038
rect -422 -3042 -420 -3038
rect -418 -3042 -412 -3038
rect -410 -3042 -409 -3038
rect -397 -3042 -396 -3038
rect -394 -3042 -388 -3038
rect -386 -3042 -385 -3038
rect -325 -3042 -324 -3038
rect -322 -3042 -321 -3038
rect -215 -3042 -214 -3038
rect -212 -3042 -210 -3038
rect -206 -3042 -204 -3038
rect -202 -3042 -201 -3038
rect -189 -3042 -188 -3038
rect -186 -3042 -180 -3038
rect -178 -3042 -177 -3038
rect -165 -3042 -164 -3038
rect -162 -3042 -156 -3038
rect -154 -3042 -152 -3038
rect -148 -3042 -146 -3038
rect -144 -3042 -138 -3038
rect -136 -3042 -135 -3038
rect -123 -3042 -122 -3038
rect -120 -3042 -114 -3038
rect -112 -3042 -110 -3038
rect -106 -3042 -104 -3038
rect -102 -3042 -96 -3038
rect -94 -3042 -93 -3038
rect -81 -3042 -80 -3038
rect -78 -3042 -72 -3038
rect -70 -3042 -68 -3038
rect -64 -3042 -62 -3038
rect -60 -3042 -54 -3038
rect -52 -3042 -51 -3038
rect -39 -3042 -38 -3038
rect -36 -3042 -30 -3038
rect -28 -3042 -27 -3038
rect 213 -3042 214 -3038
rect 216 -3042 218 -3038
rect 222 -3042 224 -3038
rect 226 -3042 227 -3038
rect 239 -3042 240 -3038
rect 242 -3042 248 -3038
rect 250 -3042 251 -3038
rect 263 -3042 264 -3038
rect 266 -3042 272 -3038
rect 274 -3042 276 -3038
rect 280 -3042 282 -3038
rect 284 -3042 290 -3038
rect 292 -3042 293 -3038
rect 305 -3042 306 -3038
rect 308 -3042 314 -3038
rect 316 -3042 318 -3038
rect 322 -3042 324 -3038
rect 326 -3042 332 -3038
rect 334 -3042 335 -3038
rect 347 -3042 348 -3038
rect 350 -3042 356 -3038
rect 358 -3042 360 -3038
rect 364 -3042 366 -3038
rect 368 -3042 374 -3038
rect 376 -3042 377 -3038
rect 389 -3042 390 -3038
rect 392 -3042 398 -3038
rect 400 -3042 401 -3038
rect 476 -3042 477 -3038
rect 479 -3042 480 -3038
rect 845 -3042 846 -3034
rect 848 -3042 849 -3034
rect 1203 -3042 1204 -3038
rect 1206 -3042 1207 -3038
rect -1260 -3158 -1259 -3154
rect -1257 -3158 -1255 -3154
rect -1251 -3158 -1249 -3154
rect -1247 -3158 -1246 -3154
rect -1234 -3158 -1233 -3154
rect -1231 -3158 -1225 -3154
rect -1223 -3158 -1222 -3154
rect -1210 -3158 -1209 -3154
rect -1207 -3158 -1201 -3154
rect -1199 -3158 -1197 -3154
rect -1193 -3158 -1191 -3154
rect -1189 -3158 -1183 -3154
rect -1181 -3158 -1180 -3154
rect -1168 -3158 -1167 -3154
rect -1165 -3158 -1159 -3154
rect -1157 -3158 -1155 -3154
rect -1151 -3158 -1149 -3154
rect -1147 -3158 -1141 -3154
rect -1139 -3158 -1138 -3154
rect -1126 -3158 -1125 -3154
rect -1123 -3158 -1117 -3154
rect -1115 -3158 -1113 -3154
rect -1109 -3158 -1107 -3154
rect -1105 -3158 -1099 -3154
rect -1097 -3158 -1096 -3154
rect -1084 -3158 -1083 -3154
rect -1081 -3158 -1075 -3154
rect -1073 -3158 -1072 -3154
rect -1022 -3158 -1021 -3154
rect -1019 -3158 -1018 -3154
rect -931 -3158 -930 -3154
rect -928 -3158 -926 -3154
rect -922 -3158 -920 -3154
rect -918 -3158 -917 -3154
rect -905 -3158 -904 -3154
rect -902 -3158 -896 -3154
rect -894 -3158 -893 -3154
rect -881 -3158 -880 -3154
rect -878 -3158 -872 -3154
rect -870 -3158 -868 -3154
rect -864 -3158 -862 -3154
rect -860 -3158 -854 -3154
rect -852 -3158 -851 -3154
rect -839 -3158 -838 -3154
rect -836 -3158 -830 -3154
rect -828 -3158 -826 -3154
rect -822 -3158 -820 -3154
rect -818 -3158 -812 -3154
rect -810 -3158 -809 -3154
rect -797 -3158 -796 -3154
rect -794 -3158 -788 -3154
rect -786 -3158 -784 -3154
rect -780 -3158 -778 -3154
rect -776 -3158 -770 -3154
rect -768 -3158 -767 -3154
rect -755 -3158 -754 -3154
rect -752 -3158 -746 -3154
rect -744 -3158 -743 -3154
rect -573 -3158 -572 -3154
rect -570 -3158 -568 -3154
rect -564 -3158 -562 -3154
rect -560 -3158 -559 -3154
rect -547 -3158 -546 -3154
rect -544 -3158 -538 -3154
rect -536 -3158 -535 -3154
rect -523 -3158 -522 -3154
rect -520 -3158 -514 -3154
rect -512 -3158 -510 -3154
rect -506 -3158 -504 -3154
rect -502 -3158 -496 -3154
rect -494 -3158 -493 -3154
rect -481 -3158 -480 -3154
rect -478 -3158 -472 -3154
rect -470 -3158 -468 -3154
rect -464 -3158 -462 -3154
rect -460 -3158 -454 -3154
rect -452 -3158 -451 -3154
rect -439 -3158 -438 -3154
rect -436 -3158 -430 -3154
rect -428 -3158 -426 -3154
rect -422 -3158 -420 -3154
rect -418 -3158 -412 -3154
rect -410 -3158 -409 -3154
rect -397 -3158 -396 -3154
rect -394 -3158 -388 -3154
rect -386 -3158 -385 -3154
rect -325 -3158 -324 -3154
rect -322 -3158 -321 -3154
rect -215 -3158 -214 -3154
rect -212 -3158 -210 -3154
rect -206 -3158 -204 -3154
rect -202 -3158 -201 -3154
rect -189 -3158 -188 -3154
rect -186 -3158 -180 -3154
rect -178 -3158 -177 -3154
rect -165 -3158 -164 -3154
rect -162 -3158 -156 -3154
rect -154 -3158 -152 -3154
rect -148 -3158 -146 -3154
rect -144 -3158 -138 -3154
rect -136 -3158 -135 -3154
rect -123 -3158 -122 -3154
rect -120 -3158 -114 -3154
rect -112 -3158 -110 -3154
rect -106 -3158 -104 -3154
rect -102 -3158 -96 -3154
rect -94 -3158 -93 -3154
rect -81 -3158 -80 -3154
rect -78 -3158 -72 -3154
rect -70 -3158 -68 -3154
rect -64 -3158 -62 -3154
rect -60 -3158 -54 -3154
rect -52 -3158 -51 -3154
rect -39 -3158 -38 -3154
rect -36 -3158 -30 -3154
rect -28 -3158 -27 -3154
rect 213 -3158 214 -3154
rect 216 -3158 218 -3154
rect 222 -3158 224 -3154
rect 226 -3158 227 -3154
rect 239 -3158 240 -3154
rect 242 -3158 248 -3154
rect 250 -3158 251 -3154
rect 263 -3158 264 -3154
rect 266 -3158 272 -3154
rect 274 -3158 276 -3154
rect 280 -3158 282 -3154
rect 284 -3158 290 -3154
rect 292 -3158 293 -3154
rect 305 -3158 306 -3154
rect 308 -3158 314 -3154
rect 316 -3158 318 -3154
rect 322 -3158 324 -3154
rect 326 -3158 332 -3154
rect 334 -3158 335 -3154
rect 347 -3158 348 -3154
rect 350 -3158 356 -3154
rect 358 -3158 360 -3154
rect 364 -3158 366 -3154
rect 368 -3158 374 -3154
rect 376 -3158 377 -3154
rect 389 -3158 390 -3154
rect 392 -3158 398 -3154
rect 400 -3158 401 -3154
rect 476 -3158 477 -3154
rect 479 -3158 480 -3154
rect 569 -3158 570 -3154
rect 572 -3158 574 -3154
rect 578 -3158 580 -3154
rect 582 -3158 583 -3154
rect 595 -3158 596 -3154
rect 598 -3158 604 -3154
rect 606 -3158 607 -3154
rect 619 -3158 620 -3154
rect 622 -3158 628 -3154
rect 630 -3158 632 -3154
rect 636 -3158 638 -3154
rect 640 -3158 646 -3154
rect 648 -3158 649 -3154
rect 661 -3158 662 -3154
rect 664 -3158 670 -3154
rect 672 -3158 674 -3154
rect 678 -3158 680 -3154
rect 682 -3158 688 -3154
rect 690 -3158 691 -3154
rect 703 -3158 704 -3154
rect 706 -3158 712 -3154
rect 714 -3158 716 -3154
rect 720 -3158 722 -3154
rect 724 -3158 730 -3154
rect 732 -3158 733 -3154
rect 745 -3158 746 -3154
rect 748 -3158 754 -3154
rect 756 -3158 757 -3154
rect 967 -3158 968 -3154
rect 970 -3158 972 -3154
rect 976 -3158 978 -3154
rect 980 -3158 981 -3154
rect 993 -3158 994 -3154
rect 996 -3158 1002 -3154
rect 1004 -3158 1005 -3154
rect 1017 -3158 1018 -3154
rect 1020 -3158 1026 -3154
rect 1028 -3158 1030 -3154
rect 1034 -3158 1036 -3154
rect 1038 -3158 1044 -3154
rect 1046 -3158 1047 -3154
rect 1059 -3158 1060 -3154
rect 1062 -3158 1068 -3154
rect 1070 -3158 1072 -3154
rect 1076 -3158 1078 -3154
rect 1080 -3158 1086 -3154
rect 1088 -3158 1089 -3154
rect 1101 -3158 1102 -3154
rect 1104 -3158 1110 -3154
rect 1112 -3158 1114 -3154
rect 1118 -3158 1120 -3154
rect 1122 -3158 1128 -3154
rect 1130 -3158 1131 -3154
rect 1143 -3158 1144 -3154
rect 1146 -3158 1152 -3154
rect 1154 -3158 1155 -3154
rect 1203 -3158 1204 -3154
rect 1206 -3158 1207 -3154
rect 1325 -3158 1326 -3154
rect 1328 -3158 1330 -3154
rect 1334 -3158 1336 -3154
rect 1338 -3158 1339 -3154
rect 1351 -3158 1352 -3154
rect 1354 -3158 1360 -3154
rect 1362 -3158 1363 -3154
rect 1375 -3158 1376 -3154
rect 1378 -3158 1384 -3154
rect 1386 -3158 1388 -3154
rect 1392 -3158 1394 -3154
rect 1396 -3158 1402 -3154
rect 1404 -3158 1405 -3154
rect 1417 -3158 1418 -3154
rect 1420 -3158 1426 -3154
rect 1428 -3158 1430 -3154
rect 1434 -3158 1436 -3154
rect 1438 -3158 1444 -3154
rect 1446 -3158 1447 -3154
rect 1459 -3158 1460 -3154
rect 1462 -3158 1468 -3154
rect 1470 -3158 1472 -3154
rect 1476 -3158 1478 -3154
rect 1480 -3158 1486 -3154
rect 1488 -3158 1489 -3154
rect 1501 -3158 1502 -3154
rect 1504 -3158 1510 -3154
rect 1512 -3158 1513 -3154
rect -1260 -3279 -1259 -3275
rect -1257 -3279 -1255 -3275
rect -1251 -3279 -1249 -3275
rect -1247 -3279 -1246 -3275
rect -1234 -3279 -1233 -3275
rect -1231 -3279 -1225 -3275
rect -1223 -3279 -1222 -3275
rect -1210 -3279 -1209 -3275
rect -1207 -3279 -1201 -3275
rect -1199 -3279 -1197 -3275
rect -1193 -3279 -1191 -3275
rect -1189 -3279 -1183 -3275
rect -1181 -3279 -1180 -3275
rect -1168 -3279 -1167 -3275
rect -1165 -3279 -1159 -3275
rect -1157 -3279 -1155 -3275
rect -1151 -3279 -1149 -3275
rect -1147 -3279 -1141 -3275
rect -1139 -3279 -1138 -3275
rect -1126 -3279 -1125 -3275
rect -1123 -3279 -1117 -3275
rect -1115 -3279 -1113 -3275
rect -1109 -3279 -1107 -3275
rect -1105 -3279 -1099 -3275
rect -1097 -3279 -1096 -3275
rect -1084 -3279 -1083 -3275
rect -1081 -3279 -1075 -3275
rect -1073 -3279 -1072 -3275
rect -931 -3279 -930 -3275
rect -928 -3279 -926 -3275
rect -922 -3279 -920 -3275
rect -918 -3279 -917 -3275
rect -905 -3279 -904 -3275
rect -902 -3279 -896 -3275
rect -894 -3279 -893 -3275
rect -881 -3279 -880 -3275
rect -878 -3279 -872 -3275
rect -870 -3279 -868 -3275
rect -864 -3279 -862 -3275
rect -860 -3279 -854 -3275
rect -852 -3279 -851 -3275
rect -839 -3279 -838 -3275
rect -836 -3279 -830 -3275
rect -828 -3279 -826 -3275
rect -822 -3279 -820 -3275
rect -818 -3279 -812 -3275
rect -810 -3279 -809 -3275
rect -797 -3279 -796 -3275
rect -794 -3279 -788 -3275
rect -786 -3279 -784 -3275
rect -780 -3279 -778 -3275
rect -776 -3279 -770 -3275
rect -768 -3279 -767 -3275
rect -755 -3279 -754 -3275
rect -752 -3279 -746 -3275
rect -744 -3279 -743 -3275
rect -573 -3279 -572 -3275
rect -570 -3279 -568 -3275
rect -564 -3279 -562 -3275
rect -560 -3279 -559 -3275
rect -547 -3279 -546 -3275
rect -544 -3279 -538 -3275
rect -536 -3279 -535 -3275
rect -523 -3279 -522 -3275
rect -520 -3279 -514 -3275
rect -512 -3279 -510 -3275
rect -506 -3279 -504 -3275
rect -502 -3279 -496 -3275
rect -494 -3279 -493 -3275
rect -481 -3279 -480 -3275
rect -478 -3279 -472 -3275
rect -470 -3279 -468 -3275
rect -464 -3279 -462 -3275
rect -460 -3279 -454 -3275
rect -452 -3279 -451 -3275
rect -439 -3279 -438 -3275
rect -436 -3279 -430 -3275
rect -428 -3279 -426 -3275
rect -422 -3279 -420 -3275
rect -418 -3279 -412 -3275
rect -410 -3279 -409 -3275
rect -397 -3279 -396 -3275
rect -394 -3279 -388 -3275
rect -386 -3279 -385 -3275
rect -215 -3279 -214 -3275
rect -212 -3279 -210 -3275
rect -206 -3279 -204 -3275
rect -202 -3279 -201 -3275
rect -189 -3279 -188 -3275
rect -186 -3279 -180 -3275
rect -178 -3279 -177 -3275
rect -165 -3279 -164 -3275
rect -162 -3279 -156 -3275
rect -154 -3279 -152 -3275
rect -148 -3279 -146 -3275
rect -144 -3279 -138 -3275
rect -136 -3279 -135 -3275
rect -123 -3279 -122 -3275
rect -120 -3279 -114 -3275
rect -112 -3279 -110 -3275
rect -106 -3279 -104 -3275
rect -102 -3279 -96 -3275
rect -94 -3279 -93 -3275
rect -81 -3279 -80 -3275
rect -78 -3279 -72 -3275
rect -70 -3279 -68 -3275
rect -64 -3279 -62 -3275
rect -60 -3279 -54 -3275
rect -52 -3279 -51 -3275
rect -39 -3279 -38 -3275
rect -36 -3279 -30 -3275
rect -28 -3279 -27 -3275
rect 213 -3279 214 -3275
rect 216 -3279 218 -3275
rect 222 -3279 224 -3275
rect 226 -3279 227 -3275
rect 239 -3279 240 -3275
rect 242 -3279 248 -3275
rect 250 -3279 251 -3275
rect 263 -3279 264 -3275
rect 266 -3279 272 -3275
rect 274 -3279 276 -3275
rect 280 -3279 282 -3275
rect 284 -3279 290 -3275
rect 292 -3279 293 -3275
rect 305 -3279 306 -3275
rect 308 -3279 314 -3275
rect 316 -3279 318 -3275
rect 322 -3279 324 -3275
rect 326 -3279 332 -3275
rect 334 -3279 335 -3275
rect 347 -3279 348 -3275
rect 350 -3279 356 -3275
rect 358 -3279 360 -3275
rect 364 -3279 366 -3275
rect 368 -3279 374 -3275
rect 376 -3279 377 -3275
rect 389 -3279 390 -3275
rect 392 -3279 398 -3275
rect 400 -3279 401 -3275
rect 569 -3279 570 -3275
rect 572 -3279 574 -3275
rect 578 -3279 580 -3275
rect 582 -3279 583 -3275
rect 595 -3279 596 -3275
rect 598 -3279 604 -3275
rect 606 -3279 607 -3275
rect 619 -3279 620 -3275
rect 622 -3279 628 -3275
rect 630 -3279 632 -3275
rect 636 -3279 638 -3275
rect 640 -3279 646 -3275
rect 648 -3279 649 -3275
rect 661 -3279 662 -3275
rect 664 -3279 670 -3275
rect 672 -3279 674 -3275
rect 678 -3279 680 -3275
rect 682 -3279 688 -3275
rect 690 -3279 691 -3275
rect 703 -3279 704 -3275
rect 706 -3279 712 -3275
rect 714 -3279 716 -3275
rect 720 -3279 722 -3275
rect 724 -3279 730 -3275
rect 732 -3279 733 -3275
rect 745 -3279 746 -3275
rect 748 -3279 754 -3275
rect 756 -3279 757 -3275
rect 967 -3279 968 -3275
rect 970 -3279 972 -3275
rect 976 -3279 978 -3275
rect 980 -3279 981 -3275
rect 993 -3279 994 -3275
rect 996 -3279 1002 -3275
rect 1004 -3279 1005 -3275
rect 1017 -3279 1018 -3275
rect 1020 -3279 1026 -3275
rect 1028 -3279 1030 -3275
rect 1034 -3279 1036 -3275
rect 1038 -3279 1044 -3275
rect 1046 -3279 1047 -3275
rect 1059 -3279 1060 -3275
rect 1062 -3279 1068 -3275
rect 1070 -3279 1072 -3275
rect 1076 -3279 1078 -3275
rect 1080 -3279 1086 -3275
rect 1088 -3279 1089 -3275
rect 1101 -3279 1102 -3275
rect 1104 -3279 1110 -3275
rect 1112 -3279 1114 -3275
rect 1118 -3279 1120 -3275
rect 1122 -3279 1128 -3275
rect 1130 -3279 1131 -3275
rect 1143 -3279 1144 -3275
rect 1146 -3279 1152 -3275
rect 1154 -3279 1155 -3275
rect 1325 -3279 1326 -3275
rect 1328 -3279 1330 -3275
rect 1334 -3279 1336 -3275
rect 1338 -3279 1339 -3275
rect 1351 -3279 1352 -3275
rect 1354 -3279 1360 -3275
rect 1362 -3279 1363 -3275
rect 1375 -3279 1376 -3275
rect 1378 -3279 1384 -3275
rect 1386 -3279 1388 -3275
rect 1392 -3279 1394 -3275
rect 1396 -3279 1402 -3275
rect 1404 -3279 1405 -3275
rect 1417 -3279 1418 -3275
rect 1420 -3279 1426 -3275
rect 1428 -3279 1430 -3275
rect 1434 -3279 1436 -3275
rect 1438 -3279 1444 -3275
rect 1446 -3279 1447 -3275
rect 1459 -3279 1460 -3275
rect 1462 -3279 1468 -3275
rect 1470 -3279 1472 -3275
rect 1476 -3279 1478 -3275
rect 1480 -3279 1486 -3275
rect 1488 -3279 1489 -3275
rect 1501 -3279 1502 -3275
rect 1504 -3279 1510 -3275
rect 1512 -3279 1513 -3275
rect -1260 -3393 -1259 -3389
rect -1257 -3393 -1255 -3389
rect -1251 -3393 -1249 -3389
rect -1247 -3393 -1246 -3389
rect -1234 -3393 -1233 -3389
rect -1231 -3393 -1225 -3389
rect -1223 -3393 -1222 -3389
rect -1210 -3393 -1209 -3389
rect -1207 -3393 -1201 -3389
rect -1199 -3393 -1197 -3389
rect -1193 -3393 -1191 -3389
rect -1189 -3393 -1183 -3389
rect -1181 -3393 -1180 -3389
rect -1168 -3393 -1167 -3389
rect -1165 -3393 -1159 -3389
rect -1157 -3393 -1155 -3389
rect -1151 -3393 -1149 -3389
rect -1147 -3393 -1141 -3389
rect -1139 -3393 -1138 -3389
rect -1126 -3393 -1125 -3389
rect -1123 -3393 -1117 -3389
rect -1115 -3393 -1113 -3389
rect -1109 -3393 -1107 -3389
rect -1105 -3393 -1099 -3389
rect -1097 -3393 -1096 -3389
rect -1084 -3393 -1083 -3389
rect -1081 -3393 -1075 -3389
rect -1073 -3393 -1072 -3389
rect -931 -3393 -930 -3389
rect -928 -3393 -926 -3389
rect -922 -3393 -920 -3389
rect -918 -3393 -917 -3389
rect -905 -3393 -904 -3389
rect -902 -3393 -896 -3389
rect -894 -3393 -893 -3389
rect -881 -3393 -880 -3389
rect -878 -3393 -872 -3389
rect -870 -3393 -868 -3389
rect -864 -3393 -862 -3389
rect -860 -3393 -854 -3389
rect -852 -3393 -851 -3389
rect -839 -3393 -838 -3389
rect -836 -3393 -830 -3389
rect -828 -3393 -826 -3389
rect -822 -3393 -820 -3389
rect -818 -3393 -812 -3389
rect -810 -3393 -809 -3389
rect -797 -3393 -796 -3389
rect -794 -3393 -788 -3389
rect -786 -3393 -784 -3389
rect -780 -3393 -778 -3389
rect -776 -3393 -770 -3389
rect -768 -3393 -767 -3389
rect -755 -3393 -754 -3389
rect -752 -3393 -746 -3389
rect -744 -3393 -743 -3389
rect -573 -3393 -572 -3389
rect -570 -3393 -568 -3389
rect -564 -3393 -562 -3389
rect -560 -3393 -559 -3389
rect -547 -3393 -546 -3389
rect -544 -3393 -538 -3389
rect -536 -3393 -535 -3389
rect -523 -3393 -522 -3389
rect -520 -3393 -514 -3389
rect -512 -3393 -510 -3389
rect -506 -3393 -504 -3389
rect -502 -3393 -496 -3389
rect -494 -3393 -493 -3389
rect -481 -3393 -480 -3389
rect -478 -3393 -472 -3389
rect -470 -3393 -468 -3389
rect -464 -3393 -462 -3389
rect -460 -3393 -454 -3389
rect -452 -3393 -451 -3389
rect -439 -3393 -438 -3389
rect -436 -3393 -430 -3389
rect -428 -3393 -426 -3389
rect -422 -3393 -420 -3389
rect -418 -3393 -412 -3389
rect -410 -3393 -409 -3389
rect -397 -3393 -396 -3389
rect -394 -3393 -388 -3389
rect -386 -3393 -385 -3389
rect -1335 -3510 -1334 -3506
rect -1332 -3510 -1326 -3506
rect -1324 -3510 -1322 -3506
rect -1318 -3510 -1316 -3506
rect -1314 -3510 -1313 -3506
rect -931 -3510 -930 -3506
rect -928 -3510 -922 -3506
rect -920 -3510 -918 -3506
rect -914 -3510 -912 -3506
rect -910 -3510 -909 -3506
rect -573 -3510 -572 -3506
rect -570 -3510 -564 -3506
rect -562 -3510 -560 -3506
rect -556 -3510 -554 -3506
rect -552 -3510 -551 -3506
rect -215 -3510 -214 -3506
rect -212 -3510 -206 -3506
rect -204 -3510 -202 -3506
rect -198 -3510 -196 -3506
rect -194 -3510 -193 -3506
rect 213 -3510 214 -3506
rect 216 -3510 222 -3506
rect 224 -3510 226 -3506
rect 230 -3510 232 -3506
rect 234 -3510 235 -3506
rect 569 -3510 570 -3506
rect 572 -3510 578 -3506
rect 580 -3510 582 -3506
rect 586 -3510 588 -3506
rect 590 -3510 591 -3506
rect 967 -3510 968 -3506
rect 970 -3510 976 -3506
rect 978 -3510 980 -3506
rect 984 -3510 986 -3506
rect 988 -3510 989 -3506
rect 1325 -3510 1326 -3506
rect 1328 -3510 1334 -3506
rect 1336 -3510 1338 -3506
rect 1342 -3510 1344 -3506
rect 1346 -3510 1347 -3506
rect -1260 -3634 -1259 -3630
rect -1257 -3634 -1255 -3630
rect -1251 -3634 -1249 -3630
rect -1247 -3634 -1246 -3630
rect -1234 -3634 -1233 -3630
rect -1231 -3634 -1229 -3630
rect -1225 -3634 -1223 -3630
rect -1221 -3634 -1215 -3630
rect -1213 -3634 -1211 -3630
rect -1207 -3634 -1205 -3630
rect -1203 -3634 -1202 -3630
rect -1190 -3634 -1189 -3630
rect -1187 -3634 -1181 -3630
rect -1179 -3634 -1177 -3630
rect -1173 -3634 -1171 -3630
rect -1169 -3634 -1168 -3630
rect -931 -3634 -930 -3630
rect -928 -3634 -926 -3630
rect -922 -3634 -920 -3630
rect -918 -3634 -917 -3630
rect -905 -3634 -904 -3630
rect -902 -3634 -900 -3630
rect -896 -3634 -894 -3630
rect -892 -3634 -891 -3630
rect -879 -3634 -878 -3630
rect -876 -3634 -875 -3630
rect -871 -3634 -868 -3630
rect -866 -3634 -860 -3630
rect -858 -3634 -857 -3630
rect -853 -3634 -850 -3630
rect -848 -3634 -847 -3630
rect -835 -3634 -834 -3630
rect -832 -3634 -826 -3630
rect -824 -3634 -822 -3630
rect -818 -3634 -816 -3630
rect -814 -3634 -813 -3630
rect -801 -3634 -800 -3630
rect -798 -3634 -796 -3630
rect -792 -3634 -790 -3630
rect -788 -3634 -782 -3630
rect -780 -3634 -778 -3630
rect -774 -3634 -772 -3630
rect -770 -3634 -769 -3630
rect -757 -3634 -756 -3630
rect -754 -3634 -748 -3630
rect -746 -3634 -745 -3630
rect -733 -3634 -732 -3630
rect -730 -3634 -725 -3630
rect -721 -3634 -716 -3630
rect -714 -3634 -713 -3630
rect -709 -3634 -708 -3630
rect -706 -3634 -704 -3630
rect -700 -3634 -698 -3630
rect -696 -3634 -695 -3630
rect -573 -3634 -572 -3630
rect -570 -3634 -568 -3630
rect -564 -3634 -562 -3630
rect -560 -3634 -559 -3630
rect -547 -3634 -546 -3630
rect -544 -3634 -542 -3630
rect -538 -3634 -536 -3630
rect -534 -3634 -533 -3630
rect -521 -3634 -520 -3630
rect -518 -3634 -517 -3630
rect -513 -3634 -510 -3630
rect -508 -3634 -502 -3630
rect -500 -3634 -499 -3630
rect -495 -3634 -492 -3630
rect -490 -3634 -489 -3630
rect -477 -3634 -476 -3630
rect -474 -3634 -468 -3630
rect -466 -3634 -464 -3630
rect -460 -3634 -458 -3630
rect -456 -3634 -455 -3630
rect -443 -3634 -442 -3630
rect -440 -3634 -438 -3630
rect -434 -3634 -432 -3630
rect -430 -3634 -424 -3630
rect -422 -3634 -420 -3630
rect -416 -3634 -414 -3630
rect -412 -3634 -411 -3630
rect -399 -3634 -398 -3630
rect -396 -3634 -390 -3630
rect -388 -3634 -387 -3630
rect -375 -3634 -374 -3630
rect -372 -3634 -367 -3630
rect -363 -3634 -358 -3630
rect -356 -3634 -355 -3630
rect -351 -3634 -350 -3630
rect -348 -3634 -346 -3630
rect -342 -3634 -340 -3630
rect -338 -3634 -337 -3630
rect -215 -3634 -214 -3630
rect -212 -3634 -210 -3630
rect -206 -3634 -204 -3630
rect -202 -3634 -201 -3630
rect -189 -3634 -188 -3630
rect -186 -3634 -184 -3630
rect -180 -3634 -178 -3630
rect -176 -3634 -175 -3630
rect -163 -3634 -162 -3630
rect -160 -3634 -159 -3630
rect -155 -3634 -152 -3630
rect -150 -3634 -144 -3630
rect -142 -3634 -141 -3630
rect -137 -3634 -134 -3630
rect -132 -3634 -131 -3630
rect -119 -3634 -118 -3630
rect -116 -3634 -110 -3630
rect -108 -3634 -106 -3630
rect -102 -3634 -100 -3630
rect -98 -3634 -97 -3630
rect -85 -3634 -84 -3630
rect -82 -3634 -80 -3630
rect -76 -3634 -74 -3630
rect -72 -3634 -66 -3630
rect -64 -3634 -62 -3630
rect -58 -3634 -56 -3630
rect -54 -3634 -53 -3630
rect -41 -3634 -40 -3630
rect -38 -3634 -32 -3630
rect -30 -3634 -29 -3630
rect -17 -3634 -16 -3630
rect -14 -3634 -9 -3630
rect -5 -3634 0 -3630
rect 2 -3634 3 -3630
rect 7 -3634 8 -3630
rect 10 -3634 12 -3630
rect 16 -3634 18 -3630
rect 20 -3634 21 -3630
rect 213 -3634 214 -3630
rect 216 -3634 218 -3630
rect 222 -3634 224 -3630
rect 226 -3634 227 -3630
rect 239 -3634 240 -3630
rect 242 -3634 244 -3630
rect 248 -3634 250 -3630
rect 252 -3634 253 -3630
rect 265 -3634 266 -3630
rect 268 -3634 269 -3630
rect 273 -3634 276 -3630
rect 278 -3634 284 -3630
rect 286 -3634 287 -3630
rect 291 -3634 294 -3630
rect 296 -3634 297 -3630
rect 309 -3634 310 -3630
rect 312 -3634 318 -3630
rect 320 -3634 322 -3630
rect 326 -3634 328 -3630
rect 330 -3634 331 -3630
rect 343 -3634 344 -3630
rect 346 -3634 348 -3630
rect 352 -3634 354 -3630
rect 356 -3634 362 -3630
rect 364 -3634 366 -3630
rect 370 -3634 372 -3630
rect 374 -3634 375 -3630
rect 387 -3634 388 -3630
rect 390 -3634 396 -3630
rect 398 -3634 399 -3630
rect 411 -3634 412 -3630
rect 414 -3634 419 -3630
rect 423 -3634 428 -3630
rect 430 -3634 431 -3630
rect 435 -3634 436 -3630
rect 438 -3634 440 -3630
rect 444 -3634 446 -3630
rect 448 -3634 449 -3630
rect 569 -3634 570 -3630
rect 572 -3634 574 -3630
rect 578 -3634 580 -3630
rect 582 -3634 583 -3630
rect 595 -3634 596 -3630
rect 598 -3634 600 -3630
rect 604 -3634 606 -3630
rect 608 -3634 609 -3630
rect 621 -3634 622 -3630
rect 624 -3634 625 -3630
rect 629 -3634 632 -3630
rect 634 -3634 640 -3630
rect 642 -3634 643 -3630
rect 647 -3634 650 -3630
rect 652 -3634 653 -3630
rect 665 -3634 666 -3630
rect 668 -3634 674 -3630
rect 676 -3634 678 -3630
rect 682 -3634 684 -3630
rect 686 -3634 687 -3630
rect 699 -3634 700 -3630
rect 702 -3634 704 -3630
rect 708 -3634 710 -3630
rect 712 -3634 718 -3630
rect 720 -3634 722 -3630
rect 726 -3634 728 -3630
rect 730 -3634 731 -3630
rect 743 -3634 744 -3630
rect 746 -3634 752 -3630
rect 754 -3634 755 -3630
rect 767 -3634 768 -3630
rect 770 -3634 775 -3630
rect 779 -3634 784 -3630
rect 786 -3634 787 -3630
rect 791 -3634 792 -3630
rect 794 -3634 796 -3630
rect 800 -3634 802 -3630
rect 804 -3634 805 -3630
rect 967 -3634 968 -3630
rect 970 -3634 972 -3630
rect 976 -3634 978 -3630
rect 980 -3634 981 -3630
rect 993 -3634 994 -3630
rect 996 -3634 998 -3630
rect 1002 -3634 1004 -3630
rect 1006 -3634 1007 -3630
rect 1019 -3634 1020 -3630
rect 1022 -3634 1023 -3630
rect 1027 -3634 1030 -3630
rect 1032 -3634 1038 -3630
rect 1040 -3634 1041 -3630
rect 1045 -3634 1048 -3630
rect 1050 -3634 1051 -3630
rect 1063 -3634 1064 -3630
rect 1066 -3634 1072 -3630
rect 1074 -3634 1076 -3630
rect 1080 -3634 1082 -3630
rect 1084 -3634 1085 -3630
rect 1097 -3634 1098 -3630
rect 1100 -3634 1102 -3630
rect 1106 -3634 1108 -3630
rect 1110 -3634 1116 -3630
rect 1118 -3634 1120 -3630
rect 1124 -3634 1126 -3630
rect 1128 -3634 1129 -3630
rect 1141 -3634 1142 -3630
rect 1144 -3634 1150 -3630
rect 1152 -3634 1153 -3630
rect 1165 -3634 1166 -3630
rect 1168 -3634 1173 -3630
rect 1177 -3634 1182 -3630
rect 1184 -3634 1185 -3630
rect 1189 -3634 1190 -3630
rect 1192 -3634 1194 -3630
rect 1198 -3634 1200 -3630
rect 1202 -3634 1203 -3630
rect 1325 -3634 1326 -3630
rect 1328 -3634 1330 -3630
rect 1334 -3634 1336 -3630
rect 1338 -3634 1339 -3630
rect 1351 -3634 1352 -3630
rect 1354 -3634 1356 -3630
rect 1360 -3634 1362 -3630
rect 1364 -3634 1365 -3630
rect 1377 -3634 1378 -3630
rect 1380 -3634 1381 -3630
rect 1385 -3634 1388 -3630
rect 1390 -3634 1396 -3630
rect 1398 -3634 1399 -3630
rect 1403 -3634 1406 -3630
rect 1408 -3634 1409 -3630
rect 1421 -3634 1422 -3630
rect 1424 -3634 1430 -3630
rect 1432 -3634 1434 -3630
rect 1438 -3634 1440 -3630
rect 1442 -3634 1443 -3630
rect 1455 -3634 1456 -3630
rect 1458 -3634 1460 -3630
rect 1464 -3634 1466 -3630
rect 1468 -3634 1474 -3630
rect 1476 -3634 1478 -3630
rect 1482 -3634 1484 -3630
rect 1486 -3634 1487 -3630
rect 1499 -3634 1500 -3630
rect 1502 -3634 1508 -3630
rect 1510 -3634 1511 -3630
rect 1523 -3634 1524 -3630
rect 1526 -3634 1531 -3630
rect 1535 -3634 1540 -3630
rect 1542 -3634 1543 -3630
rect 1547 -3634 1548 -3630
rect 1550 -3634 1552 -3630
rect 1556 -3634 1558 -3630
rect 1560 -3634 1561 -3630
rect -1260 -3764 -1259 -3760
rect -1257 -3764 -1255 -3760
rect -1251 -3764 -1249 -3760
rect -1247 -3764 -1246 -3760
rect -1234 -3764 -1233 -3760
rect -1231 -3764 -1225 -3760
rect -1223 -3764 -1222 -3760
rect -1210 -3764 -1209 -3760
rect -1207 -3764 -1201 -3760
rect -1199 -3764 -1197 -3760
rect -1193 -3764 -1191 -3760
rect -1189 -3764 -1183 -3760
rect -1181 -3764 -1180 -3760
rect -1168 -3764 -1167 -3760
rect -1165 -3764 -1159 -3760
rect -1157 -3764 -1155 -3760
rect -1151 -3764 -1149 -3760
rect -1147 -3764 -1141 -3760
rect -1139 -3764 -1138 -3760
rect -1126 -3764 -1125 -3760
rect -1123 -3764 -1117 -3760
rect -1115 -3764 -1113 -3760
rect -1109 -3764 -1107 -3760
rect -1105 -3764 -1099 -3760
rect -1097 -3764 -1096 -3760
rect -1084 -3764 -1083 -3760
rect -1081 -3764 -1075 -3760
rect -1073 -3764 -1072 -3760
rect -931 -3764 -930 -3760
rect -928 -3764 -926 -3760
rect -922 -3764 -920 -3760
rect -918 -3764 -917 -3760
rect -905 -3764 -904 -3760
rect -902 -3764 -896 -3760
rect -894 -3764 -893 -3760
rect -881 -3764 -880 -3760
rect -878 -3764 -872 -3760
rect -870 -3764 -868 -3760
rect -864 -3764 -862 -3760
rect -860 -3764 -854 -3760
rect -852 -3764 -851 -3760
rect -839 -3764 -838 -3760
rect -836 -3764 -830 -3760
rect -828 -3764 -826 -3760
rect -822 -3764 -820 -3760
rect -818 -3764 -812 -3760
rect -810 -3764 -809 -3760
rect -797 -3764 -796 -3760
rect -794 -3764 -788 -3760
rect -786 -3764 -784 -3760
rect -780 -3764 -778 -3760
rect -776 -3764 -770 -3760
rect -768 -3764 -767 -3760
rect -755 -3764 -754 -3760
rect -752 -3764 -746 -3760
rect -744 -3764 -743 -3760
rect -573 -3764 -572 -3760
rect -570 -3764 -568 -3760
rect -564 -3764 -562 -3760
rect -560 -3764 -559 -3760
rect -547 -3764 -546 -3760
rect -544 -3764 -538 -3760
rect -536 -3764 -535 -3760
rect -523 -3764 -522 -3760
rect -520 -3764 -514 -3760
rect -512 -3764 -510 -3760
rect -506 -3764 -504 -3760
rect -502 -3764 -496 -3760
rect -494 -3764 -493 -3760
rect -481 -3764 -480 -3760
rect -478 -3764 -472 -3760
rect -470 -3764 -468 -3760
rect -464 -3764 -462 -3760
rect -460 -3764 -454 -3760
rect -452 -3764 -451 -3760
rect -439 -3764 -438 -3760
rect -436 -3764 -430 -3760
rect -428 -3764 -426 -3760
rect -422 -3764 -420 -3760
rect -418 -3764 -412 -3760
rect -410 -3764 -409 -3760
rect -397 -3764 -396 -3760
rect -394 -3764 -388 -3760
rect -386 -3764 -385 -3760
rect -215 -3764 -214 -3760
rect -212 -3764 -210 -3760
rect -206 -3764 -204 -3760
rect -202 -3764 -201 -3760
rect -189 -3764 -188 -3760
rect -186 -3764 -180 -3760
rect -178 -3764 -177 -3760
rect -165 -3764 -164 -3760
rect -162 -3764 -156 -3760
rect -154 -3764 -152 -3760
rect -148 -3764 -146 -3760
rect -144 -3764 -138 -3760
rect -136 -3764 -135 -3760
rect -123 -3764 -122 -3760
rect -120 -3764 -114 -3760
rect -112 -3764 -110 -3760
rect -106 -3764 -104 -3760
rect -102 -3764 -96 -3760
rect -94 -3764 -93 -3760
rect -81 -3764 -80 -3760
rect -78 -3764 -72 -3760
rect -70 -3764 -68 -3760
rect -64 -3764 -62 -3760
rect -60 -3764 -54 -3760
rect -52 -3764 -51 -3760
rect -39 -3764 -38 -3760
rect -36 -3764 -30 -3760
rect -28 -3764 -27 -3760
rect 72 -3879 73 -3863
rect 75 -3879 76 -3863
rect -1260 -3995 -1259 -3991
rect -1257 -3995 -1255 -3991
rect -1251 -3995 -1249 -3991
rect -1247 -3995 -1246 -3991
rect -1234 -3995 -1233 -3991
rect -1231 -3995 -1225 -3991
rect -1223 -3995 -1222 -3991
rect -1210 -3995 -1209 -3991
rect -1207 -3995 -1201 -3991
rect -1199 -3995 -1197 -3991
rect -1193 -3995 -1191 -3991
rect -1189 -3995 -1183 -3991
rect -1181 -3995 -1180 -3991
rect -1168 -3995 -1167 -3991
rect -1165 -3995 -1159 -3991
rect -1157 -3995 -1155 -3991
rect -1151 -3995 -1149 -3991
rect -1147 -3995 -1141 -3991
rect -1139 -3995 -1138 -3991
rect -1126 -3995 -1125 -3991
rect -1123 -3995 -1117 -3991
rect -1115 -3995 -1113 -3991
rect -1109 -3995 -1107 -3991
rect -1105 -3995 -1099 -3991
rect -1097 -3995 -1096 -3991
rect -1084 -3995 -1083 -3991
rect -1081 -3995 -1075 -3991
rect -1073 -3995 -1072 -3991
rect -931 -3995 -930 -3991
rect -928 -3995 -926 -3991
rect -922 -3995 -920 -3991
rect -918 -3995 -917 -3991
rect -905 -3995 -904 -3991
rect -902 -3995 -896 -3991
rect -894 -3995 -893 -3991
rect -881 -3995 -880 -3991
rect -878 -3995 -872 -3991
rect -870 -3995 -868 -3991
rect -864 -3995 -862 -3991
rect -860 -3995 -854 -3991
rect -852 -3995 -851 -3991
rect -839 -3995 -838 -3991
rect -836 -3995 -830 -3991
rect -828 -3995 -826 -3991
rect -822 -3995 -820 -3991
rect -818 -3995 -812 -3991
rect -810 -3995 -809 -3991
rect -797 -3995 -796 -3991
rect -794 -3995 -788 -3991
rect -786 -3995 -784 -3991
rect -780 -3995 -778 -3991
rect -776 -3995 -770 -3991
rect -768 -3995 -767 -3991
rect -755 -3995 -754 -3991
rect -752 -3995 -746 -3991
rect -744 -3995 -743 -3991
rect -573 -3995 -572 -3991
rect -570 -3995 -568 -3991
rect -564 -3995 -562 -3991
rect -560 -3995 -559 -3991
rect -547 -3995 -546 -3991
rect -544 -3995 -538 -3991
rect -536 -3995 -535 -3991
rect -523 -3995 -522 -3991
rect -520 -3995 -514 -3991
rect -512 -3995 -510 -3991
rect -506 -3995 -504 -3991
rect -502 -3995 -496 -3991
rect -494 -3995 -493 -3991
rect -481 -3995 -480 -3991
rect -478 -3995 -472 -3991
rect -470 -3995 -468 -3991
rect -464 -3995 -462 -3991
rect -460 -3995 -454 -3991
rect -452 -3995 -451 -3991
rect -439 -3995 -438 -3991
rect -436 -3995 -430 -3991
rect -428 -3995 -426 -3991
rect -422 -3995 -420 -3991
rect -418 -3995 -412 -3991
rect -410 -3995 -409 -3991
rect -397 -3995 -396 -3991
rect -394 -3995 -388 -3991
rect -386 -3995 -385 -3991
rect -215 -3995 -214 -3991
rect -212 -3995 -210 -3991
rect -206 -3995 -204 -3991
rect -202 -3995 -201 -3991
rect -189 -3995 -188 -3991
rect -186 -3995 -180 -3991
rect -178 -3995 -177 -3991
rect -165 -3995 -164 -3991
rect -162 -3995 -156 -3991
rect -154 -3995 -152 -3991
rect -148 -3995 -146 -3991
rect -144 -3995 -138 -3991
rect -136 -3995 -135 -3991
rect -123 -3995 -122 -3991
rect -120 -3995 -114 -3991
rect -112 -3995 -110 -3991
rect -106 -3995 -104 -3991
rect -102 -3995 -96 -3991
rect -94 -3995 -93 -3991
rect -81 -3995 -80 -3991
rect -78 -3995 -72 -3991
rect -70 -3995 -68 -3991
rect -64 -3995 -62 -3991
rect -60 -3995 -54 -3991
rect -52 -3995 -51 -3991
rect -39 -3995 -38 -3991
rect -36 -3995 -30 -3991
rect -28 -3995 -27 -3991
rect 213 -3995 214 -3991
rect 216 -3995 218 -3991
rect 222 -3995 224 -3991
rect 226 -3995 227 -3991
rect 239 -3995 240 -3991
rect 242 -3995 248 -3991
rect 250 -3995 251 -3991
rect 263 -3995 264 -3991
rect 266 -3995 272 -3991
rect 274 -3995 276 -3991
rect 280 -3995 282 -3991
rect 284 -3995 290 -3991
rect 292 -3995 293 -3991
rect 305 -3995 306 -3991
rect 308 -3995 314 -3991
rect 316 -3995 318 -3991
rect 322 -3995 324 -3991
rect 326 -3995 332 -3991
rect 334 -3995 335 -3991
rect 347 -3995 348 -3991
rect 350 -3995 356 -3991
rect 358 -3995 360 -3991
rect 364 -3995 366 -3991
rect 368 -3995 374 -3991
rect 376 -3995 377 -3991
rect 389 -3995 390 -3991
rect 392 -3995 398 -3991
rect 400 -3995 401 -3991
rect 569 -3995 570 -3991
rect 572 -3995 574 -3991
rect 578 -3995 580 -3991
rect 582 -3995 583 -3991
rect 595 -3995 596 -3991
rect 598 -3995 604 -3991
rect 606 -3995 607 -3991
rect 619 -3995 620 -3991
rect 622 -3995 628 -3991
rect 630 -3995 632 -3991
rect 636 -3995 638 -3991
rect 640 -3995 646 -3991
rect 648 -3995 649 -3991
rect 661 -3995 662 -3991
rect 664 -3995 670 -3991
rect 672 -3995 674 -3991
rect 678 -3995 680 -3991
rect 682 -3995 688 -3991
rect 690 -3995 691 -3991
rect 703 -3995 704 -3991
rect 706 -3995 712 -3991
rect 714 -3995 716 -3991
rect 720 -3995 722 -3991
rect 724 -3995 730 -3991
rect 732 -3995 733 -3991
rect 745 -3995 746 -3991
rect 748 -3995 754 -3991
rect 756 -3995 757 -3991
rect 967 -3995 968 -3991
rect 970 -3995 972 -3991
rect 976 -3995 978 -3991
rect 980 -3995 981 -3991
rect 993 -3995 994 -3991
rect 996 -3995 1002 -3991
rect 1004 -3995 1005 -3991
rect 1017 -3995 1018 -3991
rect 1020 -3995 1026 -3991
rect 1028 -3995 1030 -3991
rect 1034 -3995 1036 -3991
rect 1038 -3995 1044 -3991
rect 1046 -3995 1047 -3991
rect 1059 -3995 1060 -3991
rect 1062 -3995 1068 -3991
rect 1070 -3995 1072 -3991
rect 1076 -3995 1078 -3991
rect 1080 -3995 1086 -3991
rect 1088 -3995 1089 -3991
rect 1101 -3995 1102 -3991
rect 1104 -3995 1110 -3991
rect 1112 -3995 1114 -3991
rect 1118 -3995 1120 -3991
rect 1122 -3995 1128 -3991
rect 1130 -3995 1131 -3991
rect 1143 -3995 1144 -3991
rect 1146 -3995 1152 -3991
rect 1154 -3995 1155 -3991
rect 1325 -3995 1326 -3991
rect 1328 -3995 1330 -3991
rect 1334 -3995 1336 -3991
rect 1338 -3995 1339 -3991
rect 1351 -3995 1352 -3991
rect 1354 -3995 1360 -3991
rect 1362 -3995 1363 -3991
rect 1375 -3995 1376 -3991
rect 1378 -3995 1384 -3991
rect 1386 -3995 1388 -3991
rect 1392 -3995 1394 -3991
rect 1396 -3995 1402 -3991
rect 1404 -3995 1405 -3991
rect 1417 -3995 1418 -3991
rect 1420 -3995 1426 -3991
rect 1428 -3995 1430 -3991
rect 1434 -3995 1436 -3991
rect 1438 -3995 1444 -3991
rect 1446 -3995 1447 -3991
rect 1459 -3995 1460 -3991
rect 1462 -3995 1468 -3991
rect 1470 -3995 1472 -3991
rect 1476 -3995 1478 -3991
rect 1480 -3995 1486 -3991
rect 1488 -3995 1489 -3991
rect 1501 -3995 1502 -3991
rect 1504 -3995 1510 -3991
rect 1512 -3995 1513 -3991
rect -1260 -4120 -1259 -4116
rect -1257 -4120 -1255 -4116
rect -1251 -4120 -1249 -4116
rect -1247 -4120 -1246 -4116
rect -1234 -4120 -1233 -4116
rect -1231 -4120 -1225 -4116
rect -1223 -4120 -1222 -4116
rect -1210 -4120 -1209 -4116
rect -1207 -4120 -1201 -4116
rect -1199 -4120 -1197 -4116
rect -1193 -4120 -1191 -4116
rect -1189 -4120 -1183 -4116
rect -1181 -4120 -1180 -4116
rect -1168 -4120 -1167 -4116
rect -1165 -4120 -1159 -4116
rect -1157 -4120 -1155 -4116
rect -1151 -4120 -1149 -4116
rect -1147 -4120 -1141 -4116
rect -1139 -4120 -1138 -4116
rect -1126 -4120 -1125 -4116
rect -1123 -4120 -1117 -4116
rect -1115 -4120 -1113 -4116
rect -1109 -4120 -1107 -4116
rect -1105 -4120 -1099 -4116
rect -1097 -4120 -1096 -4116
rect -1084 -4120 -1083 -4116
rect -1081 -4120 -1075 -4116
rect -1073 -4120 -1072 -4116
rect -931 -4120 -930 -4116
rect -928 -4120 -926 -4116
rect -922 -4120 -920 -4116
rect -918 -4120 -917 -4116
rect -905 -4120 -904 -4116
rect -902 -4120 -896 -4116
rect -894 -4120 -893 -4116
rect -881 -4120 -880 -4116
rect -878 -4120 -872 -4116
rect -870 -4120 -868 -4116
rect -864 -4120 -862 -4116
rect -860 -4120 -854 -4116
rect -852 -4120 -851 -4116
rect -839 -4120 -838 -4116
rect -836 -4120 -830 -4116
rect -828 -4120 -826 -4116
rect -822 -4120 -820 -4116
rect -818 -4120 -812 -4116
rect -810 -4120 -809 -4116
rect -797 -4120 -796 -4116
rect -794 -4120 -788 -4116
rect -786 -4120 -784 -4116
rect -780 -4120 -778 -4116
rect -776 -4120 -770 -4116
rect -768 -4120 -767 -4116
rect -755 -4120 -754 -4116
rect -752 -4120 -746 -4116
rect -744 -4120 -743 -4116
rect -573 -4120 -572 -4116
rect -570 -4120 -568 -4116
rect -564 -4120 -562 -4116
rect -560 -4120 -559 -4116
rect -547 -4120 -546 -4116
rect -544 -4120 -538 -4116
rect -536 -4120 -535 -4116
rect -523 -4120 -522 -4116
rect -520 -4120 -514 -4116
rect -512 -4120 -510 -4116
rect -506 -4120 -504 -4116
rect -502 -4120 -496 -4116
rect -494 -4120 -493 -4116
rect -481 -4120 -480 -4116
rect -478 -4120 -472 -4116
rect -470 -4120 -468 -4116
rect -464 -4120 -462 -4116
rect -460 -4120 -454 -4116
rect -452 -4120 -451 -4116
rect -439 -4120 -438 -4116
rect -436 -4120 -430 -4116
rect -428 -4120 -426 -4116
rect -422 -4120 -420 -4116
rect -418 -4120 -412 -4116
rect -410 -4120 -409 -4116
rect -397 -4120 -396 -4116
rect -394 -4120 -388 -4116
rect -386 -4120 -385 -4116
rect -215 -4120 -214 -4116
rect -212 -4120 -210 -4116
rect -206 -4120 -204 -4116
rect -202 -4120 -201 -4116
rect -189 -4120 -188 -4116
rect -186 -4120 -180 -4116
rect -178 -4120 -177 -4116
rect -165 -4120 -164 -4116
rect -162 -4120 -156 -4116
rect -154 -4120 -152 -4116
rect -148 -4120 -146 -4116
rect -144 -4120 -138 -4116
rect -136 -4120 -135 -4116
rect -123 -4120 -122 -4116
rect -120 -4120 -114 -4116
rect -112 -4120 -110 -4116
rect -106 -4120 -104 -4116
rect -102 -4120 -96 -4116
rect -94 -4120 -93 -4116
rect -81 -4120 -80 -4116
rect -78 -4120 -72 -4116
rect -70 -4120 -68 -4116
rect -64 -4120 -62 -4116
rect -60 -4120 -54 -4116
rect -52 -4120 -51 -4116
rect -39 -4120 -38 -4116
rect -36 -4120 -30 -4116
rect -28 -4120 -27 -4116
rect 213 -4120 214 -4116
rect 216 -4120 218 -4116
rect 222 -4120 224 -4116
rect 226 -4120 227 -4116
rect 239 -4120 240 -4116
rect 242 -4120 248 -4116
rect 250 -4120 251 -4116
rect 263 -4120 264 -4116
rect 266 -4120 272 -4116
rect 274 -4120 276 -4116
rect 280 -4120 282 -4116
rect 284 -4120 290 -4116
rect 292 -4120 293 -4116
rect 305 -4120 306 -4116
rect 308 -4120 314 -4116
rect 316 -4120 318 -4116
rect 322 -4120 324 -4116
rect 326 -4120 332 -4116
rect 334 -4120 335 -4116
rect 347 -4120 348 -4116
rect 350 -4120 356 -4116
rect 358 -4120 360 -4116
rect 364 -4120 366 -4116
rect 368 -4120 374 -4116
rect 376 -4120 377 -4116
rect 389 -4120 390 -4116
rect 392 -4120 398 -4116
rect 400 -4120 401 -4116
rect 569 -4120 570 -4116
rect 572 -4120 574 -4116
rect 578 -4120 580 -4116
rect 582 -4120 583 -4116
rect 595 -4120 596 -4116
rect 598 -4120 604 -4116
rect 606 -4120 607 -4116
rect 619 -4120 620 -4116
rect 622 -4120 628 -4116
rect 630 -4120 632 -4116
rect 636 -4120 638 -4116
rect 640 -4120 646 -4116
rect 648 -4120 649 -4116
rect 661 -4120 662 -4116
rect 664 -4120 670 -4116
rect 672 -4120 674 -4116
rect 678 -4120 680 -4116
rect 682 -4120 688 -4116
rect 690 -4120 691 -4116
rect 703 -4120 704 -4116
rect 706 -4120 712 -4116
rect 714 -4120 716 -4116
rect 720 -4120 722 -4116
rect 724 -4120 730 -4116
rect 732 -4120 733 -4116
rect 745 -4120 746 -4116
rect 748 -4120 754 -4116
rect 756 -4120 757 -4116
rect 967 -4120 968 -4116
rect 970 -4120 972 -4116
rect 976 -4120 978 -4116
rect 980 -4120 981 -4116
rect 993 -4120 994 -4116
rect 996 -4120 1002 -4116
rect 1004 -4120 1005 -4116
rect 1017 -4120 1018 -4116
rect 1020 -4120 1026 -4116
rect 1028 -4120 1030 -4116
rect 1034 -4120 1036 -4116
rect 1038 -4120 1044 -4116
rect 1046 -4120 1047 -4116
rect 1059 -4120 1060 -4116
rect 1062 -4120 1068 -4116
rect 1070 -4120 1072 -4116
rect 1076 -4120 1078 -4116
rect 1080 -4120 1086 -4116
rect 1088 -4120 1089 -4116
rect 1101 -4120 1102 -4116
rect 1104 -4120 1110 -4116
rect 1112 -4120 1114 -4116
rect 1118 -4120 1120 -4116
rect 1122 -4120 1128 -4116
rect 1130 -4120 1131 -4116
rect 1143 -4120 1144 -4116
rect 1146 -4120 1152 -4116
rect 1154 -4120 1155 -4116
rect 1325 -4120 1326 -4116
rect 1328 -4120 1330 -4116
rect 1334 -4120 1336 -4116
rect 1338 -4120 1339 -4116
rect 1351 -4120 1352 -4116
rect 1354 -4120 1360 -4116
rect 1362 -4120 1363 -4116
rect 1375 -4120 1376 -4116
rect 1378 -4120 1384 -4116
rect 1386 -4120 1388 -4116
rect 1392 -4120 1394 -4116
rect 1396 -4120 1402 -4116
rect 1404 -4120 1405 -4116
rect 1417 -4120 1418 -4116
rect 1420 -4120 1426 -4116
rect 1428 -4120 1430 -4116
rect 1434 -4120 1436 -4116
rect 1438 -4120 1444 -4116
rect 1446 -4120 1447 -4116
rect 1459 -4120 1460 -4116
rect 1462 -4120 1468 -4116
rect 1470 -4120 1472 -4116
rect 1476 -4120 1478 -4116
rect 1480 -4120 1486 -4116
rect 1488 -4120 1489 -4116
rect 1501 -4120 1502 -4116
rect 1504 -4120 1510 -4116
rect 1512 -4120 1513 -4116
rect -1260 -4244 -1259 -4240
rect -1257 -4244 -1255 -4240
rect -1251 -4244 -1249 -4240
rect -1247 -4244 -1246 -4240
rect -1234 -4244 -1233 -4240
rect -1231 -4244 -1225 -4240
rect -1223 -4244 -1222 -4240
rect -1210 -4244 -1209 -4240
rect -1207 -4244 -1201 -4240
rect -1199 -4244 -1197 -4240
rect -1193 -4244 -1191 -4240
rect -1189 -4244 -1183 -4240
rect -1181 -4244 -1180 -4240
rect -1168 -4244 -1167 -4240
rect -1165 -4244 -1159 -4240
rect -1157 -4244 -1155 -4240
rect -1151 -4244 -1149 -4240
rect -1147 -4244 -1141 -4240
rect -1139 -4244 -1138 -4240
rect -1126 -4244 -1125 -4240
rect -1123 -4244 -1117 -4240
rect -1115 -4244 -1113 -4240
rect -1109 -4244 -1107 -4240
rect -1105 -4244 -1099 -4240
rect -1097 -4244 -1096 -4240
rect -1084 -4244 -1083 -4240
rect -1081 -4244 -1075 -4240
rect -1073 -4244 -1072 -4240
rect -1025 -4244 -1024 -4240
rect -1022 -4244 -1021 -4240
rect -931 -4244 -930 -4240
rect -928 -4244 -926 -4240
rect -922 -4244 -920 -4240
rect -918 -4244 -917 -4240
rect -905 -4244 -904 -4240
rect -902 -4244 -896 -4240
rect -894 -4244 -893 -4240
rect -881 -4244 -880 -4240
rect -878 -4244 -872 -4240
rect -870 -4244 -868 -4240
rect -864 -4244 -862 -4240
rect -860 -4244 -854 -4240
rect -852 -4244 -851 -4240
rect -839 -4244 -838 -4240
rect -836 -4244 -830 -4240
rect -828 -4244 -826 -4240
rect -822 -4244 -820 -4240
rect -818 -4244 -812 -4240
rect -810 -4244 -809 -4240
rect -797 -4244 -796 -4240
rect -794 -4244 -788 -4240
rect -786 -4244 -784 -4240
rect -780 -4244 -778 -4240
rect -776 -4244 -770 -4240
rect -768 -4244 -767 -4240
rect -755 -4244 -754 -4240
rect -752 -4244 -746 -4240
rect -744 -4244 -743 -4240
rect -573 -4244 -572 -4240
rect -570 -4244 -568 -4240
rect -564 -4244 -562 -4240
rect -560 -4244 -559 -4240
rect -547 -4244 -546 -4240
rect -544 -4244 -538 -4240
rect -536 -4244 -535 -4240
rect -523 -4244 -522 -4240
rect -520 -4244 -514 -4240
rect -512 -4244 -510 -4240
rect -506 -4244 -504 -4240
rect -502 -4244 -496 -4240
rect -494 -4244 -493 -4240
rect -481 -4244 -480 -4240
rect -478 -4244 -472 -4240
rect -470 -4244 -468 -4240
rect -464 -4244 -462 -4240
rect -460 -4244 -454 -4240
rect -452 -4244 -451 -4240
rect -439 -4244 -438 -4240
rect -436 -4244 -430 -4240
rect -428 -4244 -426 -4240
rect -422 -4244 -420 -4240
rect -418 -4244 -412 -4240
rect -410 -4244 -409 -4240
rect -397 -4244 -396 -4240
rect -394 -4244 -388 -4240
rect -386 -4244 -385 -4240
rect -328 -4244 -327 -4240
rect -325 -4244 -324 -4240
rect -215 -4244 -214 -4240
rect -212 -4244 -210 -4240
rect -206 -4244 -204 -4240
rect -202 -4244 -201 -4240
rect -189 -4244 -188 -4240
rect -186 -4244 -180 -4240
rect -178 -4244 -177 -4240
rect -165 -4244 -164 -4240
rect -162 -4244 -156 -4240
rect -154 -4244 -152 -4240
rect -148 -4244 -146 -4240
rect -144 -4244 -138 -4240
rect -136 -4244 -135 -4240
rect -123 -4244 -122 -4240
rect -120 -4244 -114 -4240
rect -112 -4244 -110 -4240
rect -106 -4244 -104 -4240
rect -102 -4244 -96 -4240
rect -94 -4244 -93 -4240
rect -81 -4244 -80 -4240
rect -78 -4244 -72 -4240
rect -70 -4244 -68 -4240
rect -64 -4244 -62 -4240
rect -60 -4244 -54 -4240
rect -52 -4244 -51 -4240
rect -39 -4244 -38 -4240
rect -36 -4244 -30 -4240
rect -28 -4244 -27 -4240
rect 460 -4244 461 -4240
rect 463 -4244 464 -4240
rect 1205 -4244 1206 -4240
rect 1208 -4244 1209 -4240
rect -1335 -4355 -1334 -4351
rect -1332 -4355 -1326 -4351
rect -1324 -4355 -1322 -4351
rect -1318 -4355 -1316 -4351
rect -1314 -4355 -1313 -4351
rect -1025 -4355 -1024 -4351
rect -1022 -4355 -1021 -4351
rect -931 -4355 -930 -4351
rect -928 -4355 -922 -4351
rect -920 -4355 -918 -4351
rect -914 -4355 -912 -4351
rect -910 -4355 -909 -4351
rect -669 -4355 -668 -4347
rect -666 -4355 -665 -4347
rect -573 -4355 -572 -4351
rect -570 -4355 -564 -4351
rect -562 -4355 -560 -4351
rect -556 -4355 -554 -4351
rect -552 -4355 -551 -4351
rect -328 -4355 -327 -4351
rect -325 -4355 -324 -4351
rect -215 -4355 -214 -4351
rect -212 -4355 -206 -4351
rect -204 -4355 -202 -4351
rect -198 -4355 -196 -4351
rect -194 -4355 -193 -4351
rect 213 -4355 214 -4351
rect 216 -4355 222 -4351
rect 224 -4355 226 -4351
rect 230 -4355 232 -4351
rect 234 -4355 235 -4351
rect 460 -4355 461 -4351
rect 463 -4355 464 -4351
rect 569 -4355 570 -4351
rect 572 -4355 578 -4351
rect 580 -4355 582 -4351
rect 586 -4355 588 -4351
rect 590 -4355 591 -4351
rect 864 -4355 865 -4347
rect 867 -4355 868 -4347
rect 967 -4355 968 -4351
rect 970 -4355 976 -4351
rect 978 -4355 980 -4351
rect 984 -4355 986 -4351
rect 988 -4355 989 -4351
rect 1205 -4355 1206 -4351
rect 1208 -4355 1209 -4351
rect 1325 -4355 1326 -4351
rect 1328 -4355 1334 -4351
rect 1336 -4355 1338 -4351
rect 1342 -4355 1344 -4351
rect 1346 -4355 1347 -4351
rect -1260 -4474 -1259 -4470
rect -1257 -4474 -1255 -4470
rect -1251 -4474 -1249 -4470
rect -1247 -4474 -1246 -4470
rect -1234 -4474 -1233 -4470
rect -1231 -4474 -1229 -4470
rect -1225 -4474 -1223 -4470
rect -1221 -4474 -1215 -4470
rect -1213 -4474 -1211 -4470
rect -1207 -4474 -1205 -4470
rect -1203 -4474 -1202 -4470
rect -1190 -4474 -1189 -4470
rect -1187 -4474 -1181 -4470
rect -1179 -4474 -1177 -4470
rect -1173 -4474 -1171 -4470
rect -1169 -4474 -1168 -4470
rect -931 -4474 -930 -4470
rect -928 -4474 -926 -4470
rect -922 -4474 -920 -4470
rect -918 -4474 -917 -4470
rect -905 -4474 -904 -4470
rect -902 -4474 -900 -4470
rect -896 -4474 -894 -4470
rect -892 -4474 -891 -4470
rect -879 -4474 -878 -4470
rect -876 -4474 -875 -4470
rect -871 -4474 -868 -4470
rect -866 -4474 -860 -4470
rect -858 -4474 -857 -4470
rect -853 -4474 -850 -4470
rect -848 -4474 -847 -4470
rect -835 -4474 -834 -4470
rect -832 -4474 -826 -4470
rect -824 -4474 -822 -4470
rect -818 -4474 -816 -4470
rect -814 -4474 -813 -4470
rect -801 -4474 -800 -4470
rect -798 -4474 -796 -4470
rect -792 -4474 -790 -4470
rect -788 -4474 -782 -4470
rect -780 -4474 -778 -4470
rect -774 -4474 -772 -4470
rect -770 -4474 -769 -4470
rect -757 -4474 -756 -4470
rect -754 -4474 -748 -4470
rect -746 -4474 -745 -4470
rect -733 -4474 -732 -4470
rect -730 -4474 -725 -4470
rect -721 -4474 -716 -4470
rect -714 -4474 -713 -4470
rect -709 -4474 -708 -4470
rect -706 -4474 -704 -4470
rect -700 -4474 -698 -4470
rect -696 -4474 -695 -4470
rect -573 -4474 -572 -4470
rect -570 -4474 -568 -4470
rect -564 -4474 -562 -4470
rect -560 -4474 -559 -4470
rect -547 -4474 -546 -4470
rect -544 -4474 -542 -4470
rect -538 -4474 -536 -4470
rect -534 -4474 -533 -4470
rect -521 -4474 -520 -4470
rect -518 -4474 -517 -4470
rect -513 -4474 -510 -4470
rect -508 -4474 -502 -4470
rect -500 -4474 -499 -4470
rect -495 -4474 -492 -4470
rect -490 -4474 -489 -4470
rect -477 -4474 -476 -4470
rect -474 -4474 -468 -4470
rect -466 -4474 -464 -4470
rect -460 -4474 -458 -4470
rect -456 -4474 -455 -4470
rect -443 -4474 -442 -4470
rect -440 -4474 -438 -4470
rect -434 -4474 -432 -4470
rect -430 -4474 -424 -4470
rect -422 -4474 -420 -4470
rect -416 -4474 -414 -4470
rect -412 -4474 -411 -4470
rect -399 -4474 -398 -4470
rect -396 -4474 -390 -4470
rect -388 -4474 -387 -4470
rect -375 -4474 -374 -4470
rect -372 -4474 -367 -4470
rect -363 -4474 -358 -4470
rect -356 -4474 -355 -4470
rect -351 -4474 -350 -4470
rect -348 -4474 -346 -4470
rect -342 -4474 -340 -4470
rect -338 -4474 -337 -4470
rect -215 -4474 -214 -4470
rect -212 -4474 -210 -4470
rect -206 -4474 -204 -4470
rect -202 -4474 -201 -4470
rect -189 -4474 -188 -4470
rect -186 -4474 -184 -4470
rect -180 -4474 -178 -4470
rect -176 -4474 -175 -4470
rect -163 -4474 -162 -4470
rect -160 -4474 -159 -4470
rect -155 -4474 -152 -4470
rect -150 -4474 -144 -4470
rect -142 -4474 -141 -4470
rect -137 -4474 -134 -4470
rect -132 -4474 -131 -4470
rect -119 -4474 -118 -4470
rect -116 -4474 -110 -4470
rect -108 -4474 -106 -4470
rect -102 -4474 -100 -4470
rect -98 -4474 -97 -4470
rect -85 -4474 -84 -4470
rect -82 -4474 -80 -4470
rect -76 -4474 -74 -4470
rect -72 -4474 -66 -4470
rect -64 -4474 -62 -4470
rect -58 -4474 -56 -4470
rect -54 -4474 -53 -4470
rect -41 -4474 -40 -4470
rect -38 -4474 -32 -4470
rect -30 -4474 -29 -4470
rect -17 -4474 -16 -4470
rect -14 -4474 -9 -4470
rect -5 -4474 0 -4470
rect 2 -4474 3 -4470
rect 7 -4474 8 -4470
rect 10 -4474 12 -4470
rect 16 -4474 18 -4470
rect 20 -4474 21 -4470
rect 213 -4474 214 -4470
rect 216 -4474 218 -4470
rect 222 -4474 224 -4470
rect 226 -4474 227 -4470
rect 239 -4474 240 -4470
rect 242 -4474 244 -4470
rect 248 -4474 250 -4470
rect 252 -4474 253 -4470
rect 265 -4474 266 -4470
rect 268 -4474 269 -4470
rect 273 -4474 276 -4470
rect 278 -4474 284 -4470
rect 286 -4474 287 -4470
rect 291 -4474 294 -4470
rect 296 -4474 297 -4470
rect 309 -4474 310 -4470
rect 312 -4474 318 -4470
rect 320 -4474 322 -4470
rect 326 -4474 328 -4470
rect 330 -4474 331 -4470
rect 343 -4474 344 -4470
rect 346 -4474 348 -4470
rect 352 -4474 354 -4470
rect 356 -4474 362 -4470
rect 364 -4474 366 -4470
rect 370 -4474 372 -4470
rect 374 -4474 375 -4470
rect 387 -4474 388 -4470
rect 390 -4474 396 -4470
rect 398 -4474 399 -4470
rect 411 -4474 412 -4470
rect 414 -4474 419 -4470
rect 423 -4474 428 -4470
rect 430 -4474 431 -4470
rect 435 -4474 436 -4470
rect 438 -4474 440 -4470
rect 444 -4474 446 -4470
rect 448 -4474 449 -4470
rect 569 -4474 570 -4470
rect 572 -4474 574 -4470
rect 578 -4474 580 -4470
rect 582 -4474 583 -4470
rect 595 -4474 596 -4470
rect 598 -4474 600 -4470
rect 604 -4474 606 -4470
rect 608 -4474 609 -4470
rect 621 -4474 622 -4470
rect 624 -4474 625 -4470
rect 629 -4474 632 -4470
rect 634 -4474 640 -4470
rect 642 -4474 643 -4470
rect 647 -4474 650 -4470
rect 652 -4474 653 -4470
rect 665 -4474 666 -4470
rect 668 -4474 674 -4470
rect 676 -4474 678 -4470
rect 682 -4474 684 -4470
rect 686 -4474 687 -4470
rect 699 -4474 700 -4470
rect 702 -4474 704 -4470
rect 708 -4474 710 -4470
rect 712 -4474 718 -4470
rect 720 -4474 722 -4470
rect 726 -4474 728 -4470
rect 730 -4474 731 -4470
rect 743 -4474 744 -4470
rect 746 -4474 752 -4470
rect 754 -4474 755 -4470
rect 767 -4474 768 -4470
rect 770 -4474 775 -4470
rect 779 -4474 784 -4470
rect 786 -4474 787 -4470
rect 791 -4474 792 -4470
rect 794 -4474 796 -4470
rect 800 -4474 802 -4470
rect 804 -4474 805 -4470
rect 967 -4474 968 -4470
rect 970 -4474 972 -4470
rect 976 -4474 978 -4470
rect 980 -4474 981 -4470
rect 993 -4474 994 -4470
rect 996 -4474 998 -4470
rect 1002 -4474 1004 -4470
rect 1006 -4474 1007 -4470
rect 1019 -4474 1020 -4470
rect 1022 -4474 1023 -4470
rect 1027 -4474 1030 -4470
rect 1032 -4474 1038 -4470
rect 1040 -4474 1041 -4470
rect 1045 -4474 1048 -4470
rect 1050 -4474 1051 -4470
rect 1063 -4474 1064 -4470
rect 1066 -4474 1072 -4470
rect 1074 -4474 1076 -4470
rect 1080 -4474 1082 -4470
rect 1084 -4474 1085 -4470
rect 1097 -4474 1098 -4470
rect 1100 -4474 1102 -4470
rect 1106 -4474 1108 -4470
rect 1110 -4474 1116 -4470
rect 1118 -4474 1120 -4470
rect 1124 -4474 1126 -4470
rect 1128 -4474 1129 -4470
rect 1141 -4474 1142 -4470
rect 1144 -4474 1150 -4470
rect 1152 -4474 1153 -4470
rect 1165 -4474 1166 -4470
rect 1168 -4474 1173 -4470
rect 1177 -4474 1182 -4470
rect 1184 -4474 1185 -4470
rect 1189 -4474 1190 -4470
rect 1192 -4474 1194 -4470
rect 1198 -4474 1200 -4470
rect 1202 -4474 1203 -4470
rect 1325 -4474 1326 -4470
rect 1328 -4474 1330 -4470
rect 1334 -4474 1336 -4470
rect 1338 -4474 1339 -4470
rect 1351 -4474 1352 -4470
rect 1354 -4474 1356 -4470
rect 1360 -4474 1362 -4470
rect 1364 -4474 1365 -4470
rect 1377 -4474 1378 -4470
rect 1380 -4474 1381 -4470
rect 1385 -4474 1388 -4470
rect 1390 -4474 1396 -4470
rect 1398 -4474 1399 -4470
rect 1403 -4474 1406 -4470
rect 1408 -4474 1409 -4470
rect 1421 -4474 1422 -4470
rect 1424 -4474 1430 -4470
rect 1432 -4474 1434 -4470
rect 1438 -4474 1440 -4470
rect 1442 -4474 1443 -4470
rect 1455 -4474 1456 -4470
rect 1458 -4474 1460 -4470
rect 1464 -4474 1466 -4470
rect 1468 -4474 1474 -4470
rect 1476 -4474 1478 -4470
rect 1482 -4474 1484 -4470
rect 1486 -4474 1487 -4470
rect 1499 -4474 1500 -4470
rect 1502 -4474 1508 -4470
rect 1510 -4474 1511 -4470
rect 1523 -4474 1524 -4470
rect 1526 -4474 1531 -4470
rect 1535 -4474 1540 -4470
rect 1542 -4474 1543 -4470
rect 1547 -4474 1548 -4470
rect 1550 -4474 1552 -4470
rect 1556 -4474 1558 -4470
rect 1560 -4474 1561 -4470
rect -1260 -4597 -1259 -4593
rect -1257 -4597 -1255 -4593
rect -1251 -4597 -1249 -4593
rect -1247 -4597 -1246 -4593
rect -1234 -4597 -1233 -4593
rect -1231 -4597 -1225 -4593
rect -1223 -4597 -1222 -4593
rect -1210 -4597 -1209 -4593
rect -1207 -4597 -1201 -4593
rect -1199 -4597 -1197 -4593
rect -1193 -4597 -1191 -4593
rect -1189 -4597 -1183 -4593
rect -1181 -4597 -1180 -4593
rect -1168 -4597 -1167 -4593
rect -1165 -4597 -1159 -4593
rect -1157 -4597 -1155 -4593
rect -1151 -4597 -1149 -4593
rect -1147 -4597 -1141 -4593
rect -1139 -4597 -1138 -4593
rect -1126 -4597 -1125 -4593
rect -1123 -4597 -1117 -4593
rect -1115 -4597 -1113 -4593
rect -1109 -4597 -1107 -4593
rect -1105 -4597 -1099 -4593
rect -1097 -4597 -1096 -4593
rect -1084 -4597 -1083 -4593
rect -1081 -4597 -1075 -4593
rect -1073 -4597 -1072 -4593
rect -931 -4597 -930 -4593
rect -928 -4597 -926 -4593
rect -922 -4597 -920 -4593
rect -918 -4597 -917 -4593
rect -905 -4597 -904 -4593
rect -902 -4597 -896 -4593
rect -894 -4597 -893 -4593
rect -881 -4597 -880 -4593
rect -878 -4597 -872 -4593
rect -870 -4597 -868 -4593
rect -864 -4597 -862 -4593
rect -860 -4597 -854 -4593
rect -852 -4597 -851 -4593
rect -839 -4597 -838 -4593
rect -836 -4597 -830 -4593
rect -828 -4597 -826 -4593
rect -822 -4597 -820 -4593
rect -818 -4597 -812 -4593
rect -810 -4597 -809 -4593
rect -797 -4597 -796 -4593
rect -794 -4597 -788 -4593
rect -786 -4597 -784 -4593
rect -780 -4597 -778 -4593
rect -776 -4597 -770 -4593
rect -768 -4597 -767 -4593
rect -755 -4597 -754 -4593
rect -752 -4597 -746 -4593
rect -744 -4597 -743 -4593
rect -573 -4597 -572 -4593
rect -570 -4597 -568 -4593
rect -564 -4597 -562 -4593
rect -560 -4597 -559 -4593
rect -547 -4597 -546 -4593
rect -544 -4597 -538 -4593
rect -536 -4597 -535 -4593
rect -523 -4597 -522 -4593
rect -520 -4597 -514 -4593
rect -512 -4597 -510 -4593
rect -506 -4597 -504 -4593
rect -502 -4597 -496 -4593
rect -494 -4597 -493 -4593
rect -481 -4597 -480 -4593
rect -478 -4597 -472 -4593
rect -470 -4597 -468 -4593
rect -464 -4597 -462 -4593
rect -460 -4597 -454 -4593
rect -452 -4597 -451 -4593
rect -439 -4597 -438 -4593
rect -436 -4597 -430 -4593
rect -428 -4597 -426 -4593
rect -422 -4597 -420 -4593
rect -418 -4597 -412 -4593
rect -410 -4597 -409 -4593
rect -397 -4597 -396 -4593
rect -394 -4597 -388 -4593
rect -386 -4597 -385 -4593
rect -1260 -4718 -1259 -4714
rect -1257 -4718 -1255 -4714
rect -1251 -4718 -1249 -4714
rect -1247 -4718 -1246 -4714
rect -1234 -4718 -1233 -4714
rect -1231 -4718 -1225 -4714
rect -1223 -4718 -1222 -4714
rect -1210 -4718 -1209 -4714
rect -1207 -4718 -1201 -4714
rect -1199 -4718 -1197 -4714
rect -1193 -4718 -1191 -4714
rect -1189 -4718 -1183 -4714
rect -1181 -4718 -1180 -4714
rect -1168 -4718 -1167 -4714
rect -1165 -4718 -1159 -4714
rect -1157 -4718 -1155 -4714
rect -1151 -4718 -1149 -4714
rect -1147 -4718 -1141 -4714
rect -1139 -4718 -1138 -4714
rect -1126 -4718 -1125 -4714
rect -1123 -4718 -1117 -4714
rect -1115 -4718 -1113 -4714
rect -1109 -4718 -1107 -4714
rect -1105 -4718 -1099 -4714
rect -1097 -4718 -1096 -4714
rect -1084 -4718 -1083 -4714
rect -1081 -4718 -1075 -4714
rect -1073 -4718 -1072 -4714
rect -931 -4718 -930 -4714
rect -928 -4718 -926 -4714
rect -922 -4718 -920 -4714
rect -918 -4718 -917 -4714
rect -905 -4718 -904 -4714
rect -902 -4718 -896 -4714
rect -894 -4718 -893 -4714
rect -881 -4718 -880 -4714
rect -878 -4718 -872 -4714
rect -870 -4718 -868 -4714
rect -864 -4718 -862 -4714
rect -860 -4718 -854 -4714
rect -852 -4718 -851 -4714
rect -839 -4718 -838 -4714
rect -836 -4718 -830 -4714
rect -828 -4718 -826 -4714
rect -822 -4718 -820 -4714
rect -818 -4718 -812 -4714
rect -810 -4718 -809 -4714
rect -797 -4718 -796 -4714
rect -794 -4718 -788 -4714
rect -786 -4718 -784 -4714
rect -780 -4718 -778 -4714
rect -776 -4718 -770 -4714
rect -768 -4718 -767 -4714
rect -755 -4718 -754 -4714
rect -752 -4718 -746 -4714
rect -744 -4718 -743 -4714
rect -573 -4718 -572 -4714
rect -570 -4718 -568 -4714
rect -564 -4718 -562 -4714
rect -560 -4718 -559 -4714
rect -547 -4718 -546 -4714
rect -544 -4718 -538 -4714
rect -536 -4718 -535 -4714
rect -523 -4718 -522 -4714
rect -520 -4718 -514 -4714
rect -512 -4718 -510 -4714
rect -506 -4718 -504 -4714
rect -502 -4718 -496 -4714
rect -494 -4718 -493 -4714
rect -481 -4718 -480 -4714
rect -478 -4718 -472 -4714
rect -470 -4718 -468 -4714
rect -464 -4718 -462 -4714
rect -460 -4718 -454 -4714
rect -452 -4718 -451 -4714
rect -439 -4718 -438 -4714
rect -436 -4718 -430 -4714
rect -428 -4718 -426 -4714
rect -422 -4718 -420 -4714
rect -418 -4718 -412 -4714
rect -410 -4718 -409 -4714
rect -397 -4718 -396 -4714
rect -394 -4718 -388 -4714
rect -386 -4718 -385 -4714
rect -215 -4718 -214 -4714
rect -212 -4718 -210 -4714
rect -206 -4718 -204 -4714
rect -202 -4718 -201 -4714
rect -189 -4718 -188 -4714
rect -186 -4718 -180 -4714
rect -178 -4718 -177 -4714
rect -165 -4718 -164 -4714
rect -162 -4718 -156 -4714
rect -154 -4718 -152 -4714
rect -148 -4718 -146 -4714
rect -144 -4718 -138 -4714
rect -136 -4718 -135 -4714
rect -123 -4718 -122 -4714
rect -120 -4718 -114 -4714
rect -112 -4718 -110 -4714
rect -106 -4718 -104 -4714
rect -102 -4718 -96 -4714
rect -94 -4718 -93 -4714
rect -81 -4718 -80 -4714
rect -78 -4718 -72 -4714
rect -70 -4718 -68 -4714
rect -64 -4718 -62 -4714
rect -60 -4718 -54 -4714
rect -52 -4718 -51 -4714
rect -39 -4718 -38 -4714
rect -36 -4718 -30 -4714
rect -28 -4718 -27 -4714
rect 213 -4718 214 -4714
rect 216 -4718 218 -4714
rect 222 -4718 224 -4714
rect 226 -4718 227 -4714
rect 239 -4718 240 -4714
rect 242 -4718 248 -4714
rect 250 -4718 251 -4714
rect 263 -4718 264 -4714
rect 266 -4718 272 -4714
rect 274 -4718 276 -4714
rect 280 -4718 282 -4714
rect 284 -4718 290 -4714
rect 292 -4718 293 -4714
rect 305 -4718 306 -4714
rect 308 -4718 314 -4714
rect 316 -4718 318 -4714
rect 322 -4718 324 -4714
rect 326 -4718 332 -4714
rect 334 -4718 335 -4714
rect 347 -4718 348 -4714
rect 350 -4718 356 -4714
rect 358 -4718 360 -4714
rect 364 -4718 366 -4714
rect 368 -4718 374 -4714
rect 376 -4718 377 -4714
rect 389 -4718 390 -4714
rect 392 -4718 398 -4714
rect 400 -4718 401 -4714
rect 569 -4718 570 -4714
rect 572 -4718 574 -4714
rect 578 -4718 580 -4714
rect 582 -4718 583 -4714
rect 595 -4718 596 -4714
rect 598 -4718 604 -4714
rect 606 -4718 607 -4714
rect 619 -4718 620 -4714
rect 622 -4718 628 -4714
rect 630 -4718 632 -4714
rect 636 -4718 638 -4714
rect 640 -4718 646 -4714
rect 648 -4718 649 -4714
rect 661 -4718 662 -4714
rect 664 -4718 670 -4714
rect 672 -4718 674 -4714
rect 678 -4718 680 -4714
rect 682 -4718 688 -4714
rect 690 -4718 691 -4714
rect 703 -4718 704 -4714
rect 706 -4718 712 -4714
rect 714 -4718 716 -4714
rect 720 -4718 722 -4714
rect 724 -4718 730 -4714
rect 732 -4718 733 -4714
rect 745 -4718 746 -4714
rect 748 -4718 754 -4714
rect 756 -4718 757 -4714
rect 967 -4718 968 -4714
rect 970 -4718 972 -4714
rect 976 -4718 978 -4714
rect 980 -4718 981 -4714
rect 993 -4718 994 -4714
rect 996 -4718 1002 -4714
rect 1004 -4718 1005 -4714
rect 1017 -4718 1018 -4714
rect 1020 -4718 1026 -4714
rect 1028 -4718 1030 -4714
rect 1034 -4718 1036 -4714
rect 1038 -4718 1044 -4714
rect 1046 -4718 1047 -4714
rect 1059 -4718 1060 -4714
rect 1062 -4718 1068 -4714
rect 1070 -4718 1072 -4714
rect 1076 -4718 1078 -4714
rect 1080 -4718 1086 -4714
rect 1088 -4718 1089 -4714
rect 1101 -4718 1102 -4714
rect 1104 -4718 1110 -4714
rect 1112 -4718 1114 -4714
rect 1118 -4718 1120 -4714
rect 1122 -4718 1128 -4714
rect 1130 -4718 1131 -4714
rect 1143 -4718 1144 -4714
rect 1146 -4718 1152 -4714
rect 1154 -4718 1155 -4714
rect 1325 -4718 1326 -4714
rect 1328 -4718 1330 -4714
rect 1334 -4718 1336 -4714
rect 1338 -4718 1339 -4714
rect 1351 -4718 1352 -4714
rect 1354 -4718 1360 -4714
rect 1362 -4718 1363 -4714
rect 1375 -4718 1376 -4714
rect 1378 -4718 1384 -4714
rect 1386 -4718 1388 -4714
rect 1392 -4718 1394 -4714
rect 1396 -4718 1402 -4714
rect 1404 -4718 1405 -4714
rect 1417 -4718 1418 -4714
rect 1420 -4718 1426 -4714
rect 1428 -4718 1430 -4714
rect 1434 -4718 1436 -4714
rect 1438 -4718 1444 -4714
rect 1446 -4718 1447 -4714
rect 1459 -4718 1460 -4714
rect 1462 -4718 1468 -4714
rect 1470 -4718 1472 -4714
rect 1476 -4718 1478 -4714
rect 1480 -4718 1486 -4714
rect 1488 -4718 1489 -4714
rect 1501 -4718 1502 -4714
rect 1504 -4718 1510 -4714
rect 1512 -4718 1513 -4714
rect -1260 -4839 -1259 -4835
rect -1257 -4839 -1255 -4835
rect -1251 -4839 -1249 -4835
rect -1247 -4839 -1246 -4835
rect -1234 -4839 -1233 -4835
rect -1231 -4839 -1225 -4835
rect -1223 -4839 -1222 -4835
rect -1210 -4839 -1209 -4835
rect -1207 -4839 -1201 -4835
rect -1199 -4839 -1197 -4835
rect -1193 -4839 -1191 -4835
rect -1189 -4839 -1183 -4835
rect -1181 -4839 -1180 -4835
rect -1168 -4839 -1167 -4835
rect -1165 -4839 -1159 -4835
rect -1157 -4839 -1155 -4835
rect -1151 -4839 -1149 -4835
rect -1147 -4839 -1141 -4835
rect -1139 -4839 -1138 -4835
rect -1126 -4839 -1125 -4835
rect -1123 -4839 -1117 -4835
rect -1115 -4839 -1113 -4835
rect -1109 -4839 -1107 -4835
rect -1105 -4839 -1099 -4835
rect -1097 -4839 -1096 -4835
rect -1084 -4839 -1083 -4835
rect -1081 -4839 -1075 -4835
rect -1073 -4839 -1072 -4835
rect -931 -4839 -930 -4835
rect -928 -4839 -926 -4835
rect -922 -4839 -920 -4835
rect -918 -4839 -917 -4835
rect -905 -4839 -904 -4835
rect -902 -4839 -896 -4835
rect -894 -4839 -893 -4835
rect -881 -4839 -880 -4835
rect -878 -4839 -872 -4835
rect -870 -4839 -868 -4835
rect -864 -4839 -862 -4835
rect -860 -4839 -854 -4835
rect -852 -4839 -851 -4835
rect -839 -4839 -838 -4835
rect -836 -4839 -830 -4835
rect -828 -4839 -826 -4835
rect -822 -4839 -820 -4835
rect -818 -4839 -812 -4835
rect -810 -4839 -809 -4835
rect -797 -4839 -796 -4835
rect -794 -4839 -788 -4835
rect -786 -4839 -784 -4835
rect -780 -4839 -778 -4835
rect -776 -4839 -770 -4835
rect -768 -4839 -767 -4835
rect -755 -4839 -754 -4835
rect -752 -4839 -746 -4835
rect -744 -4839 -743 -4835
rect -573 -4839 -572 -4835
rect -570 -4839 -568 -4835
rect -564 -4839 -562 -4835
rect -560 -4839 -559 -4835
rect -547 -4839 -546 -4835
rect -544 -4839 -538 -4835
rect -536 -4839 -535 -4835
rect -523 -4839 -522 -4835
rect -520 -4839 -514 -4835
rect -512 -4839 -510 -4835
rect -506 -4839 -504 -4835
rect -502 -4839 -496 -4835
rect -494 -4839 -493 -4835
rect -481 -4839 -480 -4835
rect -478 -4839 -472 -4835
rect -470 -4839 -468 -4835
rect -464 -4839 -462 -4835
rect -460 -4839 -454 -4835
rect -452 -4839 -451 -4835
rect -439 -4839 -438 -4835
rect -436 -4839 -430 -4835
rect -428 -4839 -426 -4835
rect -422 -4839 -420 -4835
rect -418 -4839 -412 -4835
rect -410 -4839 -409 -4835
rect -397 -4839 -396 -4835
rect -394 -4839 -388 -4835
rect -386 -4839 -385 -4835
rect -215 -4839 -214 -4835
rect -212 -4839 -210 -4835
rect -206 -4839 -204 -4835
rect -202 -4839 -201 -4835
rect -189 -4839 -188 -4835
rect -186 -4839 -180 -4835
rect -178 -4839 -177 -4835
rect -165 -4839 -164 -4835
rect -162 -4839 -156 -4835
rect -154 -4839 -152 -4835
rect -148 -4839 -146 -4835
rect -144 -4839 -138 -4835
rect -136 -4839 -135 -4835
rect -123 -4839 -122 -4835
rect -120 -4839 -114 -4835
rect -112 -4839 -110 -4835
rect -106 -4839 -104 -4835
rect -102 -4839 -96 -4835
rect -94 -4839 -93 -4835
rect -81 -4839 -80 -4835
rect -78 -4839 -72 -4835
rect -70 -4839 -68 -4835
rect -64 -4839 -62 -4835
rect -60 -4839 -54 -4835
rect -52 -4839 -51 -4835
rect -39 -4839 -38 -4835
rect -36 -4839 -30 -4835
rect -28 -4839 -27 -4835
rect 94 -4839 95 -4823
rect 97 -4839 98 -4823
rect 213 -4839 214 -4835
rect 216 -4839 218 -4835
rect 222 -4839 224 -4835
rect 226 -4839 227 -4835
rect 239 -4839 240 -4835
rect 242 -4839 248 -4835
rect 250 -4839 251 -4835
rect 263 -4839 264 -4835
rect 266 -4839 272 -4835
rect 274 -4839 276 -4835
rect 280 -4839 282 -4835
rect 284 -4839 290 -4835
rect 292 -4839 293 -4835
rect 305 -4839 306 -4835
rect 308 -4839 314 -4835
rect 316 -4839 318 -4835
rect 322 -4839 324 -4835
rect 326 -4839 332 -4835
rect 334 -4839 335 -4835
rect 347 -4839 348 -4835
rect 350 -4839 356 -4835
rect 358 -4839 360 -4835
rect 364 -4839 366 -4835
rect 368 -4839 374 -4835
rect 376 -4839 377 -4835
rect 389 -4839 390 -4835
rect 392 -4839 398 -4835
rect 400 -4839 401 -4835
rect 569 -4839 570 -4835
rect 572 -4839 574 -4835
rect 578 -4839 580 -4835
rect 582 -4839 583 -4835
rect 595 -4839 596 -4835
rect 598 -4839 604 -4835
rect 606 -4839 607 -4835
rect 619 -4839 620 -4835
rect 622 -4839 628 -4835
rect 630 -4839 632 -4835
rect 636 -4839 638 -4835
rect 640 -4839 646 -4835
rect 648 -4839 649 -4835
rect 661 -4839 662 -4835
rect 664 -4839 670 -4835
rect 672 -4839 674 -4835
rect 678 -4839 680 -4835
rect 682 -4839 688 -4835
rect 690 -4839 691 -4835
rect 703 -4839 704 -4835
rect 706 -4839 712 -4835
rect 714 -4839 716 -4835
rect 720 -4839 722 -4835
rect 724 -4839 730 -4835
rect 732 -4839 733 -4835
rect 745 -4839 746 -4835
rect 748 -4839 754 -4835
rect 756 -4839 757 -4835
rect 967 -4839 968 -4835
rect 970 -4839 972 -4835
rect 976 -4839 978 -4835
rect 980 -4839 981 -4835
rect 993 -4839 994 -4835
rect 996 -4839 1002 -4835
rect 1004 -4839 1005 -4835
rect 1017 -4839 1018 -4835
rect 1020 -4839 1026 -4835
rect 1028 -4839 1030 -4835
rect 1034 -4839 1036 -4835
rect 1038 -4839 1044 -4835
rect 1046 -4839 1047 -4835
rect 1059 -4839 1060 -4835
rect 1062 -4839 1068 -4835
rect 1070 -4839 1072 -4835
rect 1076 -4839 1078 -4835
rect 1080 -4839 1086 -4835
rect 1088 -4839 1089 -4835
rect 1101 -4839 1102 -4835
rect 1104 -4839 1110 -4835
rect 1112 -4839 1114 -4835
rect 1118 -4839 1120 -4835
rect 1122 -4839 1128 -4835
rect 1130 -4839 1131 -4835
rect 1143 -4839 1144 -4835
rect 1146 -4839 1152 -4835
rect 1154 -4839 1155 -4835
rect 1325 -4839 1326 -4835
rect 1328 -4839 1330 -4835
rect 1334 -4839 1336 -4835
rect 1338 -4839 1339 -4835
rect 1351 -4839 1352 -4835
rect 1354 -4839 1360 -4835
rect 1362 -4839 1363 -4835
rect 1375 -4839 1376 -4835
rect 1378 -4839 1384 -4835
rect 1386 -4839 1388 -4835
rect 1392 -4839 1394 -4835
rect 1396 -4839 1402 -4835
rect 1404 -4839 1405 -4835
rect 1417 -4839 1418 -4835
rect 1420 -4839 1426 -4835
rect 1428 -4839 1430 -4835
rect 1434 -4839 1436 -4835
rect 1438 -4839 1444 -4835
rect 1446 -4839 1447 -4835
rect 1459 -4839 1460 -4835
rect 1462 -4839 1468 -4835
rect 1470 -4839 1472 -4835
rect 1476 -4839 1478 -4835
rect 1480 -4839 1486 -4835
rect 1488 -4839 1489 -4835
rect 1501 -4839 1502 -4835
rect 1504 -4839 1510 -4835
rect 1512 -4839 1513 -4835
rect -1260 -4957 -1259 -4953
rect -1257 -4957 -1255 -4953
rect -1251 -4957 -1249 -4953
rect -1247 -4957 -1246 -4953
rect -1234 -4957 -1233 -4953
rect -1231 -4957 -1225 -4953
rect -1223 -4957 -1222 -4953
rect -1210 -4957 -1209 -4953
rect -1207 -4957 -1201 -4953
rect -1199 -4957 -1197 -4953
rect -1193 -4957 -1191 -4953
rect -1189 -4957 -1183 -4953
rect -1181 -4957 -1180 -4953
rect -1168 -4957 -1167 -4953
rect -1165 -4957 -1159 -4953
rect -1157 -4957 -1155 -4953
rect -1151 -4957 -1149 -4953
rect -1147 -4957 -1141 -4953
rect -1139 -4957 -1138 -4953
rect -1126 -4957 -1125 -4953
rect -1123 -4957 -1117 -4953
rect -1115 -4957 -1113 -4953
rect -1109 -4957 -1107 -4953
rect -1105 -4957 -1099 -4953
rect -1097 -4957 -1096 -4953
rect -1084 -4957 -1083 -4953
rect -1081 -4957 -1075 -4953
rect -1073 -4957 -1072 -4953
rect -931 -4957 -930 -4953
rect -928 -4957 -926 -4953
rect -922 -4957 -920 -4953
rect -918 -4957 -917 -4953
rect -905 -4957 -904 -4953
rect -902 -4957 -896 -4953
rect -894 -4957 -893 -4953
rect -881 -4957 -880 -4953
rect -878 -4957 -872 -4953
rect -870 -4957 -868 -4953
rect -864 -4957 -862 -4953
rect -860 -4957 -854 -4953
rect -852 -4957 -851 -4953
rect -839 -4957 -838 -4953
rect -836 -4957 -830 -4953
rect -828 -4957 -826 -4953
rect -822 -4957 -820 -4953
rect -818 -4957 -812 -4953
rect -810 -4957 -809 -4953
rect -797 -4957 -796 -4953
rect -794 -4957 -788 -4953
rect -786 -4957 -784 -4953
rect -780 -4957 -778 -4953
rect -776 -4957 -770 -4953
rect -768 -4957 -767 -4953
rect -755 -4957 -754 -4953
rect -752 -4957 -746 -4953
rect -744 -4957 -743 -4953
rect -573 -4957 -572 -4953
rect -570 -4957 -568 -4953
rect -564 -4957 -562 -4953
rect -560 -4957 -559 -4953
rect -547 -4957 -546 -4953
rect -544 -4957 -538 -4953
rect -536 -4957 -535 -4953
rect -523 -4957 -522 -4953
rect -520 -4957 -514 -4953
rect -512 -4957 -510 -4953
rect -506 -4957 -504 -4953
rect -502 -4957 -496 -4953
rect -494 -4957 -493 -4953
rect -481 -4957 -480 -4953
rect -478 -4957 -472 -4953
rect -470 -4957 -468 -4953
rect -464 -4957 -462 -4953
rect -460 -4957 -454 -4953
rect -452 -4957 -451 -4953
rect -439 -4957 -438 -4953
rect -436 -4957 -430 -4953
rect -428 -4957 -426 -4953
rect -422 -4957 -420 -4953
rect -418 -4957 -412 -4953
rect -410 -4957 -409 -4953
rect -397 -4957 -396 -4953
rect -394 -4957 -388 -4953
rect -386 -4957 -385 -4953
rect -215 -4957 -214 -4953
rect -212 -4957 -210 -4953
rect -206 -4957 -204 -4953
rect -202 -4957 -201 -4953
rect -189 -4957 -188 -4953
rect -186 -4957 -180 -4953
rect -178 -4957 -177 -4953
rect -165 -4957 -164 -4953
rect -162 -4957 -156 -4953
rect -154 -4957 -152 -4953
rect -148 -4957 -146 -4953
rect -144 -4957 -138 -4953
rect -136 -4957 -135 -4953
rect -123 -4957 -122 -4953
rect -120 -4957 -114 -4953
rect -112 -4957 -110 -4953
rect -106 -4957 -104 -4953
rect -102 -4957 -96 -4953
rect -94 -4957 -93 -4953
rect -81 -4957 -80 -4953
rect -78 -4957 -72 -4953
rect -70 -4957 -68 -4953
rect -64 -4957 -62 -4953
rect -60 -4957 -54 -4953
rect -52 -4957 -51 -4953
rect -39 -4957 -38 -4953
rect -36 -4957 -30 -4953
rect -28 -4957 -27 -4953
rect 213 -4957 214 -4953
rect 216 -4957 218 -4953
rect 222 -4957 224 -4953
rect 226 -4957 227 -4953
rect 239 -4957 240 -4953
rect 242 -4957 248 -4953
rect 250 -4957 251 -4953
rect 263 -4957 264 -4953
rect 266 -4957 272 -4953
rect 274 -4957 276 -4953
rect 280 -4957 282 -4953
rect 284 -4957 290 -4953
rect 292 -4957 293 -4953
rect 305 -4957 306 -4953
rect 308 -4957 314 -4953
rect 316 -4957 318 -4953
rect 322 -4957 324 -4953
rect 326 -4957 332 -4953
rect 334 -4957 335 -4953
rect 347 -4957 348 -4953
rect 350 -4957 356 -4953
rect 358 -4957 360 -4953
rect 364 -4957 366 -4953
rect 368 -4957 374 -4953
rect 376 -4957 377 -4953
rect 389 -4957 390 -4953
rect 392 -4957 398 -4953
rect 400 -4957 401 -4953
rect -1335 -5074 -1334 -5070
rect -1332 -5074 -1326 -5070
rect -1324 -5074 -1322 -5070
rect -1318 -5074 -1316 -5070
rect -1314 -5074 -1313 -5070
rect -931 -5074 -930 -5070
rect -928 -5074 -922 -5070
rect -920 -5074 -918 -5070
rect -914 -5074 -912 -5070
rect -910 -5074 -909 -5070
rect -573 -5074 -572 -5070
rect -570 -5074 -564 -5070
rect -562 -5074 -560 -5070
rect -556 -5074 -554 -5070
rect -552 -5074 -551 -5070
rect -215 -5074 -214 -5070
rect -212 -5074 -206 -5070
rect -204 -5074 -202 -5070
rect -198 -5074 -196 -5070
rect -194 -5074 -193 -5070
rect 213 -5074 214 -5070
rect 216 -5074 222 -5070
rect 224 -5074 226 -5070
rect 230 -5074 232 -5070
rect 234 -5074 235 -5070
rect 569 -5074 570 -5070
rect 572 -5074 578 -5070
rect 580 -5074 582 -5070
rect 586 -5074 588 -5070
rect 590 -5074 591 -5070
rect 967 -5074 968 -5070
rect 970 -5074 976 -5070
rect 978 -5074 980 -5070
rect 984 -5074 986 -5070
rect 988 -5074 989 -5070
rect 1325 -5074 1326 -5070
rect 1328 -5074 1334 -5070
rect 1336 -5074 1338 -5070
rect 1342 -5074 1344 -5070
rect 1346 -5074 1347 -5070
rect -1260 -5193 -1259 -5189
rect -1257 -5193 -1255 -5189
rect -1251 -5193 -1249 -5189
rect -1247 -5193 -1246 -5189
rect -1234 -5193 -1233 -5189
rect -1231 -5193 -1229 -5189
rect -1225 -5193 -1223 -5189
rect -1221 -5193 -1215 -5189
rect -1213 -5193 -1211 -5189
rect -1207 -5193 -1205 -5189
rect -1203 -5193 -1202 -5189
rect -1190 -5193 -1189 -5189
rect -1187 -5193 -1181 -5189
rect -1179 -5193 -1177 -5189
rect -1173 -5193 -1171 -5189
rect -1169 -5193 -1168 -5189
rect -931 -5193 -930 -5189
rect -928 -5193 -926 -5189
rect -922 -5193 -920 -5189
rect -918 -5193 -917 -5189
rect -905 -5193 -904 -5189
rect -902 -5193 -900 -5189
rect -896 -5193 -894 -5189
rect -892 -5193 -891 -5189
rect -879 -5193 -878 -5189
rect -876 -5193 -875 -5189
rect -871 -5193 -868 -5189
rect -866 -5193 -860 -5189
rect -858 -5193 -857 -5189
rect -853 -5193 -850 -5189
rect -848 -5193 -847 -5189
rect -835 -5193 -834 -5189
rect -832 -5193 -826 -5189
rect -824 -5193 -822 -5189
rect -818 -5193 -816 -5189
rect -814 -5193 -813 -5189
rect -801 -5193 -800 -5189
rect -798 -5193 -796 -5189
rect -792 -5193 -790 -5189
rect -788 -5193 -782 -5189
rect -780 -5193 -778 -5189
rect -774 -5193 -772 -5189
rect -770 -5193 -769 -5189
rect -757 -5193 -756 -5189
rect -754 -5193 -748 -5189
rect -746 -5193 -745 -5189
rect -733 -5193 -732 -5189
rect -730 -5193 -725 -5189
rect -721 -5193 -716 -5189
rect -714 -5193 -713 -5189
rect -709 -5193 -708 -5189
rect -706 -5193 -704 -5189
rect -700 -5193 -698 -5189
rect -696 -5193 -695 -5189
rect -573 -5193 -572 -5189
rect -570 -5193 -568 -5189
rect -564 -5193 -562 -5189
rect -560 -5193 -559 -5189
rect -547 -5193 -546 -5189
rect -544 -5193 -542 -5189
rect -538 -5193 -536 -5189
rect -534 -5193 -533 -5189
rect -521 -5193 -520 -5189
rect -518 -5193 -517 -5189
rect -513 -5193 -510 -5189
rect -508 -5193 -502 -5189
rect -500 -5193 -499 -5189
rect -495 -5193 -492 -5189
rect -490 -5193 -489 -5189
rect -477 -5193 -476 -5189
rect -474 -5193 -468 -5189
rect -466 -5193 -464 -5189
rect -460 -5193 -458 -5189
rect -456 -5193 -455 -5189
rect -443 -5193 -442 -5189
rect -440 -5193 -438 -5189
rect -434 -5193 -432 -5189
rect -430 -5193 -424 -5189
rect -422 -5193 -420 -5189
rect -416 -5193 -414 -5189
rect -412 -5193 -411 -5189
rect -399 -5193 -398 -5189
rect -396 -5193 -390 -5189
rect -388 -5193 -387 -5189
rect -375 -5193 -374 -5189
rect -372 -5193 -367 -5189
rect -363 -5193 -358 -5189
rect -356 -5193 -355 -5189
rect -351 -5193 -350 -5189
rect -348 -5193 -346 -5189
rect -342 -5193 -340 -5189
rect -338 -5193 -337 -5189
rect -215 -5193 -214 -5189
rect -212 -5193 -210 -5189
rect -206 -5193 -204 -5189
rect -202 -5193 -201 -5189
rect -189 -5193 -188 -5189
rect -186 -5193 -184 -5189
rect -180 -5193 -178 -5189
rect -176 -5193 -175 -5189
rect -163 -5193 -162 -5189
rect -160 -5193 -159 -5189
rect -155 -5193 -152 -5189
rect -150 -5193 -144 -5189
rect -142 -5193 -141 -5189
rect -137 -5193 -134 -5189
rect -132 -5193 -131 -5189
rect -119 -5193 -118 -5189
rect -116 -5193 -110 -5189
rect -108 -5193 -106 -5189
rect -102 -5193 -100 -5189
rect -98 -5193 -97 -5189
rect -85 -5193 -84 -5189
rect -82 -5193 -80 -5189
rect -76 -5193 -74 -5189
rect -72 -5193 -66 -5189
rect -64 -5193 -62 -5189
rect -58 -5193 -56 -5189
rect -54 -5193 -53 -5189
rect -41 -5193 -40 -5189
rect -38 -5193 -32 -5189
rect -30 -5193 -29 -5189
rect -17 -5193 -16 -5189
rect -14 -5193 -9 -5189
rect -5 -5193 0 -5189
rect 2 -5193 3 -5189
rect 7 -5193 8 -5189
rect 10 -5193 12 -5189
rect 16 -5193 18 -5189
rect 20 -5193 21 -5189
rect 213 -5193 214 -5189
rect 216 -5193 218 -5189
rect 222 -5193 224 -5189
rect 226 -5193 227 -5189
rect 239 -5193 240 -5189
rect 242 -5193 244 -5189
rect 248 -5193 250 -5189
rect 252 -5193 253 -5189
rect 265 -5193 266 -5189
rect 268 -5193 269 -5189
rect 273 -5193 276 -5189
rect 278 -5193 284 -5189
rect 286 -5193 287 -5189
rect 291 -5193 294 -5189
rect 296 -5193 297 -5189
rect 309 -5193 310 -5189
rect 312 -5193 318 -5189
rect 320 -5193 322 -5189
rect 326 -5193 328 -5189
rect 330 -5193 331 -5189
rect 343 -5193 344 -5189
rect 346 -5193 348 -5189
rect 352 -5193 354 -5189
rect 356 -5193 362 -5189
rect 364 -5193 366 -5189
rect 370 -5193 372 -5189
rect 374 -5193 375 -5189
rect 387 -5193 388 -5189
rect 390 -5193 396 -5189
rect 398 -5193 399 -5189
rect 411 -5193 412 -5189
rect 414 -5193 419 -5189
rect 423 -5193 428 -5189
rect 430 -5193 431 -5189
rect 435 -5193 436 -5189
rect 438 -5193 440 -5189
rect 444 -5193 446 -5189
rect 448 -5193 449 -5189
rect 569 -5193 570 -5189
rect 572 -5193 574 -5189
rect 578 -5193 580 -5189
rect 582 -5193 583 -5189
rect 595 -5193 596 -5189
rect 598 -5193 600 -5189
rect 604 -5193 606 -5189
rect 608 -5193 609 -5189
rect 621 -5193 622 -5189
rect 624 -5193 625 -5189
rect 629 -5193 632 -5189
rect 634 -5193 640 -5189
rect 642 -5193 643 -5189
rect 647 -5193 650 -5189
rect 652 -5193 653 -5189
rect 665 -5193 666 -5189
rect 668 -5193 674 -5189
rect 676 -5193 678 -5189
rect 682 -5193 684 -5189
rect 686 -5193 687 -5189
rect 699 -5193 700 -5189
rect 702 -5193 704 -5189
rect 708 -5193 710 -5189
rect 712 -5193 718 -5189
rect 720 -5193 722 -5189
rect 726 -5193 728 -5189
rect 730 -5193 731 -5189
rect 743 -5193 744 -5189
rect 746 -5193 752 -5189
rect 754 -5193 755 -5189
rect 767 -5193 768 -5189
rect 770 -5193 775 -5189
rect 779 -5193 784 -5189
rect 786 -5193 787 -5189
rect 791 -5193 792 -5189
rect 794 -5193 796 -5189
rect 800 -5193 802 -5189
rect 804 -5193 805 -5189
rect 967 -5193 968 -5189
rect 970 -5193 972 -5189
rect 976 -5193 978 -5189
rect 980 -5193 981 -5189
rect 993 -5193 994 -5189
rect 996 -5193 998 -5189
rect 1002 -5193 1004 -5189
rect 1006 -5193 1007 -5189
rect 1019 -5193 1020 -5189
rect 1022 -5193 1023 -5189
rect 1027 -5193 1030 -5189
rect 1032 -5193 1038 -5189
rect 1040 -5193 1041 -5189
rect 1045 -5193 1048 -5189
rect 1050 -5193 1051 -5189
rect 1063 -5193 1064 -5189
rect 1066 -5193 1072 -5189
rect 1074 -5193 1076 -5189
rect 1080 -5193 1082 -5189
rect 1084 -5193 1085 -5189
rect 1097 -5193 1098 -5189
rect 1100 -5193 1102 -5189
rect 1106 -5193 1108 -5189
rect 1110 -5193 1116 -5189
rect 1118 -5193 1120 -5189
rect 1124 -5193 1126 -5189
rect 1128 -5193 1129 -5189
rect 1141 -5193 1142 -5189
rect 1144 -5193 1150 -5189
rect 1152 -5193 1153 -5189
rect 1165 -5193 1166 -5189
rect 1168 -5193 1173 -5189
rect 1177 -5193 1182 -5189
rect 1184 -5193 1185 -5189
rect 1189 -5193 1190 -5189
rect 1192 -5193 1194 -5189
rect 1198 -5193 1200 -5189
rect 1202 -5193 1203 -5189
rect 1325 -5193 1326 -5189
rect 1328 -5193 1330 -5189
rect 1334 -5193 1336 -5189
rect 1338 -5193 1339 -5189
rect 1351 -5193 1352 -5189
rect 1354 -5193 1356 -5189
rect 1360 -5193 1362 -5189
rect 1364 -5193 1365 -5189
rect 1377 -5193 1378 -5189
rect 1380 -5193 1381 -5189
rect 1385 -5193 1388 -5189
rect 1390 -5193 1396 -5189
rect 1398 -5193 1399 -5189
rect 1403 -5193 1406 -5189
rect 1408 -5193 1409 -5189
rect 1421 -5193 1422 -5189
rect 1424 -5193 1430 -5189
rect 1432 -5193 1434 -5189
rect 1438 -5193 1440 -5189
rect 1442 -5193 1443 -5189
rect 1455 -5193 1456 -5189
rect 1458 -5193 1460 -5189
rect 1464 -5193 1466 -5189
rect 1468 -5193 1474 -5189
rect 1476 -5193 1478 -5189
rect 1482 -5193 1484 -5189
rect 1486 -5193 1487 -5189
rect 1499 -5193 1500 -5189
rect 1502 -5193 1508 -5189
rect 1510 -5193 1511 -5189
rect 1523 -5193 1524 -5189
rect 1526 -5193 1531 -5189
rect 1535 -5193 1540 -5189
rect 1542 -5193 1543 -5189
rect 1547 -5193 1548 -5189
rect 1550 -5193 1552 -5189
rect 1556 -5193 1558 -5189
rect 1560 -5193 1561 -5189
rect -1260 -5312 -1259 -5308
rect -1257 -5312 -1255 -5308
rect -1251 -5312 -1249 -5308
rect -1247 -5312 -1246 -5308
rect -1234 -5312 -1233 -5308
rect -1231 -5312 -1225 -5308
rect -1223 -5312 -1222 -5308
rect -1210 -5312 -1209 -5308
rect -1207 -5312 -1201 -5308
rect -1199 -5312 -1197 -5308
rect -1193 -5312 -1191 -5308
rect -1189 -5312 -1183 -5308
rect -1181 -5312 -1180 -5308
rect -1168 -5312 -1167 -5308
rect -1165 -5312 -1159 -5308
rect -1157 -5312 -1155 -5308
rect -1151 -5312 -1149 -5308
rect -1147 -5312 -1141 -5308
rect -1139 -5312 -1138 -5308
rect -1126 -5312 -1125 -5308
rect -1123 -5312 -1117 -5308
rect -1115 -5312 -1113 -5308
rect -1109 -5312 -1107 -5308
rect -1105 -5312 -1099 -5308
rect -1097 -5312 -1096 -5308
rect -1084 -5312 -1083 -5308
rect -1081 -5312 -1075 -5308
rect -1073 -5312 -1072 -5308
rect -931 -5312 -930 -5308
rect -928 -5312 -926 -5308
rect -922 -5312 -920 -5308
rect -918 -5312 -917 -5308
rect -905 -5312 -904 -5308
rect -902 -5312 -896 -5308
rect -894 -5312 -893 -5308
rect -881 -5312 -880 -5308
rect -878 -5312 -872 -5308
rect -870 -5312 -868 -5308
rect -864 -5312 -862 -5308
rect -860 -5312 -854 -5308
rect -852 -5312 -851 -5308
rect -839 -5312 -838 -5308
rect -836 -5312 -830 -5308
rect -828 -5312 -826 -5308
rect -822 -5312 -820 -5308
rect -818 -5312 -812 -5308
rect -810 -5312 -809 -5308
rect -797 -5312 -796 -5308
rect -794 -5312 -788 -5308
rect -786 -5312 -784 -5308
rect -780 -5312 -778 -5308
rect -776 -5312 -770 -5308
rect -768 -5312 -767 -5308
rect -755 -5312 -754 -5308
rect -752 -5312 -746 -5308
rect -744 -5312 -743 -5308
rect -1260 -5433 -1259 -5429
rect -1257 -5433 -1255 -5429
rect -1251 -5433 -1249 -5429
rect -1247 -5433 -1246 -5429
rect -1234 -5433 -1233 -5429
rect -1231 -5433 -1225 -5429
rect -1223 -5433 -1222 -5429
rect -1210 -5433 -1209 -5429
rect -1207 -5433 -1201 -5429
rect -1199 -5433 -1197 -5429
rect -1193 -5433 -1191 -5429
rect -1189 -5433 -1183 -5429
rect -1181 -5433 -1180 -5429
rect -1168 -5433 -1167 -5429
rect -1165 -5433 -1159 -5429
rect -1157 -5433 -1155 -5429
rect -1151 -5433 -1149 -5429
rect -1147 -5433 -1141 -5429
rect -1139 -5433 -1138 -5429
rect -1126 -5433 -1125 -5429
rect -1123 -5433 -1117 -5429
rect -1115 -5433 -1113 -5429
rect -1109 -5433 -1107 -5429
rect -1105 -5433 -1099 -5429
rect -1097 -5433 -1096 -5429
rect -1084 -5433 -1083 -5429
rect -1081 -5433 -1075 -5429
rect -1073 -5433 -1072 -5429
rect -1022 -5433 -1021 -5429
rect -1019 -5433 -1018 -5429
rect -931 -5433 -930 -5429
rect -928 -5433 -926 -5429
rect -922 -5433 -920 -5429
rect -918 -5433 -917 -5429
rect -905 -5433 -904 -5429
rect -902 -5433 -896 -5429
rect -894 -5433 -893 -5429
rect -881 -5433 -880 -5429
rect -878 -5433 -872 -5429
rect -870 -5433 -868 -5429
rect -864 -5433 -862 -5429
rect -860 -5433 -854 -5429
rect -852 -5433 -851 -5429
rect -839 -5433 -838 -5429
rect -836 -5433 -830 -5429
rect -828 -5433 -826 -5429
rect -822 -5433 -820 -5429
rect -818 -5433 -812 -5429
rect -810 -5433 -809 -5429
rect -797 -5433 -796 -5429
rect -794 -5433 -788 -5429
rect -786 -5433 -784 -5429
rect -780 -5433 -778 -5429
rect -776 -5433 -770 -5429
rect -768 -5433 -767 -5429
rect -755 -5433 -754 -5429
rect -752 -5433 -746 -5429
rect -744 -5433 -743 -5429
rect -669 -5433 -668 -5425
rect -666 -5433 -665 -5425
rect -573 -5433 -572 -5429
rect -570 -5433 -568 -5429
rect -564 -5433 -562 -5429
rect -560 -5433 -559 -5429
rect -547 -5433 -546 -5429
rect -544 -5433 -538 -5429
rect -536 -5433 -535 -5429
rect -523 -5433 -522 -5429
rect -520 -5433 -514 -5429
rect -512 -5433 -510 -5429
rect -506 -5433 -504 -5429
rect -502 -5433 -496 -5429
rect -494 -5433 -493 -5429
rect -481 -5433 -480 -5429
rect -478 -5433 -472 -5429
rect -470 -5433 -468 -5429
rect -464 -5433 -462 -5429
rect -460 -5433 -454 -5429
rect -452 -5433 -451 -5429
rect -439 -5433 -438 -5429
rect -436 -5433 -430 -5429
rect -428 -5433 -426 -5429
rect -422 -5433 -420 -5429
rect -418 -5433 -412 -5429
rect -410 -5433 -409 -5429
rect -397 -5433 -396 -5429
rect -394 -5433 -388 -5429
rect -386 -5433 -385 -5429
rect -323 -5433 -322 -5429
rect -320 -5433 -319 -5429
rect -215 -5433 -214 -5429
rect -212 -5433 -210 -5429
rect -206 -5433 -204 -5429
rect -202 -5433 -201 -5429
rect -189 -5433 -188 -5429
rect -186 -5433 -180 -5429
rect -178 -5433 -177 -5429
rect -165 -5433 -164 -5429
rect -162 -5433 -156 -5429
rect -154 -5433 -152 -5429
rect -148 -5433 -146 -5429
rect -144 -5433 -138 -5429
rect -136 -5433 -135 -5429
rect -123 -5433 -122 -5429
rect -120 -5433 -114 -5429
rect -112 -5433 -110 -5429
rect -106 -5433 -104 -5429
rect -102 -5433 -96 -5429
rect -94 -5433 -93 -5429
rect -81 -5433 -80 -5429
rect -78 -5433 -72 -5429
rect -70 -5433 -68 -5429
rect -64 -5433 -62 -5429
rect -60 -5433 -54 -5429
rect -52 -5433 -51 -5429
rect -39 -5433 -38 -5429
rect -36 -5433 -30 -5429
rect -28 -5433 -27 -5429
rect 213 -5433 214 -5429
rect 216 -5433 218 -5429
rect 222 -5433 224 -5429
rect 226 -5433 227 -5429
rect 239 -5433 240 -5429
rect 242 -5433 248 -5429
rect 250 -5433 251 -5429
rect 263 -5433 264 -5429
rect 266 -5433 272 -5429
rect 274 -5433 276 -5429
rect 280 -5433 282 -5429
rect 284 -5433 290 -5429
rect 292 -5433 293 -5429
rect 305 -5433 306 -5429
rect 308 -5433 314 -5429
rect 316 -5433 318 -5429
rect 322 -5433 324 -5429
rect 326 -5433 332 -5429
rect 334 -5433 335 -5429
rect 347 -5433 348 -5429
rect 350 -5433 356 -5429
rect 358 -5433 360 -5429
rect 364 -5433 366 -5429
rect 368 -5433 374 -5429
rect 376 -5433 377 -5429
rect 389 -5433 390 -5429
rect 392 -5433 398 -5429
rect 400 -5433 401 -5429
rect 470 -5433 471 -5429
rect 473 -5433 474 -5429
rect 569 -5433 570 -5429
rect 572 -5433 574 -5429
rect 578 -5433 580 -5429
rect 582 -5433 583 -5429
rect 595 -5433 596 -5429
rect 598 -5433 604 -5429
rect 606 -5433 607 -5429
rect 619 -5433 620 -5429
rect 622 -5433 628 -5429
rect 630 -5433 632 -5429
rect 636 -5433 638 -5429
rect 640 -5433 646 -5429
rect 648 -5433 649 -5429
rect 661 -5433 662 -5429
rect 664 -5433 670 -5429
rect 672 -5433 674 -5429
rect 678 -5433 680 -5429
rect 682 -5433 688 -5429
rect 690 -5433 691 -5429
rect 703 -5433 704 -5429
rect 706 -5433 712 -5429
rect 714 -5433 716 -5429
rect 720 -5433 722 -5429
rect 724 -5433 730 -5429
rect 732 -5433 733 -5429
rect 745 -5433 746 -5429
rect 748 -5433 754 -5429
rect 756 -5433 757 -5429
rect 871 -5433 872 -5425
rect 874 -5433 875 -5425
rect 967 -5433 968 -5429
rect 970 -5433 972 -5429
rect 976 -5433 978 -5429
rect 980 -5433 981 -5429
rect 993 -5433 994 -5429
rect 996 -5433 1002 -5429
rect 1004 -5433 1005 -5429
rect 1017 -5433 1018 -5429
rect 1020 -5433 1026 -5429
rect 1028 -5433 1030 -5429
rect 1034 -5433 1036 -5429
rect 1038 -5433 1044 -5429
rect 1046 -5433 1047 -5429
rect 1059 -5433 1060 -5429
rect 1062 -5433 1068 -5429
rect 1070 -5433 1072 -5429
rect 1076 -5433 1078 -5429
rect 1080 -5433 1086 -5429
rect 1088 -5433 1089 -5429
rect 1101 -5433 1102 -5429
rect 1104 -5433 1110 -5429
rect 1112 -5433 1114 -5429
rect 1118 -5433 1120 -5429
rect 1122 -5433 1128 -5429
rect 1130 -5433 1131 -5429
rect 1143 -5433 1144 -5429
rect 1146 -5433 1152 -5429
rect 1154 -5433 1155 -5429
rect 1214 -5433 1215 -5429
rect 1217 -5433 1218 -5429
rect 1325 -5433 1326 -5429
rect 1328 -5433 1330 -5429
rect 1334 -5433 1336 -5429
rect 1338 -5433 1339 -5429
rect 1351 -5433 1352 -5429
rect 1354 -5433 1360 -5429
rect 1362 -5433 1363 -5429
rect 1375 -5433 1376 -5429
rect 1378 -5433 1384 -5429
rect 1386 -5433 1388 -5429
rect 1392 -5433 1394 -5429
rect 1396 -5433 1402 -5429
rect 1404 -5433 1405 -5429
rect 1417 -5433 1418 -5429
rect 1420 -5433 1426 -5429
rect 1428 -5433 1430 -5429
rect 1434 -5433 1436 -5429
rect 1438 -5433 1444 -5429
rect 1446 -5433 1447 -5429
rect 1459 -5433 1460 -5429
rect 1462 -5433 1468 -5429
rect 1470 -5433 1472 -5429
rect 1476 -5433 1478 -5429
rect 1480 -5433 1486 -5429
rect 1488 -5433 1489 -5429
rect 1501 -5433 1502 -5429
rect 1504 -5433 1510 -5429
rect 1512 -5433 1513 -5429
rect -1260 -5553 -1259 -5549
rect -1257 -5553 -1255 -5549
rect -1251 -5553 -1249 -5549
rect -1247 -5553 -1246 -5549
rect -1234 -5553 -1233 -5549
rect -1231 -5553 -1225 -5549
rect -1223 -5553 -1222 -5549
rect -1210 -5553 -1209 -5549
rect -1207 -5553 -1201 -5549
rect -1199 -5553 -1197 -5549
rect -1193 -5553 -1191 -5549
rect -1189 -5553 -1183 -5549
rect -1181 -5553 -1180 -5549
rect -1168 -5553 -1167 -5549
rect -1165 -5553 -1159 -5549
rect -1157 -5553 -1155 -5549
rect -1151 -5553 -1149 -5549
rect -1147 -5553 -1141 -5549
rect -1139 -5553 -1138 -5549
rect -1126 -5553 -1125 -5549
rect -1123 -5553 -1117 -5549
rect -1115 -5553 -1113 -5549
rect -1109 -5553 -1107 -5549
rect -1105 -5553 -1099 -5549
rect -1097 -5553 -1096 -5549
rect -1084 -5553 -1083 -5549
rect -1081 -5553 -1075 -5549
rect -1073 -5553 -1072 -5549
rect -1022 -5553 -1021 -5549
rect -1019 -5553 -1018 -5549
rect -931 -5553 -930 -5549
rect -928 -5553 -926 -5549
rect -922 -5553 -920 -5549
rect -918 -5553 -917 -5549
rect -905 -5553 -904 -5549
rect -902 -5553 -896 -5549
rect -894 -5553 -893 -5549
rect -881 -5553 -880 -5549
rect -878 -5553 -872 -5549
rect -870 -5553 -868 -5549
rect -864 -5553 -862 -5549
rect -860 -5553 -854 -5549
rect -852 -5553 -851 -5549
rect -839 -5553 -838 -5549
rect -836 -5553 -830 -5549
rect -828 -5553 -826 -5549
rect -822 -5553 -820 -5549
rect -818 -5553 -812 -5549
rect -810 -5553 -809 -5549
rect -797 -5553 -796 -5549
rect -794 -5553 -788 -5549
rect -786 -5553 -784 -5549
rect -780 -5553 -778 -5549
rect -776 -5553 -770 -5549
rect -768 -5553 -767 -5549
rect -755 -5553 -754 -5549
rect -752 -5553 -746 -5549
rect -744 -5553 -743 -5549
rect -573 -5553 -572 -5549
rect -570 -5553 -568 -5549
rect -564 -5553 -562 -5549
rect -560 -5553 -559 -5549
rect -547 -5553 -546 -5549
rect -544 -5553 -538 -5549
rect -536 -5553 -535 -5549
rect -523 -5553 -522 -5549
rect -520 -5553 -514 -5549
rect -512 -5553 -510 -5549
rect -506 -5553 -504 -5549
rect -502 -5553 -496 -5549
rect -494 -5553 -493 -5549
rect -481 -5553 -480 -5549
rect -478 -5553 -472 -5549
rect -470 -5553 -468 -5549
rect -464 -5553 -462 -5549
rect -460 -5553 -454 -5549
rect -452 -5553 -451 -5549
rect -439 -5553 -438 -5549
rect -436 -5553 -430 -5549
rect -428 -5553 -426 -5549
rect -422 -5553 -420 -5549
rect -418 -5553 -412 -5549
rect -410 -5553 -409 -5549
rect -397 -5553 -396 -5549
rect -394 -5553 -388 -5549
rect -386 -5553 -385 -5549
rect -323 -5553 -322 -5549
rect -320 -5553 -319 -5549
rect -215 -5553 -214 -5549
rect -212 -5553 -210 -5549
rect -206 -5553 -204 -5549
rect -202 -5553 -201 -5549
rect -189 -5553 -188 -5549
rect -186 -5553 -180 -5549
rect -178 -5553 -177 -5549
rect -165 -5553 -164 -5549
rect -162 -5553 -156 -5549
rect -154 -5553 -152 -5549
rect -148 -5553 -146 -5549
rect -144 -5553 -138 -5549
rect -136 -5553 -135 -5549
rect -123 -5553 -122 -5549
rect -120 -5553 -114 -5549
rect -112 -5553 -110 -5549
rect -106 -5553 -104 -5549
rect -102 -5553 -96 -5549
rect -94 -5553 -93 -5549
rect -81 -5553 -80 -5549
rect -78 -5553 -72 -5549
rect -70 -5553 -68 -5549
rect -64 -5553 -62 -5549
rect -60 -5553 -54 -5549
rect -52 -5553 -51 -5549
rect -39 -5553 -38 -5549
rect -36 -5553 -30 -5549
rect -28 -5553 -27 -5549
rect 213 -5553 214 -5549
rect 216 -5553 218 -5549
rect 222 -5553 224 -5549
rect 226 -5553 227 -5549
rect 239 -5553 240 -5549
rect 242 -5553 248 -5549
rect 250 -5553 251 -5549
rect 263 -5553 264 -5549
rect 266 -5553 272 -5549
rect 274 -5553 276 -5549
rect 280 -5553 282 -5549
rect 284 -5553 290 -5549
rect 292 -5553 293 -5549
rect 305 -5553 306 -5549
rect 308 -5553 314 -5549
rect 316 -5553 318 -5549
rect 322 -5553 324 -5549
rect 326 -5553 332 -5549
rect 334 -5553 335 -5549
rect 347 -5553 348 -5549
rect 350 -5553 356 -5549
rect 358 -5553 360 -5549
rect 364 -5553 366 -5549
rect 368 -5553 374 -5549
rect 376 -5553 377 -5549
rect 389 -5553 390 -5549
rect 392 -5553 398 -5549
rect 400 -5553 401 -5549
rect 470 -5553 471 -5549
rect 473 -5553 474 -5549
rect 569 -5553 570 -5549
rect 572 -5553 574 -5549
rect 578 -5553 580 -5549
rect 582 -5553 583 -5549
rect 595 -5553 596 -5549
rect 598 -5553 604 -5549
rect 606 -5553 607 -5549
rect 619 -5553 620 -5549
rect 622 -5553 628 -5549
rect 630 -5553 632 -5549
rect 636 -5553 638 -5549
rect 640 -5553 646 -5549
rect 648 -5553 649 -5549
rect 661 -5553 662 -5549
rect 664 -5553 670 -5549
rect 672 -5553 674 -5549
rect 678 -5553 680 -5549
rect 682 -5553 688 -5549
rect 690 -5553 691 -5549
rect 703 -5553 704 -5549
rect 706 -5553 712 -5549
rect 714 -5553 716 -5549
rect 720 -5553 722 -5549
rect 724 -5553 730 -5549
rect 732 -5553 733 -5549
rect 745 -5553 746 -5549
rect 748 -5553 754 -5549
rect 756 -5553 757 -5549
rect 967 -5553 968 -5549
rect 970 -5553 972 -5549
rect 976 -5553 978 -5549
rect 980 -5553 981 -5549
rect 993 -5553 994 -5549
rect 996 -5553 1002 -5549
rect 1004 -5553 1005 -5549
rect 1017 -5553 1018 -5549
rect 1020 -5553 1026 -5549
rect 1028 -5553 1030 -5549
rect 1034 -5553 1036 -5549
rect 1038 -5553 1044 -5549
rect 1046 -5553 1047 -5549
rect 1059 -5553 1060 -5549
rect 1062 -5553 1068 -5549
rect 1070 -5553 1072 -5549
rect 1076 -5553 1078 -5549
rect 1080 -5553 1086 -5549
rect 1088 -5553 1089 -5549
rect 1101 -5553 1102 -5549
rect 1104 -5553 1110 -5549
rect 1112 -5553 1114 -5549
rect 1118 -5553 1120 -5549
rect 1122 -5553 1128 -5549
rect 1130 -5553 1131 -5549
rect 1143 -5553 1144 -5549
rect 1146 -5553 1152 -5549
rect 1154 -5553 1155 -5549
rect 1214 -5553 1215 -5549
rect 1217 -5553 1218 -5549
rect 1325 -5553 1326 -5549
rect 1328 -5553 1330 -5549
rect 1334 -5553 1336 -5549
rect 1338 -5553 1339 -5549
rect 1351 -5553 1352 -5549
rect 1354 -5553 1360 -5549
rect 1362 -5553 1363 -5549
rect 1375 -5553 1376 -5549
rect 1378 -5553 1384 -5549
rect 1386 -5553 1388 -5549
rect 1392 -5553 1394 -5549
rect 1396 -5553 1402 -5549
rect 1404 -5553 1405 -5549
rect 1417 -5553 1418 -5549
rect 1420 -5553 1426 -5549
rect 1428 -5553 1430 -5549
rect 1434 -5553 1436 -5549
rect 1438 -5553 1444 -5549
rect 1446 -5553 1447 -5549
rect 1459 -5553 1460 -5549
rect 1462 -5553 1468 -5549
rect 1470 -5553 1472 -5549
rect 1476 -5553 1478 -5549
rect 1480 -5553 1486 -5549
rect 1488 -5553 1489 -5549
rect 1501 -5553 1502 -5549
rect 1504 -5553 1510 -5549
rect 1512 -5553 1513 -5549
rect -1260 -5670 -1259 -5666
rect -1257 -5670 -1255 -5666
rect -1251 -5670 -1249 -5666
rect -1247 -5670 -1246 -5666
rect -1234 -5670 -1233 -5666
rect -1231 -5670 -1225 -5666
rect -1223 -5670 -1222 -5666
rect -1210 -5670 -1209 -5666
rect -1207 -5670 -1201 -5666
rect -1199 -5670 -1197 -5666
rect -1193 -5670 -1191 -5666
rect -1189 -5670 -1183 -5666
rect -1181 -5670 -1180 -5666
rect -1168 -5670 -1167 -5666
rect -1165 -5670 -1159 -5666
rect -1157 -5670 -1155 -5666
rect -1151 -5670 -1149 -5666
rect -1147 -5670 -1141 -5666
rect -1139 -5670 -1138 -5666
rect -1126 -5670 -1125 -5666
rect -1123 -5670 -1117 -5666
rect -1115 -5670 -1113 -5666
rect -1109 -5670 -1107 -5666
rect -1105 -5670 -1099 -5666
rect -1097 -5670 -1096 -5666
rect -1084 -5670 -1083 -5666
rect -1081 -5670 -1075 -5666
rect -1073 -5670 -1072 -5666
rect -931 -5670 -930 -5666
rect -928 -5670 -926 -5666
rect -922 -5670 -920 -5666
rect -918 -5670 -917 -5666
rect -905 -5670 -904 -5666
rect -902 -5670 -896 -5666
rect -894 -5670 -893 -5666
rect -881 -5670 -880 -5666
rect -878 -5670 -872 -5666
rect -870 -5670 -868 -5666
rect -864 -5670 -862 -5666
rect -860 -5670 -854 -5666
rect -852 -5670 -851 -5666
rect -839 -5670 -838 -5666
rect -836 -5670 -830 -5666
rect -828 -5670 -826 -5666
rect -822 -5670 -820 -5666
rect -818 -5670 -812 -5666
rect -810 -5670 -809 -5666
rect -797 -5670 -796 -5666
rect -794 -5670 -788 -5666
rect -786 -5670 -784 -5666
rect -780 -5670 -778 -5666
rect -776 -5670 -770 -5666
rect -768 -5670 -767 -5666
rect -755 -5670 -754 -5666
rect -752 -5670 -746 -5666
rect -744 -5670 -743 -5666
rect -573 -5670 -572 -5666
rect -570 -5670 -568 -5666
rect -564 -5670 -562 -5666
rect -560 -5670 -559 -5666
rect -547 -5670 -546 -5666
rect -544 -5670 -538 -5666
rect -536 -5670 -535 -5666
rect -523 -5670 -522 -5666
rect -520 -5670 -514 -5666
rect -512 -5670 -510 -5666
rect -506 -5670 -504 -5666
rect -502 -5670 -496 -5666
rect -494 -5670 -493 -5666
rect -481 -5670 -480 -5666
rect -478 -5670 -472 -5666
rect -470 -5670 -468 -5666
rect -464 -5670 -462 -5666
rect -460 -5670 -454 -5666
rect -452 -5670 -451 -5666
rect -439 -5670 -438 -5666
rect -436 -5670 -430 -5666
rect -428 -5670 -426 -5666
rect -422 -5670 -420 -5666
rect -418 -5670 -412 -5666
rect -410 -5670 -409 -5666
rect -397 -5670 -396 -5666
rect -394 -5670 -388 -5666
rect -386 -5670 -385 -5666
rect -215 -5670 -214 -5666
rect -212 -5670 -210 -5666
rect -206 -5670 -204 -5666
rect -202 -5670 -201 -5666
rect -189 -5670 -188 -5666
rect -186 -5670 -180 -5666
rect -178 -5670 -177 -5666
rect -165 -5670 -164 -5666
rect -162 -5670 -156 -5666
rect -154 -5670 -152 -5666
rect -148 -5670 -146 -5666
rect -144 -5670 -138 -5666
rect -136 -5670 -135 -5666
rect -123 -5670 -122 -5666
rect -120 -5670 -114 -5666
rect -112 -5670 -110 -5666
rect -106 -5670 -104 -5666
rect -102 -5670 -96 -5666
rect -94 -5670 -93 -5666
rect -81 -5670 -80 -5666
rect -78 -5670 -72 -5666
rect -70 -5670 -68 -5666
rect -64 -5670 -62 -5666
rect -60 -5670 -54 -5666
rect -52 -5670 -51 -5666
rect -39 -5670 -38 -5666
rect -36 -5670 -30 -5666
rect -28 -5670 -27 -5666
rect 213 -5670 214 -5666
rect 216 -5670 218 -5666
rect 222 -5670 224 -5666
rect 226 -5670 227 -5666
rect 239 -5670 240 -5666
rect 242 -5670 248 -5666
rect 250 -5670 251 -5666
rect 263 -5670 264 -5666
rect 266 -5670 272 -5666
rect 274 -5670 276 -5666
rect 280 -5670 282 -5666
rect 284 -5670 290 -5666
rect 292 -5670 293 -5666
rect 305 -5670 306 -5666
rect 308 -5670 314 -5666
rect 316 -5670 318 -5666
rect 322 -5670 324 -5666
rect 326 -5670 332 -5666
rect 334 -5670 335 -5666
rect 347 -5670 348 -5666
rect 350 -5670 356 -5666
rect 358 -5670 360 -5666
rect 364 -5670 366 -5666
rect 368 -5670 374 -5666
rect 376 -5670 377 -5666
rect 389 -5670 390 -5666
rect 392 -5670 398 -5666
rect 400 -5670 401 -5666
rect 569 -5670 570 -5666
rect 572 -5670 574 -5666
rect 578 -5670 580 -5666
rect 582 -5670 583 -5666
rect 595 -5670 596 -5666
rect 598 -5670 604 -5666
rect 606 -5670 607 -5666
rect 619 -5670 620 -5666
rect 622 -5670 628 -5666
rect 630 -5670 632 -5666
rect 636 -5670 638 -5666
rect 640 -5670 646 -5666
rect 648 -5670 649 -5666
rect 661 -5670 662 -5666
rect 664 -5670 670 -5666
rect 672 -5670 674 -5666
rect 678 -5670 680 -5666
rect 682 -5670 688 -5666
rect 690 -5670 691 -5666
rect 703 -5670 704 -5666
rect 706 -5670 712 -5666
rect 714 -5670 716 -5666
rect 720 -5670 722 -5666
rect 724 -5670 730 -5666
rect 732 -5670 733 -5666
rect 745 -5670 746 -5666
rect 748 -5670 754 -5666
rect 756 -5670 757 -5666
rect -1335 -5787 -1334 -5783
rect -1332 -5787 -1326 -5783
rect -1324 -5787 -1322 -5783
rect -1318 -5787 -1316 -5783
rect -1314 -5787 -1313 -5783
rect -931 -5787 -930 -5783
rect -928 -5787 -922 -5783
rect -920 -5787 -918 -5783
rect -914 -5787 -912 -5783
rect -910 -5787 -909 -5783
rect -573 -5787 -572 -5783
rect -570 -5787 -564 -5783
rect -562 -5787 -560 -5783
rect -556 -5787 -554 -5783
rect -552 -5787 -551 -5783
rect -215 -5787 -214 -5783
rect -212 -5787 -206 -5783
rect -204 -5787 -202 -5783
rect -198 -5787 -196 -5783
rect -194 -5787 -193 -5783
rect 213 -5787 214 -5783
rect 216 -5787 222 -5783
rect 224 -5787 226 -5783
rect 230 -5787 232 -5783
rect 234 -5787 235 -5783
rect 569 -5787 570 -5783
rect 572 -5787 578 -5783
rect 580 -5787 582 -5783
rect 586 -5787 588 -5783
rect 590 -5787 591 -5783
rect 967 -5787 968 -5783
rect 970 -5787 976 -5783
rect 978 -5787 980 -5783
rect 984 -5787 986 -5783
rect 988 -5787 989 -5783
rect 1325 -5787 1326 -5783
rect 1328 -5787 1334 -5783
rect 1336 -5787 1338 -5783
rect 1342 -5787 1344 -5783
rect 1346 -5787 1347 -5783
rect -1260 -5906 -1259 -5902
rect -1257 -5906 -1255 -5902
rect -1251 -5906 -1249 -5902
rect -1247 -5906 -1246 -5902
rect -1234 -5906 -1233 -5902
rect -1231 -5906 -1229 -5902
rect -1225 -5906 -1223 -5902
rect -1221 -5906 -1215 -5902
rect -1213 -5906 -1211 -5902
rect -1207 -5906 -1205 -5902
rect -1203 -5906 -1202 -5902
rect -1190 -5906 -1189 -5902
rect -1187 -5906 -1181 -5902
rect -1179 -5906 -1177 -5902
rect -1173 -5906 -1171 -5902
rect -1169 -5906 -1168 -5902
rect -931 -5906 -930 -5902
rect -928 -5906 -926 -5902
rect -922 -5906 -920 -5902
rect -918 -5906 -917 -5902
rect -905 -5906 -904 -5902
rect -902 -5906 -900 -5902
rect -896 -5906 -894 -5902
rect -892 -5906 -891 -5902
rect -879 -5906 -878 -5902
rect -876 -5906 -875 -5902
rect -871 -5906 -868 -5902
rect -866 -5906 -860 -5902
rect -858 -5906 -857 -5902
rect -853 -5906 -850 -5902
rect -848 -5906 -847 -5902
rect -835 -5906 -834 -5902
rect -832 -5906 -826 -5902
rect -824 -5906 -822 -5902
rect -818 -5906 -816 -5902
rect -814 -5906 -813 -5902
rect -801 -5906 -800 -5902
rect -798 -5906 -796 -5902
rect -792 -5906 -790 -5902
rect -788 -5906 -782 -5902
rect -780 -5906 -778 -5902
rect -774 -5906 -772 -5902
rect -770 -5906 -769 -5902
rect -757 -5906 -756 -5902
rect -754 -5906 -748 -5902
rect -746 -5906 -745 -5902
rect -733 -5906 -732 -5902
rect -730 -5906 -725 -5902
rect -721 -5906 -716 -5902
rect -714 -5906 -713 -5902
rect -709 -5906 -708 -5902
rect -706 -5906 -704 -5902
rect -700 -5906 -698 -5902
rect -696 -5906 -695 -5902
rect -573 -5906 -572 -5902
rect -570 -5906 -568 -5902
rect -564 -5906 -562 -5902
rect -560 -5906 -559 -5902
rect -547 -5906 -546 -5902
rect -544 -5906 -542 -5902
rect -538 -5906 -536 -5902
rect -534 -5906 -533 -5902
rect -521 -5906 -520 -5902
rect -518 -5906 -517 -5902
rect -513 -5906 -510 -5902
rect -508 -5906 -502 -5902
rect -500 -5906 -499 -5902
rect -495 -5906 -492 -5902
rect -490 -5906 -489 -5902
rect -477 -5906 -476 -5902
rect -474 -5906 -468 -5902
rect -466 -5906 -464 -5902
rect -460 -5906 -458 -5902
rect -456 -5906 -455 -5902
rect -443 -5906 -442 -5902
rect -440 -5906 -438 -5902
rect -434 -5906 -432 -5902
rect -430 -5906 -424 -5902
rect -422 -5906 -420 -5902
rect -416 -5906 -414 -5902
rect -412 -5906 -411 -5902
rect -399 -5906 -398 -5902
rect -396 -5906 -390 -5902
rect -388 -5906 -387 -5902
rect -375 -5906 -374 -5902
rect -372 -5906 -367 -5902
rect -363 -5906 -358 -5902
rect -356 -5906 -355 -5902
rect -351 -5906 -350 -5902
rect -348 -5906 -346 -5902
rect -342 -5906 -340 -5902
rect -338 -5906 -337 -5902
rect -215 -5906 -214 -5902
rect -212 -5906 -210 -5902
rect -206 -5906 -204 -5902
rect -202 -5906 -201 -5902
rect -189 -5906 -188 -5902
rect -186 -5906 -184 -5902
rect -180 -5906 -178 -5902
rect -176 -5906 -175 -5902
rect -163 -5906 -162 -5902
rect -160 -5906 -159 -5902
rect -155 -5906 -152 -5902
rect -150 -5906 -144 -5902
rect -142 -5906 -141 -5902
rect -137 -5906 -134 -5902
rect -132 -5906 -131 -5902
rect -119 -5906 -118 -5902
rect -116 -5906 -110 -5902
rect -108 -5906 -106 -5902
rect -102 -5906 -100 -5902
rect -98 -5906 -97 -5902
rect -85 -5906 -84 -5902
rect -82 -5906 -80 -5902
rect -76 -5906 -74 -5902
rect -72 -5906 -66 -5902
rect -64 -5906 -62 -5902
rect -58 -5906 -56 -5902
rect -54 -5906 -53 -5902
rect -41 -5906 -40 -5902
rect -38 -5906 -32 -5902
rect -30 -5906 -29 -5902
rect -17 -5906 -16 -5902
rect -14 -5906 -9 -5902
rect -5 -5906 0 -5902
rect 2 -5906 3 -5902
rect 7 -5906 8 -5902
rect 10 -5906 12 -5902
rect 16 -5906 18 -5902
rect 20 -5906 21 -5902
rect 213 -5906 214 -5902
rect 216 -5906 218 -5902
rect 222 -5906 224 -5902
rect 226 -5906 227 -5902
rect 239 -5906 240 -5902
rect 242 -5906 244 -5902
rect 248 -5906 250 -5902
rect 252 -5906 253 -5902
rect 265 -5906 266 -5902
rect 268 -5906 269 -5902
rect 273 -5906 276 -5902
rect 278 -5906 284 -5902
rect 286 -5906 287 -5902
rect 291 -5906 294 -5902
rect 296 -5906 297 -5902
rect 309 -5906 310 -5902
rect 312 -5906 318 -5902
rect 320 -5906 322 -5902
rect 326 -5906 328 -5902
rect 330 -5906 331 -5902
rect 343 -5906 344 -5902
rect 346 -5906 348 -5902
rect 352 -5906 354 -5902
rect 356 -5906 362 -5902
rect 364 -5906 366 -5902
rect 370 -5906 372 -5902
rect 374 -5906 375 -5902
rect 387 -5906 388 -5902
rect 390 -5906 396 -5902
rect 398 -5906 399 -5902
rect 411 -5906 412 -5902
rect 414 -5906 419 -5902
rect 423 -5906 428 -5902
rect 430 -5906 431 -5902
rect 435 -5906 436 -5902
rect 438 -5906 440 -5902
rect 444 -5906 446 -5902
rect 448 -5906 449 -5902
rect 569 -5906 570 -5902
rect 572 -5906 574 -5902
rect 578 -5906 580 -5902
rect 582 -5906 583 -5902
rect 595 -5906 596 -5902
rect 598 -5906 600 -5902
rect 604 -5906 606 -5902
rect 608 -5906 609 -5902
rect 621 -5906 622 -5902
rect 624 -5906 625 -5902
rect 629 -5906 632 -5902
rect 634 -5906 640 -5902
rect 642 -5906 643 -5902
rect 647 -5906 650 -5902
rect 652 -5906 653 -5902
rect 665 -5906 666 -5902
rect 668 -5906 674 -5902
rect 676 -5906 678 -5902
rect 682 -5906 684 -5902
rect 686 -5906 687 -5902
rect 699 -5906 700 -5902
rect 702 -5906 704 -5902
rect 708 -5906 710 -5902
rect 712 -5906 718 -5902
rect 720 -5906 722 -5902
rect 726 -5906 728 -5902
rect 730 -5906 731 -5902
rect 743 -5906 744 -5902
rect 746 -5906 752 -5902
rect 754 -5906 755 -5902
rect 767 -5906 768 -5902
rect 770 -5906 775 -5902
rect 779 -5906 784 -5902
rect 786 -5906 787 -5902
rect 791 -5906 792 -5902
rect 794 -5906 796 -5902
rect 800 -5906 802 -5902
rect 804 -5906 805 -5902
rect 967 -5906 968 -5902
rect 970 -5906 972 -5902
rect 976 -5906 978 -5902
rect 980 -5906 981 -5902
rect 993 -5906 994 -5902
rect 996 -5906 998 -5902
rect 1002 -5906 1004 -5902
rect 1006 -5906 1007 -5902
rect 1019 -5906 1020 -5902
rect 1022 -5906 1023 -5902
rect 1027 -5906 1030 -5902
rect 1032 -5906 1038 -5902
rect 1040 -5906 1041 -5902
rect 1045 -5906 1048 -5902
rect 1050 -5906 1051 -5902
rect 1063 -5906 1064 -5902
rect 1066 -5906 1072 -5902
rect 1074 -5906 1076 -5902
rect 1080 -5906 1082 -5902
rect 1084 -5906 1085 -5902
rect 1097 -5906 1098 -5902
rect 1100 -5906 1102 -5902
rect 1106 -5906 1108 -5902
rect 1110 -5906 1116 -5902
rect 1118 -5906 1120 -5902
rect 1124 -5906 1126 -5902
rect 1128 -5906 1129 -5902
rect 1141 -5906 1142 -5902
rect 1144 -5906 1150 -5902
rect 1152 -5906 1153 -5902
rect 1165 -5906 1166 -5902
rect 1168 -5906 1173 -5902
rect 1177 -5906 1182 -5902
rect 1184 -5906 1185 -5902
rect 1189 -5906 1190 -5902
rect 1192 -5906 1194 -5902
rect 1198 -5906 1200 -5902
rect 1202 -5906 1203 -5902
rect 1325 -5906 1326 -5902
rect 1328 -5906 1330 -5902
rect 1334 -5906 1336 -5902
rect 1338 -5906 1339 -5902
rect 1351 -5906 1352 -5902
rect 1354 -5906 1356 -5902
rect 1360 -5906 1362 -5902
rect 1364 -5906 1365 -5902
rect 1377 -5906 1378 -5902
rect 1380 -5906 1381 -5902
rect 1385 -5906 1388 -5902
rect 1390 -5906 1396 -5902
rect 1398 -5906 1399 -5902
rect 1403 -5906 1406 -5902
rect 1408 -5906 1409 -5902
rect 1421 -5906 1422 -5902
rect 1424 -5906 1430 -5902
rect 1432 -5906 1434 -5902
rect 1438 -5906 1440 -5902
rect 1442 -5906 1443 -5902
rect 1455 -5906 1456 -5902
rect 1458 -5906 1460 -5902
rect 1464 -5906 1466 -5902
rect 1468 -5906 1474 -5902
rect 1476 -5906 1478 -5902
rect 1482 -5906 1484 -5902
rect 1486 -5906 1487 -5902
rect 1499 -5906 1500 -5902
rect 1502 -5906 1508 -5902
rect 1510 -5906 1511 -5902
rect 1523 -5906 1524 -5902
rect 1526 -5906 1531 -5902
rect 1535 -5906 1540 -5902
rect 1542 -5906 1543 -5902
rect 1547 -5906 1548 -5902
rect 1550 -5906 1552 -5902
rect 1556 -5906 1558 -5902
rect 1560 -5906 1561 -5902
rect -1260 -6029 -1259 -6025
rect -1257 -6029 -1255 -6025
rect -1251 -6029 -1249 -6025
rect -1247 -6029 -1246 -6025
rect -1234 -6029 -1233 -6025
rect -1231 -6029 -1225 -6025
rect -1223 -6029 -1222 -6025
rect -1210 -6029 -1209 -6025
rect -1207 -6029 -1201 -6025
rect -1199 -6029 -1197 -6025
rect -1193 -6029 -1191 -6025
rect -1189 -6029 -1183 -6025
rect -1181 -6029 -1180 -6025
rect -1168 -6029 -1167 -6025
rect -1165 -6029 -1159 -6025
rect -1157 -6029 -1155 -6025
rect -1151 -6029 -1149 -6025
rect -1147 -6029 -1141 -6025
rect -1139 -6029 -1138 -6025
rect -1126 -6029 -1125 -6025
rect -1123 -6029 -1117 -6025
rect -1115 -6029 -1113 -6025
rect -1109 -6029 -1107 -6025
rect -1105 -6029 -1099 -6025
rect -1097 -6029 -1096 -6025
rect -1084 -6029 -1083 -6025
rect -1081 -6029 -1075 -6025
rect -1073 -6029 -1072 -6025
rect -931 -6029 -930 -6025
rect -928 -6029 -926 -6025
rect -922 -6029 -920 -6025
rect -918 -6029 -917 -6025
rect -905 -6029 -904 -6025
rect -902 -6029 -896 -6025
rect -894 -6029 -893 -6025
rect -881 -6029 -880 -6025
rect -878 -6029 -872 -6025
rect -870 -6029 -868 -6025
rect -864 -6029 -862 -6025
rect -860 -6029 -854 -6025
rect -852 -6029 -851 -6025
rect -839 -6029 -838 -6025
rect -836 -6029 -830 -6025
rect -828 -6029 -826 -6025
rect -822 -6029 -820 -6025
rect -818 -6029 -812 -6025
rect -810 -6029 -809 -6025
rect -797 -6029 -796 -6025
rect -794 -6029 -788 -6025
rect -786 -6029 -784 -6025
rect -780 -6029 -778 -6025
rect -776 -6029 -770 -6025
rect -768 -6029 -767 -6025
rect -755 -6029 -754 -6025
rect -752 -6029 -746 -6025
rect -744 -6029 -743 -6025
rect -573 -6029 -572 -6025
rect -570 -6029 -568 -6025
rect -564 -6029 -562 -6025
rect -560 -6029 -559 -6025
rect -547 -6029 -546 -6025
rect -544 -6029 -538 -6025
rect -536 -6029 -535 -6025
rect -523 -6029 -522 -6025
rect -520 -6029 -514 -6025
rect -512 -6029 -510 -6025
rect -506 -6029 -504 -6025
rect -502 -6029 -496 -6025
rect -494 -6029 -493 -6025
rect -481 -6029 -480 -6025
rect -478 -6029 -472 -6025
rect -470 -6029 -468 -6025
rect -464 -6029 -462 -6025
rect -460 -6029 -454 -6025
rect -452 -6029 -451 -6025
rect -439 -6029 -438 -6025
rect -436 -6029 -430 -6025
rect -428 -6029 -426 -6025
rect -422 -6029 -420 -6025
rect -418 -6029 -412 -6025
rect -410 -6029 -409 -6025
rect -397 -6029 -396 -6025
rect -394 -6029 -388 -6025
rect -386 -6029 -385 -6025
rect -215 -6029 -214 -6025
rect -212 -6029 -210 -6025
rect -206 -6029 -204 -6025
rect -202 -6029 -201 -6025
rect -189 -6029 -188 -6025
rect -186 -6029 -180 -6025
rect -178 -6029 -177 -6025
rect -165 -6029 -164 -6025
rect -162 -6029 -156 -6025
rect -154 -6029 -152 -6025
rect -148 -6029 -146 -6025
rect -144 -6029 -138 -6025
rect -136 -6029 -135 -6025
rect -123 -6029 -122 -6025
rect -120 -6029 -114 -6025
rect -112 -6029 -110 -6025
rect -106 -6029 -104 -6025
rect -102 -6029 -96 -6025
rect -94 -6029 -93 -6025
rect -81 -6029 -80 -6025
rect -78 -6029 -72 -6025
rect -70 -6029 -68 -6025
rect -64 -6029 -62 -6025
rect -60 -6029 -54 -6025
rect -52 -6029 -51 -6025
rect -39 -6029 -38 -6025
rect -36 -6029 -30 -6025
rect -28 -6029 -27 -6025
rect 213 -6029 214 -6025
rect 216 -6029 218 -6025
rect 222 -6029 224 -6025
rect 226 -6029 227 -6025
rect 239 -6029 240 -6025
rect 242 -6029 248 -6025
rect 250 -6029 251 -6025
rect 263 -6029 264 -6025
rect 266 -6029 272 -6025
rect 274 -6029 276 -6025
rect 280 -6029 282 -6025
rect 284 -6029 290 -6025
rect 292 -6029 293 -6025
rect 305 -6029 306 -6025
rect 308 -6029 314 -6025
rect 316 -6029 318 -6025
rect 322 -6029 324 -6025
rect 326 -6029 332 -6025
rect 334 -6029 335 -6025
rect 347 -6029 348 -6025
rect 350 -6029 356 -6025
rect 358 -6029 360 -6025
rect 364 -6029 366 -6025
rect 368 -6029 374 -6025
rect 376 -6029 377 -6025
rect 389 -6029 390 -6025
rect 392 -6029 398 -6025
rect 400 -6029 401 -6025
rect 569 -6029 570 -6025
rect 572 -6029 574 -6025
rect 578 -6029 580 -6025
rect 582 -6029 583 -6025
rect 595 -6029 596 -6025
rect 598 -6029 604 -6025
rect 606 -6029 607 -6025
rect 619 -6029 620 -6025
rect 622 -6029 628 -6025
rect 630 -6029 632 -6025
rect 636 -6029 638 -6025
rect 640 -6029 646 -6025
rect 648 -6029 649 -6025
rect 661 -6029 662 -6025
rect 664 -6029 670 -6025
rect 672 -6029 674 -6025
rect 678 -6029 680 -6025
rect 682 -6029 688 -6025
rect 690 -6029 691 -6025
rect 703 -6029 704 -6025
rect 706 -6029 712 -6025
rect 714 -6029 716 -6025
rect 720 -6029 722 -6025
rect 724 -6029 730 -6025
rect 732 -6029 733 -6025
rect 745 -6029 746 -6025
rect 748 -6029 754 -6025
rect 756 -6029 757 -6025
rect 967 -6029 968 -6025
rect 970 -6029 972 -6025
rect 976 -6029 978 -6025
rect 980 -6029 981 -6025
rect 993 -6029 994 -6025
rect 996 -6029 1002 -6025
rect 1004 -6029 1005 -6025
rect 1017 -6029 1018 -6025
rect 1020 -6029 1026 -6025
rect 1028 -6029 1030 -6025
rect 1034 -6029 1036 -6025
rect 1038 -6029 1044 -6025
rect 1046 -6029 1047 -6025
rect 1059 -6029 1060 -6025
rect 1062 -6029 1068 -6025
rect 1070 -6029 1072 -6025
rect 1076 -6029 1078 -6025
rect 1080 -6029 1086 -6025
rect 1088 -6029 1089 -6025
rect 1101 -6029 1102 -6025
rect 1104 -6029 1110 -6025
rect 1112 -6029 1114 -6025
rect 1118 -6029 1120 -6025
rect 1122 -6029 1128 -6025
rect 1130 -6029 1131 -6025
rect 1143 -6029 1144 -6025
rect 1146 -6029 1152 -6025
rect 1154 -6029 1155 -6025
rect 1325 -6029 1326 -6025
rect 1328 -6029 1330 -6025
rect 1334 -6029 1336 -6025
rect 1338 -6029 1339 -6025
rect 1351 -6029 1352 -6025
rect 1354 -6029 1360 -6025
rect 1362 -6029 1363 -6025
rect 1375 -6029 1376 -6025
rect 1378 -6029 1384 -6025
rect 1386 -6029 1388 -6025
rect 1392 -6029 1394 -6025
rect 1396 -6029 1402 -6025
rect 1404 -6029 1405 -6025
rect 1417 -6029 1418 -6025
rect 1420 -6029 1426 -6025
rect 1428 -6029 1430 -6025
rect 1434 -6029 1436 -6025
rect 1438 -6029 1444 -6025
rect 1446 -6029 1447 -6025
rect 1459 -6029 1460 -6025
rect 1462 -6029 1468 -6025
rect 1470 -6029 1472 -6025
rect 1476 -6029 1478 -6025
rect 1480 -6029 1486 -6025
rect 1488 -6029 1489 -6025
rect 1501 -6029 1502 -6025
rect 1504 -6029 1510 -6025
rect 1512 -6029 1513 -6025
rect 1325 -6147 1326 -6143
rect 1328 -6147 1330 -6143
rect 1334 -6147 1336 -6143
rect 1338 -6147 1339 -6143
rect 1351 -6147 1352 -6143
rect 1354 -6147 1360 -6143
rect 1362 -6147 1363 -6143
rect 1375 -6147 1376 -6143
rect 1378 -6147 1384 -6143
rect 1386 -6147 1388 -6143
rect 1392 -6147 1394 -6143
rect 1396 -6147 1402 -6143
rect 1404 -6147 1405 -6143
rect 1417 -6147 1418 -6143
rect 1420 -6147 1426 -6143
rect 1428 -6147 1430 -6143
rect 1434 -6147 1436 -6143
rect 1438 -6147 1444 -6143
rect 1446 -6147 1447 -6143
rect 1459 -6147 1460 -6143
rect 1462 -6147 1468 -6143
rect 1470 -6147 1472 -6143
rect 1476 -6147 1478 -6143
rect 1480 -6147 1486 -6143
rect 1488 -6147 1489 -6143
rect 1501 -6147 1502 -6143
rect 1504 -6147 1510 -6143
rect 1512 -6147 1513 -6143
<< pdiffusion >>
rect -1333 -1046 -1332 -1038
rect -1330 -1046 -1329 -1038
rect -1325 -1046 -1324 -1038
rect -1322 -1046 -1320 -1038
rect -1316 -1046 -1314 -1038
rect -1312 -1046 -1311 -1038
rect -932 -1046 -931 -1038
rect -929 -1046 -928 -1038
rect -924 -1046 -923 -1038
rect -921 -1046 -919 -1038
rect -915 -1046 -913 -1038
rect -911 -1046 -910 -1038
rect -573 -1046 -572 -1038
rect -570 -1046 -569 -1038
rect -565 -1046 -564 -1038
rect -562 -1046 -560 -1038
rect -556 -1046 -554 -1038
rect -552 -1046 -551 -1038
rect -215 -1046 -214 -1038
rect -212 -1046 -211 -1038
rect -207 -1046 -206 -1038
rect -204 -1046 -202 -1038
rect -198 -1046 -196 -1038
rect -194 -1046 -193 -1038
rect 213 -1046 214 -1038
rect 216 -1046 217 -1038
rect 221 -1046 222 -1038
rect 224 -1046 226 -1038
rect 230 -1046 232 -1038
rect 234 -1046 235 -1038
rect 569 -1046 570 -1038
rect 572 -1046 573 -1038
rect 577 -1046 578 -1038
rect 580 -1046 582 -1038
rect 586 -1046 588 -1038
rect 590 -1046 591 -1038
rect 967 -1046 968 -1038
rect 970 -1046 971 -1038
rect 975 -1046 976 -1038
rect 978 -1046 980 -1038
rect 984 -1046 986 -1038
rect 988 -1046 989 -1038
rect 1325 -1046 1326 -1038
rect 1328 -1046 1329 -1038
rect 1333 -1046 1334 -1038
rect 1336 -1046 1338 -1038
rect 1342 -1046 1344 -1038
rect 1346 -1046 1347 -1038
rect -1256 -1160 -1255 -1152
rect -1253 -1160 -1251 -1152
rect -1247 -1160 -1245 -1152
rect -1243 -1160 -1242 -1152
rect -1230 -1160 -1229 -1152
rect -1227 -1160 -1226 -1152
rect -1222 -1160 -1221 -1152
rect -1219 -1160 -1214 -1152
rect -1210 -1160 -1205 -1152
rect -1203 -1160 -1202 -1152
rect -1198 -1160 -1197 -1152
rect -1195 -1160 -1193 -1152
rect -1189 -1160 -1187 -1152
rect -1185 -1160 -1184 -1152
rect -1180 -1160 -1179 -1152
rect -1177 -1160 -1172 -1152
rect -1168 -1160 -1163 -1152
rect -1161 -1160 -1160 -1152
rect -1156 -1160 -1155 -1152
rect -1153 -1160 -1151 -1152
rect -1147 -1160 -1145 -1152
rect -1143 -1160 -1142 -1152
rect -1138 -1160 -1137 -1152
rect -1135 -1160 -1130 -1152
rect -1126 -1160 -1121 -1152
rect -1119 -1160 -1118 -1152
rect -1114 -1160 -1113 -1152
rect -1111 -1160 -1109 -1152
rect -1105 -1160 -1103 -1152
rect -1101 -1160 -1100 -1152
rect -1096 -1160 -1095 -1152
rect -1093 -1160 -1088 -1152
rect -1084 -1160 -1079 -1152
rect -1077 -1160 -1076 -1152
rect -1072 -1160 -1071 -1152
rect -1069 -1160 -1068 -1152
rect -931 -1160 -930 -1152
rect -928 -1160 -926 -1152
rect -922 -1160 -920 -1152
rect -918 -1160 -917 -1152
rect -905 -1160 -904 -1152
rect -902 -1160 -901 -1152
rect -897 -1160 -896 -1152
rect -894 -1160 -889 -1152
rect -885 -1160 -880 -1152
rect -878 -1160 -877 -1152
rect -873 -1160 -872 -1152
rect -870 -1160 -868 -1152
rect -864 -1160 -862 -1152
rect -860 -1160 -859 -1152
rect -855 -1160 -854 -1152
rect -852 -1160 -847 -1152
rect -843 -1160 -838 -1152
rect -836 -1160 -835 -1152
rect -831 -1160 -830 -1152
rect -828 -1160 -826 -1152
rect -822 -1160 -820 -1152
rect -818 -1160 -817 -1152
rect -813 -1160 -812 -1152
rect -810 -1160 -805 -1152
rect -801 -1160 -796 -1152
rect -794 -1160 -793 -1152
rect -789 -1160 -788 -1152
rect -786 -1160 -784 -1152
rect -780 -1160 -778 -1152
rect -776 -1160 -775 -1152
rect -771 -1160 -770 -1152
rect -768 -1160 -763 -1152
rect -759 -1160 -754 -1152
rect -752 -1160 -751 -1152
rect -747 -1160 -746 -1152
rect -744 -1160 -743 -1152
rect -573 -1160 -572 -1152
rect -570 -1160 -568 -1152
rect -564 -1160 -562 -1152
rect -560 -1160 -559 -1152
rect -547 -1160 -546 -1152
rect -544 -1160 -543 -1152
rect -539 -1160 -538 -1152
rect -536 -1160 -531 -1152
rect -527 -1160 -522 -1152
rect -520 -1160 -519 -1152
rect -515 -1160 -514 -1152
rect -512 -1160 -510 -1152
rect -506 -1160 -504 -1152
rect -502 -1160 -501 -1152
rect -497 -1160 -496 -1152
rect -494 -1160 -489 -1152
rect -485 -1160 -480 -1152
rect -478 -1160 -477 -1152
rect -473 -1160 -472 -1152
rect -470 -1160 -468 -1152
rect -464 -1160 -462 -1152
rect -460 -1160 -459 -1152
rect -455 -1160 -454 -1152
rect -452 -1160 -447 -1152
rect -443 -1160 -438 -1152
rect -436 -1160 -435 -1152
rect -431 -1160 -430 -1152
rect -428 -1160 -426 -1152
rect -422 -1160 -420 -1152
rect -418 -1160 -417 -1152
rect -413 -1160 -412 -1152
rect -410 -1160 -405 -1152
rect -401 -1160 -396 -1152
rect -394 -1160 -393 -1152
rect -389 -1160 -388 -1152
rect -386 -1160 -385 -1152
rect -215 -1160 -214 -1152
rect -212 -1160 -210 -1152
rect -206 -1160 -204 -1152
rect -202 -1160 -201 -1152
rect -189 -1160 -188 -1152
rect -186 -1160 -185 -1152
rect -181 -1160 -180 -1152
rect -178 -1160 -173 -1152
rect -169 -1160 -164 -1152
rect -162 -1160 -161 -1152
rect -157 -1160 -156 -1152
rect -154 -1160 -152 -1152
rect -148 -1160 -146 -1152
rect -144 -1160 -143 -1152
rect -139 -1160 -138 -1152
rect -136 -1160 -131 -1152
rect -127 -1160 -122 -1152
rect -120 -1160 -119 -1152
rect -115 -1160 -114 -1152
rect -112 -1160 -110 -1152
rect -106 -1160 -104 -1152
rect -102 -1160 -101 -1152
rect -97 -1160 -96 -1152
rect -94 -1160 -89 -1152
rect -85 -1160 -80 -1152
rect -78 -1160 -77 -1152
rect -73 -1160 -72 -1152
rect -70 -1160 -68 -1152
rect -64 -1160 -62 -1152
rect -60 -1160 -59 -1152
rect -55 -1160 -54 -1152
rect -52 -1160 -47 -1152
rect -43 -1160 -38 -1152
rect -36 -1160 -35 -1152
rect -31 -1160 -30 -1152
rect -28 -1160 -27 -1152
rect 213 -1160 214 -1152
rect 216 -1160 218 -1152
rect 222 -1160 224 -1152
rect 226 -1160 227 -1152
rect 239 -1160 240 -1152
rect 242 -1160 243 -1152
rect 247 -1160 248 -1152
rect 250 -1160 255 -1152
rect 259 -1160 264 -1152
rect 266 -1160 267 -1152
rect 271 -1160 272 -1152
rect 274 -1160 276 -1152
rect 280 -1160 282 -1152
rect 284 -1160 285 -1152
rect 289 -1160 290 -1152
rect 292 -1160 297 -1152
rect 301 -1160 306 -1152
rect 308 -1160 309 -1152
rect 313 -1160 314 -1152
rect 316 -1160 318 -1152
rect 322 -1160 324 -1152
rect 326 -1160 327 -1152
rect 331 -1160 332 -1152
rect 334 -1160 339 -1152
rect 343 -1160 348 -1152
rect 350 -1160 351 -1152
rect 355 -1160 356 -1152
rect 358 -1160 360 -1152
rect 364 -1160 366 -1152
rect 368 -1160 369 -1152
rect 373 -1160 374 -1152
rect 376 -1160 381 -1152
rect 385 -1160 390 -1152
rect 392 -1160 393 -1152
rect 397 -1160 398 -1152
rect 400 -1160 401 -1152
rect 569 -1160 570 -1152
rect 572 -1160 574 -1152
rect 578 -1160 580 -1152
rect 582 -1160 583 -1152
rect 595 -1160 596 -1152
rect 598 -1160 599 -1152
rect 603 -1160 604 -1152
rect 606 -1160 611 -1152
rect 615 -1160 620 -1152
rect 622 -1160 623 -1152
rect 627 -1160 628 -1152
rect 630 -1160 632 -1152
rect 636 -1160 638 -1152
rect 640 -1160 641 -1152
rect 645 -1160 646 -1152
rect 648 -1160 653 -1152
rect 657 -1160 662 -1152
rect 664 -1160 665 -1152
rect 669 -1160 670 -1152
rect 672 -1160 674 -1152
rect 678 -1160 680 -1152
rect 682 -1160 683 -1152
rect 687 -1160 688 -1152
rect 690 -1160 695 -1152
rect 699 -1160 704 -1152
rect 706 -1160 707 -1152
rect 711 -1160 712 -1152
rect 714 -1160 716 -1152
rect 720 -1160 722 -1152
rect 724 -1160 725 -1152
rect 729 -1160 730 -1152
rect 732 -1160 737 -1152
rect 741 -1160 746 -1152
rect 748 -1160 749 -1152
rect 753 -1160 754 -1152
rect 756 -1160 757 -1152
rect 967 -1160 968 -1152
rect 970 -1160 972 -1152
rect 976 -1160 978 -1152
rect 980 -1160 981 -1152
rect 993 -1160 994 -1152
rect 996 -1160 997 -1152
rect 1001 -1160 1002 -1152
rect 1004 -1160 1009 -1152
rect 1013 -1160 1018 -1152
rect 1020 -1160 1021 -1152
rect 1025 -1160 1026 -1152
rect 1028 -1160 1030 -1152
rect 1034 -1160 1036 -1152
rect 1038 -1160 1039 -1152
rect 1043 -1160 1044 -1152
rect 1046 -1160 1051 -1152
rect 1055 -1160 1060 -1152
rect 1062 -1160 1063 -1152
rect 1067 -1160 1068 -1152
rect 1070 -1160 1072 -1152
rect 1076 -1160 1078 -1152
rect 1080 -1160 1081 -1152
rect 1085 -1160 1086 -1152
rect 1088 -1160 1093 -1152
rect 1097 -1160 1102 -1152
rect 1104 -1160 1105 -1152
rect 1109 -1160 1110 -1152
rect 1112 -1160 1114 -1152
rect 1118 -1160 1120 -1152
rect 1122 -1160 1123 -1152
rect 1127 -1160 1128 -1152
rect 1130 -1160 1135 -1152
rect 1139 -1160 1144 -1152
rect 1146 -1160 1147 -1152
rect 1151 -1160 1152 -1152
rect 1154 -1160 1155 -1152
rect -1335 -1276 -1334 -1268
rect -1332 -1276 -1331 -1268
rect -1327 -1276 -1326 -1268
rect -1324 -1276 -1322 -1268
rect -1318 -1276 -1316 -1268
rect -1314 -1276 -1313 -1268
rect -931 -1276 -930 -1268
rect -928 -1276 -927 -1268
rect -923 -1276 -922 -1268
rect -920 -1276 -918 -1268
rect -914 -1276 -912 -1268
rect -910 -1276 -909 -1268
rect -573 -1276 -572 -1268
rect -570 -1276 -569 -1268
rect -565 -1276 -564 -1268
rect -562 -1276 -560 -1268
rect -556 -1276 -554 -1268
rect -552 -1276 -551 -1268
rect -215 -1276 -214 -1268
rect -212 -1276 -211 -1268
rect -207 -1276 -206 -1268
rect -204 -1276 -202 -1268
rect -198 -1276 -196 -1268
rect -194 -1276 -193 -1268
rect 213 -1276 214 -1268
rect 216 -1276 217 -1268
rect 221 -1276 222 -1268
rect 224 -1276 226 -1268
rect 230 -1276 232 -1268
rect 234 -1276 235 -1268
rect 569 -1276 570 -1268
rect 572 -1276 573 -1268
rect 577 -1276 578 -1268
rect 580 -1276 582 -1268
rect 586 -1276 588 -1268
rect 590 -1276 591 -1268
rect 967 -1276 968 -1268
rect 970 -1276 971 -1268
rect 975 -1276 976 -1268
rect 978 -1276 980 -1268
rect 984 -1276 986 -1268
rect 988 -1276 989 -1268
rect 1325 -1276 1326 -1268
rect 1328 -1276 1329 -1268
rect 1333 -1276 1334 -1268
rect 1336 -1276 1338 -1268
rect 1342 -1276 1344 -1268
rect 1346 -1276 1347 -1268
rect -1256 -1390 -1255 -1382
rect -1253 -1390 -1251 -1382
rect -1247 -1390 -1245 -1382
rect -1243 -1390 -1242 -1382
rect -1230 -1390 -1229 -1382
rect -1227 -1390 -1219 -1382
rect -1217 -1390 -1216 -1382
rect -1212 -1390 -1211 -1382
rect -1209 -1390 -1201 -1382
rect -1199 -1390 -1194 -1382
rect -1190 -1390 -1185 -1382
rect -1183 -1390 -1182 -1382
rect -1178 -1390 -1177 -1382
rect -1175 -1390 -1173 -1382
rect -1169 -1390 -1167 -1382
rect -1165 -1390 -1164 -1382
rect -931 -1390 -930 -1382
rect -928 -1390 -926 -1382
rect -922 -1390 -920 -1382
rect -918 -1390 -917 -1382
rect -905 -1390 -904 -1382
rect -902 -1390 -900 -1382
rect -896 -1390 -894 -1382
rect -892 -1390 -891 -1382
rect -879 -1390 -878 -1382
rect -876 -1390 -868 -1382
rect -866 -1390 -865 -1382
rect -861 -1390 -860 -1382
rect -858 -1390 -850 -1382
rect -848 -1390 -843 -1382
rect -839 -1390 -834 -1382
rect -832 -1390 -831 -1382
rect -827 -1390 -826 -1382
rect -824 -1390 -822 -1382
rect -818 -1390 -816 -1382
rect -814 -1390 -813 -1382
rect -801 -1390 -800 -1382
rect -798 -1390 -790 -1382
rect -788 -1390 -787 -1382
rect -783 -1390 -782 -1382
rect -780 -1390 -772 -1382
rect -770 -1390 -765 -1382
rect -761 -1390 -756 -1382
rect -754 -1390 -753 -1382
rect -749 -1390 -748 -1382
rect -746 -1390 -741 -1382
rect -737 -1390 -732 -1382
rect -730 -1390 -729 -1382
rect -717 -1390 -716 -1382
rect -714 -1390 -708 -1382
rect -706 -1390 -704 -1382
rect -700 -1390 -698 -1382
rect -696 -1390 -695 -1382
rect -573 -1390 -572 -1382
rect -570 -1390 -568 -1382
rect -564 -1390 -562 -1382
rect -560 -1390 -559 -1382
rect -547 -1390 -546 -1382
rect -544 -1390 -542 -1382
rect -538 -1390 -536 -1382
rect -534 -1390 -533 -1382
rect -521 -1390 -520 -1382
rect -518 -1390 -510 -1382
rect -508 -1390 -507 -1382
rect -503 -1390 -502 -1382
rect -500 -1390 -492 -1382
rect -490 -1390 -485 -1382
rect -481 -1390 -476 -1382
rect -474 -1390 -473 -1382
rect -469 -1390 -468 -1382
rect -466 -1390 -464 -1382
rect -460 -1390 -458 -1382
rect -456 -1390 -455 -1382
rect -443 -1390 -442 -1382
rect -440 -1390 -432 -1382
rect -430 -1390 -429 -1382
rect -425 -1390 -424 -1382
rect -422 -1390 -414 -1382
rect -412 -1390 -407 -1382
rect -403 -1390 -398 -1382
rect -396 -1390 -395 -1382
rect -391 -1390 -390 -1382
rect -388 -1390 -383 -1382
rect -379 -1390 -374 -1382
rect -372 -1390 -371 -1382
rect -359 -1390 -358 -1382
rect -356 -1390 -350 -1382
rect -348 -1390 -346 -1382
rect -342 -1390 -340 -1382
rect -338 -1390 -337 -1382
rect -215 -1390 -214 -1382
rect -212 -1390 -210 -1382
rect -206 -1390 -204 -1382
rect -202 -1390 -201 -1382
rect -189 -1390 -188 -1382
rect -186 -1390 -184 -1382
rect -180 -1390 -178 -1382
rect -176 -1390 -175 -1382
rect -163 -1390 -162 -1382
rect -160 -1390 -152 -1382
rect -150 -1390 -149 -1382
rect -145 -1390 -144 -1382
rect -142 -1390 -134 -1382
rect -132 -1390 -127 -1382
rect -123 -1390 -118 -1382
rect -116 -1390 -115 -1382
rect -111 -1390 -110 -1382
rect -108 -1390 -106 -1382
rect -102 -1390 -100 -1382
rect -98 -1390 -97 -1382
rect -85 -1390 -84 -1382
rect -82 -1390 -74 -1382
rect -72 -1390 -71 -1382
rect -67 -1390 -66 -1382
rect -64 -1390 -56 -1382
rect -54 -1390 -49 -1382
rect -45 -1390 -40 -1382
rect -38 -1390 -37 -1382
rect -33 -1390 -32 -1382
rect -30 -1390 -25 -1382
rect -21 -1390 -16 -1382
rect -14 -1390 -13 -1382
rect -1 -1390 0 -1382
rect 2 -1390 8 -1382
rect 10 -1390 12 -1382
rect 16 -1390 18 -1382
rect 20 -1390 21 -1382
rect 213 -1390 214 -1382
rect 216 -1390 218 -1382
rect 222 -1390 224 -1382
rect 226 -1390 227 -1382
rect 239 -1390 240 -1382
rect 242 -1390 244 -1382
rect 248 -1390 250 -1382
rect 252 -1390 253 -1382
rect 265 -1390 266 -1382
rect 268 -1390 276 -1382
rect 278 -1390 279 -1382
rect 283 -1390 284 -1382
rect 286 -1390 294 -1382
rect 296 -1390 301 -1382
rect 305 -1390 310 -1382
rect 312 -1390 313 -1382
rect 317 -1390 318 -1382
rect 320 -1390 322 -1382
rect 326 -1390 328 -1382
rect 330 -1390 331 -1382
rect 343 -1390 344 -1382
rect 346 -1390 354 -1382
rect 356 -1390 357 -1382
rect 361 -1390 362 -1382
rect 364 -1390 372 -1382
rect 374 -1390 379 -1382
rect 383 -1390 388 -1382
rect 390 -1390 391 -1382
rect 395 -1390 396 -1382
rect 398 -1390 403 -1382
rect 407 -1390 412 -1382
rect 414 -1390 415 -1382
rect 427 -1390 428 -1382
rect 430 -1390 436 -1382
rect 438 -1390 440 -1382
rect 444 -1390 446 -1382
rect 448 -1390 449 -1382
rect 569 -1390 570 -1382
rect 572 -1390 574 -1382
rect 578 -1390 580 -1382
rect 582 -1390 583 -1382
rect 595 -1390 596 -1382
rect 598 -1390 600 -1382
rect 604 -1390 606 -1382
rect 608 -1390 609 -1382
rect 621 -1390 622 -1382
rect 624 -1390 632 -1382
rect 634 -1390 635 -1382
rect 639 -1390 640 -1382
rect 642 -1390 650 -1382
rect 652 -1390 657 -1382
rect 661 -1390 666 -1382
rect 668 -1390 669 -1382
rect 673 -1390 674 -1382
rect 676 -1390 678 -1382
rect 682 -1390 684 -1382
rect 686 -1390 687 -1382
rect 699 -1390 700 -1382
rect 702 -1390 710 -1382
rect 712 -1390 713 -1382
rect 717 -1390 718 -1382
rect 720 -1390 728 -1382
rect 730 -1390 735 -1382
rect 739 -1390 744 -1382
rect 746 -1390 747 -1382
rect 751 -1390 752 -1382
rect 754 -1390 759 -1382
rect 763 -1390 768 -1382
rect 770 -1390 771 -1382
rect 783 -1390 784 -1382
rect 786 -1390 792 -1382
rect 794 -1390 796 -1382
rect 800 -1390 802 -1382
rect 804 -1390 805 -1382
rect 967 -1390 968 -1382
rect 970 -1390 972 -1382
rect 976 -1390 978 -1382
rect 980 -1390 981 -1382
rect 993 -1390 994 -1382
rect 996 -1390 998 -1382
rect 1002 -1390 1004 -1382
rect 1006 -1390 1007 -1382
rect 1019 -1390 1020 -1382
rect 1022 -1390 1030 -1382
rect 1032 -1390 1033 -1382
rect 1037 -1390 1038 -1382
rect 1040 -1390 1048 -1382
rect 1050 -1390 1055 -1382
rect 1059 -1390 1064 -1382
rect 1066 -1390 1067 -1382
rect 1071 -1390 1072 -1382
rect 1074 -1390 1076 -1382
rect 1080 -1390 1082 -1382
rect 1084 -1390 1085 -1382
rect 1097 -1390 1098 -1382
rect 1100 -1390 1108 -1382
rect 1110 -1390 1111 -1382
rect 1115 -1390 1116 -1382
rect 1118 -1390 1126 -1382
rect 1128 -1390 1133 -1382
rect 1137 -1390 1142 -1382
rect 1144 -1390 1145 -1382
rect 1149 -1390 1150 -1382
rect 1152 -1390 1157 -1382
rect 1161 -1390 1166 -1382
rect 1168 -1390 1169 -1382
rect 1181 -1390 1182 -1382
rect 1184 -1390 1190 -1382
rect 1192 -1390 1194 -1382
rect 1198 -1390 1200 -1382
rect 1202 -1390 1203 -1382
rect 1325 -1390 1326 -1382
rect 1328 -1390 1330 -1382
rect 1334 -1390 1336 -1382
rect 1338 -1390 1339 -1382
rect 1351 -1390 1352 -1382
rect 1354 -1390 1362 -1382
rect 1364 -1390 1365 -1382
rect 1369 -1390 1370 -1382
rect 1372 -1390 1380 -1382
rect 1382 -1390 1387 -1382
rect 1391 -1390 1396 -1382
rect 1398 -1390 1399 -1382
rect 1403 -1390 1404 -1382
rect 1406 -1390 1408 -1382
rect 1412 -1390 1414 -1382
rect 1416 -1390 1417 -1382
rect -1256 -1513 -1255 -1505
rect -1253 -1513 -1251 -1505
rect -1247 -1513 -1245 -1505
rect -1243 -1513 -1242 -1505
rect -1230 -1513 -1229 -1505
rect -1227 -1513 -1226 -1505
rect -1222 -1513 -1221 -1505
rect -1219 -1513 -1214 -1505
rect -1210 -1513 -1205 -1505
rect -1203 -1513 -1202 -1505
rect -1198 -1513 -1197 -1505
rect -1195 -1513 -1193 -1505
rect -1189 -1513 -1187 -1505
rect -1185 -1513 -1184 -1505
rect -1180 -1513 -1179 -1505
rect -1177 -1513 -1172 -1505
rect -1168 -1513 -1163 -1505
rect -1161 -1513 -1160 -1505
rect -1156 -1513 -1155 -1505
rect -1153 -1513 -1151 -1505
rect -1147 -1513 -1145 -1505
rect -1143 -1513 -1142 -1505
rect -1138 -1513 -1137 -1505
rect -1135 -1513 -1130 -1505
rect -1126 -1513 -1121 -1505
rect -1119 -1513 -1118 -1505
rect -1114 -1513 -1113 -1505
rect -1111 -1513 -1109 -1505
rect -1105 -1513 -1103 -1505
rect -1101 -1513 -1100 -1505
rect -1096 -1513 -1095 -1505
rect -1093 -1513 -1088 -1505
rect -1084 -1513 -1079 -1505
rect -1077 -1513 -1076 -1505
rect -1072 -1513 -1071 -1505
rect -1069 -1513 -1068 -1505
rect -931 -1513 -930 -1505
rect -928 -1513 -926 -1505
rect -922 -1513 -920 -1505
rect -918 -1513 -917 -1505
rect -905 -1513 -904 -1505
rect -902 -1513 -901 -1505
rect -897 -1513 -896 -1505
rect -894 -1513 -889 -1505
rect -885 -1513 -880 -1505
rect -878 -1513 -877 -1505
rect -873 -1513 -872 -1505
rect -870 -1513 -868 -1505
rect -864 -1513 -862 -1505
rect -860 -1513 -859 -1505
rect -855 -1513 -854 -1505
rect -852 -1513 -847 -1505
rect -843 -1513 -838 -1505
rect -836 -1513 -835 -1505
rect -831 -1513 -830 -1505
rect -828 -1513 -826 -1505
rect -822 -1513 -820 -1505
rect -818 -1513 -817 -1505
rect -813 -1513 -812 -1505
rect -810 -1513 -805 -1505
rect -801 -1513 -796 -1505
rect -794 -1513 -793 -1505
rect -789 -1513 -788 -1505
rect -786 -1513 -784 -1505
rect -780 -1513 -778 -1505
rect -776 -1513 -775 -1505
rect -771 -1513 -770 -1505
rect -768 -1513 -763 -1505
rect -759 -1513 -754 -1505
rect -752 -1513 -751 -1505
rect -747 -1513 -746 -1505
rect -744 -1513 -743 -1505
rect -573 -1513 -572 -1505
rect -570 -1513 -568 -1505
rect -564 -1513 -562 -1505
rect -560 -1513 -559 -1505
rect -547 -1513 -546 -1505
rect -544 -1513 -543 -1505
rect -539 -1513 -538 -1505
rect -536 -1513 -531 -1505
rect -527 -1513 -522 -1505
rect -520 -1513 -519 -1505
rect -515 -1513 -514 -1505
rect -512 -1513 -510 -1505
rect -506 -1513 -504 -1505
rect -502 -1513 -501 -1505
rect -497 -1513 -496 -1505
rect -494 -1513 -489 -1505
rect -485 -1513 -480 -1505
rect -478 -1513 -477 -1505
rect -473 -1513 -472 -1505
rect -470 -1513 -468 -1505
rect -464 -1513 -462 -1505
rect -460 -1513 -459 -1505
rect -455 -1513 -454 -1505
rect -452 -1513 -447 -1505
rect -443 -1513 -438 -1505
rect -436 -1513 -435 -1505
rect -431 -1513 -430 -1505
rect -428 -1513 -426 -1505
rect -422 -1513 -420 -1505
rect -418 -1513 -417 -1505
rect -413 -1513 -412 -1505
rect -410 -1513 -405 -1505
rect -401 -1513 -396 -1505
rect -394 -1513 -393 -1505
rect -389 -1513 -388 -1505
rect -386 -1513 -385 -1505
rect -215 -1513 -214 -1505
rect -212 -1513 -210 -1505
rect -206 -1513 -204 -1505
rect -202 -1513 -201 -1505
rect -189 -1513 -188 -1505
rect -186 -1513 -185 -1505
rect -181 -1513 -180 -1505
rect -178 -1513 -173 -1505
rect -169 -1513 -164 -1505
rect -162 -1513 -161 -1505
rect -157 -1513 -156 -1505
rect -154 -1513 -152 -1505
rect -148 -1513 -146 -1505
rect -144 -1513 -143 -1505
rect -139 -1513 -138 -1505
rect -136 -1513 -131 -1505
rect -127 -1513 -122 -1505
rect -120 -1513 -119 -1505
rect -115 -1513 -114 -1505
rect -112 -1513 -110 -1505
rect -106 -1513 -104 -1505
rect -102 -1513 -101 -1505
rect -97 -1513 -96 -1505
rect -94 -1513 -89 -1505
rect -85 -1513 -80 -1505
rect -78 -1513 -77 -1505
rect -73 -1513 -72 -1505
rect -70 -1513 -68 -1505
rect -64 -1513 -62 -1505
rect -60 -1513 -59 -1505
rect -55 -1513 -54 -1505
rect -52 -1513 -47 -1505
rect -43 -1513 -38 -1505
rect -36 -1513 -35 -1505
rect -31 -1513 -30 -1505
rect -28 -1513 -27 -1505
rect 213 -1513 214 -1505
rect 216 -1513 218 -1505
rect 222 -1513 224 -1505
rect 226 -1513 227 -1505
rect 239 -1513 240 -1505
rect 242 -1513 243 -1505
rect 247 -1513 248 -1505
rect 250 -1513 255 -1505
rect 259 -1513 264 -1505
rect 266 -1513 267 -1505
rect 271 -1513 272 -1505
rect 274 -1513 276 -1505
rect 280 -1513 282 -1505
rect 284 -1513 285 -1505
rect 289 -1513 290 -1505
rect 292 -1513 297 -1505
rect 301 -1513 306 -1505
rect 308 -1513 309 -1505
rect 313 -1513 314 -1505
rect 316 -1513 318 -1505
rect 322 -1513 324 -1505
rect 326 -1513 327 -1505
rect 331 -1513 332 -1505
rect 334 -1513 339 -1505
rect 343 -1513 348 -1505
rect 350 -1513 351 -1505
rect 355 -1513 356 -1505
rect 358 -1513 360 -1505
rect 364 -1513 366 -1505
rect 368 -1513 369 -1505
rect 373 -1513 374 -1505
rect 376 -1513 381 -1505
rect 385 -1513 390 -1505
rect 392 -1513 393 -1505
rect 397 -1513 398 -1505
rect 400 -1513 401 -1505
rect 569 -1513 570 -1505
rect 572 -1513 574 -1505
rect 578 -1513 580 -1505
rect 582 -1513 583 -1505
rect 595 -1513 596 -1505
rect 598 -1513 599 -1505
rect 603 -1513 604 -1505
rect 606 -1513 611 -1505
rect 615 -1513 620 -1505
rect 622 -1513 623 -1505
rect 627 -1513 628 -1505
rect 630 -1513 632 -1505
rect 636 -1513 638 -1505
rect 640 -1513 641 -1505
rect 645 -1513 646 -1505
rect 648 -1513 653 -1505
rect 657 -1513 662 -1505
rect 664 -1513 665 -1505
rect 669 -1513 670 -1505
rect 672 -1513 674 -1505
rect 678 -1513 680 -1505
rect 682 -1513 683 -1505
rect 687 -1513 688 -1505
rect 690 -1513 695 -1505
rect 699 -1513 704 -1505
rect 706 -1513 707 -1505
rect 711 -1513 712 -1505
rect 714 -1513 716 -1505
rect 720 -1513 722 -1505
rect 724 -1513 725 -1505
rect 729 -1513 730 -1505
rect 732 -1513 737 -1505
rect 741 -1513 746 -1505
rect 748 -1513 749 -1505
rect 753 -1513 754 -1505
rect 756 -1513 757 -1505
rect 967 -1513 968 -1505
rect 970 -1513 972 -1505
rect 976 -1513 978 -1505
rect 980 -1513 981 -1505
rect 993 -1513 994 -1505
rect 996 -1513 997 -1505
rect 1001 -1513 1002 -1505
rect 1004 -1513 1009 -1505
rect 1013 -1513 1018 -1505
rect 1020 -1513 1021 -1505
rect 1025 -1513 1026 -1505
rect 1028 -1513 1030 -1505
rect 1034 -1513 1036 -1505
rect 1038 -1513 1039 -1505
rect 1043 -1513 1044 -1505
rect 1046 -1513 1051 -1505
rect 1055 -1513 1060 -1505
rect 1062 -1513 1063 -1505
rect 1067 -1513 1068 -1505
rect 1070 -1513 1072 -1505
rect 1076 -1513 1078 -1505
rect 1080 -1513 1081 -1505
rect 1085 -1513 1086 -1505
rect 1088 -1513 1093 -1505
rect 1097 -1513 1102 -1505
rect 1104 -1513 1105 -1505
rect 1109 -1513 1110 -1505
rect 1112 -1513 1114 -1505
rect 1118 -1513 1120 -1505
rect 1122 -1513 1123 -1505
rect 1127 -1513 1128 -1505
rect 1130 -1513 1135 -1505
rect 1139 -1513 1144 -1505
rect 1146 -1513 1147 -1505
rect 1151 -1513 1152 -1505
rect 1154 -1513 1155 -1505
rect -1256 -1634 -1255 -1626
rect -1253 -1634 -1251 -1626
rect -1247 -1634 -1245 -1626
rect -1243 -1634 -1242 -1626
rect -1230 -1634 -1229 -1626
rect -1227 -1634 -1226 -1626
rect -1222 -1634 -1221 -1626
rect -1219 -1634 -1214 -1626
rect -1210 -1634 -1205 -1626
rect -1203 -1634 -1202 -1626
rect -1198 -1634 -1197 -1626
rect -1195 -1634 -1193 -1626
rect -1189 -1634 -1187 -1626
rect -1185 -1634 -1184 -1626
rect -1180 -1634 -1179 -1626
rect -1177 -1634 -1172 -1626
rect -1168 -1634 -1163 -1626
rect -1161 -1634 -1160 -1626
rect -1156 -1634 -1155 -1626
rect -1153 -1634 -1151 -1626
rect -1147 -1634 -1145 -1626
rect -1143 -1634 -1142 -1626
rect -1138 -1634 -1137 -1626
rect -1135 -1634 -1130 -1626
rect -1126 -1634 -1121 -1626
rect -1119 -1634 -1118 -1626
rect -1114 -1634 -1113 -1626
rect -1111 -1634 -1109 -1626
rect -1105 -1634 -1103 -1626
rect -1101 -1634 -1100 -1626
rect -1096 -1634 -1095 -1626
rect -1093 -1634 -1088 -1626
rect -1084 -1634 -1079 -1626
rect -1077 -1634 -1076 -1626
rect -1072 -1634 -1071 -1626
rect -1069 -1634 -1068 -1626
rect -931 -1634 -930 -1626
rect -928 -1634 -926 -1626
rect -922 -1634 -920 -1626
rect -918 -1634 -917 -1626
rect -905 -1634 -904 -1626
rect -902 -1634 -901 -1626
rect -897 -1634 -896 -1626
rect -894 -1634 -889 -1626
rect -885 -1634 -880 -1626
rect -878 -1634 -877 -1626
rect -873 -1634 -872 -1626
rect -870 -1634 -868 -1626
rect -864 -1634 -862 -1626
rect -860 -1634 -859 -1626
rect -855 -1634 -854 -1626
rect -852 -1634 -847 -1626
rect -843 -1634 -838 -1626
rect -836 -1634 -835 -1626
rect -831 -1634 -830 -1626
rect -828 -1634 -826 -1626
rect -822 -1634 -820 -1626
rect -818 -1634 -817 -1626
rect -813 -1634 -812 -1626
rect -810 -1634 -805 -1626
rect -801 -1634 -796 -1626
rect -794 -1634 -793 -1626
rect -789 -1634 -788 -1626
rect -786 -1634 -784 -1626
rect -780 -1634 -778 -1626
rect -776 -1634 -775 -1626
rect -771 -1634 -770 -1626
rect -768 -1634 -763 -1626
rect -759 -1634 -754 -1626
rect -752 -1634 -751 -1626
rect -747 -1634 -746 -1626
rect -744 -1634 -743 -1626
rect -573 -1634 -572 -1626
rect -570 -1634 -568 -1626
rect -564 -1634 -562 -1626
rect -560 -1634 -559 -1626
rect -547 -1634 -546 -1626
rect -544 -1634 -543 -1626
rect -539 -1634 -538 -1626
rect -536 -1634 -531 -1626
rect -527 -1634 -522 -1626
rect -520 -1634 -519 -1626
rect -515 -1634 -514 -1626
rect -512 -1634 -510 -1626
rect -506 -1634 -504 -1626
rect -502 -1634 -501 -1626
rect -497 -1634 -496 -1626
rect -494 -1634 -489 -1626
rect -485 -1634 -480 -1626
rect -478 -1634 -477 -1626
rect -473 -1634 -472 -1626
rect -470 -1634 -468 -1626
rect -464 -1634 -462 -1626
rect -460 -1634 -459 -1626
rect -455 -1634 -454 -1626
rect -452 -1634 -447 -1626
rect -443 -1634 -438 -1626
rect -436 -1634 -435 -1626
rect -431 -1634 -430 -1626
rect -428 -1634 -426 -1626
rect -422 -1634 -420 -1626
rect -418 -1634 -417 -1626
rect -413 -1634 -412 -1626
rect -410 -1634 -405 -1626
rect -401 -1634 -396 -1626
rect -394 -1634 -393 -1626
rect -389 -1634 -388 -1626
rect -386 -1634 -385 -1626
rect -215 -1634 -214 -1626
rect -212 -1634 -210 -1626
rect -206 -1634 -204 -1626
rect -202 -1634 -201 -1626
rect -189 -1634 -188 -1626
rect -186 -1634 -185 -1626
rect -181 -1634 -180 -1626
rect -178 -1634 -173 -1626
rect -169 -1634 -164 -1626
rect -162 -1634 -161 -1626
rect -157 -1634 -156 -1626
rect -154 -1634 -152 -1626
rect -148 -1634 -146 -1626
rect -144 -1634 -143 -1626
rect -139 -1634 -138 -1626
rect -136 -1634 -131 -1626
rect -127 -1634 -122 -1626
rect -120 -1634 -119 -1626
rect -115 -1634 -114 -1626
rect -112 -1634 -110 -1626
rect -106 -1634 -104 -1626
rect -102 -1634 -101 -1626
rect -97 -1634 -96 -1626
rect -94 -1634 -89 -1626
rect -85 -1634 -80 -1626
rect -78 -1634 -77 -1626
rect -73 -1634 -72 -1626
rect -70 -1634 -68 -1626
rect -64 -1634 -62 -1626
rect -60 -1634 -59 -1626
rect -55 -1634 -54 -1626
rect -52 -1634 -47 -1626
rect -43 -1634 -38 -1626
rect -36 -1634 -35 -1626
rect -31 -1634 -30 -1626
rect -28 -1634 -27 -1626
rect 213 -1634 214 -1626
rect 216 -1634 218 -1626
rect 222 -1634 224 -1626
rect 226 -1634 227 -1626
rect 239 -1634 240 -1626
rect 242 -1634 243 -1626
rect 247 -1634 248 -1626
rect 250 -1634 255 -1626
rect 259 -1634 264 -1626
rect 266 -1634 267 -1626
rect 271 -1634 272 -1626
rect 274 -1634 276 -1626
rect 280 -1634 282 -1626
rect 284 -1634 285 -1626
rect 289 -1634 290 -1626
rect 292 -1634 297 -1626
rect 301 -1634 306 -1626
rect 308 -1634 309 -1626
rect 313 -1634 314 -1626
rect 316 -1634 318 -1626
rect 322 -1634 324 -1626
rect 326 -1634 327 -1626
rect 331 -1634 332 -1626
rect 334 -1634 339 -1626
rect 343 -1634 348 -1626
rect 350 -1634 351 -1626
rect 355 -1634 356 -1626
rect 358 -1634 360 -1626
rect 364 -1634 366 -1626
rect 368 -1634 369 -1626
rect 373 -1634 374 -1626
rect 376 -1634 381 -1626
rect 385 -1634 390 -1626
rect 392 -1634 393 -1626
rect 397 -1634 398 -1626
rect 400 -1634 401 -1626
rect 569 -1634 570 -1626
rect 572 -1634 574 -1626
rect 578 -1634 580 -1626
rect 582 -1634 583 -1626
rect 595 -1634 596 -1626
rect 598 -1634 599 -1626
rect 603 -1634 604 -1626
rect 606 -1634 611 -1626
rect 615 -1634 620 -1626
rect 622 -1634 623 -1626
rect 627 -1634 628 -1626
rect 630 -1634 632 -1626
rect 636 -1634 638 -1626
rect 640 -1634 641 -1626
rect 645 -1634 646 -1626
rect 648 -1634 653 -1626
rect 657 -1634 662 -1626
rect 664 -1634 665 -1626
rect 669 -1634 670 -1626
rect 672 -1634 674 -1626
rect 678 -1634 680 -1626
rect 682 -1634 683 -1626
rect 687 -1634 688 -1626
rect 690 -1634 695 -1626
rect 699 -1634 704 -1626
rect 706 -1634 707 -1626
rect 711 -1634 712 -1626
rect 714 -1634 716 -1626
rect 720 -1634 722 -1626
rect 724 -1634 725 -1626
rect 729 -1634 730 -1626
rect 732 -1634 737 -1626
rect 741 -1634 746 -1626
rect 748 -1634 749 -1626
rect 753 -1634 754 -1626
rect 756 -1634 757 -1626
rect 967 -1634 968 -1626
rect 970 -1634 972 -1626
rect 976 -1634 978 -1626
rect 980 -1634 981 -1626
rect 993 -1634 994 -1626
rect 996 -1634 997 -1626
rect 1001 -1634 1002 -1626
rect 1004 -1634 1009 -1626
rect 1013 -1634 1018 -1626
rect 1020 -1634 1021 -1626
rect 1025 -1634 1026 -1626
rect 1028 -1634 1030 -1626
rect 1034 -1634 1036 -1626
rect 1038 -1634 1039 -1626
rect 1043 -1634 1044 -1626
rect 1046 -1634 1051 -1626
rect 1055 -1634 1060 -1626
rect 1062 -1634 1063 -1626
rect 1067 -1634 1068 -1626
rect 1070 -1634 1072 -1626
rect 1076 -1634 1078 -1626
rect 1080 -1634 1081 -1626
rect 1085 -1634 1086 -1626
rect 1088 -1634 1093 -1626
rect 1097 -1634 1102 -1626
rect 1104 -1634 1105 -1626
rect 1109 -1634 1110 -1626
rect 1112 -1634 1114 -1626
rect 1118 -1634 1120 -1626
rect 1122 -1634 1123 -1626
rect 1127 -1634 1128 -1626
rect 1130 -1634 1135 -1626
rect 1139 -1634 1144 -1626
rect 1146 -1634 1147 -1626
rect 1151 -1634 1152 -1626
rect 1154 -1634 1155 -1626
rect 1325 -1634 1326 -1626
rect 1328 -1634 1330 -1626
rect 1334 -1634 1336 -1626
rect 1338 -1634 1339 -1626
rect 1351 -1634 1352 -1626
rect 1354 -1634 1355 -1626
rect 1359 -1634 1360 -1626
rect 1362 -1634 1367 -1626
rect 1371 -1634 1376 -1626
rect 1378 -1634 1379 -1626
rect 1383 -1634 1384 -1626
rect 1386 -1634 1388 -1626
rect 1392 -1634 1394 -1626
rect 1396 -1634 1397 -1626
rect 1401 -1634 1402 -1626
rect 1404 -1634 1409 -1626
rect 1413 -1634 1418 -1626
rect 1420 -1634 1421 -1626
rect 1425 -1634 1426 -1626
rect 1428 -1634 1430 -1626
rect 1434 -1634 1436 -1626
rect 1438 -1634 1439 -1626
rect 1443 -1634 1444 -1626
rect 1446 -1634 1451 -1626
rect 1455 -1634 1460 -1626
rect 1462 -1634 1463 -1626
rect 1467 -1634 1468 -1626
rect 1470 -1634 1472 -1626
rect 1476 -1634 1478 -1626
rect 1480 -1634 1481 -1626
rect 1485 -1634 1486 -1626
rect 1488 -1634 1493 -1626
rect 1497 -1634 1502 -1626
rect 1504 -1634 1505 -1626
rect 1509 -1634 1510 -1626
rect 1512 -1634 1513 -1626
rect -1256 -1755 -1255 -1747
rect -1253 -1755 -1251 -1747
rect -1247 -1755 -1245 -1747
rect -1243 -1755 -1242 -1747
rect -1230 -1755 -1229 -1747
rect -1227 -1755 -1226 -1747
rect -1222 -1755 -1221 -1747
rect -1219 -1755 -1214 -1747
rect -1210 -1755 -1205 -1747
rect -1203 -1755 -1202 -1747
rect -1198 -1755 -1197 -1747
rect -1195 -1755 -1193 -1747
rect -1189 -1755 -1187 -1747
rect -1185 -1755 -1184 -1747
rect -1180 -1755 -1179 -1747
rect -1177 -1755 -1172 -1747
rect -1168 -1755 -1163 -1747
rect -1161 -1755 -1160 -1747
rect -1156 -1755 -1155 -1747
rect -1153 -1755 -1151 -1747
rect -1147 -1755 -1145 -1747
rect -1143 -1755 -1142 -1747
rect -1138 -1755 -1137 -1747
rect -1135 -1755 -1130 -1747
rect -1126 -1755 -1121 -1747
rect -1119 -1755 -1118 -1747
rect -1114 -1755 -1113 -1747
rect -1111 -1755 -1109 -1747
rect -1105 -1755 -1103 -1747
rect -1101 -1755 -1100 -1747
rect -1096 -1755 -1095 -1747
rect -1093 -1755 -1088 -1747
rect -1084 -1755 -1079 -1747
rect -1077 -1755 -1076 -1747
rect -1072 -1755 -1071 -1747
rect -1069 -1755 -1068 -1747
rect -1025 -1755 -1024 -1747
rect -1022 -1755 -1021 -1747
rect -931 -1755 -930 -1747
rect -928 -1755 -926 -1747
rect -922 -1755 -920 -1747
rect -918 -1755 -917 -1747
rect -905 -1755 -904 -1747
rect -902 -1755 -901 -1747
rect -897 -1755 -896 -1747
rect -894 -1755 -889 -1747
rect -885 -1755 -880 -1747
rect -878 -1755 -877 -1747
rect -873 -1755 -872 -1747
rect -870 -1755 -868 -1747
rect -864 -1755 -862 -1747
rect -860 -1755 -859 -1747
rect -855 -1755 -854 -1747
rect -852 -1755 -847 -1747
rect -843 -1755 -838 -1747
rect -836 -1755 -835 -1747
rect -831 -1755 -830 -1747
rect -828 -1755 -826 -1747
rect -822 -1755 -820 -1747
rect -818 -1755 -817 -1747
rect -813 -1755 -812 -1747
rect -810 -1755 -805 -1747
rect -801 -1755 -796 -1747
rect -794 -1755 -793 -1747
rect -789 -1755 -788 -1747
rect -786 -1755 -784 -1747
rect -780 -1755 -778 -1747
rect -776 -1755 -775 -1747
rect -771 -1755 -770 -1747
rect -768 -1755 -763 -1747
rect -759 -1755 -754 -1747
rect -752 -1755 -751 -1747
rect -747 -1755 -746 -1747
rect -744 -1755 -743 -1747
rect -573 -1755 -572 -1747
rect -570 -1755 -568 -1747
rect -564 -1755 -562 -1747
rect -560 -1755 -559 -1747
rect -547 -1755 -546 -1747
rect -544 -1755 -543 -1747
rect -539 -1755 -538 -1747
rect -536 -1755 -531 -1747
rect -527 -1755 -522 -1747
rect -520 -1755 -519 -1747
rect -515 -1755 -514 -1747
rect -512 -1755 -510 -1747
rect -506 -1755 -504 -1747
rect -502 -1755 -501 -1747
rect -497 -1755 -496 -1747
rect -494 -1755 -489 -1747
rect -485 -1755 -480 -1747
rect -478 -1755 -477 -1747
rect -473 -1755 -472 -1747
rect -470 -1755 -468 -1747
rect -464 -1755 -462 -1747
rect -460 -1755 -459 -1747
rect -455 -1755 -454 -1747
rect -452 -1755 -447 -1747
rect -443 -1755 -438 -1747
rect -436 -1755 -435 -1747
rect -431 -1755 -430 -1747
rect -428 -1755 -426 -1747
rect -422 -1755 -420 -1747
rect -418 -1755 -417 -1747
rect -413 -1755 -412 -1747
rect -410 -1755 -405 -1747
rect -401 -1755 -396 -1747
rect -394 -1755 -393 -1747
rect -389 -1755 -388 -1747
rect -386 -1755 -385 -1747
rect -328 -1755 -327 -1747
rect -325 -1755 -324 -1747
rect -215 -1755 -214 -1747
rect -212 -1755 -210 -1747
rect -206 -1755 -204 -1747
rect -202 -1755 -201 -1747
rect -189 -1755 -188 -1747
rect -186 -1755 -185 -1747
rect -181 -1755 -180 -1747
rect -178 -1755 -173 -1747
rect -169 -1755 -164 -1747
rect -162 -1755 -161 -1747
rect -157 -1755 -156 -1747
rect -154 -1755 -152 -1747
rect -148 -1755 -146 -1747
rect -144 -1755 -143 -1747
rect -139 -1755 -138 -1747
rect -136 -1755 -131 -1747
rect -127 -1755 -122 -1747
rect -120 -1755 -119 -1747
rect -115 -1755 -114 -1747
rect -112 -1755 -110 -1747
rect -106 -1755 -104 -1747
rect -102 -1755 -101 -1747
rect -97 -1755 -96 -1747
rect -94 -1755 -89 -1747
rect -85 -1755 -80 -1747
rect -78 -1755 -77 -1747
rect -73 -1755 -72 -1747
rect -70 -1755 -68 -1747
rect -64 -1755 -62 -1747
rect -60 -1755 -59 -1747
rect -55 -1755 -54 -1747
rect -52 -1755 -47 -1747
rect -43 -1755 -38 -1747
rect -36 -1755 -35 -1747
rect -31 -1755 -30 -1747
rect -28 -1755 -27 -1747
rect 213 -1755 214 -1747
rect 216 -1755 218 -1747
rect 222 -1755 224 -1747
rect 226 -1755 227 -1747
rect 239 -1755 240 -1747
rect 242 -1755 243 -1747
rect 247 -1755 248 -1747
rect 250 -1755 255 -1747
rect 259 -1755 264 -1747
rect 266 -1755 267 -1747
rect 271 -1755 272 -1747
rect 274 -1755 276 -1747
rect 280 -1755 282 -1747
rect 284 -1755 285 -1747
rect 289 -1755 290 -1747
rect 292 -1755 297 -1747
rect 301 -1755 306 -1747
rect 308 -1755 309 -1747
rect 313 -1755 314 -1747
rect 316 -1755 318 -1747
rect 322 -1755 324 -1747
rect 326 -1755 327 -1747
rect 331 -1755 332 -1747
rect 334 -1755 339 -1747
rect 343 -1755 348 -1747
rect 350 -1755 351 -1747
rect 355 -1755 356 -1747
rect 358 -1755 360 -1747
rect 364 -1755 366 -1747
rect 368 -1755 369 -1747
rect 373 -1755 374 -1747
rect 376 -1755 381 -1747
rect 385 -1755 390 -1747
rect 392 -1755 393 -1747
rect 397 -1755 398 -1747
rect 400 -1755 401 -1747
rect 468 -1755 469 -1747
rect 471 -1755 472 -1747
rect 569 -1755 570 -1747
rect 572 -1755 574 -1747
rect 578 -1755 580 -1747
rect 582 -1755 583 -1747
rect 595 -1755 596 -1747
rect 598 -1755 599 -1747
rect 603 -1755 604 -1747
rect 606 -1755 611 -1747
rect 615 -1755 620 -1747
rect 622 -1755 623 -1747
rect 627 -1755 628 -1747
rect 630 -1755 632 -1747
rect 636 -1755 638 -1747
rect 640 -1755 641 -1747
rect 645 -1755 646 -1747
rect 648 -1755 653 -1747
rect 657 -1755 662 -1747
rect 664 -1755 665 -1747
rect 669 -1755 670 -1747
rect 672 -1755 674 -1747
rect 678 -1755 680 -1747
rect 682 -1755 683 -1747
rect 687 -1755 688 -1747
rect 690 -1755 695 -1747
rect 699 -1755 704 -1747
rect 706 -1755 707 -1747
rect 711 -1755 712 -1747
rect 714 -1755 716 -1747
rect 720 -1755 722 -1747
rect 724 -1755 725 -1747
rect 729 -1755 730 -1747
rect 732 -1755 737 -1747
rect 741 -1755 746 -1747
rect 748 -1755 749 -1747
rect 753 -1755 754 -1747
rect 756 -1755 757 -1747
rect 967 -1755 968 -1747
rect 970 -1755 972 -1747
rect 976 -1755 978 -1747
rect 980 -1755 981 -1747
rect 993 -1755 994 -1747
rect 996 -1755 997 -1747
rect 1001 -1755 1002 -1747
rect 1004 -1755 1009 -1747
rect 1013 -1755 1018 -1747
rect 1020 -1755 1021 -1747
rect 1025 -1755 1026 -1747
rect 1028 -1755 1030 -1747
rect 1034 -1755 1036 -1747
rect 1038 -1755 1039 -1747
rect 1043 -1755 1044 -1747
rect 1046 -1755 1051 -1747
rect 1055 -1755 1060 -1747
rect 1062 -1755 1063 -1747
rect 1067 -1755 1068 -1747
rect 1070 -1755 1072 -1747
rect 1076 -1755 1078 -1747
rect 1080 -1755 1081 -1747
rect 1085 -1755 1086 -1747
rect 1088 -1755 1093 -1747
rect 1097 -1755 1102 -1747
rect 1104 -1755 1105 -1747
rect 1109 -1755 1110 -1747
rect 1112 -1755 1114 -1747
rect 1118 -1755 1120 -1747
rect 1122 -1755 1123 -1747
rect 1127 -1755 1128 -1747
rect 1130 -1755 1135 -1747
rect 1139 -1755 1144 -1747
rect 1146 -1755 1147 -1747
rect 1151 -1755 1152 -1747
rect 1154 -1755 1155 -1747
rect 1207 -1755 1208 -1747
rect 1210 -1755 1211 -1747
rect 1325 -1755 1326 -1747
rect 1328 -1755 1330 -1747
rect 1334 -1755 1336 -1747
rect 1338 -1755 1339 -1747
rect 1351 -1755 1352 -1747
rect 1354 -1755 1355 -1747
rect 1359 -1755 1360 -1747
rect 1362 -1755 1367 -1747
rect 1371 -1755 1376 -1747
rect 1378 -1755 1379 -1747
rect 1383 -1755 1384 -1747
rect 1386 -1755 1388 -1747
rect 1392 -1755 1394 -1747
rect 1396 -1755 1397 -1747
rect 1401 -1755 1402 -1747
rect 1404 -1755 1409 -1747
rect 1413 -1755 1418 -1747
rect 1420 -1755 1421 -1747
rect 1425 -1755 1426 -1747
rect 1428 -1755 1430 -1747
rect 1434 -1755 1436 -1747
rect 1438 -1755 1439 -1747
rect 1443 -1755 1444 -1747
rect 1446 -1755 1451 -1747
rect 1455 -1755 1460 -1747
rect 1462 -1755 1463 -1747
rect 1467 -1755 1468 -1747
rect 1470 -1755 1472 -1747
rect 1476 -1755 1478 -1747
rect 1480 -1755 1481 -1747
rect 1485 -1755 1486 -1747
rect 1488 -1755 1493 -1747
rect 1497 -1755 1502 -1747
rect 1504 -1755 1505 -1747
rect 1509 -1755 1510 -1747
rect 1512 -1755 1513 -1747
rect -1256 -1870 -1255 -1862
rect -1253 -1870 -1251 -1862
rect -1247 -1870 -1245 -1862
rect -1243 -1870 -1242 -1862
rect -1230 -1870 -1229 -1862
rect -1227 -1870 -1226 -1862
rect -1222 -1870 -1221 -1862
rect -1219 -1870 -1214 -1862
rect -1210 -1870 -1205 -1862
rect -1203 -1870 -1202 -1862
rect -1198 -1870 -1197 -1862
rect -1195 -1870 -1193 -1862
rect -1189 -1870 -1187 -1862
rect -1185 -1870 -1184 -1862
rect -1180 -1870 -1179 -1862
rect -1177 -1870 -1172 -1862
rect -1168 -1870 -1163 -1862
rect -1161 -1870 -1160 -1862
rect -1156 -1870 -1155 -1862
rect -1153 -1870 -1151 -1862
rect -1147 -1870 -1145 -1862
rect -1143 -1870 -1142 -1862
rect -1138 -1870 -1137 -1862
rect -1135 -1870 -1130 -1862
rect -1126 -1870 -1121 -1862
rect -1119 -1870 -1118 -1862
rect -1114 -1870 -1113 -1862
rect -1111 -1870 -1109 -1862
rect -1105 -1870 -1103 -1862
rect -1101 -1870 -1100 -1862
rect -1096 -1870 -1095 -1862
rect -1093 -1870 -1088 -1862
rect -1084 -1870 -1079 -1862
rect -1077 -1870 -1076 -1862
rect -1072 -1870 -1071 -1862
rect -1069 -1870 -1068 -1862
rect -1025 -1870 -1024 -1862
rect -1022 -1870 -1021 -1862
rect -669 -1878 -668 -1862
rect -666 -1878 -665 -1862
rect -328 -1870 -327 -1862
rect -325 -1870 -324 -1862
rect 468 -1870 469 -1862
rect 471 -1870 472 -1862
rect 845 -1878 846 -1862
rect 848 -1878 849 -1862
rect 1207 -1870 1208 -1862
rect 1210 -1870 1211 -1862
rect -1335 -1982 -1334 -1974
rect -1332 -1982 -1331 -1974
rect -1327 -1982 -1326 -1974
rect -1324 -1982 -1322 -1974
rect -1318 -1982 -1316 -1974
rect -1314 -1982 -1313 -1974
rect -931 -1982 -930 -1974
rect -928 -1982 -927 -1974
rect -923 -1982 -922 -1974
rect -920 -1982 -918 -1974
rect -914 -1982 -912 -1974
rect -910 -1982 -909 -1974
rect -573 -1982 -572 -1974
rect -570 -1982 -569 -1974
rect -565 -1982 -564 -1974
rect -562 -1982 -560 -1974
rect -556 -1982 -554 -1974
rect -552 -1982 -551 -1974
rect -215 -1982 -214 -1974
rect -212 -1982 -211 -1974
rect -207 -1982 -206 -1974
rect -204 -1982 -202 -1974
rect -198 -1982 -196 -1974
rect -194 -1982 -193 -1974
rect 213 -1982 214 -1974
rect 216 -1982 217 -1974
rect 221 -1982 222 -1974
rect 224 -1982 226 -1974
rect 230 -1982 232 -1974
rect 234 -1982 235 -1974
rect 569 -1982 570 -1974
rect 572 -1982 573 -1974
rect 577 -1982 578 -1974
rect 580 -1982 582 -1974
rect 586 -1982 588 -1974
rect 590 -1982 591 -1974
rect 967 -1982 968 -1974
rect 970 -1982 971 -1974
rect 975 -1982 976 -1974
rect 978 -1982 980 -1974
rect 984 -1982 986 -1974
rect 988 -1982 989 -1974
rect 1325 -1982 1326 -1974
rect 1328 -1982 1329 -1974
rect 1333 -1982 1334 -1974
rect 1336 -1982 1338 -1974
rect 1342 -1982 1344 -1974
rect 1346 -1982 1347 -1974
rect -1256 -2101 -1255 -2093
rect -1253 -2101 -1251 -2093
rect -1247 -2101 -1245 -2093
rect -1243 -2101 -1242 -2093
rect -1230 -2101 -1229 -2093
rect -1227 -2101 -1219 -2093
rect -1217 -2101 -1216 -2093
rect -1212 -2101 -1211 -2093
rect -1209 -2101 -1201 -2093
rect -1199 -2101 -1194 -2093
rect -1190 -2101 -1185 -2093
rect -1183 -2101 -1182 -2093
rect -1178 -2101 -1177 -2093
rect -1175 -2101 -1173 -2093
rect -1169 -2101 -1167 -2093
rect -1165 -2101 -1164 -2093
rect -931 -2101 -930 -2093
rect -928 -2101 -926 -2093
rect -922 -2101 -920 -2093
rect -918 -2101 -917 -2093
rect -905 -2101 -904 -2093
rect -902 -2101 -900 -2093
rect -896 -2101 -894 -2093
rect -892 -2101 -891 -2093
rect -879 -2101 -878 -2093
rect -876 -2101 -868 -2093
rect -866 -2101 -865 -2093
rect -861 -2101 -860 -2093
rect -858 -2101 -850 -2093
rect -848 -2101 -843 -2093
rect -839 -2101 -834 -2093
rect -832 -2101 -831 -2093
rect -827 -2101 -826 -2093
rect -824 -2101 -822 -2093
rect -818 -2101 -816 -2093
rect -814 -2101 -813 -2093
rect -801 -2101 -800 -2093
rect -798 -2101 -790 -2093
rect -788 -2101 -787 -2093
rect -783 -2101 -782 -2093
rect -780 -2101 -772 -2093
rect -770 -2101 -765 -2093
rect -761 -2101 -756 -2093
rect -754 -2101 -753 -2093
rect -749 -2101 -748 -2093
rect -746 -2101 -741 -2093
rect -737 -2101 -732 -2093
rect -730 -2101 -729 -2093
rect -717 -2101 -716 -2093
rect -714 -2101 -708 -2093
rect -706 -2101 -704 -2093
rect -700 -2101 -698 -2093
rect -696 -2101 -695 -2093
rect -573 -2101 -572 -2093
rect -570 -2101 -568 -2093
rect -564 -2101 -562 -2093
rect -560 -2101 -559 -2093
rect -547 -2101 -546 -2093
rect -544 -2101 -542 -2093
rect -538 -2101 -536 -2093
rect -534 -2101 -533 -2093
rect -521 -2101 -520 -2093
rect -518 -2101 -510 -2093
rect -508 -2101 -507 -2093
rect -503 -2101 -502 -2093
rect -500 -2101 -492 -2093
rect -490 -2101 -485 -2093
rect -481 -2101 -476 -2093
rect -474 -2101 -473 -2093
rect -469 -2101 -468 -2093
rect -466 -2101 -464 -2093
rect -460 -2101 -458 -2093
rect -456 -2101 -455 -2093
rect -443 -2101 -442 -2093
rect -440 -2101 -432 -2093
rect -430 -2101 -429 -2093
rect -425 -2101 -424 -2093
rect -422 -2101 -414 -2093
rect -412 -2101 -407 -2093
rect -403 -2101 -398 -2093
rect -396 -2101 -395 -2093
rect -391 -2101 -390 -2093
rect -388 -2101 -383 -2093
rect -379 -2101 -374 -2093
rect -372 -2101 -371 -2093
rect -359 -2101 -358 -2093
rect -356 -2101 -350 -2093
rect -348 -2101 -346 -2093
rect -342 -2101 -340 -2093
rect -338 -2101 -337 -2093
rect -215 -2101 -214 -2093
rect -212 -2101 -210 -2093
rect -206 -2101 -204 -2093
rect -202 -2101 -201 -2093
rect -189 -2101 -188 -2093
rect -186 -2101 -184 -2093
rect -180 -2101 -178 -2093
rect -176 -2101 -175 -2093
rect -163 -2101 -162 -2093
rect -160 -2101 -152 -2093
rect -150 -2101 -149 -2093
rect -145 -2101 -144 -2093
rect -142 -2101 -134 -2093
rect -132 -2101 -127 -2093
rect -123 -2101 -118 -2093
rect -116 -2101 -115 -2093
rect -111 -2101 -110 -2093
rect -108 -2101 -106 -2093
rect -102 -2101 -100 -2093
rect -98 -2101 -97 -2093
rect -85 -2101 -84 -2093
rect -82 -2101 -74 -2093
rect -72 -2101 -71 -2093
rect -67 -2101 -66 -2093
rect -64 -2101 -56 -2093
rect -54 -2101 -49 -2093
rect -45 -2101 -40 -2093
rect -38 -2101 -37 -2093
rect -33 -2101 -32 -2093
rect -30 -2101 -25 -2093
rect -21 -2101 -16 -2093
rect -14 -2101 -13 -2093
rect -1 -2101 0 -2093
rect 2 -2101 8 -2093
rect 10 -2101 12 -2093
rect 16 -2101 18 -2093
rect 20 -2101 21 -2093
rect 213 -2101 214 -2093
rect 216 -2101 218 -2093
rect 222 -2101 224 -2093
rect 226 -2101 227 -2093
rect 239 -2101 240 -2093
rect 242 -2101 244 -2093
rect 248 -2101 250 -2093
rect 252 -2101 253 -2093
rect 265 -2101 266 -2093
rect 268 -2101 276 -2093
rect 278 -2101 279 -2093
rect 283 -2101 284 -2093
rect 286 -2101 294 -2093
rect 296 -2101 301 -2093
rect 305 -2101 310 -2093
rect 312 -2101 313 -2093
rect 317 -2101 318 -2093
rect 320 -2101 322 -2093
rect 326 -2101 328 -2093
rect 330 -2101 331 -2093
rect 343 -2101 344 -2093
rect 346 -2101 354 -2093
rect 356 -2101 357 -2093
rect 361 -2101 362 -2093
rect 364 -2101 372 -2093
rect 374 -2101 379 -2093
rect 383 -2101 388 -2093
rect 390 -2101 391 -2093
rect 395 -2101 396 -2093
rect 398 -2101 403 -2093
rect 407 -2101 412 -2093
rect 414 -2101 415 -2093
rect 427 -2101 428 -2093
rect 430 -2101 436 -2093
rect 438 -2101 440 -2093
rect 444 -2101 446 -2093
rect 448 -2101 449 -2093
rect 569 -2101 570 -2093
rect 572 -2101 574 -2093
rect 578 -2101 580 -2093
rect 582 -2101 583 -2093
rect 595 -2101 596 -2093
rect 598 -2101 600 -2093
rect 604 -2101 606 -2093
rect 608 -2101 609 -2093
rect 621 -2101 622 -2093
rect 624 -2101 632 -2093
rect 634 -2101 635 -2093
rect 639 -2101 640 -2093
rect 642 -2101 650 -2093
rect 652 -2101 657 -2093
rect 661 -2101 666 -2093
rect 668 -2101 669 -2093
rect 673 -2101 674 -2093
rect 676 -2101 678 -2093
rect 682 -2101 684 -2093
rect 686 -2101 687 -2093
rect 699 -2101 700 -2093
rect 702 -2101 710 -2093
rect 712 -2101 713 -2093
rect 717 -2101 718 -2093
rect 720 -2101 728 -2093
rect 730 -2101 735 -2093
rect 739 -2101 744 -2093
rect 746 -2101 747 -2093
rect 751 -2101 752 -2093
rect 754 -2101 759 -2093
rect 763 -2101 768 -2093
rect 770 -2101 771 -2093
rect 783 -2101 784 -2093
rect 786 -2101 792 -2093
rect 794 -2101 796 -2093
rect 800 -2101 802 -2093
rect 804 -2101 805 -2093
rect 967 -2101 968 -2093
rect 970 -2101 972 -2093
rect 976 -2101 978 -2093
rect 980 -2101 981 -2093
rect 993 -2101 994 -2093
rect 996 -2101 998 -2093
rect 1002 -2101 1004 -2093
rect 1006 -2101 1007 -2093
rect 1019 -2101 1020 -2093
rect 1022 -2101 1030 -2093
rect 1032 -2101 1033 -2093
rect 1037 -2101 1038 -2093
rect 1040 -2101 1048 -2093
rect 1050 -2101 1055 -2093
rect 1059 -2101 1064 -2093
rect 1066 -2101 1067 -2093
rect 1071 -2101 1072 -2093
rect 1074 -2101 1076 -2093
rect 1080 -2101 1082 -2093
rect 1084 -2101 1085 -2093
rect 1097 -2101 1098 -2093
rect 1100 -2101 1108 -2093
rect 1110 -2101 1111 -2093
rect 1115 -2101 1116 -2093
rect 1118 -2101 1126 -2093
rect 1128 -2101 1133 -2093
rect 1137 -2101 1142 -2093
rect 1144 -2101 1145 -2093
rect 1149 -2101 1150 -2093
rect 1152 -2101 1157 -2093
rect 1161 -2101 1166 -2093
rect 1168 -2101 1169 -2093
rect 1181 -2101 1182 -2093
rect 1184 -2101 1190 -2093
rect 1192 -2101 1194 -2093
rect 1198 -2101 1200 -2093
rect 1202 -2101 1203 -2093
rect 1325 -2101 1326 -2093
rect 1328 -2101 1330 -2093
rect 1334 -2101 1336 -2093
rect 1338 -2101 1339 -2093
rect 1351 -2101 1352 -2093
rect 1354 -2101 1356 -2093
rect 1360 -2101 1362 -2093
rect 1364 -2101 1365 -2093
rect 1377 -2101 1378 -2093
rect 1380 -2101 1388 -2093
rect 1390 -2101 1391 -2093
rect 1395 -2101 1396 -2093
rect 1398 -2101 1406 -2093
rect 1408 -2101 1413 -2093
rect 1417 -2101 1422 -2093
rect 1424 -2101 1425 -2093
rect 1429 -2101 1430 -2093
rect 1432 -2101 1434 -2093
rect 1438 -2101 1440 -2093
rect 1442 -2101 1443 -2093
rect 1455 -2101 1456 -2093
rect 1458 -2101 1466 -2093
rect 1468 -2101 1469 -2093
rect 1473 -2101 1474 -2093
rect 1476 -2101 1484 -2093
rect 1486 -2101 1491 -2093
rect 1495 -2101 1500 -2093
rect 1502 -2101 1503 -2093
rect 1507 -2101 1508 -2093
rect 1510 -2101 1515 -2093
rect 1519 -2101 1524 -2093
rect 1526 -2101 1527 -2093
rect 1539 -2101 1540 -2093
rect 1542 -2101 1548 -2093
rect 1550 -2101 1552 -2093
rect 1556 -2101 1558 -2093
rect 1560 -2101 1561 -2093
rect -1260 -2245 -1259 -2237
rect -1257 -2245 -1255 -2237
rect -1251 -2245 -1249 -2237
rect -1247 -2245 -1246 -2237
rect -1234 -2245 -1233 -2237
rect -1231 -2245 -1230 -2237
rect -1226 -2245 -1225 -2237
rect -1223 -2245 -1218 -2237
rect -1214 -2245 -1209 -2237
rect -1207 -2245 -1206 -2237
rect -1202 -2245 -1201 -2237
rect -1199 -2245 -1197 -2237
rect -1193 -2245 -1191 -2237
rect -1189 -2245 -1188 -2237
rect -1184 -2245 -1183 -2237
rect -1181 -2245 -1176 -2237
rect -1172 -2245 -1167 -2237
rect -1165 -2245 -1164 -2237
rect -1160 -2245 -1159 -2237
rect -1157 -2245 -1155 -2237
rect -1151 -2245 -1149 -2237
rect -1147 -2245 -1146 -2237
rect -1142 -2245 -1141 -2237
rect -1139 -2245 -1134 -2237
rect -1130 -2245 -1125 -2237
rect -1123 -2245 -1122 -2237
rect -1118 -2245 -1117 -2237
rect -1115 -2245 -1113 -2237
rect -1109 -2245 -1107 -2237
rect -1105 -2245 -1104 -2237
rect -1100 -2245 -1099 -2237
rect -1097 -2245 -1092 -2237
rect -1088 -2245 -1083 -2237
rect -1081 -2245 -1080 -2237
rect -1076 -2245 -1075 -2237
rect -1073 -2245 -1072 -2237
rect -931 -2245 -930 -2237
rect -928 -2245 -926 -2237
rect -922 -2245 -920 -2237
rect -918 -2245 -917 -2237
rect -905 -2245 -904 -2237
rect -902 -2245 -901 -2237
rect -897 -2245 -896 -2237
rect -894 -2245 -889 -2237
rect -885 -2245 -880 -2237
rect -878 -2245 -877 -2237
rect -873 -2245 -872 -2237
rect -870 -2245 -868 -2237
rect -864 -2245 -862 -2237
rect -860 -2245 -859 -2237
rect -855 -2245 -854 -2237
rect -852 -2245 -847 -2237
rect -843 -2245 -838 -2237
rect -836 -2245 -835 -2237
rect -831 -2245 -830 -2237
rect -828 -2245 -826 -2237
rect -822 -2245 -820 -2237
rect -818 -2245 -817 -2237
rect -813 -2245 -812 -2237
rect -810 -2245 -805 -2237
rect -801 -2245 -796 -2237
rect -794 -2245 -793 -2237
rect -789 -2245 -788 -2237
rect -786 -2245 -784 -2237
rect -780 -2245 -778 -2237
rect -776 -2245 -775 -2237
rect -771 -2245 -770 -2237
rect -768 -2245 -763 -2237
rect -759 -2245 -754 -2237
rect -752 -2245 -751 -2237
rect -747 -2245 -746 -2237
rect -744 -2245 -743 -2237
rect -573 -2245 -572 -2237
rect -570 -2245 -568 -2237
rect -564 -2245 -562 -2237
rect -560 -2245 -559 -2237
rect -547 -2245 -546 -2237
rect -544 -2245 -543 -2237
rect -539 -2245 -538 -2237
rect -536 -2245 -531 -2237
rect -527 -2245 -522 -2237
rect -520 -2245 -519 -2237
rect -515 -2245 -514 -2237
rect -512 -2245 -510 -2237
rect -506 -2245 -504 -2237
rect -502 -2245 -501 -2237
rect -497 -2245 -496 -2237
rect -494 -2245 -489 -2237
rect -485 -2245 -480 -2237
rect -478 -2245 -477 -2237
rect -473 -2245 -472 -2237
rect -470 -2245 -468 -2237
rect -464 -2245 -462 -2237
rect -460 -2245 -459 -2237
rect -455 -2245 -454 -2237
rect -452 -2245 -447 -2237
rect -443 -2245 -438 -2237
rect -436 -2245 -435 -2237
rect -431 -2245 -430 -2237
rect -428 -2245 -426 -2237
rect -422 -2245 -420 -2237
rect -418 -2245 -417 -2237
rect -413 -2245 -412 -2237
rect -410 -2245 -405 -2237
rect -401 -2245 -396 -2237
rect -394 -2245 -393 -2237
rect -389 -2245 -388 -2237
rect -386 -2245 -385 -2237
rect -215 -2245 -214 -2237
rect -212 -2245 -210 -2237
rect -206 -2245 -204 -2237
rect -202 -2245 -201 -2237
rect -189 -2245 -188 -2237
rect -186 -2245 -185 -2237
rect -181 -2245 -180 -2237
rect -178 -2245 -173 -2237
rect -169 -2245 -164 -2237
rect -162 -2245 -161 -2237
rect -157 -2245 -156 -2237
rect -154 -2245 -152 -2237
rect -148 -2245 -146 -2237
rect -144 -2245 -143 -2237
rect -139 -2245 -138 -2237
rect -136 -2245 -131 -2237
rect -127 -2245 -122 -2237
rect -120 -2245 -119 -2237
rect -115 -2245 -114 -2237
rect -112 -2245 -110 -2237
rect -106 -2245 -104 -2237
rect -102 -2245 -101 -2237
rect -97 -2245 -96 -2237
rect -94 -2245 -89 -2237
rect -85 -2245 -80 -2237
rect -78 -2245 -77 -2237
rect -73 -2245 -72 -2237
rect -70 -2245 -68 -2237
rect -64 -2245 -62 -2237
rect -60 -2245 -59 -2237
rect -55 -2245 -54 -2237
rect -52 -2245 -47 -2237
rect -43 -2245 -38 -2237
rect -36 -2245 -35 -2237
rect -31 -2245 -30 -2237
rect -28 -2245 -27 -2237
rect 213 -2245 214 -2237
rect 216 -2245 218 -2237
rect 222 -2245 224 -2237
rect 226 -2245 227 -2237
rect 239 -2245 240 -2237
rect 242 -2245 243 -2237
rect 247 -2245 248 -2237
rect 250 -2245 255 -2237
rect 259 -2245 264 -2237
rect 266 -2245 267 -2237
rect 271 -2245 272 -2237
rect 274 -2245 276 -2237
rect 280 -2245 282 -2237
rect 284 -2245 285 -2237
rect 289 -2245 290 -2237
rect 292 -2245 297 -2237
rect 301 -2245 306 -2237
rect 308 -2245 309 -2237
rect 313 -2245 314 -2237
rect 316 -2245 318 -2237
rect 322 -2245 324 -2237
rect 326 -2245 327 -2237
rect 331 -2245 332 -2237
rect 334 -2245 339 -2237
rect 343 -2245 348 -2237
rect 350 -2245 351 -2237
rect 355 -2245 356 -2237
rect 358 -2245 360 -2237
rect 364 -2245 366 -2237
rect 368 -2245 369 -2237
rect 373 -2245 374 -2237
rect 376 -2245 381 -2237
rect 385 -2245 390 -2237
rect 392 -2245 393 -2237
rect 397 -2245 398 -2237
rect 400 -2245 401 -2237
rect 569 -2245 570 -2237
rect 572 -2245 574 -2237
rect 578 -2245 580 -2237
rect 582 -2245 583 -2237
rect 595 -2245 596 -2237
rect 598 -2245 599 -2237
rect 603 -2245 604 -2237
rect 606 -2245 611 -2237
rect 615 -2245 620 -2237
rect 622 -2245 623 -2237
rect 627 -2245 628 -2237
rect 630 -2245 632 -2237
rect 636 -2245 638 -2237
rect 640 -2245 641 -2237
rect 645 -2245 646 -2237
rect 648 -2245 653 -2237
rect 657 -2245 662 -2237
rect 664 -2245 665 -2237
rect 669 -2245 670 -2237
rect 672 -2245 674 -2237
rect 678 -2245 680 -2237
rect 682 -2245 683 -2237
rect 687 -2245 688 -2237
rect 690 -2245 695 -2237
rect 699 -2245 704 -2237
rect 706 -2245 707 -2237
rect 711 -2245 712 -2237
rect 714 -2245 716 -2237
rect 720 -2245 722 -2237
rect 724 -2245 725 -2237
rect 729 -2245 730 -2237
rect 732 -2245 737 -2237
rect 741 -2245 746 -2237
rect 748 -2245 749 -2237
rect 753 -2245 754 -2237
rect 756 -2245 757 -2237
rect -1260 -2376 -1259 -2368
rect -1257 -2376 -1255 -2368
rect -1251 -2376 -1249 -2368
rect -1247 -2376 -1246 -2368
rect -1234 -2376 -1233 -2368
rect -1231 -2376 -1230 -2368
rect -1226 -2376 -1225 -2368
rect -1223 -2376 -1218 -2368
rect -1214 -2376 -1209 -2368
rect -1207 -2376 -1206 -2368
rect -1202 -2376 -1201 -2368
rect -1199 -2376 -1197 -2368
rect -1193 -2376 -1191 -2368
rect -1189 -2376 -1188 -2368
rect -1184 -2376 -1183 -2368
rect -1181 -2376 -1176 -2368
rect -1172 -2376 -1167 -2368
rect -1165 -2376 -1164 -2368
rect -1160 -2376 -1159 -2368
rect -1157 -2376 -1155 -2368
rect -1151 -2376 -1149 -2368
rect -1147 -2376 -1146 -2368
rect -1142 -2376 -1141 -2368
rect -1139 -2376 -1134 -2368
rect -1130 -2376 -1125 -2368
rect -1123 -2376 -1122 -2368
rect -1118 -2376 -1117 -2368
rect -1115 -2376 -1113 -2368
rect -1109 -2376 -1107 -2368
rect -1105 -2376 -1104 -2368
rect -1100 -2376 -1099 -2368
rect -1097 -2376 -1092 -2368
rect -1088 -2376 -1083 -2368
rect -1081 -2376 -1080 -2368
rect -1076 -2376 -1075 -2368
rect -1073 -2376 -1072 -2368
rect -931 -2376 -930 -2368
rect -928 -2376 -926 -2368
rect -922 -2376 -920 -2368
rect -918 -2376 -917 -2368
rect -905 -2376 -904 -2368
rect -902 -2376 -901 -2368
rect -897 -2376 -896 -2368
rect -894 -2376 -889 -2368
rect -885 -2376 -880 -2368
rect -878 -2376 -877 -2368
rect -873 -2376 -872 -2368
rect -870 -2376 -868 -2368
rect -864 -2376 -862 -2368
rect -860 -2376 -859 -2368
rect -855 -2376 -854 -2368
rect -852 -2376 -847 -2368
rect -843 -2376 -838 -2368
rect -836 -2376 -835 -2368
rect -831 -2376 -830 -2368
rect -828 -2376 -826 -2368
rect -822 -2376 -820 -2368
rect -818 -2376 -817 -2368
rect -813 -2376 -812 -2368
rect -810 -2376 -805 -2368
rect -801 -2376 -796 -2368
rect -794 -2376 -793 -2368
rect -789 -2376 -788 -2368
rect -786 -2376 -784 -2368
rect -780 -2376 -778 -2368
rect -776 -2376 -775 -2368
rect -771 -2376 -770 -2368
rect -768 -2376 -763 -2368
rect -759 -2376 -754 -2368
rect -752 -2376 -751 -2368
rect -747 -2376 -746 -2368
rect -744 -2376 -743 -2368
rect -573 -2376 -572 -2368
rect -570 -2376 -568 -2368
rect -564 -2376 -562 -2368
rect -560 -2376 -559 -2368
rect -547 -2376 -546 -2368
rect -544 -2376 -543 -2368
rect -539 -2376 -538 -2368
rect -536 -2376 -531 -2368
rect -527 -2376 -522 -2368
rect -520 -2376 -519 -2368
rect -515 -2376 -514 -2368
rect -512 -2376 -510 -2368
rect -506 -2376 -504 -2368
rect -502 -2376 -501 -2368
rect -497 -2376 -496 -2368
rect -494 -2376 -489 -2368
rect -485 -2376 -480 -2368
rect -478 -2376 -477 -2368
rect -473 -2376 -472 -2368
rect -470 -2376 -468 -2368
rect -464 -2376 -462 -2368
rect -460 -2376 -459 -2368
rect -455 -2376 -454 -2368
rect -452 -2376 -447 -2368
rect -443 -2376 -438 -2368
rect -436 -2376 -435 -2368
rect -431 -2376 -430 -2368
rect -428 -2376 -426 -2368
rect -422 -2376 -420 -2368
rect -418 -2376 -417 -2368
rect -413 -2376 -412 -2368
rect -410 -2376 -405 -2368
rect -401 -2376 -396 -2368
rect -394 -2376 -393 -2368
rect -389 -2376 -388 -2368
rect -386 -2376 -385 -2368
rect -215 -2376 -214 -2368
rect -212 -2376 -210 -2368
rect -206 -2376 -204 -2368
rect -202 -2376 -201 -2368
rect -189 -2376 -188 -2368
rect -186 -2376 -185 -2368
rect -181 -2376 -180 -2368
rect -178 -2376 -173 -2368
rect -169 -2376 -164 -2368
rect -162 -2376 -161 -2368
rect -157 -2376 -156 -2368
rect -154 -2376 -152 -2368
rect -148 -2376 -146 -2368
rect -144 -2376 -143 -2368
rect -139 -2376 -138 -2368
rect -136 -2376 -131 -2368
rect -127 -2376 -122 -2368
rect -120 -2376 -119 -2368
rect -115 -2376 -114 -2368
rect -112 -2376 -110 -2368
rect -106 -2376 -104 -2368
rect -102 -2376 -101 -2368
rect -97 -2376 -96 -2368
rect -94 -2376 -89 -2368
rect -85 -2376 -80 -2368
rect -78 -2376 -77 -2368
rect -73 -2376 -72 -2368
rect -70 -2376 -68 -2368
rect -64 -2376 -62 -2368
rect -60 -2376 -59 -2368
rect -55 -2376 -54 -2368
rect -52 -2376 -47 -2368
rect -43 -2376 -38 -2368
rect -36 -2376 -35 -2368
rect -31 -2376 -30 -2368
rect -28 -2376 -27 -2368
rect 213 -2376 214 -2368
rect 216 -2376 218 -2368
rect 222 -2376 224 -2368
rect 226 -2376 227 -2368
rect 239 -2376 240 -2368
rect 242 -2376 243 -2368
rect 247 -2376 248 -2368
rect 250 -2376 255 -2368
rect 259 -2376 264 -2368
rect 266 -2376 267 -2368
rect 271 -2376 272 -2368
rect 274 -2376 276 -2368
rect 280 -2376 282 -2368
rect 284 -2376 285 -2368
rect 289 -2376 290 -2368
rect 292 -2376 297 -2368
rect 301 -2376 306 -2368
rect 308 -2376 309 -2368
rect 313 -2376 314 -2368
rect 316 -2376 318 -2368
rect 322 -2376 324 -2368
rect 326 -2376 327 -2368
rect 331 -2376 332 -2368
rect 334 -2376 339 -2368
rect 343 -2376 348 -2368
rect 350 -2376 351 -2368
rect 355 -2376 356 -2368
rect 358 -2376 360 -2368
rect 364 -2376 366 -2368
rect 368 -2376 369 -2368
rect 373 -2376 374 -2368
rect 376 -2376 381 -2368
rect 385 -2376 390 -2368
rect 392 -2376 393 -2368
rect 397 -2376 398 -2368
rect 400 -2376 401 -2368
rect 569 -2376 570 -2368
rect 572 -2376 574 -2368
rect 578 -2376 580 -2368
rect 582 -2376 583 -2368
rect 595 -2376 596 -2368
rect 598 -2376 599 -2368
rect 603 -2376 604 -2368
rect 606 -2376 611 -2368
rect 615 -2376 620 -2368
rect 622 -2376 623 -2368
rect 627 -2376 628 -2368
rect 630 -2376 632 -2368
rect 636 -2376 638 -2368
rect 640 -2376 641 -2368
rect 645 -2376 646 -2368
rect 648 -2376 653 -2368
rect 657 -2376 662 -2368
rect 664 -2376 665 -2368
rect 669 -2376 670 -2368
rect 672 -2376 674 -2368
rect 678 -2376 680 -2368
rect 682 -2376 683 -2368
rect 687 -2376 688 -2368
rect 690 -2376 695 -2368
rect 699 -2376 704 -2368
rect 706 -2376 707 -2368
rect 711 -2376 712 -2368
rect 714 -2376 716 -2368
rect 720 -2376 722 -2368
rect 724 -2376 725 -2368
rect 729 -2376 730 -2368
rect 732 -2376 737 -2368
rect 741 -2376 746 -2368
rect 748 -2376 749 -2368
rect 753 -2376 754 -2368
rect 756 -2376 757 -2368
rect 967 -2376 968 -2368
rect 970 -2376 972 -2368
rect 976 -2376 978 -2368
rect 980 -2376 981 -2368
rect 993 -2376 994 -2368
rect 996 -2376 997 -2368
rect 1001 -2376 1002 -2368
rect 1004 -2376 1009 -2368
rect 1013 -2376 1018 -2368
rect 1020 -2376 1021 -2368
rect 1025 -2376 1026 -2368
rect 1028 -2376 1030 -2368
rect 1034 -2376 1036 -2368
rect 1038 -2376 1039 -2368
rect 1043 -2376 1044 -2368
rect 1046 -2376 1051 -2368
rect 1055 -2376 1060 -2368
rect 1062 -2376 1063 -2368
rect 1067 -2376 1068 -2368
rect 1070 -2376 1072 -2368
rect 1076 -2376 1078 -2368
rect 1080 -2376 1081 -2368
rect 1085 -2376 1086 -2368
rect 1088 -2376 1093 -2368
rect 1097 -2376 1102 -2368
rect 1104 -2376 1105 -2368
rect 1109 -2376 1110 -2368
rect 1112 -2376 1114 -2368
rect 1118 -2376 1120 -2368
rect 1122 -2376 1123 -2368
rect 1127 -2376 1128 -2368
rect 1130 -2376 1135 -2368
rect 1139 -2376 1144 -2368
rect 1146 -2376 1147 -2368
rect 1151 -2376 1152 -2368
rect 1154 -2376 1155 -2368
rect 1325 -2376 1326 -2368
rect 1328 -2376 1330 -2368
rect 1334 -2376 1336 -2368
rect 1338 -2376 1339 -2368
rect 1351 -2376 1352 -2368
rect 1354 -2376 1355 -2368
rect 1359 -2376 1360 -2368
rect 1362 -2376 1367 -2368
rect 1371 -2376 1376 -2368
rect 1378 -2376 1379 -2368
rect 1383 -2376 1384 -2368
rect 1386 -2376 1388 -2368
rect 1392 -2376 1394 -2368
rect 1396 -2376 1397 -2368
rect 1401 -2376 1402 -2368
rect 1404 -2376 1409 -2368
rect 1413 -2376 1418 -2368
rect 1420 -2376 1421 -2368
rect 1425 -2376 1426 -2368
rect 1428 -2376 1430 -2368
rect 1434 -2376 1436 -2368
rect 1438 -2376 1439 -2368
rect 1443 -2376 1444 -2368
rect 1446 -2376 1451 -2368
rect 1455 -2376 1460 -2368
rect 1462 -2376 1463 -2368
rect 1467 -2376 1468 -2368
rect 1470 -2376 1472 -2368
rect 1476 -2376 1478 -2368
rect 1480 -2376 1481 -2368
rect 1485 -2376 1486 -2368
rect 1488 -2376 1493 -2368
rect 1497 -2376 1502 -2368
rect 1504 -2376 1505 -2368
rect 1509 -2376 1510 -2368
rect 1512 -2376 1513 -2368
rect -1260 -2507 -1259 -2499
rect -1257 -2507 -1255 -2499
rect -1251 -2507 -1249 -2499
rect -1247 -2507 -1246 -2499
rect -1234 -2507 -1233 -2499
rect -1231 -2507 -1230 -2499
rect -1226 -2507 -1225 -2499
rect -1223 -2507 -1218 -2499
rect -1214 -2507 -1209 -2499
rect -1207 -2507 -1206 -2499
rect -1202 -2507 -1201 -2499
rect -1199 -2507 -1197 -2499
rect -1193 -2507 -1191 -2499
rect -1189 -2507 -1188 -2499
rect -1184 -2507 -1183 -2499
rect -1181 -2507 -1176 -2499
rect -1172 -2507 -1167 -2499
rect -1165 -2507 -1164 -2499
rect -1160 -2507 -1159 -2499
rect -1157 -2507 -1155 -2499
rect -1151 -2507 -1149 -2499
rect -1147 -2507 -1146 -2499
rect -1142 -2507 -1141 -2499
rect -1139 -2507 -1134 -2499
rect -1130 -2507 -1125 -2499
rect -1123 -2507 -1122 -2499
rect -1118 -2507 -1117 -2499
rect -1115 -2507 -1113 -2499
rect -1109 -2507 -1107 -2499
rect -1105 -2507 -1104 -2499
rect -1100 -2507 -1099 -2499
rect -1097 -2507 -1092 -2499
rect -1088 -2507 -1083 -2499
rect -1081 -2507 -1080 -2499
rect -1076 -2507 -1075 -2499
rect -1073 -2507 -1072 -2499
rect -931 -2507 -930 -2499
rect -928 -2507 -926 -2499
rect -922 -2507 -920 -2499
rect -918 -2507 -917 -2499
rect -905 -2507 -904 -2499
rect -902 -2507 -901 -2499
rect -897 -2507 -896 -2499
rect -894 -2507 -889 -2499
rect -885 -2507 -880 -2499
rect -878 -2507 -877 -2499
rect -873 -2507 -872 -2499
rect -870 -2507 -868 -2499
rect -864 -2507 -862 -2499
rect -860 -2507 -859 -2499
rect -855 -2507 -854 -2499
rect -852 -2507 -847 -2499
rect -843 -2507 -838 -2499
rect -836 -2507 -835 -2499
rect -831 -2507 -830 -2499
rect -828 -2507 -826 -2499
rect -822 -2507 -820 -2499
rect -818 -2507 -817 -2499
rect -813 -2507 -812 -2499
rect -810 -2507 -805 -2499
rect -801 -2507 -796 -2499
rect -794 -2507 -793 -2499
rect -789 -2507 -788 -2499
rect -786 -2507 -784 -2499
rect -780 -2507 -778 -2499
rect -776 -2507 -775 -2499
rect -771 -2507 -770 -2499
rect -768 -2507 -763 -2499
rect -759 -2507 -754 -2499
rect -752 -2507 -751 -2499
rect -747 -2507 -746 -2499
rect -744 -2507 -743 -2499
rect -573 -2507 -572 -2499
rect -570 -2507 -568 -2499
rect -564 -2507 -562 -2499
rect -560 -2507 -559 -2499
rect -547 -2507 -546 -2499
rect -544 -2507 -543 -2499
rect -539 -2507 -538 -2499
rect -536 -2507 -531 -2499
rect -527 -2507 -522 -2499
rect -520 -2507 -519 -2499
rect -515 -2507 -514 -2499
rect -512 -2507 -510 -2499
rect -506 -2507 -504 -2499
rect -502 -2507 -501 -2499
rect -497 -2507 -496 -2499
rect -494 -2507 -489 -2499
rect -485 -2507 -480 -2499
rect -478 -2507 -477 -2499
rect -473 -2507 -472 -2499
rect -470 -2507 -468 -2499
rect -464 -2507 -462 -2499
rect -460 -2507 -459 -2499
rect -455 -2507 -454 -2499
rect -452 -2507 -447 -2499
rect -443 -2507 -438 -2499
rect -436 -2507 -435 -2499
rect -431 -2507 -430 -2499
rect -428 -2507 -426 -2499
rect -422 -2507 -420 -2499
rect -418 -2507 -417 -2499
rect -413 -2507 -412 -2499
rect -410 -2507 -405 -2499
rect -401 -2507 -396 -2499
rect -394 -2507 -393 -2499
rect -389 -2507 -388 -2499
rect -386 -2507 -385 -2499
rect -215 -2507 -214 -2499
rect -212 -2507 -210 -2499
rect -206 -2507 -204 -2499
rect -202 -2507 -201 -2499
rect -189 -2507 -188 -2499
rect -186 -2507 -185 -2499
rect -181 -2507 -180 -2499
rect -178 -2507 -173 -2499
rect -169 -2507 -164 -2499
rect -162 -2507 -161 -2499
rect -157 -2507 -156 -2499
rect -154 -2507 -152 -2499
rect -148 -2507 -146 -2499
rect -144 -2507 -143 -2499
rect -139 -2507 -138 -2499
rect -136 -2507 -131 -2499
rect -127 -2507 -122 -2499
rect -120 -2507 -119 -2499
rect -115 -2507 -114 -2499
rect -112 -2507 -110 -2499
rect -106 -2507 -104 -2499
rect -102 -2507 -101 -2499
rect -97 -2507 -96 -2499
rect -94 -2507 -89 -2499
rect -85 -2507 -80 -2499
rect -78 -2507 -77 -2499
rect -73 -2507 -72 -2499
rect -70 -2507 -68 -2499
rect -64 -2507 -62 -2499
rect -60 -2507 -59 -2499
rect -55 -2507 -54 -2499
rect -52 -2507 -47 -2499
rect -43 -2507 -38 -2499
rect -36 -2507 -35 -2499
rect -31 -2507 -30 -2499
rect -28 -2507 -27 -2499
rect 94 -2531 95 -2499
rect 97 -2531 98 -2499
rect 213 -2507 214 -2499
rect 216 -2507 218 -2499
rect 222 -2507 224 -2499
rect 226 -2507 227 -2499
rect 239 -2507 240 -2499
rect 242 -2507 243 -2499
rect 247 -2507 248 -2499
rect 250 -2507 255 -2499
rect 259 -2507 264 -2499
rect 266 -2507 267 -2499
rect 271 -2507 272 -2499
rect 274 -2507 276 -2499
rect 280 -2507 282 -2499
rect 284 -2507 285 -2499
rect 289 -2507 290 -2499
rect 292 -2507 297 -2499
rect 301 -2507 306 -2499
rect 308 -2507 309 -2499
rect 313 -2507 314 -2499
rect 316 -2507 318 -2499
rect 322 -2507 324 -2499
rect 326 -2507 327 -2499
rect 331 -2507 332 -2499
rect 334 -2507 339 -2499
rect 343 -2507 348 -2499
rect 350 -2507 351 -2499
rect 355 -2507 356 -2499
rect 358 -2507 360 -2499
rect 364 -2507 366 -2499
rect 368 -2507 369 -2499
rect 373 -2507 374 -2499
rect 376 -2507 381 -2499
rect 385 -2507 390 -2499
rect 392 -2507 393 -2499
rect 397 -2507 398 -2499
rect 400 -2507 401 -2499
rect 569 -2507 570 -2499
rect 572 -2507 574 -2499
rect 578 -2507 580 -2499
rect 582 -2507 583 -2499
rect 595 -2507 596 -2499
rect 598 -2507 599 -2499
rect 603 -2507 604 -2499
rect 606 -2507 611 -2499
rect 615 -2507 620 -2499
rect 622 -2507 623 -2499
rect 627 -2507 628 -2499
rect 630 -2507 632 -2499
rect 636 -2507 638 -2499
rect 640 -2507 641 -2499
rect 645 -2507 646 -2499
rect 648 -2507 653 -2499
rect 657 -2507 662 -2499
rect 664 -2507 665 -2499
rect 669 -2507 670 -2499
rect 672 -2507 674 -2499
rect 678 -2507 680 -2499
rect 682 -2507 683 -2499
rect 687 -2507 688 -2499
rect 690 -2507 695 -2499
rect 699 -2507 704 -2499
rect 706 -2507 707 -2499
rect 711 -2507 712 -2499
rect 714 -2507 716 -2499
rect 720 -2507 722 -2499
rect 724 -2507 725 -2499
rect 729 -2507 730 -2499
rect 732 -2507 737 -2499
rect 741 -2507 746 -2499
rect 748 -2507 749 -2499
rect 753 -2507 754 -2499
rect 756 -2507 757 -2499
rect 967 -2507 968 -2499
rect 970 -2507 972 -2499
rect 976 -2507 978 -2499
rect 980 -2507 981 -2499
rect 993 -2507 994 -2499
rect 996 -2507 997 -2499
rect 1001 -2507 1002 -2499
rect 1004 -2507 1009 -2499
rect 1013 -2507 1018 -2499
rect 1020 -2507 1021 -2499
rect 1025 -2507 1026 -2499
rect 1028 -2507 1030 -2499
rect 1034 -2507 1036 -2499
rect 1038 -2507 1039 -2499
rect 1043 -2507 1044 -2499
rect 1046 -2507 1051 -2499
rect 1055 -2507 1060 -2499
rect 1062 -2507 1063 -2499
rect 1067 -2507 1068 -2499
rect 1070 -2507 1072 -2499
rect 1076 -2507 1078 -2499
rect 1080 -2507 1081 -2499
rect 1085 -2507 1086 -2499
rect 1088 -2507 1093 -2499
rect 1097 -2507 1102 -2499
rect 1104 -2507 1105 -2499
rect 1109 -2507 1110 -2499
rect 1112 -2507 1114 -2499
rect 1118 -2507 1120 -2499
rect 1122 -2507 1123 -2499
rect 1127 -2507 1128 -2499
rect 1130 -2507 1135 -2499
rect 1139 -2507 1144 -2499
rect 1146 -2507 1147 -2499
rect 1151 -2507 1152 -2499
rect 1154 -2507 1155 -2499
rect 1325 -2507 1326 -2499
rect 1328 -2507 1330 -2499
rect 1334 -2507 1336 -2499
rect 1338 -2507 1339 -2499
rect 1351 -2507 1352 -2499
rect 1354 -2507 1355 -2499
rect 1359 -2507 1360 -2499
rect 1362 -2507 1367 -2499
rect 1371 -2507 1376 -2499
rect 1378 -2507 1379 -2499
rect 1383 -2507 1384 -2499
rect 1386 -2507 1388 -2499
rect 1392 -2507 1394 -2499
rect 1396 -2507 1397 -2499
rect 1401 -2507 1402 -2499
rect 1404 -2507 1409 -2499
rect 1413 -2507 1418 -2499
rect 1420 -2507 1421 -2499
rect 1425 -2507 1426 -2499
rect 1428 -2507 1430 -2499
rect 1434 -2507 1436 -2499
rect 1438 -2507 1439 -2499
rect 1443 -2507 1444 -2499
rect 1446 -2507 1451 -2499
rect 1455 -2507 1460 -2499
rect 1462 -2507 1463 -2499
rect 1467 -2507 1468 -2499
rect 1470 -2507 1472 -2499
rect 1476 -2507 1478 -2499
rect 1480 -2507 1481 -2499
rect 1485 -2507 1486 -2499
rect 1488 -2507 1493 -2499
rect 1497 -2507 1502 -2499
rect 1504 -2507 1505 -2499
rect 1509 -2507 1510 -2499
rect 1512 -2507 1513 -2499
rect -1260 -2619 -1259 -2611
rect -1257 -2619 -1255 -2611
rect -1251 -2619 -1249 -2611
rect -1247 -2619 -1246 -2611
rect -1234 -2619 -1233 -2611
rect -1231 -2619 -1230 -2611
rect -1226 -2619 -1225 -2611
rect -1223 -2619 -1218 -2611
rect -1214 -2619 -1209 -2611
rect -1207 -2619 -1206 -2611
rect -1202 -2619 -1201 -2611
rect -1199 -2619 -1197 -2611
rect -1193 -2619 -1191 -2611
rect -1189 -2619 -1188 -2611
rect -1184 -2619 -1183 -2611
rect -1181 -2619 -1176 -2611
rect -1172 -2619 -1167 -2611
rect -1165 -2619 -1164 -2611
rect -1160 -2619 -1159 -2611
rect -1157 -2619 -1155 -2611
rect -1151 -2619 -1149 -2611
rect -1147 -2619 -1146 -2611
rect -1142 -2619 -1141 -2611
rect -1139 -2619 -1134 -2611
rect -1130 -2619 -1125 -2611
rect -1123 -2619 -1122 -2611
rect -1118 -2619 -1117 -2611
rect -1115 -2619 -1113 -2611
rect -1109 -2619 -1107 -2611
rect -1105 -2619 -1104 -2611
rect -1100 -2619 -1099 -2611
rect -1097 -2619 -1092 -2611
rect -1088 -2619 -1083 -2611
rect -1081 -2619 -1080 -2611
rect -1076 -2619 -1075 -2611
rect -1073 -2619 -1072 -2611
rect -931 -2619 -930 -2611
rect -928 -2619 -926 -2611
rect -922 -2619 -920 -2611
rect -918 -2619 -917 -2611
rect -905 -2619 -904 -2611
rect -902 -2619 -901 -2611
rect -897 -2619 -896 -2611
rect -894 -2619 -889 -2611
rect -885 -2619 -880 -2611
rect -878 -2619 -877 -2611
rect -873 -2619 -872 -2611
rect -870 -2619 -868 -2611
rect -864 -2619 -862 -2611
rect -860 -2619 -859 -2611
rect -855 -2619 -854 -2611
rect -852 -2619 -847 -2611
rect -843 -2619 -838 -2611
rect -836 -2619 -835 -2611
rect -831 -2619 -830 -2611
rect -828 -2619 -826 -2611
rect -822 -2619 -820 -2611
rect -818 -2619 -817 -2611
rect -813 -2619 -812 -2611
rect -810 -2619 -805 -2611
rect -801 -2619 -796 -2611
rect -794 -2619 -793 -2611
rect -789 -2619 -788 -2611
rect -786 -2619 -784 -2611
rect -780 -2619 -778 -2611
rect -776 -2619 -775 -2611
rect -771 -2619 -770 -2611
rect -768 -2619 -763 -2611
rect -759 -2619 -754 -2611
rect -752 -2619 -751 -2611
rect -747 -2619 -746 -2611
rect -744 -2619 -743 -2611
rect -1335 -2732 -1334 -2724
rect -1332 -2732 -1331 -2724
rect -1327 -2732 -1326 -2724
rect -1324 -2732 -1322 -2724
rect -1318 -2732 -1316 -2724
rect -1314 -2732 -1313 -2724
rect -931 -2732 -930 -2724
rect -928 -2732 -927 -2724
rect -923 -2732 -922 -2724
rect -920 -2732 -918 -2724
rect -914 -2732 -912 -2724
rect -910 -2732 -909 -2724
rect -573 -2732 -572 -2724
rect -570 -2732 -569 -2724
rect -565 -2732 -564 -2724
rect -562 -2732 -560 -2724
rect -556 -2732 -554 -2724
rect -552 -2732 -551 -2724
rect -215 -2732 -214 -2724
rect -212 -2732 -211 -2724
rect -207 -2732 -206 -2724
rect -204 -2732 -202 -2724
rect -198 -2732 -196 -2724
rect -194 -2732 -193 -2724
rect 213 -2732 214 -2724
rect 216 -2732 217 -2724
rect 221 -2732 222 -2724
rect 224 -2732 226 -2724
rect 230 -2732 232 -2724
rect 234 -2732 235 -2724
rect 569 -2732 570 -2724
rect 572 -2732 573 -2724
rect 577 -2732 578 -2724
rect 580 -2732 582 -2724
rect 586 -2732 588 -2724
rect 590 -2732 591 -2724
rect 967 -2732 968 -2724
rect 970 -2732 971 -2724
rect 975 -2732 976 -2724
rect 978 -2732 980 -2724
rect 984 -2732 986 -2724
rect 988 -2732 989 -2724
rect 1325 -2732 1326 -2724
rect 1328 -2732 1329 -2724
rect 1333 -2732 1334 -2724
rect 1336 -2732 1338 -2724
rect 1342 -2732 1344 -2724
rect 1346 -2732 1347 -2724
rect -1260 -2851 -1259 -2843
rect -1257 -2851 -1255 -2843
rect -1251 -2851 -1249 -2843
rect -1247 -2851 -1246 -2843
rect -1234 -2851 -1233 -2843
rect -1231 -2851 -1223 -2843
rect -1221 -2851 -1220 -2843
rect -1216 -2851 -1215 -2843
rect -1213 -2851 -1205 -2843
rect -1203 -2851 -1198 -2843
rect -1194 -2851 -1189 -2843
rect -1187 -2851 -1186 -2843
rect -1182 -2851 -1181 -2843
rect -1179 -2851 -1177 -2843
rect -1173 -2851 -1171 -2843
rect -1169 -2851 -1168 -2843
rect -931 -2851 -930 -2843
rect -928 -2851 -926 -2843
rect -922 -2851 -920 -2843
rect -918 -2851 -917 -2843
rect -905 -2851 -904 -2843
rect -902 -2851 -900 -2843
rect -896 -2851 -894 -2843
rect -892 -2851 -891 -2843
rect -879 -2851 -878 -2843
rect -876 -2851 -868 -2843
rect -866 -2851 -865 -2843
rect -861 -2851 -860 -2843
rect -858 -2851 -850 -2843
rect -848 -2851 -843 -2843
rect -839 -2851 -834 -2843
rect -832 -2851 -831 -2843
rect -827 -2851 -826 -2843
rect -824 -2851 -822 -2843
rect -818 -2851 -816 -2843
rect -814 -2851 -813 -2843
rect -801 -2851 -800 -2843
rect -798 -2851 -790 -2843
rect -788 -2851 -787 -2843
rect -783 -2851 -782 -2843
rect -780 -2851 -772 -2843
rect -770 -2851 -765 -2843
rect -761 -2851 -756 -2843
rect -754 -2851 -753 -2843
rect -749 -2851 -748 -2843
rect -746 -2851 -741 -2843
rect -737 -2851 -732 -2843
rect -730 -2851 -729 -2843
rect -717 -2851 -716 -2843
rect -714 -2851 -708 -2843
rect -706 -2851 -704 -2843
rect -700 -2851 -698 -2843
rect -696 -2851 -695 -2843
rect -573 -2851 -572 -2843
rect -570 -2851 -568 -2843
rect -564 -2851 -562 -2843
rect -560 -2851 -559 -2843
rect -547 -2851 -546 -2843
rect -544 -2851 -542 -2843
rect -538 -2851 -536 -2843
rect -534 -2851 -533 -2843
rect -521 -2851 -520 -2843
rect -518 -2851 -510 -2843
rect -508 -2851 -507 -2843
rect -503 -2851 -502 -2843
rect -500 -2851 -492 -2843
rect -490 -2851 -485 -2843
rect -481 -2851 -476 -2843
rect -474 -2851 -473 -2843
rect -469 -2851 -468 -2843
rect -466 -2851 -464 -2843
rect -460 -2851 -458 -2843
rect -456 -2851 -455 -2843
rect -443 -2851 -442 -2843
rect -440 -2851 -432 -2843
rect -430 -2851 -429 -2843
rect -425 -2851 -424 -2843
rect -422 -2851 -414 -2843
rect -412 -2851 -407 -2843
rect -403 -2851 -398 -2843
rect -396 -2851 -395 -2843
rect -391 -2851 -390 -2843
rect -388 -2851 -383 -2843
rect -379 -2851 -374 -2843
rect -372 -2851 -371 -2843
rect -359 -2851 -358 -2843
rect -356 -2851 -350 -2843
rect -348 -2851 -346 -2843
rect -342 -2851 -340 -2843
rect -338 -2851 -337 -2843
rect -215 -2851 -214 -2843
rect -212 -2851 -210 -2843
rect -206 -2851 -204 -2843
rect -202 -2851 -201 -2843
rect -189 -2851 -188 -2843
rect -186 -2851 -184 -2843
rect -180 -2851 -178 -2843
rect -176 -2851 -175 -2843
rect -163 -2851 -162 -2843
rect -160 -2851 -152 -2843
rect -150 -2851 -149 -2843
rect -145 -2851 -144 -2843
rect -142 -2851 -134 -2843
rect -132 -2851 -127 -2843
rect -123 -2851 -118 -2843
rect -116 -2851 -115 -2843
rect -111 -2851 -110 -2843
rect -108 -2851 -106 -2843
rect -102 -2851 -100 -2843
rect -98 -2851 -97 -2843
rect -85 -2851 -84 -2843
rect -82 -2851 -74 -2843
rect -72 -2851 -71 -2843
rect -67 -2851 -66 -2843
rect -64 -2851 -56 -2843
rect -54 -2851 -49 -2843
rect -45 -2851 -40 -2843
rect -38 -2851 -37 -2843
rect -33 -2851 -32 -2843
rect -30 -2851 -25 -2843
rect -21 -2851 -16 -2843
rect -14 -2851 -13 -2843
rect -1 -2851 0 -2843
rect 2 -2851 8 -2843
rect 10 -2851 12 -2843
rect 16 -2851 18 -2843
rect 20 -2851 21 -2843
rect 213 -2851 214 -2843
rect 216 -2851 218 -2843
rect 222 -2851 224 -2843
rect 226 -2851 227 -2843
rect 239 -2851 240 -2843
rect 242 -2851 244 -2843
rect 248 -2851 250 -2843
rect 252 -2851 253 -2843
rect 265 -2851 266 -2843
rect 268 -2851 276 -2843
rect 278 -2851 279 -2843
rect 283 -2851 284 -2843
rect 286 -2851 294 -2843
rect 296 -2851 301 -2843
rect 305 -2851 310 -2843
rect 312 -2851 313 -2843
rect 317 -2851 318 -2843
rect 320 -2851 322 -2843
rect 326 -2851 328 -2843
rect 330 -2851 331 -2843
rect 343 -2851 344 -2843
rect 346 -2851 354 -2843
rect 356 -2851 357 -2843
rect 361 -2851 362 -2843
rect 364 -2851 372 -2843
rect 374 -2851 379 -2843
rect 383 -2851 388 -2843
rect 390 -2851 391 -2843
rect 395 -2851 396 -2843
rect 398 -2851 403 -2843
rect 407 -2851 412 -2843
rect 414 -2851 415 -2843
rect 427 -2851 428 -2843
rect 430 -2851 436 -2843
rect 438 -2851 440 -2843
rect 444 -2851 446 -2843
rect 448 -2851 449 -2843
rect 569 -2851 570 -2843
rect 572 -2851 574 -2843
rect 578 -2851 580 -2843
rect 582 -2851 583 -2843
rect 595 -2851 596 -2843
rect 598 -2851 600 -2843
rect 604 -2851 606 -2843
rect 608 -2851 609 -2843
rect 621 -2851 622 -2843
rect 624 -2851 632 -2843
rect 634 -2851 635 -2843
rect 639 -2851 640 -2843
rect 642 -2851 650 -2843
rect 652 -2851 657 -2843
rect 661 -2851 666 -2843
rect 668 -2851 669 -2843
rect 673 -2851 674 -2843
rect 676 -2851 678 -2843
rect 682 -2851 684 -2843
rect 686 -2851 687 -2843
rect 699 -2851 700 -2843
rect 702 -2851 710 -2843
rect 712 -2851 713 -2843
rect 717 -2851 718 -2843
rect 720 -2851 728 -2843
rect 730 -2851 735 -2843
rect 739 -2851 744 -2843
rect 746 -2851 747 -2843
rect 751 -2851 752 -2843
rect 754 -2851 759 -2843
rect 763 -2851 768 -2843
rect 770 -2851 771 -2843
rect 783 -2851 784 -2843
rect 786 -2851 792 -2843
rect 794 -2851 796 -2843
rect 800 -2851 802 -2843
rect 804 -2851 805 -2843
rect 967 -2851 968 -2843
rect 970 -2851 972 -2843
rect 976 -2851 978 -2843
rect 980 -2851 981 -2843
rect 993 -2851 994 -2843
rect 996 -2851 998 -2843
rect 1002 -2851 1004 -2843
rect 1006 -2851 1007 -2843
rect 1019 -2851 1020 -2843
rect 1022 -2851 1030 -2843
rect 1032 -2851 1033 -2843
rect 1037 -2851 1038 -2843
rect 1040 -2851 1048 -2843
rect 1050 -2851 1055 -2843
rect 1059 -2851 1064 -2843
rect 1066 -2851 1067 -2843
rect 1071 -2851 1072 -2843
rect 1074 -2851 1076 -2843
rect 1080 -2851 1082 -2843
rect 1084 -2851 1085 -2843
rect 1097 -2851 1098 -2843
rect 1100 -2851 1108 -2843
rect 1110 -2851 1111 -2843
rect 1115 -2851 1116 -2843
rect 1118 -2851 1126 -2843
rect 1128 -2851 1133 -2843
rect 1137 -2851 1142 -2843
rect 1144 -2851 1145 -2843
rect 1149 -2851 1150 -2843
rect 1152 -2851 1157 -2843
rect 1161 -2851 1166 -2843
rect 1168 -2851 1169 -2843
rect 1181 -2851 1182 -2843
rect 1184 -2851 1190 -2843
rect 1192 -2851 1194 -2843
rect 1198 -2851 1200 -2843
rect 1202 -2851 1203 -2843
rect 1325 -2851 1326 -2843
rect 1328 -2851 1330 -2843
rect 1334 -2851 1336 -2843
rect 1338 -2851 1339 -2843
rect 1351 -2851 1352 -2843
rect 1354 -2851 1356 -2843
rect 1360 -2851 1362 -2843
rect 1364 -2851 1365 -2843
rect 1377 -2851 1378 -2843
rect 1380 -2851 1388 -2843
rect 1390 -2851 1391 -2843
rect 1395 -2851 1396 -2843
rect 1398 -2851 1406 -2843
rect 1408 -2851 1413 -2843
rect 1417 -2851 1422 -2843
rect 1424 -2851 1425 -2843
rect 1429 -2851 1430 -2843
rect 1432 -2851 1434 -2843
rect 1438 -2851 1440 -2843
rect 1442 -2851 1443 -2843
rect 1455 -2851 1456 -2843
rect 1458 -2851 1466 -2843
rect 1468 -2851 1469 -2843
rect 1473 -2851 1474 -2843
rect 1476 -2851 1484 -2843
rect 1486 -2851 1491 -2843
rect 1495 -2851 1500 -2843
rect 1502 -2851 1503 -2843
rect 1507 -2851 1508 -2843
rect 1510 -2851 1515 -2843
rect 1519 -2851 1524 -2843
rect 1526 -2851 1527 -2843
rect 1539 -2851 1540 -2843
rect 1542 -2851 1548 -2843
rect 1550 -2851 1552 -2843
rect 1556 -2851 1558 -2843
rect 1560 -2851 1561 -2843
rect -1260 -2970 -1259 -2962
rect -1257 -2970 -1255 -2962
rect -1251 -2970 -1249 -2962
rect -1247 -2970 -1246 -2962
rect -1234 -2970 -1233 -2962
rect -1231 -2970 -1230 -2962
rect -1226 -2970 -1225 -2962
rect -1223 -2970 -1218 -2962
rect -1214 -2970 -1209 -2962
rect -1207 -2970 -1206 -2962
rect -1202 -2970 -1201 -2962
rect -1199 -2970 -1197 -2962
rect -1193 -2970 -1191 -2962
rect -1189 -2970 -1188 -2962
rect -1184 -2970 -1183 -2962
rect -1181 -2970 -1176 -2962
rect -1172 -2970 -1167 -2962
rect -1165 -2970 -1164 -2962
rect -1160 -2970 -1159 -2962
rect -1157 -2970 -1155 -2962
rect -1151 -2970 -1149 -2962
rect -1147 -2970 -1146 -2962
rect -1142 -2970 -1141 -2962
rect -1139 -2970 -1134 -2962
rect -1130 -2970 -1125 -2962
rect -1123 -2970 -1122 -2962
rect -1118 -2970 -1117 -2962
rect -1115 -2970 -1113 -2962
rect -1109 -2970 -1107 -2962
rect -1105 -2970 -1104 -2962
rect -1100 -2970 -1099 -2962
rect -1097 -2970 -1092 -2962
rect -1088 -2970 -1083 -2962
rect -1081 -2970 -1080 -2962
rect -1076 -2970 -1075 -2962
rect -1073 -2970 -1072 -2962
rect -1022 -2970 -1021 -2962
rect -1019 -2970 -1018 -2962
rect -931 -2970 -930 -2962
rect -928 -2970 -926 -2962
rect -922 -2970 -920 -2962
rect -918 -2970 -917 -2962
rect -905 -2970 -904 -2962
rect -902 -2970 -901 -2962
rect -897 -2970 -896 -2962
rect -894 -2970 -889 -2962
rect -885 -2970 -880 -2962
rect -878 -2970 -877 -2962
rect -873 -2970 -872 -2962
rect -870 -2970 -868 -2962
rect -864 -2970 -862 -2962
rect -860 -2970 -859 -2962
rect -855 -2970 -854 -2962
rect -852 -2970 -847 -2962
rect -843 -2970 -838 -2962
rect -836 -2970 -835 -2962
rect -831 -2970 -830 -2962
rect -828 -2970 -826 -2962
rect -822 -2970 -820 -2962
rect -818 -2970 -817 -2962
rect -813 -2970 -812 -2962
rect -810 -2970 -805 -2962
rect -801 -2970 -796 -2962
rect -794 -2970 -793 -2962
rect -789 -2970 -788 -2962
rect -786 -2970 -784 -2962
rect -780 -2970 -778 -2962
rect -776 -2970 -775 -2962
rect -771 -2970 -770 -2962
rect -768 -2970 -763 -2962
rect -759 -2970 -754 -2962
rect -752 -2970 -751 -2962
rect -747 -2970 -746 -2962
rect -744 -2970 -743 -2962
rect -668 -2978 -667 -2962
rect -665 -2978 -664 -2962
rect -573 -2970 -572 -2962
rect -570 -2970 -568 -2962
rect -564 -2970 -562 -2962
rect -560 -2970 -559 -2962
rect -547 -2970 -546 -2962
rect -544 -2970 -543 -2962
rect -539 -2970 -538 -2962
rect -536 -2970 -531 -2962
rect -527 -2970 -522 -2962
rect -520 -2970 -519 -2962
rect -515 -2970 -514 -2962
rect -512 -2970 -510 -2962
rect -506 -2970 -504 -2962
rect -502 -2970 -501 -2962
rect -497 -2970 -496 -2962
rect -494 -2970 -489 -2962
rect -485 -2970 -480 -2962
rect -478 -2970 -477 -2962
rect -473 -2970 -472 -2962
rect -470 -2970 -468 -2962
rect -464 -2970 -462 -2962
rect -460 -2970 -459 -2962
rect -455 -2970 -454 -2962
rect -452 -2970 -447 -2962
rect -443 -2970 -438 -2962
rect -436 -2970 -435 -2962
rect -431 -2970 -430 -2962
rect -428 -2970 -426 -2962
rect -422 -2970 -420 -2962
rect -418 -2970 -417 -2962
rect -413 -2970 -412 -2962
rect -410 -2970 -405 -2962
rect -401 -2970 -396 -2962
rect -394 -2970 -393 -2962
rect -389 -2970 -388 -2962
rect -386 -2970 -385 -2962
rect -325 -2970 -324 -2962
rect -322 -2970 -321 -2962
rect -215 -2970 -214 -2962
rect -212 -2970 -210 -2962
rect -206 -2970 -204 -2962
rect -202 -2970 -201 -2962
rect -189 -2970 -188 -2962
rect -186 -2970 -185 -2962
rect -181 -2970 -180 -2962
rect -178 -2970 -173 -2962
rect -169 -2970 -164 -2962
rect -162 -2970 -161 -2962
rect -157 -2970 -156 -2962
rect -154 -2970 -152 -2962
rect -148 -2970 -146 -2962
rect -144 -2970 -143 -2962
rect -139 -2970 -138 -2962
rect -136 -2970 -131 -2962
rect -127 -2970 -122 -2962
rect -120 -2970 -119 -2962
rect -115 -2970 -114 -2962
rect -112 -2970 -110 -2962
rect -106 -2970 -104 -2962
rect -102 -2970 -101 -2962
rect -97 -2970 -96 -2962
rect -94 -2970 -89 -2962
rect -85 -2970 -80 -2962
rect -78 -2970 -77 -2962
rect -73 -2970 -72 -2962
rect -70 -2970 -68 -2962
rect -64 -2970 -62 -2962
rect -60 -2970 -59 -2962
rect -55 -2970 -54 -2962
rect -52 -2970 -47 -2962
rect -43 -2970 -38 -2962
rect -36 -2970 -35 -2962
rect -31 -2970 -30 -2962
rect -28 -2970 -27 -2962
rect 213 -2970 214 -2962
rect 216 -2970 218 -2962
rect 222 -2970 224 -2962
rect 226 -2970 227 -2962
rect 239 -2970 240 -2962
rect 242 -2970 243 -2962
rect 247 -2970 248 -2962
rect 250 -2970 255 -2962
rect 259 -2970 264 -2962
rect 266 -2970 267 -2962
rect 271 -2970 272 -2962
rect 274 -2970 276 -2962
rect 280 -2970 282 -2962
rect 284 -2970 285 -2962
rect 289 -2970 290 -2962
rect 292 -2970 297 -2962
rect 301 -2970 306 -2962
rect 308 -2970 309 -2962
rect 313 -2970 314 -2962
rect 316 -2970 318 -2962
rect 322 -2970 324 -2962
rect 326 -2970 327 -2962
rect 331 -2970 332 -2962
rect 334 -2970 339 -2962
rect 343 -2970 348 -2962
rect 350 -2970 351 -2962
rect 355 -2970 356 -2962
rect 358 -2970 360 -2962
rect 364 -2970 366 -2962
rect 368 -2970 369 -2962
rect 373 -2970 374 -2962
rect 376 -2970 381 -2962
rect 385 -2970 390 -2962
rect 392 -2970 393 -2962
rect 397 -2970 398 -2962
rect 400 -2970 401 -2962
rect 476 -2970 477 -2962
rect 479 -2970 480 -2962
rect 845 -2978 846 -2962
rect 848 -2978 849 -2962
rect 1203 -2970 1204 -2962
rect 1206 -2970 1207 -2962
rect -1260 -3086 -1259 -3078
rect -1257 -3086 -1255 -3078
rect -1251 -3086 -1249 -3078
rect -1247 -3086 -1246 -3078
rect -1234 -3086 -1233 -3078
rect -1231 -3086 -1230 -3078
rect -1226 -3086 -1225 -3078
rect -1223 -3086 -1218 -3078
rect -1214 -3086 -1209 -3078
rect -1207 -3086 -1206 -3078
rect -1202 -3086 -1201 -3078
rect -1199 -3086 -1197 -3078
rect -1193 -3086 -1191 -3078
rect -1189 -3086 -1188 -3078
rect -1184 -3086 -1183 -3078
rect -1181 -3086 -1176 -3078
rect -1172 -3086 -1167 -3078
rect -1165 -3086 -1164 -3078
rect -1160 -3086 -1159 -3078
rect -1157 -3086 -1155 -3078
rect -1151 -3086 -1149 -3078
rect -1147 -3086 -1146 -3078
rect -1142 -3086 -1141 -3078
rect -1139 -3086 -1134 -3078
rect -1130 -3086 -1125 -3078
rect -1123 -3086 -1122 -3078
rect -1118 -3086 -1117 -3078
rect -1115 -3086 -1113 -3078
rect -1109 -3086 -1107 -3078
rect -1105 -3086 -1104 -3078
rect -1100 -3086 -1099 -3078
rect -1097 -3086 -1092 -3078
rect -1088 -3086 -1083 -3078
rect -1081 -3086 -1080 -3078
rect -1076 -3086 -1075 -3078
rect -1073 -3086 -1072 -3078
rect -1022 -3086 -1021 -3078
rect -1019 -3086 -1018 -3078
rect -931 -3086 -930 -3078
rect -928 -3086 -926 -3078
rect -922 -3086 -920 -3078
rect -918 -3086 -917 -3078
rect -905 -3086 -904 -3078
rect -902 -3086 -901 -3078
rect -897 -3086 -896 -3078
rect -894 -3086 -889 -3078
rect -885 -3086 -880 -3078
rect -878 -3086 -877 -3078
rect -873 -3086 -872 -3078
rect -870 -3086 -868 -3078
rect -864 -3086 -862 -3078
rect -860 -3086 -859 -3078
rect -855 -3086 -854 -3078
rect -852 -3086 -847 -3078
rect -843 -3086 -838 -3078
rect -836 -3086 -835 -3078
rect -831 -3086 -830 -3078
rect -828 -3086 -826 -3078
rect -822 -3086 -820 -3078
rect -818 -3086 -817 -3078
rect -813 -3086 -812 -3078
rect -810 -3086 -805 -3078
rect -801 -3086 -796 -3078
rect -794 -3086 -793 -3078
rect -789 -3086 -788 -3078
rect -786 -3086 -784 -3078
rect -780 -3086 -778 -3078
rect -776 -3086 -775 -3078
rect -771 -3086 -770 -3078
rect -768 -3086 -763 -3078
rect -759 -3086 -754 -3078
rect -752 -3086 -751 -3078
rect -747 -3086 -746 -3078
rect -744 -3086 -743 -3078
rect -573 -3086 -572 -3078
rect -570 -3086 -568 -3078
rect -564 -3086 -562 -3078
rect -560 -3086 -559 -3078
rect -547 -3086 -546 -3078
rect -544 -3086 -543 -3078
rect -539 -3086 -538 -3078
rect -536 -3086 -531 -3078
rect -527 -3086 -522 -3078
rect -520 -3086 -519 -3078
rect -515 -3086 -514 -3078
rect -512 -3086 -510 -3078
rect -506 -3086 -504 -3078
rect -502 -3086 -501 -3078
rect -497 -3086 -496 -3078
rect -494 -3086 -489 -3078
rect -485 -3086 -480 -3078
rect -478 -3086 -477 -3078
rect -473 -3086 -472 -3078
rect -470 -3086 -468 -3078
rect -464 -3086 -462 -3078
rect -460 -3086 -459 -3078
rect -455 -3086 -454 -3078
rect -452 -3086 -447 -3078
rect -443 -3086 -438 -3078
rect -436 -3086 -435 -3078
rect -431 -3086 -430 -3078
rect -428 -3086 -426 -3078
rect -422 -3086 -420 -3078
rect -418 -3086 -417 -3078
rect -413 -3086 -412 -3078
rect -410 -3086 -405 -3078
rect -401 -3086 -396 -3078
rect -394 -3086 -393 -3078
rect -389 -3086 -388 -3078
rect -386 -3086 -385 -3078
rect -325 -3086 -324 -3078
rect -322 -3086 -321 -3078
rect -215 -3086 -214 -3078
rect -212 -3086 -210 -3078
rect -206 -3086 -204 -3078
rect -202 -3086 -201 -3078
rect -189 -3086 -188 -3078
rect -186 -3086 -185 -3078
rect -181 -3086 -180 -3078
rect -178 -3086 -173 -3078
rect -169 -3086 -164 -3078
rect -162 -3086 -161 -3078
rect -157 -3086 -156 -3078
rect -154 -3086 -152 -3078
rect -148 -3086 -146 -3078
rect -144 -3086 -143 -3078
rect -139 -3086 -138 -3078
rect -136 -3086 -131 -3078
rect -127 -3086 -122 -3078
rect -120 -3086 -119 -3078
rect -115 -3086 -114 -3078
rect -112 -3086 -110 -3078
rect -106 -3086 -104 -3078
rect -102 -3086 -101 -3078
rect -97 -3086 -96 -3078
rect -94 -3086 -89 -3078
rect -85 -3086 -80 -3078
rect -78 -3086 -77 -3078
rect -73 -3086 -72 -3078
rect -70 -3086 -68 -3078
rect -64 -3086 -62 -3078
rect -60 -3086 -59 -3078
rect -55 -3086 -54 -3078
rect -52 -3086 -47 -3078
rect -43 -3086 -38 -3078
rect -36 -3086 -35 -3078
rect -31 -3086 -30 -3078
rect -28 -3086 -27 -3078
rect 213 -3086 214 -3078
rect 216 -3086 218 -3078
rect 222 -3086 224 -3078
rect 226 -3086 227 -3078
rect 239 -3086 240 -3078
rect 242 -3086 243 -3078
rect 247 -3086 248 -3078
rect 250 -3086 255 -3078
rect 259 -3086 264 -3078
rect 266 -3086 267 -3078
rect 271 -3086 272 -3078
rect 274 -3086 276 -3078
rect 280 -3086 282 -3078
rect 284 -3086 285 -3078
rect 289 -3086 290 -3078
rect 292 -3086 297 -3078
rect 301 -3086 306 -3078
rect 308 -3086 309 -3078
rect 313 -3086 314 -3078
rect 316 -3086 318 -3078
rect 322 -3086 324 -3078
rect 326 -3086 327 -3078
rect 331 -3086 332 -3078
rect 334 -3086 339 -3078
rect 343 -3086 348 -3078
rect 350 -3086 351 -3078
rect 355 -3086 356 -3078
rect 358 -3086 360 -3078
rect 364 -3086 366 -3078
rect 368 -3086 369 -3078
rect 373 -3086 374 -3078
rect 376 -3086 381 -3078
rect 385 -3086 390 -3078
rect 392 -3086 393 -3078
rect 397 -3086 398 -3078
rect 400 -3086 401 -3078
rect 476 -3086 477 -3078
rect 479 -3086 480 -3078
rect 569 -3086 570 -3078
rect 572 -3086 574 -3078
rect 578 -3086 580 -3078
rect 582 -3086 583 -3078
rect 595 -3086 596 -3078
rect 598 -3086 599 -3078
rect 603 -3086 604 -3078
rect 606 -3086 611 -3078
rect 615 -3086 620 -3078
rect 622 -3086 623 -3078
rect 627 -3086 628 -3078
rect 630 -3086 632 -3078
rect 636 -3086 638 -3078
rect 640 -3086 641 -3078
rect 645 -3086 646 -3078
rect 648 -3086 653 -3078
rect 657 -3086 662 -3078
rect 664 -3086 665 -3078
rect 669 -3086 670 -3078
rect 672 -3086 674 -3078
rect 678 -3086 680 -3078
rect 682 -3086 683 -3078
rect 687 -3086 688 -3078
rect 690 -3086 695 -3078
rect 699 -3086 704 -3078
rect 706 -3086 707 -3078
rect 711 -3086 712 -3078
rect 714 -3086 716 -3078
rect 720 -3086 722 -3078
rect 724 -3086 725 -3078
rect 729 -3086 730 -3078
rect 732 -3086 737 -3078
rect 741 -3086 746 -3078
rect 748 -3086 749 -3078
rect 753 -3086 754 -3078
rect 756 -3086 757 -3078
rect 967 -3086 968 -3078
rect 970 -3086 972 -3078
rect 976 -3086 978 -3078
rect 980 -3086 981 -3078
rect 993 -3086 994 -3078
rect 996 -3086 997 -3078
rect 1001 -3086 1002 -3078
rect 1004 -3086 1009 -3078
rect 1013 -3086 1018 -3078
rect 1020 -3086 1021 -3078
rect 1025 -3086 1026 -3078
rect 1028 -3086 1030 -3078
rect 1034 -3086 1036 -3078
rect 1038 -3086 1039 -3078
rect 1043 -3086 1044 -3078
rect 1046 -3086 1051 -3078
rect 1055 -3086 1060 -3078
rect 1062 -3086 1063 -3078
rect 1067 -3086 1068 -3078
rect 1070 -3086 1072 -3078
rect 1076 -3086 1078 -3078
rect 1080 -3086 1081 -3078
rect 1085 -3086 1086 -3078
rect 1088 -3086 1093 -3078
rect 1097 -3086 1102 -3078
rect 1104 -3086 1105 -3078
rect 1109 -3086 1110 -3078
rect 1112 -3086 1114 -3078
rect 1118 -3086 1120 -3078
rect 1122 -3086 1123 -3078
rect 1127 -3086 1128 -3078
rect 1130 -3086 1135 -3078
rect 1139 -3086 1144 -3078
rect 1146 -3086 1147 -3078
rect 1151 -3086 1152 -3078
rect 1154 -3086 1155 -3078
rect 1203 -3086 1204 -3078
rect 1206 -3086 1207 -3078
rect 1325 -3086 1326 -3078
rect 1328 -3086 1330 -3078
rect 1334 -3086 1336 -3078
rect 1338 -3086 1339 -3078
rect 1351 -3086 1352 -3078
rect 1354 -3086 1355 -3078
rect 1359 -3086 1360 -3078
rect 1362 -3086 1367 -3078
rect 1371 -3086 1376 -3078
rect 1378 -3086 1379 -3078
rect 1383 -3086 1384 -3078
rect 1386 -3086 1388 -3078
rect 1392 -3086 1394 -3078
rect 1396 -3086 1397 -3078
rect 1401 -3086 1402 -3078
rect 1404 -3086 1409 -3078
rect 1413 -3086 1418 -3078
rect 1420 -3086 1421 -3078
rect 1425 -3086 1426 -3078
rect 1428 -3086 1430 -3078
rect 1434 -3086 1436 -3078
rect 1438 -3086 1439 -3078
rect 1443 -3086 1444 -3078
rect 1446 -3086 1451 -3078
rect 1455 -3086 1460 -3078
rect 1462 -3086 1463 -3078
rect 1467 -3086 1468 -3078
rect 1470 -3086 1472 -3078
rect 1476 -3086 1478 -3078
rect 1480 -3086 1481 -3078
rect 1485 -3086 1486 -3078
rect 1488 -3086 1493 -3078
rect 1497 -3086 1502 -3078
rect 1504 -3086 1505 -3078
rect 1509 -3086 1510 -3078
rect 1512 -3086 1513 -3078
rect -1260 -3207 -1259 -3199
rect -1257 -3207 -1255 -3199
rect -1251 -3207 -1249 -3199
rect -1247 -3207 -1246 -3199
rect -1234 -3207 -1233 -3199
rect -1231 -3207 -1230 -3199
rect -1226 -3207 -1225 -3199
rect -1223 -3207 -1218 -3199
rect -1214 -3207 -1209 -3199
rect -1207 -3207 -1206 -3199
rect -1202 -3207 -1201 -3199
rect -1199 -3207 -1197 -3199
rect -1193 -3207 -1191 -3199
rect -1189 -3207 -1188 -3199
rect -1184 -3207 -1183 -3199
rect -1181 -3207 -1176 -3199
rect -1172 -3207 -1167 -3199
rect -1165 -3207 -1164 -3199
rect -1160 -3207 -1159 -3199
rect -1157 -3207 -1155 -3199
rect -1151 -3207 -1149 -3199
rect -1147 -3207 -1146 -3199
rect -1142 -3207 -1141 -3199
rect -1139 -3207 -1134 -3199
rect -1130 -3207 -1125 -3199
rect -1123 -3207 -1122 -3199
rect -1118 -3207 -1117 -3199
rect -1115 -3207 -1113 -3199
rect -1109 -3207 -1107 -3199
rect -1105 -3207 -1104 -3199
rect -1100 -3207 -1099 -3199
rect -1097 -3207 -1092 -3199
rect -1088 -3207 -1083 -3199
rect -1081 -3207 -1080 -3199
rect -1076 -3207 -1075 -3199
rect -1073 -3207 -1072 -3199
rect -931 -3207 -930 -3199
rect -928 -3207 -926 -3199
rect -922 -3207 -920 -3199
rect -918 -3207 -917 -3199
rect -905 -3207 -904 -3199
rect -902 -3207 -901 -3199
rect -897 -3207 -896 -3199
rect -894 -3207 -889 -3199
rect -885 -3207 -880 -3199
rect -878 -3207 -877 -3199
rect -873 -3207 -872 -3199
rect -870 -3207 -868 -3199
rect -864 -3207 -862 -3199
rect -860 -3207 -859 -3199
rect -855 -3207 -854 -3199
rect -852 -3207 -847 -3199
rect -843 -3207 -838 -3199
rect -836 -3207 -835 -3199
rect -831 -3207 -830 -3199
rect -828 -3207 -826 -3199
rect -822 -3207 -820 -3199
rect -818 -3207 -817 -3199
rect -813 -3207 -812 -3199
rect -810 -3207 -805 -3199
rect -801 -3207 -796 -3199
rect -794 -3207 -793 -3199
rect -789 -3207 -788 -3199
rect -786 -3207 -784 -3199
rect -780 -3207 -778 -3199
rect -776 -3207 -775 -3199
rect -771 -3207 -770 -3199
rect -768 -3207 -763 -3199
rect -759 -3207 -754 -3199
rect -752 -3207 -751 -3199
rect -747 -3207 -746 -3199
rect -744 -3207 -743 -3199
rect -573 -3207 -572 -3199
rect -570 -3207 -568 -3199
rect -564 -3207 -562 -3199
rect -560 -3207 -559 -3199
rect -547 -3207 -546 -3199
rect -544 -3207 -543 -3199
rect -539 -3207 -538 -3199
rect -536 -3207 -531 -3199
rect -527 -3207 -522 -3199
rect -520 -3207 -519 -3199
rect -515 -3207 -514 -3199
rect -512 -3207 -510 -3199
rect -506 -3207 -504 -3199
rect -502 -3207 -501 -3199
rect -497 -3207 -496 -3199
rect -494 -3207 -489 -3199
rect -485 -3207 -480 -3199
rect -478 -3207 -477 -3199
rect -473 -3207 -472 -3199
rect -470 -3207 -468 -3199
rect -464 -3207 -462 -3199
rect -460 -3207 -459 -3199
rect -455 -3207 -454 -3199
rect -452 -3207 -447 -3199
rect -443 -3207 -438 -3199
rect -436 -3207 -435 -3199
rect -431 -3207 -430 -3199
rect -428 -3207 -426 -3199
rect -422 -3207 -420 -3199
rect -418 -3207 -417 -3199
rect -413 -3207 -412 -3199
rect -410 -3207 -405 -3199
rect -401 -3207 -396 -3199
rect -394 -3207 -393 -3199
rect -389 -3207 -388 -3199
rect -386 -3207 -385 -3199
rect -215 -3207 -214 -3199
rect -212 -3207 -210 -3199
rect -206 -3207 -204 -3199
rect -202 -3207 -201 -3199
rect -189 -3207 -188 -3199
rect -186 -3207 -185 -3199
rect -181 -3207 -180 -3199
rect -178 -3207 -173 -3199
rect -169 -3207 -164 -3199
rect -162 -3207 -161 -3199
rect -157 -3207 -156 -3199
rect -154 -3207 -152 -3199
rect -148 -3207 -146 -3199
rect -144 -3207 -143 -3199
rect -139 -3207 -138 -3199
rect -136 -3207 -131 -3199
rect -127 -3207 -122 -3199
rect -120 -3207 -119 -3199
rect -115 -3207 -114 -3199
rect -112 -3207 -110 -3199
rect -106 -3207 -104 -3199
rect -102 -3207 -101 -3199
rect -97 -3207 -96 -3199
rect -94 -3207 -89 -3199
rect -85 -3207 -80 -3199
rect -78 -3207 -77 -3199
rect -73 -3207 -72 -3199
rect -70 -3207 -68 -3199
rect -64 -3207 -62 -3199
rect -60 -3207 -59 -3199
rect -55 -3207 -54 -3199
rect -52 -3207 -47 -3199
rect -43 -3207 -38 -3199
rect -36 -3207 -35 -3199
rect -31 -3207 -30 -3199
rect -28 -3207 -27 -3199
rect 213 -3207 214 -3199
rect 216 -3207 218 -3199
rect 222 -3207 224 -3199
rect 226 -3207 227 -3199
rect 239 -3207 240 -3199
rect 242 -3207 243 -3199
rect 247 -3207 248 -3199
rect 250 -3207 255 -3199
rect 259 -3207 264 -3199
rect 266 -3207 267 -3199
rect 271 -3207 272 -3199
rect 274 -3207 276 -3199
rect 280 -3207 282 -3199
rect 284 -3207 285 -3199
rect 289 -3207 290 -3199
rect 292 -3207 297 -3199
rect 301 -3207 306 -3199
rect 308 -3207 309 -3199
rect 313 -3207 314 -3199
rect 316 -3207 318 -3199
rect 322 -3207 324 -3199
rect 326 -3207 327 -3199
rect 331 -3207 332 -3199
rect 334 -3207 339 -3199
rect 343 -3207 348 -3199
rect 350 -3207 351 -3199
rect 355 -3207 356 -3199
rect 358 -3207 360 -3199
rect 364 -3207 366 -3199
rect 368 -3207 369 -3199
rect 373 -3207 374 -3199
rect 376 -3207 381 -3199
rect 385 -3207 390 -3199
rect 392 -3207 393 -3199
rect 397 -3207 398 -3199
rect 400 -3207 401 -3199
rect 569 -3207 570 -3199
rect 572 -3207 574 -3199
rect 578 -3207 580 -3199
rect 582 -3207 583 -3199
rect 595 -3207 596 -3199
rect 598 -3207 599 -3199
rect 603 -3207 604 -3199
rect 606 -3207 611 -3199
rect 615 -3207 620 -3199
rect 622 -3207 623 -3199
rect 627 -3207 628 -3199
rect 630 -3207 632 -3199
rect 636 -3207 638 -3199
rect 640 -3207 641 -3199
rect 645 -3207 646 -3199
rect 648 -3207 653 -3199
rect 657 -3207 662 -3199
rect 664 -3207 665 -3199
rect 669 -3207 670 -3199
rect 672 -3207 674 -3199
rect 678 -3207 680 -3199
rect 682 -3207 683 -3199
rect 687 -3207 688 -3199
rect 690 -3207 695 -3199
rect 699 -3207 704 -3199
rect 706 -3207 707 -3199
rect 711 -3207 712 -3199
rect 714 -3207 716 -3199
rect 720 -3207 722 -3199
rect 724 -3207 725 -3199
rect 729 -3207 730 -3199
rect 732 -3207 737 -3199
rect 741 -3207 746 -3199
rect 748 -3207 749 -3199
rect 753 -3207 754 -3199
rect 756 -3207 757 -3199
rect 967 -3207 968 -3199
rect 970 -3207 972 -3199
rect 976 -3207 978 -3199
rect 980 -3207 981 -3199
rect 993 -3207 994 -3199
rect 996 -3207 997 -3199
rect 1001 -3207 1002 -3199
rect 1004 -3207 1009 -3199
rect 1013 -3207 1018 -3199
rect 1020 -3207 1021 -3199
rect 1025 -3207 1026 -3199
rect 1028 -3207 1030 -3199
rect 1034 -3207 1036 -3199
rect 1038 -3207 1039 -3199
rect 1043 -3207 1044 -3199
rect 1046 -3207 1051 -3199
rect 1055 -3207 1060 -3199
rect 1062 -3207 1063 -3199
rect 1067 -3207 1068 -3199
rect 1070 -3207 1072 -3199
rect 1076 -3207 1078 -3199
rect 1080 -3207 1081 -3199
rect 1085 -3207 1086 -3199
rect 1088 -3207 1093 -3199
rect 1097 -3207 1102 -3199
rect 1104 -3207 1105 -3199
rect 1109 -3207 1110 -3199
rect 1112 -3207 1114 -3199
rect 1118 -3207 1120 -3199
rect 1122 -3207 1123 -3199
rect 1127 -3207 1128 -3199
rect 1130 -3207 1135 -3199
rect 1139 -3207 1144 -3199
rect 1146 -3207 1147 -3199
rect 1151 -3207 1152 -3199
rect 1154 -3207 1155 -3199
rect 1325 -3207 1326 -3199
rect 1328 -3207 1330 -3199
rect 1334 -3207 1336 -3199
rect 1338 -3207 1339 -3199
rect 1351 -3207 1352 -3199
rect 1354 -3207 1355 -3199
rect 1359 -3207 1360 -3199
rect 1362 -3207 1367 -3199
rect 1371 -3207 1376 -3199
rect 1378 -3207 1379 -3199
rect 1383 -3207 1384 -3199
rect 1386 -3207 1388 -3199
rect 1392 -3207 1394 -3199
rect 1396 -3207 1397 -3199
rect 1401 -3207 1402 -3199
rect 1404 -3207 1409 -3199
rect 1413 -3207 1418 -3199
rect 1420 -3207 1421 -3199
rect 1425 -3207 1426 -3199
rect 1428 -3207 1430 -3199
rect 1434 -3207 1436 -3199
rect 1438 -3207 1439 -3199
rect 1443 -3207 1444 -3199
rect 1446 -3207 1451 -3199
rect 1455 -3207 1460 -3199
rect 1462 -3207 1463 -3199
rect 1467 -3207 1468 -3199
rect 1470 -3207 1472 -3199
rect 1476 -3207 1478 -3199
rect 1480 -3207 1481 -3199
rect 1485 -3207 1486 -3199
rect 1488 -3207 1493 -3199
rect 1497 -3207 1502 -3199
rect 1504 -3207 1505 -3199
rect 1509 -3207 1510 -3199
rect 1512 -3207 1513 -3199
rect -1260 -3321 -1259 -3313
rect -1257 -3321 -1255 -3313
rect -1251 -3321 -1249 -3313
rect -1247 -3321 -1246 -3313
rect -1234 -3321 -1233 -3313
rect -1231 -3321 -1230 -3313
rect -1226 -3321 -1225 -3313
rect -1223 -3321 -1218 -3313
rect -1214 -3321 -1209 -3313
rect -1207 -3321 -1206 -3313
rect -1202 -3321 -1201 -3313
rect -1199 -3321 -1197 -3313
rect -1193 -3321 -1191 -3313
rect -1189 -3321 -1188 -3313
rect -1184 -3321 -1183 -3313
rect -1181 -3321 -1176 -3313
rect -1172 -3321 -1167 -3313
rect -1165 -3321 -1164 -3313
rect -1160 -3321 -1159 -3313
rect -1157 -3321 -1155 -3313
rect -1151 -3321 -1149 -3313
rect -1147 -3321 -1146 -3313
rect -1142 -3321 -1141 -3313
rect -1139 -3321 -1134 -3313
rect -1130 -3321 -1125 -3313
rect -1123 -3321 -1122 -3313
rect -1118 -3321 -1117 -3313
rect -1115 -3321 -1113 -3313
rect -1109 -3321 -1107 -3313
rect -1105 -3321 -1104 -3313
rect -1100 -3321 -1099 -3313
rect -1097 -3321 -1092 -3313
rect -1088 -3321 -1083 -3313
rect -1081 -3321 -1080 -3313
rect -1076 -3321 -1075 -3313
rect -1073 -3321 -1072 -3313
rect -931 -3321 -930 -3313
rect -928 -3321 -926 -3313
rect -922 -3321 -920 -3313
rect -918 -3321 -917 -3313
rect -905 -3321 -904 -3313
rect -902 -3321 -901 -3313
rect -897 -3321 -896 -3313
rect -894 -3321 -889 -3313
rect -885 -3321 -880 -3313
rect -878 -3321 -877 -3313
rect -873 -3321 -872 -3313
rect -870 -3321 -868 -3313
rect -864 -3321 -862 -3313
rect -860 -3321 -859 -3313
rect -855 -3321 -854 -3313
rect -852 -3321 -847 -3313
rect -843 -3321 -838 -3313
rect -836 -3321 -835 -3313
rect -831 -3321 -830 -3313
rect -828 -3321 -826 -3313
rect -822 -3321 -820 -3313
rect -818 -3321 -817 -3313
rect -813 -3321 -812 -3313
rect -810 -3321 -805 -3313
rect -801 -3321 -796 -3313
rect -794 -3321 -793 -3313
rect -789 -3321 -788 -3313
rect -786 -3321 -784 -3313
rect -780 -3321 -778 -3313
rect -776 -3321 -775 -3313
rect -771 -3321 -770 -3313
rect -768 -3321 -763 -3313
rect -759 -3321 -754 -3313
rect -752 -3321 -751 -3313
rect -747 -3321 -746 -3313
rect -744 -3321 -743 -3313
rect -573 -3321 -572 -3313
rect -570 -3321 -568 -3313
rect -564 -3321 -562 -3313
rect -560 -3321 -559 -3313
rect -547 -3321 -546 -3313
rect -544 -3321 -543 -3313
rect -539 -3321 -538 -3313
rect -536 -3321 -531 -3313
rect -527 -3321 -522 -3313
rect -520 -3321 -519 -3313
rect -515 -3321 -514 -3313
rect -512 -3321 -510 -3313
rect -506 -3321 -504 -3313
rect -502 -3321 -501 -3313
rect -497 -3321 -496 -3313
rect -494 -3321 -489 -3313
rect -485 -3321 -480 -3313
rect -478 -3321 -477 -3313
rect -473 -3321 -472 -3313
rect -470 -3321 -468 -3313
rect -464 -3321 -462 -3313
rect -460 -3321 -459 -3313
rect -455 -3321 -454 -3313
rect -452 -3321 -447 -3313
rect -443 -3321 -438 -3313
rect -436 -3321 -435 -3313
rect -431 -3321 -430 -3313
rect -428 -3321 -426 -3313
rect -422 -3321 -420 -3313
rect -418 -3321 -417 -3313
rect -413 -3321 -412 -3313
rect -410 -3321 -405 -3313
rect -401 -3321 -396 -3313
rect -394 -3321 -393 -3313
rect -389 -3321 -388 -3313
rect -386 -3321 -385 -3313
rect -1335 -3438 -1334 -3430
rect -1332 -3438 -1331 -3430
rect -1327 -3438 -1326 -3430
rect -1324 -3438 -1322 -3430
rect -1318 -3438 -1316 -3430
rect -1314 -3438 -1313 -3430
rect -931 -3438 -930 -3430
rect -928 -3438 -927 -3430
rect -923 -3438 -922 -3430
rect -920 -3438 -918 -3430
rect -914 -3438 -912 -3430
rect -910 -3438 -909 -3430
rect -573 -3438 -572 -3430
rect -570 -3438 -569 -3430
rect -565 -3438 -564 -3430
rect -562 -3438 -560 -3430
rect -556 -3438 -554 -3430
rect -552 -3438 -551 -3430
rect -215 -3438 -214 -3430
rect -212 -3438 -211 -3430
rect -207 -3438 -206 -3430
rect -204 -3438 -202 -3430
rect -198 -3438 -196 -3430
rect -194 -3438 -193 -3430
rect 213 -3438 214 -3430
rect 216 -3438 217 -3430
rect 221 -3438 222 -3430
rect 224 -3438 226 -3430
rect 230 -3438 232 -3430
rect 234 -3438 235 -3430
rect 569 -3438 570 -3430
rect 572 -3438 573 -3430
rect 577 -3438 578 -3430
rect 580 -3438 582 -3430
rect 586 -3438 588 -3430
rect 590 -3438 591 -3430
rect 967 -3438 968 -3430
rect 970 -3438 971 -3430
rect 975 -3438 976 -3430
rect 978 -3438 980 -3430
rect 984 -3438 986 -3430
rect 988 -3438 989 -3430
rect 1325 -3438 1326 -3430
rect 1328 -3438 1329 -3430
rect 1333 -3438 1334 -3430
rect 1336 -3438 1338 -3430
rect 1342 -3438 1344 -3430
rect 1346 -3438 1347 -3430
rect -1260 -3562 -1259 -3554
rect -1257 -3562 -1255 -3554
rect -1251 -3562 -1249 -3554
rect -1247 -3562 -1246 -3554
rect -1234 -3562 -1233 -3554
rect -1231 -3562 -1223 -3554
rect -1221 -3562 -1220 -3554
rect -1216 -3562 -1215 -3554
rect -1213 -3562 -1205 -3554
rect -1203 -3562 -1198 -3554
rect -1194 -3562 -1189 -3554
rect -1187 -3562 -1186 -3554
rect -1182 -3562 -1181 -3554
rect -1179 -3562 -1177 -3554
rect -1173 -3562 -1171 -3554
rect -1169 -3562 -1168 -3554
rect -931 -3562 -930 -3554
rect -928 -3562 -926 -3554
rect -922 -3562 -920 -3554
rect -918 -3562 -917 -3554
rect -905 -3562 -904 -3554
rect -902 -3562 -900 -3554
rect -896 -3562 -894 -3554
rect -892 -3562 -891 -3554
rect -879 -3562 -878 -3554
rect -876 -3562 -868 -3554
rect -866 -3562 -865 -3554
rect -861 -3562 -860 -3554
rect -858 -3562 -850 -3554
rect -848 -3562 -843 -3554
rect -839 -3562 -834 -3554
rect -832 -3562 -831 -3554
rect -827 -3562 -826 -3554
rect -824 -3562 -822 -3554
rect -818 -3562 -816 -3554
rect -814 -3562 -813 -3554
rect -801 -3562 -800 -3554
rect -798 -3562 -790 -3554
rect -788 -3562 -787 -3554
rect -783 -3562 -782 -3554
rect -780 -3562 -772 -3554
rect -770 -3562 -765 -3554
rect -761 -3562 -756 -3554
rect -754 -3562 -753 -3554
rect -749 -3562 -748 -3554
rect -746 -3562 -741 -3554
rect -737 -3562 -732 -3554
rect -730 -3562 -729 -3554
rect -717 -3562 -716 -3554
rect -714 -3562 -708 -3554
rect -706 -3562 -704 -3554
rect -700 -3562 -698 -3554
rect -696 -3562 -695 -3554
rect -573 -3562 -572 -3554
rect -570 -3562 -568 -3554
rect -564 -3562 -562 -3554
rect -560 -3562 -559 -3554
rect -547 -3562 -546 -3554
rect -544 -3562 -542 -3554
rect -538 -3562 -536 -3554
rect -534 -3562 -533 -3554
rect -521 -3562 -520 -3554
rect -518 -3562 -510 -3554
rect -508 -3562 -507 -3554
rect -503 -3562 -502 -3554
rect -500 -3562 -492 -3554
rect -490 -3562 -485 -3554
rect -481 -3562 -476 -3554
rect -474 -3562 -473 -3554
rect -469 -3562 -468 -3554
rect -466 -3562 -464 -3554
rect -460 -3562 -458 -3554
rect -456 -3562 -455 -3554
rect -443 -3562 -442 -3554
rect -440 -3562 -432 -3554
rect -430 -3562 -429 -3554
rect -425 -3562 -424 -3554
rect -422 -3562 -414 -3554
rect -412 -3562 -407 -3554
rect -403 -3562 -398 -3554
rect -396 -3562 -395 -3554
rect -391 -3562 -390 -3554
rect -388 -3562 -383 -3554
rect -379 -3562 -374 -3554
rect -372 -3562 -371 -3554
rect -359 -3562 -358 -3554
rect -356 -3562 -350 -3554
rect -348 -3562 -346 -3554
rect -342 -3562 -340 -3554
rect -338 -3562 -337 -3554
rect -215 -3562 -214 -3554
rect -212 -3562 -210 -3554
rect -206 -3562 -204 -3554
rect -202 -3562 -201 -3554
rect -189 -3562 -188 -3554
rect -186 -3562 -184 -3554
rect -180 -3562 -178 -3554
rect -176 -3562 -175 -3554
rect -163 -3562 -162 -3554
rect -160 -3562 -152 -3554
rect -150 -3562 -149 -3554
rect -145 -3562 -144 -3554
rect -142 -3562 -134 -3554
rect -132 -3562 -127 -3554
rect -123 -3562 -118 -3554
rect -116 -3562 -115 -3554
rect -111 -3562 -110 -3554
rect -108 -3562 -106 -3554
rect -102 -3562 -100 -3554
rect -98 -3562 -97 -3554
rect -85 -3562 -84 -3554
rect -82 -3562 -74 -3554
rect -72 -3562 -71 -3554
rect -67 -3562 -66 -3554
rect -64 -3562 -56 -3554
rect -54 -3562 -49 -3554
rect -45 -3562 -40 -3554
rect -38 -3562 -37 -3554
rect -33 -3562 -32 -3554
rect -30 -3562 -25 -3554
rect -21 -3562 -16 -3554
rect -14 -3562 -13 -3554
rect -1 -3562 0 -3554
rect 2 -3562 8 -3554
rect 10 -3562 12 -3554
rect 16 -3562 18 -3554
rect 20 -3562 21 -3554
rect 213 -3562 214 -3554
rect 216 -3562 218 -3554
rect 222 -3562 224 -3554
rect 226 -3562 227 -3554
rect 239 -3562 240 -3554
rect 242 -3562 244 -3554
rect 248 -3562 250 -3554
rect 252 -3562 253 -3554
rect 265 -3562 266 -3554
rect 268 -3562 276 -3554
rect 278 -3562 279 -3554
rect 283 -3562 284 -3554
rect 286 -3562 294 -3554
rect 296 -3562 301 -3554
rect 305 -3562 310 -3554
rect 312 -3562 313 -3554
rect 317 -3562 318 -3554
rect 320 -3562 322 -3554
rect 326 -3562 328 -3554
rect 330 -3562 331 -3554
rect 343 -3562 344 -3554
rect 346 -3562 354 -3554
rect 356 -3562 357 -3554
rect 361 -3562 362 -3554
rect 364 -3562 372 -3554
rect 374 -3562 379 -3554
rect 383 -3562 388 -3554
rect 390 -3562 391 -3554
rect 395 -3562 396 -3554
rect 398 -3562 403 -3554
rect 407 -3562 412 -3554
rect 414 -3562 415 -3554
rect 427 -3562 428 -3554
rect 430 -3562 436 -3554
rect 438 -3562 440 -3554
rect 444 -3562 446 -3554
rect 448 -3562 449 -3554
rect 569 -3562 570 -3554
rect 572 -3562 574 -3554
rect 578 -3562 580 -3554
rect 582 -3562 583 -3554
rect 595 -3562 596 -3554
rect 598 -3562 600 -3554
rect 604 -3562 606 -3554
rect 608 -3562 609 -3554
rect 621 -3562 622 -3554
rect 624 -3562 632 -3554
rect 634 -3562 635 -3554
rect 639 -3562 640 -3554
rect 642 -3562 650 -3554
rect 652 -3562 657 -3554
rect 661 -3562 666 -3554
rect 668 -3562 669 -3554
rect 673 -3562 674 -3554
rect 676 -3562 678 -3554
rect 682 -3562 684 -3554
rect 686 -3562 687 -3554
rect 699 -3562 700 -3554
rect 702 -3562 710 -3554
rect 712 -3562 713 -3554
rect 717 -3562 718 -3554
rect 720 -3562 728 -3554
rect 730 -3562 735 -3554
rect 739 -3562 744 -3554
rect 746 -3562 747 -3554
rect 751 -3562 752 -3554
rect 754 -3562 759 -3554
rect 763 -3562 768 -3554
rect 770 -3562 771 -3554
rect 783 -3562 784 -3554
rect 786 -3562 792 -3554
rect 794 -3562 796 -3554
rect 800 -3562 802 -3554
rect 804 -3562 805 -3554
rect 967 -3562 968 -3554
rect 970 -3562 972 -3554
rect 976 -3562 978 -3554
rect 980 -3562 981 -3554
rect 993 -3562 994 -3554
rect 996 -3562 998 -3554
rect 1002 -3562 1004 -3554
rect 1006 -3562 1007 -3554
rect 1019 -3562 1020 -3554
rect 1022 -3562 1030 -3554
rect 1032 -3562 1033 -3554
rect 1037 -3562 1038 -3554
rect 1040 -3562 1048 -3554
rect 1050 -3562 1055 -3554
rect 1059 -3562 1064 -3554
rect 1066 -3562 1067 -3554
rect 1071 -3562 1072 -3554
rect 1074 -3562 1076 -3554
rect 1080 -3562 1082 -3554
rect 1084 -3562 1085 -3554
rect 1097 -3562 1098 -3554
rect 1100 -3562 1108 -3554
rect 1110 -3562 1111 -3554
rect 1115 -3562 1116 -3554
rect 1118 -3562 1126 -3554
rect 1128 -3562 1133 -3554
rect 1137 -3562 1142 -3554
rect 1144 -3562 1145 -3554
rect 1149 -3562 1150 -3554
rect 1152 -3562 1157 -3554
rect 1161 -3562 1166 -3554
rect 1168 -3562 1169 -3554
rect 1181 -3562 1182 -3554
rect 1184 -3562 1190 -3554
rect 1192 -3562 1194 -3554
rect 1198 -3562 1200 -3554
rect 1202 -3562 1203 -3554
rect 1325 -3562 1326 -3554
rect 1328 -3562 1330 -3554
rect 1334 -3562 1336 -3554
rect 1338 -3562 1339 -3554
rect 1351 -3562 1352 -3554
rect 1354 -3562 1356 -3554
rect 1360 -3562 1362 -3554
rect 1364 -3562 1365 -3554
rect 1377 -3562 1378 -3554
rect 1380 -3562 1388 -3554
rect 1390 -3562 1391 -3554
rect 1395 -3562 1396 -3554
rect 1398 -3562 1406 -3554
rect 1408 -3562 1413 -3554
rect 1417 -3562 1422 -3554
rect 1424 -3562 1425 -3554
rect 1429 -3562 1430 -3554
rect 1432 -3562 1434 -3554
rect 1438 -3562 1440 -3554
rect 1442 -3562 1443 -3554
rect 1455 -3562 1456 -3554
rect 1458 -3562 1466 -3554
rect 1468 -3562 1469 -3554
rect 1473 -3562 1474 -3554
rect 1476 -3562 1484 -3554
rect 1486 -3562 1491 -3554
rect 1495 -3562 1500 -3554
rect 1502 -3562 1503 -3554
rect 1507 -3562 1508 -3554
rect 1510 -3562 1515 -3554
rect 1519 -3562 1524 -3554
rect 1526 -3562 1527 -3554
rect 1539 -3562 1540 -3554
rect 1542 -3562 1548 -3554
rect 1550 -3562 1552 -3554
rect 1556 -3562 1558 -3554
rect 1560 -3562 1561 -3554
rect -1260 -3692 -1259 -3684
rect -1257 -3692 -1255 -3684
rect -1251 -3692 -1249 -3684
rect -1247 -3692 -1246 -3684
rect -1234 -3692 -1233 -3684
rect -1231 -3692 -1230 -3684
rect -1226 -3692 -1225 -3684
rect -1223 -3692 -1218 -3684
rect -1214 -3692 -1209 -3684
rect -1207 -3692 -1206 -3684
rect -1202 -3692 -1201 -3684
rect -1199 -3692 -1197 -3684
rect -1193 -3692 -1191 -3684
rect -1189 -3692 -1188 -3684
rect -1184 -3692 -1183 -3684
rect -1181 -3692 -1176 -3684
rect -1172 -3692 -1167 -3684
rect -1165 -3692 -1164 -3684
rect -1160 -3692 -1159 -3684
rect -1157 -3692 -1155 -3684
rect -1151 -3692 -1149 -3684
rect -1147 -3692 -1146 -3684
rect -1142 -3692 -1141 -3684
rect -1139 -3692 -1134 -3684
rect -1130 -3692 -1125 -3684
rect -1123 -3692 -1122 -3684
rect -1118 -3692 -1117 -3684
rect -1115 -3692 -1113 -3684
rect -1109 -3692 -1107 -3684
rect -1105 -3692 -1104 -3684
rect -1100 -3692 -1099 -3684
rect -1097 -3692 -1092 -3684
rect -1088 -3692 -1083 -3684
rect -1081 -3692 -1080 -3684
rect -1076 -3692 -1075 -3684
rect -1073 -3692 -1072 -3684
rect -931 -3692 -930 -3684
rect -928 -3692 -926 -3684
rect -922 -3692 -920 -3684
rect -918 -3692 -917 -3684
rect -905 -3692 -904 -3684
rect -902 -3692 -901 -3684
rect -897 -3692 -896 -3684
rect -894 -3692 -889 -3684
rect -885 -3692 -880 -3684
rect -878 -3692 -877 -3684
rect -873 -3692 -872 -3684
rect -870 -3692 -868 -3684
rect -864 -3692 -862 -3684
rect -860 -3692 -859 -3684
rect -855 -3692 -854 -3684
rect -852 -3692 -847 -3684
rect -843 -3692 -838 -3684
rect -836 -3692 -835 -3684
rect -831 -3692 -830 -3684
rect -828 -3692 -826 -3684
rect -822 -3692 -820 -3684
rect -818 -3692 -817 -3684
rect -813 -3692 -812 -3684
rect -810 -3692 -805 -3684
rect -801 -3692 -796 -3684
rect -794 -3692 -793 -3684
rect -789 -3692 -788 -3684
rect -786 -3692 -784 -3684
rect -780 -3692 -778 -3684
rect -776 -3692 -775 -3684
rect -771 -3692 -770 -3684
rect -768 -3692 -763 -3684
rect -759 -3692 -754 -3684
rect -752 -3692 -751 -3684
rect -747 -3692 -746 -3684
rect -744 -3692 -743 -3684
rect -573 -3692 -572 -3684
rect -570 -3692 -568 -3684
rect -564 -3692 -562 -3684
rect -560 -3692 -559 -3684
rect -547 -3692 -546 -3684
rect -544 -3692 -543 -3684
rect -539 -3692 -538 -3684
rect -536 -3692 -531 -3684
rect -527 -3692 -522 -3684
rect -520 -3692 -519 -3684
rect -515 -3692 -514 -3684
rect -512 -3692 -510 -3684
rect -506 -3692 -504 -3684
rect -502 -3692 -501 -3684
rect -497 -3692 -496 -3684
rect -494 -3692 -489 -3684
rect -485 -3692 -480 -3684
rect -478 -3692 -477 -3684
rect -473 -3692 -472 -3684
rect -470 -3692 -468 -3684
rect -464 -3692 -462 -3684
rect -460 -3692 -459 -3684
rect -455 -3692 -454 -3684
rect -452 -3692 -447 -3684
rect -443 -3692 -438 -3684
rect -436 -3692 -435 -3684
rect -431 -3692 -430 -3684
rect -428 -3692 -426 -3684
rect -422 -3692 -420 -3684
rect -418 -3692 -417 -3684
rect -413 -3692 -412 -3684
rect -410 -3692 -405 -3684
rect -401 -3692 -396 -3684
rect -394 -3692 -393 -3684
rect -389 -3692 -388 -3684
rect -386 -3692 -385 -3684
rect -215 -3692 -214 -3684
rect -212 -3692 -210 -3684
rect -206 -3692 -204 -3684
rect -202 -3692 -201 -3684
rect -189 -3692 -188 -3684
rect -186 -3692 -185 -3684
rect -181 -3692 -180 -3684
rect -178 -3692 -173 -3684
rect -169 -3692 -164 -3684
rect -162 -3692 -161 -3684
rect -157 -3692 -156 -3684
rect -154 -3692 -152 -3684
rect -148 -3692 -146 -3684
rect -144 -3692 -143 -3684
rect -139 -3692 -138 -3684
rect -136 -3692 -131 -3684
rect -127 -3692 -122 -3684
rect -120 -3692 -119 -3684
rect -115 -3692 -114 -3684
rect -112 -3692 -110 -3684
rect -106 -3692 -104 -3684
rect -102 -3692 -101 -3684
rect -97 -3692 -96 -3684
rect -94 -3692 -89 -3684
rect -85 -3692 -80 -3684
rect -78 -3692 -77 -3684
rect -73 -3692 -72 -3684
rect -70 -3692 -68 -3684
rect -64 -3692 -62 -3684
rect -60 -3692 -59 -3684
rect -55 -3692 -54 -3684
rect -52 -3692 -47 -3684
rect -43 -3692 -38 -3684
rect -36 -3692 -35 -3684
rect -31 -3692 -30 -3684
rect -28 -3692 -27 -3684
rect 72 -3831 73 -3799
rect 75 -3831 76 -3799
rect -1260 -3923 -1259 -3915
rect -1257 -3923 -1255 -3915
rect -1251 -3923 -1249 -3915
rect -1247 -3923 -1246 -3915
rect -1234 -3923 -1233 -3915
rect -1231 -3923 -1230 -3915
rect -1226 -3923 -1225 -3915
rect -1223 -3923 -1218 -3915
rect -1214 -3923 -1209 -3915
rect -1207 -3923 -1206 -3915
rect -1202 -3923 -1201 -3915
rect -1199 -3923 -1197 -3915
rect -1193 -3923 -1191 -3915
rect -1189 -3923 -1188 -3915
rect -1184 -3923 -1183 -3915
rect -1181 -3923 -1176 -3915
rect -1172 -3923 -1167 -3915
rect -1165 -3923 -1164 -3915
rect -1160 -3923 -1159 -3915
rect -1157 -3923 -1155 -3915
rect -1151 -3923 -1149 -3915
rect -1147 -3923 -1146 -3915
rect -1142 -3923 -1141 -3915
rect -1139 -3923 -1134 -3915
rect -1130 -3923 -1125 -3915
rect -1123 -3923 -1122 -3915
rect -1118 -3923 -1117 -3915
rect -1115 -3923 -1113 -3915
rect -1109 -3923 -1107 -3915
rect -1105 -3923 -1104 -3915
rect -1100 -3923 -1099 -3915
rect -1097 -3923 -1092 -3915
rect -1088 -3923 -1083 -3915
rect -1081 -3923 -1080 -3915
rect -1076 -3923 -1075 -3915
rect -1073 -3923 -1072 -3915
rect -931 -3923 -930 -3915
rect -928 -3923 -926 -3915
rect -922 -3923 -920 -3915
rect -918 -3923 -917 -3915
rect -905 -3923 -904 -3915
rect -902 -3923 -901 -3915
rect -897 -3923 -896 -3915
rect -894 -3923 -889 -3915
rect -885 -3923 -880 -3915
rect -878 -3923 -877 -3915
rect -873 -3923 -872 -3915
rect -870 -3923 -868 -3915
rect -864 -3923 -862 -3915
rect -860 -3923 -859 -3915
rect -855 -3923 -854 -3915
rect -852 -3923 -847 -3915
rect -843 -3923 -838 -3915
rect -836 -3923 -835 -3915
rect -831 -3923 -830 -3915
rect -828 -3923 -826 -3915
rect -822 -3923 -820 -3915
rect -818 -3923 -817 -3915
rect -813 -3923 -812 -3915
rect -810 -3923 -805 -3915
rect -801 -3923 -796 -3915
rect -794 -3923 -793 -3915
rect -789 -3923 -788 -3915
rect -786 -3923 -784 -3915
rect -780 -3923 -778 -3915
rect -776 -3923 -775 -3915
rect -771 -3923 -770 -3915
rect -768 -3923 -763 -3915
rect -759 -3923 -754 -3915
rect -752 -3923 -751 -3915
rect -747 -3923 -746 -3915
rect -744 -3923 -743 -3915
rect -573 -3923 -572 -3915
rect -570 -3923 -568 -3915
rect -564 -3923 -562 -3915
rect -560 -3923 -559 -3915
rect -547 -3923 -546 -3915
rect -544 -3923 -543 -3915
rect -539 -3923 -538 -3915
rect -536 -3923 -531 -3915
rect -527 -3923 -522 -3915
rect -520 -3923 -519 -3915
rect -515 -3923 -514 -3915
rect -512 -3923 -510 -3915
rect -506 -3923 -504 -3915
rect -502 -3923 -501 -3915
rect -497 -3923 -496 -3915
rect -494 -3923 -489 -3915
rect -485 -3923 -480 -3915
rect -478 -3923 -477 -3915
rect -473 -3923 -472 -3915
rect -470 -3923 -468 -3915
rect -464 -3923 -462 -3915
rect -460 -3923 -459 -3915
rect -455 -3923 -454 -3915
rect -452 -3923 -447 -3915
rect -443 -3923 -438 -3915
rect -436 -3923 -435 -3915
rect -431 -3923 -430 -3915
rect -428 -3923 -426 -3915
rect -422 -3923 -420 -3915
rect -418 -3923 -417 -3915
rect -413 -3923 -412 -3915
rect -410 -3923 -405 -3915
rect -401 -3923 -396 -3915
rect -394 -3923 -393 -3915
rect -389 -3923 -388 -3915
rect -386 -3923 -385 -3915
rect -215 -3923 -214 -3915
rect -212 -3923 -210 -3915
rect -206 -3923 -204 -3915
rect -202 -3923 -201 -3915
rect -189 -3923 -188 -3915
rect -186 -3923 -185 -3915
rect -181 -3923 -180 -3915
rect -178 -3923 -173 -3915
rect -169 -3923 -164 -3915
rect -162 -3923 -161 -3915
rect -157 -3923 -156 -3915
rect -154 -3923 -152 -3915
rect -148 -3923 -146 -3915
rect -144 -3923 -143 -3915
rect -139 -3923 -138 -3915
rect -136 -3923 -131 -3915
rect -127 -3923 -122 -3915
rect -120 -3923 -119 -3915
rect -115 -3923 -114 -3915
rect -112 -3923 -110 -3915
rect -106 -3923 -104 -3915
rect -102 -3923 -101 -3915
rect -97 -3923 -96 -3915
rect -94 -3923 -89 -3915
rect -85 -3923 -80 -3915
rect -78 -3923 -77 -3915
rect -73 -3923 -72 -3915
rect -70 -3923 -68 -3915
rect -64 -3923 -62 -3915
rect -60 -3923 -59 -3915
rect -55 -3923 -54 -3915
rect -52 -3923 -47 -3915
rect -43 -3923 -38 -3915
rect -36 -3923 -35 -3915
rect -31 -3923 -30 -3915
rect -28 -3923 -27 -3915
rect 213 -3923 214 -3915
rect 216 -3923 218 -3915
rect 222 -3923 224 -3915
rect 226 -3923 227 -3915
rect 239 -3923 240 -3915
rect 242 -3923 243 -3915
rect 247 -3923 248 -3915
rect 250 -3923 255 -3915
rect 259 -3923 264 -3915
rect 266 -3923 267 -3915
rect 271 -3923 272 -3915
rect 274 -3923 276 -3915
rect 280 -3923 282 -3915
rect 284 -3923 285 -3915
rect 289 -3923 290 -3915
rect 292 -3923 297 -3915
rect 301 -3923 306 -3915
rect 308 -3923 309 -3915
rect 313 -3923 314 -3915
rect 316 -3923 318 -3915
rect 322 -3923 324 -3915
rect 326 -3923 327 -3915
rect 331 -3923 332 -3915
rect 334 -3923 339 -3915
rect 343 -3923 348 -3915
rect 350 -3923 351 -3915
rect 355 -3923 356 -3915
rect 358 -3923 360 -3915
rect 364 -3923 366 -3915
rect 368 -3923 369 -3915
rect 373 -3923 374 -3915
rect 376 -3923 381 -3915
rect 385 -3923 390 -3915
rect 392 -3923 393 -3915
rect 397 -3923 398 -3915
rect 400 -3923 401 -3915
rect 569 -3923 570 -3915
rect 572 -3923 574 -3915
rect 578 -3923 580 -3915
rect 582 -3923 583 -3915
rect 595 -3923 596 -3915
rect 598 -3923 599 -3915
rect 603 -3923 604 -3915
rect 606 -3923 611 -3915
rect 615 -3923 620 -3915
rect 622 -3923 623 -3915
rect 627 -3923 628 -3915
rect 630 -3923 632 -3915
rect 636 -3923 638 -3915
rect 640 -3923 641 -3915
rect 645 -3923 646 -3915
rect 648 -3923 653 -3915
rect 657 -3923 662 -3915
rect 664 -3923 665 -3915
rect 669 -3923 670 -3915
rect 672 -3923 674 -3915
rect 678 -3923 680 -3915
rect 682 -3923 683 -3915
rect 687 -3923 688 -3915
rect 690 -3923 695 -3915
rect 699 -3923 704 -3915
rect 706 -3923 707 -3915
rect 711 -3923 712 -3915
rect 714 -3923 716 -3915
rect 720 -3923 722 -3915
rect 724 -3923 725 -3915
rect 729 -3923 730 -3915
rect 732 -3923 737 -3915
rect 741 -3923 746 -3915
rect 748 -3923 749 -3915
rect 753 -3923 754 -3915
rect 756 -3923 757 -3915
rect 967 -3923 968 -3915
rect 970 -3923 972 -3915
rect 976 -3923 978 -3915
rect 980 -3923 981 -3915
rect 993 -3923 994 -3915
rect 996 -3923 997 -3915
rect 1001 -3923 1002 -3915
rect 1004 -3923 1009 -3915
rect 1013 -3923 1018 -3915
rect 1020 -3923 1021 -3915
rect 1025 -3923 1026 -3915
rect 1028 -3923 1030 -3915
rect 1034 -3923 1036 -3915
rect 1038 -3923 1039 -3915
rect 1043 -3923 1044 -3915
rect 1046 -3923 1051 -3915
rect 1055 -3923 1060 -3915
rect 1062 -3923 1063 -3915
rect 1067 -3923 1068 -3915
rect 1070 -3923 1072 -3915
rect 1076 -3923 1078 -3915
rect 1080 -3923 1081 -3915
rect 1085 -3923 1086 -3915
rect 1088 -3923 1093 -3915
rect 1097 -3923 1102 -3915
rect 1104 -3923 1105 -3915
rect 1109 -3923 1110 -3915
rect 1112 -3923 1114 -3915
rect 1118 -3923 1120 -3915
rect 1122 -3923 1123 -3915
rect 1127 -3923 1128 -3915
rect 1130 -3923 1135 -3915
rect 1139 -3923 1144 -3915
rect 1146 -3923 1147 -3915
rect 1151 -3923 1152 -3915
rect 1154 -3923 1155 -3915
rect 1325 -3923 1326 -3915
rect 1328 -3923 1330 -3915
rect 1334 -3923 1336 -3915
rect 1338 -3923 1339 -3915
rect 1351 -3923 1352 -3915
rect 1354 -3923 1355 -3915
rect 1359 -3923 1360 -3915
rect 1362 -3923 1367 -3915
rect 1371 -3923 1376 -3915
rect 1378 -3923 1379 -3915
rect 1383 -3923 1384 -3915
rect 1386 -3923 1388 -3915
rect 1392 -3923 1394 -3915
rect 1396 -3923 1397 -3915
rect 1401 -3923 1402 -3915
rect 1404 -3923 1409 -3915
rect 1413 -3923 1418 -3915
rect 1420 -3923 1421 -3915
rect 1425 -3923 1426 -3915
rect 1428 -3923 1430 -3915
rect 1434 -3923 1436 -3915
rect 1438 -3923 1439 -3915
rect 1443 -3923 1444 -3915
rect 1446 -3923 1451 -3915
rect 1455 -3923 1460 -3915
rect 1462 -3923 1463 -3915
rect 1467 -3923 1468 -3915
rect 1470 -3923 1472 -3915
rect 1476 -3923 1478 -3915
rect 1480 -3923 1481 -3915
rect 1485 -3923 1486 -3915
rect 1488 -3923 1493 -3915
rect 1497 -3923 1502 -3915
rect 1504 -3923 1505 -3915
rect 1509 -3923 1510 -3915
rect 1512 -3923 1513 -3915
rect -1260 -4048 -1259 -4040
rect -1257 -4048 -1255 -4040
rect -1251 -4048 -1249 -4040
rect -1247 -4048 -1246 -4040
rect -1234 -4048 -1233 -4040
rect -1231 -4048 -1230 -4040
rect -1226 -4048 -1225 -4040
rect -1223 -4048 -1218 -4040
rect -1214 -4048 -1209 -4040
rect -1207 -4048 -1206 -4040
rect -1202 -4048 -1201 -4040
rect -1199 -4048 -1197 -4040
rect -1193 -4048 -1191 -4040
rect -1189 -4048 -1188 -4040
rect -1184 -4048 -1183 -4040
rect -1181 -4048 -1176 -4040
rect -1172 -4048 -1167 -4040
rect -1165 -4048 -1164 -4040
rect -1160 -4048 -1159 -4040
rect -1157 -4048 -1155 -4040
rect -1151 -4048 -1149 -4040
rect -1147 -4048 -1146 -4040
rect -1142 -4048 -1141 -4040
rect -1139 -4048 -1134 -4040
rect -1130 -4048 -1125 -4040
rect -1123 -4048 -1122 -4040
rect -1118 -4048 -1117 -4040
rect -1115 -4048 -1113 -4040
rect -1109 -4048 -1107 -4040
rect -1105 -4048 -1104 -4040
rect -1100 -4048 -1099 -4040
rect -1097 -4048 -1092 -4040
rect -1088 -4048 -1083 -4040
rect -1081 -4048 -1080 -4040
rect -1076 -4048 -1075 -4040
rect -1073 -4048 -1072 -4040
rect -931 -4048 -930 -4040
rect -928 -4048 -926 -4040
rect -922 -4048 -920 -4040
rect -918 -4048 -917 -4040
rect -905 -4048 -904 -4040
rect -902 -4048 -901 -4040
rect -897 -4048 -896 -4040
rect -894 -4048 -889 -4040
rect -885 -4048 -880 -4040
rect -878 -4048 -877 -4040
rect -873 -4048 -872 -4040
rect -870 -4048 -868 -4040
rect -864 -4048 -862 -4040
rect -860 -4048 -859 -4040
rect -855 -4048 -854 -4040
rect -852 -4048 -847 -4040
rect -843 -4048 -838 -4040
rect -836 -4048 -835 -4040
rect -831 -4048 -830 -4040
rect -828 -4048 -826 -4040
rect -822 -4048 -820 -4040
rect -818 -4048 -817 -4040
rect -813 -4048 -812 -4040
rect -810 -4048 -805 -4040
rect -801 -4048 -796 -4040
rect -794 -4048 -793 -4040
rect -789 -4048 -788 -4040
rect -786 -4048 -784 -4040
rect -780 -4048 -778 -4040
rect -776 -4048 -775 -4040
rect -771 -4048 -770 -4040
rect -768 -4048 -763 -4040
rect -759 -4048 -754 -4040
rect -752 -4048 -751 -4040
rect -747 -4048 -746 -4040
rect -744 -4048 -743 -4040
rect -573 -4048 -572 -4040
rect -570 -4048 -568 -4040
rect -564 -4048 -562 -4040
rect -560 -4048 -559 -4040
rect -547 -4048 -546 -4040
rect -544 -4048 -543 -4040
rect -539 -4048 -538 -4040
rect -536 -4048 -531 -4040
rect -527 -4048 -522 -4040
rect -520 -4048 -519 -4040
rect -515 -4048 -514 -4040
rect -512 -4048 -510 -4040
rect -506 -4048 -504 -4040
rect -502 -4048 -501 -4040
rect -497 -4048 -496 -4040
rect -494 -4048 -489 -4040
rect -485 -4048 -480 -4040
rect -478 -4048 -477 -4040
rect -473 -4048 -472 -4040
rect -470 -4048 -468 -4040
rect -464 -4048 -462 -4040
rect -460 -4048 -459 -4040
rect -455 -4048 -454 -4040
rect -452 -4048 -447 -4040
rect -443 -4048 -438 -4040
rect -436 -4048 -435 -4040
rect -431 -4048 -430 -4040
rect -428 -4048 -426 -4040
rect -422 -4048 -420 -4040
rect -418 -4048 -417 -4040
rect -413 -4048 -412 -4040
rect -410 -4048 -405 -4040
rect -401 -4048 -396 -4040
rect -394 -4048 -393 -4040
rect -389 -4048 -388 -4040
rect -386 -4048 -385 -4040
rect -215 -4048 -214 -4040
rect -212 -4048 -210 -4040
rect -206 -4048 -204 -4040
rect -202 -4048 -201 -4040
rect -189 -4048 -188 -4040
rect -186 -4048 -185 -4040
rect -181 -4048 -180 -4040
rect -178 -4048 -173 -4040
rect -169 -4048 -164 -4040
rect -162 -4048 -161 -4040
rect -157 -4048 -156 -4040
rect -154 -4048 -152 -4040
rect -148 -4048 -146 -4040
rect -144 -4048 -143 -4040
rect -139 -4048 -138 -4040
rect -136 -4048 -131 -4040
rect -127 -4048 -122 -4040
rect -120 -4048 -119 -4040
rect -115 -4048 -114 -4040
rect -112 -4048 -110 -4040
rect -106 -4048 -104 -4040
rect -102 -4048 -101 -4040
rect -97 -4048 -96 -4040
rect -94 -4048 -89 -4040
rect -85 -4048 -80 -4040
rect -78 -4048 -77 -4040
rect -73 -4048 -72 -4040
rect -70 -4048 -68 -4040
rect -64 -4048 -62 -4040
rect -60 -4048 -59 -4040
rect -55 -4048 -54 -4040
rect -52 -4048 -47 -4040
rect -43 -4048 -38 -4040
rect -36 -4048 -35 -4040
rect -31 -4048 -30 -4040
rect -28 -4048 -27 -4040
rect 213 -4048 214 -4040
rect 216 -4048 218 -4040
rect 222 -4048 224 -4040
rect 226 -4048 227 -4040
rect 239 -4048 240 -4040
rect 242 -4048 243 -4040
rect 247 -4048 248 -4040
rect 250 -4048 255 -4040
rect 259 -4048 264 -4040
rect 266 -4048 267 -4040
rect 271 -4048 272 -4040
rect 274 -4048 276 -4040
rect 280 -4048 282 -4040
rect 284 -4048 285 -4040
rect 289 -4048 290 -4040
rect 292 -4048 297 -4040
rect 301 -4048 306 -4040
rect 308 -4048 309 -4040
rect 313 -4048 314 -4040
rect 316 -4048 318 -4040
rect 322 -4048 324 -4040
rect 326 -4048 327 -4040
rect 331 -4048 332 -4040
rect 334 -4048 339 -4040
rect 343 -4048 348 -4040
rect 350 -4048 351 -4040
rect 355 -4048 356 -4040
rect 358 -4048 360 -4040
rect 364 -4048 366 -4040
rect 368 -4048 369 -4040
rect 373 -4048 374 -4040
rect 376 -4048 381 -4040
rect 385 -4048 390 -4040
rect 392 -4048 393 -4040
rect 397 -4048 398 -4040
rect 400 -4048 401 -4040
rect 569 -4048 570 -4040
rect 572 -4048 574 -4040
rect 578 -4048 580 -4040
rect 582 -4048 583 -4040
rect 595 -4048 596 -4040
rect 598 -4048 599 -4040
rect 603 -4048 604 -4040
rect 606 -4048 611 -4040
rect 615 -4048 620 -4040
rect 622 -4048 623 -4040
rect 627 -4048 628 -4040
rect 630 -4048 632 -4040
rect 636 -4048 638 -4040
rect 640 -4048 641 -4040
rect 645 -4048 646 -4040
rect 648 -4048 653 -4040
rect 657 -4048 662 -4040
rect 664 -4048 665 -4040
rect 669 -4048 670 -4040
rect 672 -4048 674 -4040
rect 678 -4048 680 -4040
rect 682 -4048 683 -4040
rect 687 -4048 688 -4040
rect 690 -4048 695 -4040
rect 699 -4048 704 -4040
rect 706 -4048 707 -4040
rect 711 -4048 712 -4040
rect 714 -4048 716 -4040
rect 720 -4048 722 -4040
rect 724 -4048 725 -4040
rect 729 -4048 730 -4040
rect 732 -4048 737 -4040
rect 741 -4048 746 -4040
rect 748 -4048 749 -4040
rect 753 -4048 754 -4040
rect 756 -4048 757 -4040
rect 967 -4048 968 -4040
rect 970 -4048 972 -4040
rect 976 -4048 978 -4040
rect 980 -4048 981 -4040
rect 993 -4048 994 -4040
rect 996 -4048 997 -4040
rect 1001 -4048 1002 -4040
rect 1004 -4048 1009 -4040
rect 1013 -4048 1018 -4040
rect 1020 -4048 1021 -4040
rect 1025 -4048 1026 -4040
rect 1028 -4048 1030 -4040
rect 1034 -4048 1036 -4040
rect 1038 -4048 1039 -4040
rect 1043 -4048 1044 -4040
rect 1046 -4048 1051 -4040
rect 1055 -4048 1060 -4040
rect 1062 -4048 1063 -4040
rect 1067 -4048 1068 -4040
rect 1070 -4048 1072 -4040
rect 1076 -4048 1078 -4040
rect 1080 -4048 1081 -4040
rect 1085 -4048 1086 -4040
rect 1088 -4048 1093 -4040
rect 1097 -4048 1102 -4040
rect 1104 -4048 1105 -4040
rect 1109 -4048 1110 -4040
rect 1112 -4048 1114 -4040
rect 1118 -4048 1120 -4040
rect 1122 -4048 1123 -4040
rect 1127 -4048 1128 -4040
rect 1130 -4048 1135 -4040
rect 1139 -4048 1144 -4040
rect 1146 -4048 1147 -4040
rect 1151 -4048 1152 -4040
rect 1154 -4048 1155 -4040
rect 1325 -4048 1326 -4040
rect 1328 -4048 1330 -4040
rect 1334 -4048 1336 -4040
rect 1338 -4048 1339 -4040
rect 1351 -4048 1352 -4040
rect 1354 -4048 1355 -4040
rect 1359 -4048 1360 -4040
rect 1362 -4048 1367 -4040
rect 1371 -4048 1376 -4040
rect 1378 -4048 1379 -4040
rect 1383 -4048 1384 -4040
rect 1386 -4048 1388 -4040
rect 1392 -4048 1394 -4040
rect 1396 -4048 1397 -4040
rect 1401 -4048 1402 -4040
rect 1404 -4048 1409 -4040
rect 1413 -4048 1418 -4040
rect 1420 -4048 1421 -4040
rect 1425 -4048 1426 -4040
rect 1428 -4048 1430 -4040
rect 1434 -4048 1436 -4040
rect 1438 -4048 1439 -4040
rect 1443 -4048 1444 -4040
rect 1446 -4048 1451 -4040
rect 1455 -4048 1460 -4040
rect 1462 -4048 1463 -4040
rect 1467 -4048 1468 -4040
rect 1470 -4048 1472 -4040
rect 1476 -4048 1478 -4040
rect 1480 -4048 1481 -4040
rect 1485 -4048 1486 -4040
rect 1488 -4048 1493 -4040
rect 1497 -4048 1502 -4040
rect 1504 -4048 1505 -4040
rect 1509 -4048 1510 -4040
rect 1512 -4048 1513 -4040
rect -1260 -4172 -1259 -4164
rect -1257 -4172 -1255 -4164
rect -1251 -4172 -1249 -4164
rect -1247 -4172 -1246 -4164
rect -1234 -4172 -1233 -4164
rect -1231 -4172 -1230 -4164
rect -1226 -4172 -1225 -4164
rect -1223 -4172 -1218 -4164
rect -1214 -4172 -1209 -4164
rect -1207 -4172 -1206 -4164
rect -1202 -4172 -1201 -4164
rect -1199 -4172 -1197 -4164
rect -1193 -4172 -1191 -4164
rect -1189 -4172 -1188 -4164
rect -1184 -4172 -1183 -4164
rect -1181 -4172 -1176 -4164
rect -1172 -4172 -1167 -4164
rect -1165 -4172 -1164 -4164
rect -1160 -4172 -1159 -4164
rect -1157 -4172 -1155 -4164
rect -1151 -4172 -1149 -4164
rect -1147 -4172 -1146 -4164
rect -1142 -4172 -1141 -4164
rect -1139 -4172 -1134 -4164
rect -1130 -4172 -1125 -4164
rect -1123 -4172 -1122 -4164
rect -1118 -4172 -1117 -4164
rect -1115 -4172 -1113 -4164
rect -1109 -4172 -1107 -4164
rect -1105 -4172 -1104 -4164
rect -1100 -4172 -1099 -4164
rect -1097 -4172 -1092 -4164
rect -1088 -4172 -1083 -4164
rect -1081 -4172 -1080 -4164
rect -1076 -4172 -1075 -4164
rect -1073 -4172 -1072 -4164
rect -1025 -4172 -1024 -4164
rect -1022 -4172 -1021 -4164
rect -931 -4172 -930 -4164
rect -928 -4172 -926 -4164
rect -922 -4172 -920 -4164
rect -918 -4172 -917 -4164
rect -905 -4172 -904 -4164
rect -902 -4172 -901 -4164
rect -897 -4172 -896 -4164
rect -894 -4172 -889 -4164
rect -885 -4172 -880 -4164
rect -878 -4172 -877 -4164
rect -873 -4172 -872 -4164
rect -870 -4172 -868 -4164
rect -864 -4172 -862 -4164
rect -860 -4172 -859 -4164
rect -855 -4172 -854 -4164
rect -852 -4172 -847 -4164
rect -843 -4172 -838 -4164
rect -836 -4172 -835 -4164
rect -831 -4172 -830 -4164
rect -828 -4172 -826 -4164
rect -822 -4172 -820 -4164
rect -818 -4172 -817 -4164
rect -813 -4172 -812 -4164
rect -810 -4172 -805 -4164
rect -801 -4172 -796 -4164
rect -794 -4172 -793 -4164
rect -789 -4172 -788 -4164
rect -786 -4172 -784 -4164
rect -780 -4172 -778 -4164
rect -776 -4172 -775 -4164
rect -771 -4172 -770 -4164
rect -768 -4172 -763 -4164
rect -759 -4172 -754 -4164
rect -752 -4172 -751 -4164
rect -747 -4172 -746 -4164
rect -744 -4172 -743 -4164
rect -573 -4172 -572 -4164
rect -570 -4172 -568 -4164
rect -564 -4172 -562 -4164
rect -560 -4172 -559 -4164
rect -547 -4172 -546 -4164
rect -544 -4172 -543 -4164
rect -539 -4172 -538 -4164
rect -536 -4172 -531 -4164
rect -527 -4172 -522 -4164
rect -520 -4172 -519 -4164
rect -515 -4172 -514 -4164
rect -512 -4172 -510 -4164
rect -506 -4172 -504 -4164
rect -502 -4172 -501 -4164
rect -497 -4172 -496 -4164
rect -494 -4172 -489 -4164
rect -485 -4172 -480 -4164
rect -478 -4172 -477 -4164
rect -473 -4172 -472 -4164
rect -470 -4172 -468 -4164
rect -464 -4172 -462 -4164
rect -460 -4172 -459 -4164
rect -455 -4172 -454 -4164
rect -452 -4172 -447 -4164
rect -443 -4172 -438 -4164
rect -436 -4172 -435 -4164
rect -431 -4172 -430 -4164
rect -428 -4172 -426 -4164
rect -422 -4172 -420 -4164
rect -418 -4172 -417 -4164
rect -413 -4172 -412 -4164
rect -410 -4172 -405 -4164
rect -401 -4172 -396 -4164
rect -394 -4172 -393 -4164
rect -389 -4172 -388 -4164
rect -386 -4172 -385 -4164
rect -328 -4172 -327 -4164
rect -325 -4172 -324 -4164
rect -215 -4172 -214 -4164
rect -212 -4172 -210 -4164
rect -206 -4172 -204 -4164
rect -202 -4172 -201 -4164
rect -189 -4172 -188 -4164
rect -186 -4172 -185 -4164
rect -181 -4172 -180 -4164
rect -178 -4172 -173 -4164
rect -169 -4172 -164 -4164
rect -162 -4172 -161 -4164
rect -157 -4172 -156 -4164
rect -154 -4172 -152 -4164
rect -148 -4172 -146 -4164
rect -144 -4172 -143 -4164
rect -139 -4172 -138 -4164
rect -136 -4172 -131 -4164
rect -127 -4172 -122 -4164
rect -120 -4172 -119 -4164
rect -115 -4172 -114 -4164
rect -112 -4172 -110 -4164
rect -106 -4172 -104 -4164
rect -102 -4172 -101 -4164
rect -97 -4172 -96 -4164
rect -94 -4172 -89 -4164
rect -85 -4172 -80 -4164
rect -78 -4172 -77 -4164
rect -73 -4172 -72 -4164
rect -70 -4172 -68 -4164
rect -64 -4172 -62 -4164
rect -60 -4172 -59 -4164
rect -55 -4172 -54 -4164
rect -52 -4172 -47 -4164
rect -43 -4172 -38 -4164
rect -36 -4172 -35 -4164
rect -31 -4172 -30 -4164
rect -28 -4172 -27 -4164
rect 460 -4172 461 -4164
rect 463 -4172 464 -4164
rect 1205 -4172 1206 -4164
rect 1208 -4172 1209 -4164
rect -1335 -4283 -1334 -4275
rect -1332 -4283 -1331 -4275
rect -1327 -4283 -1326 -4275
rect -1324 -4283 -1322 -4275
rect -1318 -4283 -1316 -4275
rect -1314 -4283 -1313 -4275
rect -1025 -4283 -1024 -4275
rect -1022 -4283 -1021 -4275
rect -931 -4283 -930 -4275
rect -928 -4283 -927 -4275
rect -923 -4283 -922 -4275
rect -920 -4283 -918 -4275
rect -914 -4283 -912 -4275
rect -910 -4283 -909 -4275
rect -669 -4291 -668 -4275
rect -666 -4291 -665 -4275
rect -573 -4283 -572 -4275
rect -570 -4283 -569 -4275
rect -565 -4283 -564 -4275
rect -562 -4283 -560 -4275
rect -556 -4283 -554 -4275
rect -552 -4283 -551 -4275
rect -328 -4283 -327 -4275
rect -325 -4283 -324 -4275
rect -215 -4283 -214 -4275
rect -212 -4283 -211 -4275
rect -207 -4283 -206 -4275
rect -204 -4283 -202 -4275
rect -198 -4283 -196 -4275
rect -194 -4283 -193 -4275
rect 213 -4283 214 -4275
rect 216 -4283 217 -4275
rect 221 -4283 222 -4275
rect 224 -4283 226 -4275
rect 230 -4283 232 -4275
rect 234 -4283 235 -4275
rect 460 -4283 461 -4275
rect 463 -4283 464 -4275
rect 569 -4283 570 -4275
rect 572 -4283 573 -4275
rect 577 -4283 578 -4275
rect 580 -4283 582 -4275
rect 586 -4283 588 -4275
rect 590 -4283 591 -4275
rect 864 -4291 865 -4275
rect 867 -4291 868 -4275
rect 967 -4283 968 -4275
rect 970 -4283 971 -4275
rect 975 -4283 976 -4275
rect 978 -4283 980 -4275
rect 984 -4283 986 -4275
rect 988 -4283 989 -4275
rect 1205 -4283 1206 -4275
rect 1208 -4283 1209 -4275
rect 1325 -4283 1326 -4275
rect 1328 -4283 1329 -4275
rect 1333 -4283 1334 -4275
rect 1336 -4283 1338 -4275
rect 1342 -4283 1344 -4275
rect 1346 -4283 1347 -4275
rect -1260 -4402 -1259 -4394
rect -1257 -4402 -1255 -4394
rect -1251 -4402 -1249 -4394
rect -1247 -4402 -1246 -4394
rect -1234 -4402 -1233 -4394
rect -1231 -4402 -1223 -4394
rect -1221 -4402 -1220 -4394
rect -1216 -4402 -1215 -4394
rect -1213 -4402 -1205 -4394
rect -1203 -4402 -1198 -4394
rect -1194 -4402 -1189 -4394
rect -1187 -4402 -1186 -4394
rect -1182 -4402 -1181 -4394
rect -1179 -4402 -1177 -4394
rect -1173 -4402 -1171 -4394
rect -1169 -4402 -1168 -4394
rect -931 -4402 -930 -4394
rect -928 -4402 -926 -4394
rect -922 -4402 -920 -4394
rect -918 -4402 -917 -4394
rect -905 -4402 -904 -4394
rect -902 -4402 -900 -4394
rect -896 -4402 -894 -4394
rect -892 -4402 -891 -4394
rect -879 -4402 -878 -4394
rect -876 -4402 -868 -4394
rect -866 -4402 -865 -4394
rect -861 -4402 -860 -4394
rect -858 -4402 -850 -4394
rect -848 -4402 -843 -4394
rect -839 -4402 -834 -4394
rect -832 -4402 -831 -4394
rect -827 -4402 -826 -4394
rect -824 -4402 -822 -4394
rect -818 -4402 -816 -4394
rect -814 -4402 -813 -4394
rect -801 -4402 -800 -4394
rect -798 -4402 -790 -4394
rect -788 -4402 -787 -4394
rect -783 -4402 -782 -4394
rect -780 -4402 -772 -4394
rect -770 -4402 -765 -4394
rect -761 -4402 -756 -4394
rect -754 -4402 -753 -4394
rect -749 -4402 -748 -4394
rect -746 -4402 -741 -4394
rect -737 -4402 -732 -4394
rect -730 -4402 -729 -4394
rect -717 -4402 -716 -4394
rect -714 -4402 -708 -4394
rect -706 -4402 -704 -4394
rect -700 -4402 -698 -4394
rect -696 -4402 -695 -4394
rect -573 -4402 -572 -4394
rect -570 -4402 -568 -4394
rect -564 -4402 -562 -4394
rect -560 -4402 -559 -4394
rect -547 -4402 -546 -4394
rect -544 -4402 -542 -4394
rect -538 -4402 -536 -4394
rect -534 -4402 -533 -4394
rect -521 -4402 -520 -4394
rect -518 -4402 -510 -4394
rect -508 -4402 -507 -4394
rect -503 -4402 -502 -4394
rect -500 -4402 -492 -4394
rect -490 -4402 -485 -4394
rect -481 -4402 -476 -4394
rect -474 -4402 -473 -4394
rect -469 -4402 -468 -4394
rect -466 -4402 -464 -4394
rect -460 -4402 -458 -4394
rect -456 -4402 -455 -4394
rect -443 -4402 -442 -4394
rect -440 -4402 -432 -4394
rect -430 -4402 -429 -4394
rect -425 -4402 -424 -4394
rect -422 -4402 -414 -4394
rect -412 -4402 -407 -4394
rect -403 -4402 -398 -4394
rect -396 -4402 -395 -4394
rect -391 -4402 -390 -4394
rect -388 -4402 -383 -4394
rect -379 -4402 -374 -4394
rect -372 -4402 -371 -4394
rect -359 -4402 -358 -4394
rect -356 -4402 -350 -4394
rect -348 -4402 -346 -4394
rect -342 -4402 -340 -4394
rect -338 -4402 -337 -4394
rect -215 -4402 -214 -4394
rect -212 -4402 -210 -4394
rect -206 -4402 -204 -4394
rect -202 -4402 -201 -4394
rect -189 -4402 -188 -4394
rect -186 -4402 -184 -4394
rect -180 -4402 -178 -4394
rect -176 -4402 -175 -4394
rect -163 -4402 -162 -4394
rect -160 -4402 -152 -4394
rect -150 -4402 -149 -4394
rect -145 -4402 -144 -4394
rect -142 -4402 -134 -4394
rect -132 -4402 -127 -4394
rect -123 -4402 -118 -4394
rect -116 -4402 -115 -4394
rect -111 -4402 -110 -4394
rect -108 -4402 -106 -4394
rect -102 -4402 -100 -4394
rect -98 -4402 -97 -4394
rect -85 -4402 -84 -4394
rect -82 -4402 -74 -4394
rect -72 -4402 -71 -4394
rect -67 -4402 -66 -4394
rect -64 -4402 -56 -4394
rect -54 -4402 -49 -4394
rect -45 -4402 -40 -4394
rect -38 -4402 -37 -4394
rect -33 -4402 -32 -4394
rect -30 -4402 -25 -4394
rect -21 -4402 -16 -4394
rect -14 -4402 -13 -4394
rect -1 -4402 0 -4394
rect 2 -4402 8 -4394
rect 10 -4402 12 -4394
rect 16 -4402 18 -4394
rect 20 -4402 21 -4394
rect 213 -4402 214 -4394
rect 216 -4402 218 -4394
rect 222 -4402 224 -4394
rect 226 -4402 227 -4394
rect 239 -4402 240 -4394
rect 242 -4402 244 -4394
rect 248 -4402 250 -4394
rect 252 -4402 253 -4394
rect 265 -4402 266 -4394
rect 268 -4402 276 -4394
rect 278 -4402 279 -4394
rect 283 -4402 284 -4394
rect 286 -4402 294 -4394
rect 296 -4402 301 -4394
rect 305 -4402 310 -4394
rect 312 -4402 313 -4394
rect 317 -4402 318 -4394
rect 320 -4402 322 -4394
rect 326 -4402 328 -4394
rect 330 -4402 331 -4394
rect 343 -4402 344 -4394
rect 346 -4402 354 -4394
rect 356 -4402 357 -4394
rect 361 -4402 362 -4394
rect 364 -4402 372 -4394
rect 374 -4402 379 -4394
rect 383 -4402 388 -4394
rect 390 -4402 391 -4394
rect 395 -4402 396 -4394
rect 398 -4402 403 -4394
rect 407 -4402 412 -4394
rect 414 -4402 415 -4394
rect 427 -4402 428 -4394
rect 430 -4402 436 -4394
rect 438 -4402 440 -4394
rect 444 -4402 446 -4394
rect 448 -4402 449 -4394
rect 569 -4402 570 -4394
rect 572 -4402 574 -4394
rect 578 -4402 580 -4394
rect 582 -4402 583 -4394
rect 595 -4402 596 -4394
rect 598 -4402 600 -4394
rect 604 -4402 606 -4394
rect 608 -4402 609 -4394
rect 621 -4402 622 -4394
rect 624 -4402 632 -4394
rect 634 -4402 635 -4394
rect 639 -4402 640 -4394
rect 642 -4402 650 -4394
rect 652 -4402 657 -4394
rect 661 -4402 666 -4394
rect 668 -4402 669 -4394
rect 673 -4402 674 -4394
rect 676 -4402 678 -4394
rect 682 -4402 684 -4394
rect 686 -4402 687 -4394
rect 699 -4402 700 -4394
rect 702 -4402 710 -4394
rect 712 -4402 713 -4394
rect 717 -4402 718 -4394
rect 720 -4402 728 -4394
rect 730 -4402 735 -4394
rect 739 -4402 744 -4394
rect 746 -4402 747 -4394
rect 751 -4402 752 -4394
rect 754 -4402 759 -4394
rect 763 -4402 768 -4394
rect 770 -4402 771 -4394
rect 783 -4402 784 -4394
rect 786 -4402 792 -4394
rect 794 -4402 796 -4394
rect 800 -4402 802 -4394
rect 804 -4402 805 -4394
rect 967 -4402 968 -4394
rect 970 -4402 972 -4394
rect 976 -4402 978 -4394
rect 980 -4402 981 -4394
rect 993 -4402 994 -4394
rect 996 -4402 998 -4394
rect 1002 -4402 1004 -4394
rect 1006 -4402 1007 -4394
rect 1019 -4402 1020 -4394
rect 1022 -4402 1030 -4394
rect 1032 -4402 1033 -4394
rect 1037 -4402 1038 -4394
rect 1040 -4402 1048 -4394
rect 1050 -4402 1055 -4394
rect 1059 -4402 1064 -4394
rect 1066 -4402 1067 -4394
rect 1071 -4402 1072 -4394
rect 1074 -4402 1076 -4394
rect 1080 -4402 1082 -4394
rect 1084 -4402 1085 -4394
rect 1097 -4402 1098 -4394
rect 1100 -4402 1108 -4394
rect 1110 -4402 1111 -4394
rect 1115 -4402 1116 -4394
rect 1118 -4402 1126 -4394
rect 1128 -4402 1133 -4394
rect 1137 -4402 1142 -4394
rect 1144 -4402 1145 -4394
rect 1149 -4402 1150 -4394
rect 1152 -4402 1157 -4394
rect 1161 -4402 1166 -4394
rect 1168 -4402 1169 -4394
rect 1181 -4402 1182 -4394
rect 1184 -4402 1190 -4394
rect 1192 -4402 1194 -4394
rect 1198 -4402 1200 -4394
rect 1202 -4402 1203 -4394
rect 1325 -4402 1326 -4394
rect 1328 -4402 1330 -4394
rect 1334 -4402 1336 -4394
rect 1338 -4402 1339 -4394
rect 1351 -4402 1352 -4394
rect 1354 -4402 1356 -4394
rect 1360 -4402 1362 -4394
rect 1364 -4402 1365 -4394
rect 1377 -4402 1378 -4394
rect 1380 -4402 1388 -4394
rect 1390 -4402 1391 -4394
rect 1395 -4402 1396 -4394
rect 1398 -4402 1406 -4394
rect 1408 -4402 1413 -4394
rect 1417 -4402 1422 -4394
rect 1424 -4402 1425 -4394
rect 1429 -4402 1430 -4394
rect 1432 -4402 1434 -4394
rect 1438 -4402 1440 -4394
rect 1442 -4402 1443 -4394
rect 1455 -4402 1456 -4394
rect 1458 -4402 1466 -4394
rect 1468 -4402 1469 -4394
rect 1473 -4402 1474 -4394
rect 1476 -4402 1484 -4394
rect 1486 -4402 1491 -4394
rect 1495 -4402 1500 -4394
rect 1502 -4402 1503 -4394
rect 1507 -4402 1508 -4394
rect 1510 -4402 1515 -4394
rect 1519 -4402 1524 -4394
rect 1526 -4402 1527 -4394
rect 1539 -4402 1540 -4394
rect 1542 -4402 1548 -4394
rect 1550 -4402 1552 -4394
rect 1556 -4402 1558 -4394
rect 1560 -4402 1561 -4394
rect -1260 -4525 -1259 -4517
rect -1257 -4525 -1255 -4517
rect -1251 -4525 -1249 -4517
rect -1247 -4525 -1246 -4517
rect -1234 -4525 -1233 -4517
rect -1231 -4525 -1230 -4517
rect -1226 -4525 -1225 -4517
rect -1223 -4525 -1218 -4517
rect -1214 -4525 -1209 -4517
rect -1207 -4525 -1206 -4517
rect -1202 -4525 -1201 -4517
rect -1199 -4525 -1197 -4517
rect -1193 -4525 -1191 -4517
rect -1189 -4525 -1188 -4517
rect -1184 -4525 -1183 -4517
rect -1181 -4525 -1176 -4517
rect -1172 -4525 -1167 -4517
rect -1165 -4525 -1164 -4517
rect -1160 -4525 -1159 -4517
rect -1157 -4525 -1155 -4517
rect -1151 -4525 -1149 -4517
rect -1147 -4525 -1146 -4517
rect -1142 -4525 -1141 -4517
rect -1139 -4525 -1134 -4517
rect -1130 -4525 -1125 -4517
rect -1123 -4525 -1122 -4517
rect -1118 -4525 -1117 -4517
rect -1115 -4525 -1113 -4517
rect -1109 -4525 -1107 -4517
rect -1105 -4525 -1104 -4517
rect -1100 -4525 -1099 -4517
rect -1097 -4525 -1092 -4517
rect -1088 -4525 -1083 -4517
rect -1081 -4525 -1080 -4517
rect -1076 -4525 -1075 -4517
rect -1073 -4525 -1072 -4517
rect -931 -4525 -930 -4517
rect -928 -4525 -926 -4517
rect -922 -4525 -920 -4517
rect -918 -4525 -917 -4517
rect -905 -4525 -904 -4517
rect -902 -4525 -901 -4517
rect -897 -4525 -896 -4517
rect -894 -4525 -889 -4517
rect -885 -4525 -880 -4517
rect -878 -4525 -877 -4517
rect -873 -4525 -872 -4517
rect -870 -4525 -868 -4517
rect -864 -4525 -862 -4517
rect -860 -4525 -859 -4517
rect -855 -4525 -854 -4517
rect -852 -4525 -847 -4517
rect -843 -4525 -838 -4517
rect -836 -4525 -835 -4517
rect -831 -4525 -830 -4517
rect -828 -4525 -826 -4517
rect -822 -4525 -820 -4517
rect -818 -4525 -817 -4517
rect -813 -4525 -812 -4517
rect -810 -4525 -805 -4517
rect -801 -4525 -796 -4517
rect -794 -4525 -793 -4517
rect -789 -4525 -788 -4517
rect -786 -4525 -784 -4517
rect -780 -4525 -778 -4517
rect -776 -4525 -775 -4517
rect -771 -4525 -770 -4517
rect -768 -4525 -763 -4517
rect -759 -4525 -754 -4517
rect -752 -4525 -751 -4517
rect -747 -4525 -746 -4517
rect -744 -4525 -743 -4517
rect -573 -4525 -572 -4517
rect -570 -4525 -568 -4517
rect -564 -4525 -562 -4517
rect -560 -4525 -559 -4517
rect -547 -4525 -546 -4517
rect -544 -4525 -543 -4517
rect -539 -4525 -538 -4517
rect -536 -4525 -531 -4517
rect -527 -4525 -522 -4517
rect -520 -4525 -519 -4517
rect -515 -4525 -514 -4517
rect -512 -4525 -510 -4517
rect -506 -4525 -504 -4517
rect -502 -4525 -501 -4517
rect -497 -4525 -496 -4517
rect -494 -4525 -489 -4517
rect -485 -4525 -480 -4517
rect -478 -4525 -477 -4517
rect -473 -4525 -472 -4517
rect -470 -4525 -468 -4517
rect -464 -4525 -462 -4517
rect -460 -4525 -459 -4517
rect -455 -4525 -454 -4517
rect -452 -4525 -447 -4517
rect -443 -4525 -438 -4517
rect -436 -4525 -435 -4517
rect -431 -4525 -430 -4517
rect -428 -4525 -426 -4517
rect -422 -4525 -420 -4517
rect -418 -4525 -417 -4517
rect -413 -4525 -412 -4517
rect -410 -4525 -405 -4517
rect -401 -4525 -396 -4517
rect -394 -4525 -393 -4517
rect -389 -4525 -388 -4517
rect -386 -4525 -385 -4517
rect -1260 -4646 -1259 -4638
rect -1257 -4646 -1255 -4638
rect -1251 -4646 -1249 -4638
rect -1247 -4646 -1246 -4638
rect -1234 -4646 -1233 -4638
rect -1231 -4646 -1230 -4638
rect -1226 -4646 -1225 -4638
rect -1223 -4646 -1218 -4638
rect -1214 -4646 -1209 -4638
rect -1207 -4646 -1206 -4638
rect -1202 -4646 -1201 -4638
rect -1199 -4646 -1197 -4638
rect -1193 -4646 -1191 -4638
rect -1189 -4646 -1188 -4638
rect -1184 -4646 -1183 -4638
rect -1181 -4646 -1176 -4638
rect -1172 -4646 -1167 -4638
rect -1165 -4646 -1164 -4638
rect -1160 -4646 -1159 -4638
rect -1157 -4646 -1155 -4638
rect -1151 -4646 -1149 -4638
rect -1147 -4646 -1146 -4638
rect -1142 -4646 -1141 -4638
rect -1139 -4646 -1134 -4638
rect -1130 -4646 -1125 -4638
rect -1123 -4646 -1122 -4638
rect -1118 -4646 -1117 -4638
rect -1115 -4646 -1113 -4638
rect -1109 -4646 -1107 -4638
rect -1105 -4646 -1104 -4638
rect -1100 -4646 -1099 -4638
rect -1097 -4646 -1092 -4638
rect -1088 -4646 -1083 -4638
rect -1081 -4646 -1080 -4638
rect -1076 -4646 -1075 -4638
rect -1073 -4646 -1072 -4638
rect -931 -4646 -930 -4638
rect -928 -4646 -926 -4638
rect -922 -4646 -920 -4638
rect -918 -4646 -917 -4638
rect -905 -4646 -904 -4638
rect -902 -4646 -901 -4638
rect -897 -4646 -896 -4638
rect -894 -4646 -889 -4638
rect -885 -4646 -880 -4638
rect -878 -4646 -877 -4638
rect -873 -4646 -872 -4638
rect -870 -4646 -868 -4638
rect -864 -4646 -862 -4638
rect -860 -4646 -859 -4638
rect -855 -4646 -854 -4638
rect -852 -4646 -847 -4638
rect -843 -4646 -838 -4638
rect -836 -4646 -835 -4638
rect -831 -4646 -830 -4638
rect -828 -4646 -826 -4638
rect -822 -4646 -820 -4638
rect -818 -4646 -817 -4638
rect -813 -4646 -812 -4638
rect -810 -4646 -805 -4638
rect -801 -4646 -796 -4638
rect -794 -4646 -793 -4638
rect -789 -4646 -788 -4638
rect -786 -4646 -784 -4638
rect -780 -4646 -778 -4638
rect -776 -4646 -775 -4638
rect -771 -4646 -770 -4638
rect -768 -4646 -763 -4638
rect -759 -4646 -754 -4638
rect -752 -4646 -751 -4638
rect -747 -4646 -746 -4638
rect -744 -4646 -743 -4638
rect -573 -4646 -572 -4638
rect -570 -4646 -568 -4638
rect -564 -4646 -562 -4638
rect -560 -4646 -559 -4638
rect -547 -4646 -546 -4638
rect -544 -4646 -543 -4638
rect -539 -4646 -538 -4638
rect -536 -4646 -531 -4638
rect -527 -4646 -522 -4638
rect -520 -4646 -519 -4638
rect -515 -4646 -514 -4638
rect -512 -4646 -510 -4638
rect -506 -4646 -504 -4638
rect -502 -4646 -501 -4638
rect -497 -4646 -496 -4638
rect -494 -4646 -489 -4638
rect -485 -4646 -480 -4638
rect -478 -4646 -477 -4638
rect -473 -4646 -472 -4638
rect -470 -4646 -468 -4638
rect -464 -4646 -462 -4638
rect -460 -4646 -459 -4638
rect -455 -4646 -454 -4638
rect -452 -4646 -447 -4638
rect -443 -4646 -438 -4638
rect -436 -4646 -435 -4638
rect -431 -4646 -430 -4638
rect -428 -4646 -426 -4638
rect -422 -4646 -420 -4638
rect -418 -4646 -417 -4638
rect -413 -4646 -412 -4638
rect -410 -4646 -405 -4638
rect -401 -4646 -396 -4638
rect -394 -4646 -393 -4638
rect -389 -4646 -388 -4638
rect -386 -4646 -385 -4638
rect -215 -4646 -214 -4638
rect -212 -4646 -210 -4638
rect -206 -4646 -204 -4638
rect -202 -4646 -201 -4638
rect -189 -4646 -188 -4638
rect -186 -4646 -185 -4638
rect -181 -4646 -180 -4638
rect -178 -4646 -173 -4638
rect -169 -4646 -164 -4638
rect -162 -4646 -161 -4638
rect -157 -4646 -156 -4638
rect -154 -4646 -152 -4638
rect -148 -4646 -146 -4638
rect -144 -4646 -143 -4638
rect -139 -4646 -138 -4638
rect -136 -4646 -131 -4638
rect -127 -4646 -122 -4638
rect -120 -4646 -119 -4638
rect -115 -4646 -114 -4638
rect -112 -4646 -110 -4638
rect -106 -4646 -104 -4638
rect -102 -4646 -101 -4638
rect -97 -4646 -96 -4638
rect -94 -4646 -89 -4638
rect -85 -4646 -80 -4638
rect -78 -4646 -77 -4638
rect -73 -4646 -72 -4638
rect -70 -4646 -68 -4638
rect -64 -4646 -62 -4638
rect -60 -4646 -59 -4638
rect -55 -4646 -54 -4638
rect -52 -4646 -47 -4638
rect -43 -4646 -38 -4638
rect -36 -4646 -35 -4638
rect -31 -4646 -30 -4638
rect -28 -4646 -27 -4638
rect 213 -4646 214 -4638
rect 216 -4646 218 -4638
rect 222 -4646 224 -4638
rect 226 -4646 227 -4638
rect 239 -4646 240 -4638
rect 242 -4646 243 -4638
rect 247 -4646 248 -4638
rect 250 -4646 255 -4638
rect 259 -4646 264 -4638
rect 266 -4646 267 -4638
rect 271 -4646 272 -4638
rect 274 -4646 276 -4638
rect 280 -4646 282 -4638
rect 284 -4646 285 -4638
rect 289 -4646 290 -4638
rect 292 -4646 297 -4638
rect 301 -4646 306 -4638
rect 308 -4646 309 -4638
rect 313 -4646 314 -4638
rect 316 -4646 318 -4638
rect 322 -4646 324 -4638
rect 326 -4646 327 -4638
rect 331 -4646 332 -4638
rect 334 -4646 339 -4638
rect 343 -4646 348 -4638
rect 350 -4646 351 -4638
rect 355 -4646 356 -4638
rect 358 -4646 360 -4638
rect 364 -4646 366 -4638
rect 368 -4646 369 -4638
rect 373 -4646 374 -4638
rect 376 -4646 381 -4638
rect 385 -4646 390 -4638
rect 392 -4646 393 -4638
rect 397 -4646 398 -4638
rect 400 -4646 401 -4638
rect 569 -4646 570 -4638
rect 572 -4646 574 -4638
rect 578 -4646 580 -4638
rect 582 -4646 583 -4638
rect 595 -4646 596 -4638
rect 598 -4646 599 -4638
rect 603 -4646 604 -4638
rect 606 -4646 611 -4638
rect 615 -4646 620 -4638
rect 622 -4646 623 -4638
rect 627 -4646 628 -4638
rect 630 -4646 632 -4638
rect 636 -4646 638 -4638
rect 640 -4646 641 -4638
rect 645 -4646 646 -4638
rect 648 -4646 653 -4638
rect 657 -4646 662 -4638
rect 664 -4646 665 -4638
rect 669 -4646 670 -4638
rect 672 -4646 674 -4638
rect 678 -4646 680 -4638
rect 682 -4646 683 -4638
rect 687 -4646 688 -4638
rect 690 -4646 695 -4638
rect 699 -4646 704 -4638
rect 706 -4646 707 -4638
rect 711 -4646 712 -4638
rect 714 -4646 716 -4638
rect 720 -4646 722 -4638
rect 724 -4646 725 -4638
rect 729 -4646 730 -4638
rect 732 -4646 737 -4638
rect 741 -4646 746 -4638
rect 748 -4646 749 -4638
rect 753 -4646 754 -4638
rect 756 -4646 757 -4638
rect 967 -4646 968 -4638
rect 970 -4646 972 -4638
rect 976 -4646 978 -4638
rect 980 -4646 981 -4638
rect 993 -4646 994 -4638
rect 996 -4646 997 -4638
rect 1001 -4646 1002 -4638
rect 1004 -4646 1009 -4638
rect 1013 -4646 1018 -4638
rect 1020 -4646 1021 -4638
rect 1025 -4646 1026 -4638
rect 1028 -4646 1030 -4638
rect 1034 -4646 1036 -4638
rect 1038 -4646 1039 -4638
rect 1043 -4646 1044 -4638
rect 1046 -4646 1051 -4638
rect 1055 -4646 1060 -4638
rect 1062 -4646 1063 -4638
rect 1067 -4646 1068 -4638
rect 1070 -4646 1072 -4638
rect 1076 -4646 1078 -4638
rect 1080 -4646 1081 -4638
rect 1085 -4646 1086 -4638
rect 1088 -4646 1093 -4638
rect 1097 -4646 1102 -4638
rect 1104 -4646 1105 -4638
rect 1109 -4646 1110 -4638
rect 1112 -4646 1114 -4638
rect 1118 -4646 1120 -4638
rect 1122 -4646 1123 -4638
rect 1127 -4646 1128 -4638
rect 1130 -4646 1135 -4638
rect 1139 -4646 1144 -4638
rect 1146 -4646 1147 -4638
rect 1151 -4646 1152 -4638
rect 1154 -4646 1155 -4638
rect 1325 -4646 1326 -4638
rect 1328 -4646 1330 -4638
rect 1334 -4646 1336 -4638
rect 1338 -4646 1339 -4638
rect 1351 -4646 1352 -4638
rect 1354 -4646 1355 -4638
rect 1359 -4646 1360 -4638
rect 1362 -4646 1367 -4638
rect 1371 -4646 1376 -4638
rect 1378 -4646 1379 -4638
rect 1383 -4646 1384 -4638
rect 1386 -4646 1388 -4638
rect 1392 -4646 1394 -4638
rect 1396 -4646 1397 -4638
rect 1401 -4646 1402 -4638
rect 1404 -4646 1409 -4638
rect 1413 -4646 1418 -4638
rect 1420 -4646 1421 -4638
rect 1425 -4646 1426 -4638
rect 1428 -4646 1430 -4638
rect 1434 -4646 1436 -4638
rect 1438 -4646 1439 -4638
rect 1443 -4646 1444 -4638
rect 1446 -4646 1451 -4638
rect 1455 -4646 1460 -4638
rect 1462 -4646 1463 -4638
rect 1467 -4646 1468 -4638
rect 1470 -4646 1472 -4638
rect 1476 -4646 1478 -4638
rect 1480 -4646 1481 -4638
rect 1485 -4646 1486 -4638
rect 1488 -4646 1493 -4638
rect 1497 -4646 1502 -4638
rect 1504 -4646 1505 -4638
rect 1509 -4646 1510 -4638
rect 1512 -4646 1513 -4638
rect -1260 -4767 -1259 -4759
rect -1257 -4767 -1255 -4759
rect -1251 -4767 -1249 -4759
rect -1247 -4767 -1246 -4759
rect -1234 -4767 -1233 -4759
rect -1231 -4767 -1230 -4759
rect -1226 -4767 -1225 -4759
rect -1223 -4767 -1218 -4759
rect -1214 -4767 -1209 -4759
rect -1207 -4767 -1206 -4759
rect -1202 -4767 -1201 -4759
rect -1199 -4767 -1197 -4759
rect -1193 -4767 -1191 -4759
rect -1189 -4767 -1188 -4759
rect -1184 -4767 -1183 -4759
rect -1181 -4767 -1176 -4759
rect -1172 -4767 -1167 -4759
rect -1165 -4767 -1164 -4759
rect -1160 -4767 -1159 -4759
rect -1157 -4767 -1155 -4759
rect -1151 -4767 -1149 -4759
rect -1147 -4767 -1146 -4759
rect -1142 -4767 -1141 -4759
rect -1139 -4767 -1134 -4759
rect -1130 -4767 -1125 -4759
rect -1123 -4767 -1122 -4759
rect -1118 -4767 -1117 -4759
rect -1115 -4767 -1113 -4759
rect -1109 -4767 -1107 -4759
rect -1105 -4767 -1104 -4759
rect -1100 -4767 -1099 -4759
rect -1097 -4767 -1092 -4759
rect -1088 -4767 -1083 -4759
rect -1081 -4767 -1080 -4759
rect -1076 -4767 -1075 -4759
rect -1073 -4767 -1072 -4759
rect -931 -4767 -930 -4759
rect -928 -4767 -926 -4759
rect -922 -4767 -920 -4759
rect -918 -4767 -917 -4759
rect -905 -4767 -904 -4759
rect -902 -4767 -901 -4759
rect -897 -4767 -896 -4759
rect -894 -4767 -889 -4759
rect -885 -4767 -880 -4759
rect -878 -4767 -877 -4759
rect -873 -4767 -872 -4759
rect -870 -4767 -868 -4759
rect -864 -4767 -862 -4759
rect -860 -4767 -859 -4759
rect -855 -4767 -854 -4759
rect -852 -4767 -847 -4759
rect -843 -4767 -838 -4759
rect -836 -4767 -835 -4759
rect -831 -4767 -830 -4759
rect -828 -4767 -826 -4759
rect -822 -4767 -820 -4759
rect -818 -4767 -817 -4759
rect -813 -4767 -812 -4759
rect -810 -4767 -805 -4759
rect -801 -4767 -796 -4759
rect -794 -4767 -793 -4759
rect -789 -4767 -788 -4759
rect -786 -4767 -784 -4759
rect -780 -4767 -778 -4759
rect -776 -4767 -775 -4759
rect -771 -4767 -770 -4759
rect -768 -4767 -763 -4759
rect -759 -4767 -754 -4759
rect -752 -4767 -751 -4759
rect -747 -4767 -746 -4759
rect -744 -4767 -743 -4759
rect -573 -4767 -572 -4759
rect -570 -4767 -568 -4759
rect -564 -4767 -562 -4759
rect -560 -4767 -559 -4759
rect -547 -4767 -546 -4759
rect -544 -4767 -543 -4759
rect -539 -4767 -538 -4759
rect -536 -4767 -531 -4759
rect -527 -4767 -522 -4759
rect -520 -4767 -519 -4759
rect -515 -4767 -514 -4759
rect -512 -4767 -510 -4759
rect -506 -4767 -504 -4759
rect -502 -4767 -501 -4759
rect -497 -4767 -496 -4759
rect -494 -4767 -489 -4759
rect -485 -4767 -480 -4759
rect -478 -4767 -477 -4759
rect -473 -4767 -472 -4759
rect -470 -4767 -468 -4759
rect -464 -4767 -462 -4759
rect -460 -4767 -459 -4759
rect -455 -4767 -454 -4759
rect -452 -4767 -447 -4759
rect -443 -4767 -438 -4759
rect -436 -4767 -435 -4759
rect -431 -4767 -430 -4759
rect -428 -4767 -426 -4759
rect -422 -4767 -420 -4759
rect -418 -4767 -417 -4759
rect -413 -4767 -412 -4759
rect -410 -4767 -405 -4759
rect -401 -4767 -396 -4759
rect -394 -4767 -393 -4759
rect -389 -4767 -388 -4759
rect -386 -4767 -385 -4759
rect -215 -4767 -214 -4759
rect -212 -4767 -210 -4759
rect -206 -4767 -204 -4759
rect -202 -4767 -201 -4759
rect -189 -4767 -188 -4759
rect -186 -4767 -185 -4759
rect -181 -4767 -180 -4759
rect -178 -4767 -173 -4759
rect -169 -4767 -164 -4759
rect -162 -4767 -161 -4759
rect -157 -4767 -156 -4759
rect -154 -4767 -152 -4759
rect -148 -4767 -146 -4759
rect -144 -4767 -143 -4759
rect -139 -4767 -138 -4759
rect -136 -4767 -131 -4759
rect -127 -4767 -122 -4759
rect -120 -4767 -119 -4759
rect -115 -4767 -114 -4759
rect -112 -4767 -110 -4759
rect -106 -4767 -104 -4759
rect -102 -4767 -101 -4759
rect -97 -4767 -96 -4759
rect -94 -4767 -89 -4759
rect -85 -4767 -80 -4759
rect -78 -4767 -77 -4759
rect -73 -4767 -72 -4759
rect -70 -4767 -68 -4759
rect -64 -4767 -62 -4759
rect -60 -4767 -59 -4759
rect -55 -4767 -54 -4759
rect -52 -4767 -47 -4759
rect -43 -4767 -38 -4759
rect -36 -4767 -35 -4759
rect -31 -4767 -30 -4759
rect -28 -4767 -27 -4759
rect 94 -4791 95 -4759
rect 97 -4791 98 -4759
rect 213 -4767 214 -4759
rect 216 -4767 218 -4759
rect 222 -4767 224 -4759
rect 226 -4767 227 -4759
rect 239 -4767 240 -4759
rect 242 -4767 243 -4759
rect 247 -4767 248 -4759
rect 250 -4767 255 -4759
rect 259 -4767 264 -4759
rect 266 -4767 267 -4759
rect 271 -4767 272 -4759
rect 274 -4767 276 -4759
rect 280 -4767 282 -4759
rect 284 -4767 285 -4759
rect 289 -4767 290 -4759
rect 292 -4767 297 -4759
rect 301 -4767 306 -4759
rect 308 -4767 309 -4759
rect 313 -4767 314 -4759
rect 316 -4767 318 -4759
rect 322 -4767 324 -4759
rect 326 -4767 327 -4759
rect 331 -4767 332 -4759
rect 334 -4767 339 -4759
rect 343 -4767 348 -4759
rect 350 -4767 351 -4759
rect 355 -4767 356 -4759
rect 358 -4767 360 -4759
rect 364 -4767 366 -4759
rect 368 -4767 369 -4759
rect 373 -4767 374 -4759
rect 376 -4767 381 -4759
rect 385 -4767 390 -4759
rect 392 -4767 393 -4759
rect 397 -4767 398 -4759
rect 400 -4767 401 -4759
rect 569 -4767 570 -4759
rect 572 -4767 574 -4759
rect 578 -4767 580 -4759
rect 582 -4767 583 -4759
rect 595 -4767 596 -4759
rect 598 -4767 599 -4759
rect 603 -4767 604 -4759
rect 606 -4767 611 -4759
rect 615 -4767 620 -4759
rect 622 -4767 623 -4759
rect 627 -4767 628 -4759
rect 630 -4767 632 -4759
rect 636 -4767 638 -4759
rect 640 -4767 641 -4759
rect 645 -4767 646 -4759
rect 648 -4767 653 -4759
rect 657 -4767 662 -4759
rect 664 -4767 665 -4759
rect 669 -4767 670 -4759
rect 672 -4767 674 -4759
rect 678 -4767 680 -4759
rect 682 -4767 683 -4759
rect 687 -4767 688 -4759
rect 690 -4767 695 -4759
rect 699 -4767 704 -4759
rect 706 -4767 707 -4759
rect 711 -4767 712 -4759
rect 714 -4767 716 -4759
rect 720 -4767 722 -4759
rect 724 -4767 725 -4759
rect 729 -4767 730 -4759
rect 732 -4767 737 -4759
rect 741 -4767 746 -4759
rect 748 -4767 749 -4759
rect 753 -4767 754 -4759
rect 756 -4767 757 -4759
rect 967 -4767 968 -4759
rect 970 -4767 972 -4759
rect 976 -4767 978 -4759
rect 980 -4767 981 -4759
rect 993 -4767 994 -4759
rect 996 -4767 997 -4759
rect 1001 -4767 1002 -4759
rect 1004 -4767 1009 -4759
rect 1013 -4767 1018 -4759
rect 1020 -4767 1021 -4759
rect 1025 -4767 1026 -4759
rect 1028 -4767 1030 -4759
rect 1034 -4767 1036 -4759
rect 1038 -4767 1039 -4759
rect 1043 -4767 1044 -4759
rect 1046 -4767 1051 -4759
rect 1055 -4767 1060 -4759
rect 1062 -4767 1063 -4759
rect 1067 -4767 1068 -4759
rect 1070 -4767 1072 -4759
rect 1076 -4767 1078 -4759
rect 1080 -4767 1081 -4759
rect 1085 -4767 1086 -4759
rect 1088 -4767 1093 -4759
rect 1097 -4767 1102 -4759
rect 1104 -4767 1105 -4759
rect 1109 -4767 1110 -4759
rect 1112 -4767 1114 -4759
rect 1118 -4767 1120 -4759
rect 1122 -4767 1123 -4759
rect 1127 -4767 1128 -4759
rect 1130 -4767 1135 -4759
rect 1139 -4767 1144 -4759
rect 1146 -4767 1147 -4759
rect 1151 -4767 1152 -4759
rect 1154 -4767 1155 -4759
rect 1325 -4767 1326 -4759
rect 1328 -4767 1330 -4759
rect 1334 -4767 1336 -4759
rect 1338 -4767 1339 -4759
rect 1351 -4767 1352 -4759
rect 1354 -4767 1355 -4759
rect 1359 -4767 1360 -4759
rect 1362 -4767 1367 -4759
rect 1371 -4767 1376 -4759
rect 1378 -4767 1379 -4759
rect 1383 -4767 1384 -4759
rect 1386 -4767 1388 -4759
rect 1392 -4767 1394 -4759
rect 1396 -4767 1397 -4759
rect 1401 -4767 1402 -4759
rect 1404 -4767 1409 -4759
rect 1413 -4767 1418 -4759
rect 1420 -4767 1421 -4759
rect 1425 -4767 1426 -4759
rect 1428 -4767 1430 -4759
rect 1434 -4767 1436 -4759
rect 1438 -4767 1439 -4759
rect 1443 -4767 1444 -4759
rect 1446 -4767 1451 -4759
rect 1455 -4767 1460 -4759
rect 1462 -4767 1463 -4759
rect 1467 -4767 1468 -4759
rect 1470 -4767 1472 -4759
rect 1476 -4767 1478 -4759
rect 1480 -4767 1481 -4759
rect 1485 -4767 1486 -4759
rect 1488 -4767 1493 -4759
rect 1497 -4767 1502 -4759
rect 1504 -4767 1505 -4759
rect 1509 -4767 1510 -4759
rect 1512 -4767 1513 -4759
rect -1260 -4885 -1259 -4877
rect -1257 -4885 -1255 -4877
rect -1251 -4885 -1249 -4877
rect -1247 -4885 -1246 -4877
rect -1234 -4885 -1233 -4877
rect -1231 -4885 -1230 -4877
rect -1226 -4885 -1225 -4877
rect -1223 -4885 -1218 -4877
rect -1214 -4885 -1209 -4877
rect -1207 -4885 -1206 -4877
rect -1202 -4885 -1201 -4877
rect -1199 -4885 -1197 -4877
rect -1193 -4885 -1191 -4877
rect -1189 -4885 -1188 -4877
rect -1184 -4885 -1183 -4877
rect -1181 -4885 -1176 -4877
rect -1172 -4885 -1167 -4877
rect -1165 -4885 -1164 -4877
rect -1160 -4885 -1159 -4877
rect -1157 -4885 -1155 -4877
rect -1151 -4885 -1149 -4877
rect -1147 -4885 -1146 -4877
rect -1142 -4885 -1141 -4877
rect -1139 -4885 -1134 -4877
rect -1130 -4885 -1125 -4877
rect -1123 -4885 -1122 -4877
rect -1118 -4885 -1117 -4877
rect -1115 -4885 -1113 -4877
rect -1109 -4885 -1107 -4877
rect -1105 -4885 -1104 -4877
rect -1100 -4885 -1099 -4877
rect -1097 -4885 -1092 -4877
rect -1088 -4885 -1083 -4877
rect -1081 -4885 -1080 -4877
rect -1076 -4885 -1075 -4877
rect -1073 -4885 -1072 -4877
rect -931 -4885 -930 -4877
rect -928 -4885 -926 -4877
rect -922 -4885 -920 -4877
rect -918 -4885 -917 -4877
rect -905 -4885 -904 -4877
rect -902 -4885 -901 -4877
rect -897 -4885 -896 -4877
rect -894 -4885 -889 -4877
rect -885 -4885 -880 -4877
rect -878 -4885 -877 -4877
rect -873 -4885 -872 -4877
rect -870 -4885 -868 -4877
rect -864 -4885 -862 -4877
rect -860 -4885 -859 -4877
rect -855 -4885 -854 -4877
rect -852 -4885 -847 -4877
rect -843 -4885 -838 -4877
rect -836 -4885 -835 -4877
rect -831 -4885 -830 -4877
rect -828 -4885 -826 -4877
rect -822 -4885 -820 -4877
rect -818 -4885 -817 -4877
rect -813 -4885 -812 -4877
rect -810 -4885 -805 -4877
rect -801 -4885 -796 -4877
rect -794 -4885 -793 -4877
rect -789 -4885 -788 -4877
rect -786 -4885 -784 -4877
rect -780 -4885 -778 -4877
rect -776 -4885 -775 -4877
rect -771 -4885 -770 -4877
rect -768 -4885 -763 -4877
rect -759 -4885 -754 -4877
rect -752 -4885 -751 -4877
rect -747 -4885 -746 -4877
rect -744 -4885 -743 -4877
rect -573 -4885 -572 -4877
rect -570 -4885 -568 -4877
rect -564 -4885 -562 -4877
rect -560 -4885 -559 -4877
rect -547 -4885 -546 -4877
rect -544 -4885 -543 -4877
rect -539 -4885 -538 -4877
rect -536 -4885 -531 -4877
rect -527 -4885 -522 -4877
rect -520 -4885 -519 -4877
rect -515 -4885 -514 -4877
rect -512 -4885 -510 -4877
rect -506 -4885 -504 -4877
rect -502 -4885 -501 -4877
rect -497 -4885 -496 -4877
rect -494 -4885 -489 -4877
rect -485 -4885 -480 -4877
rect -478 -4885 -477 -4877
rect -473 -4885 -472 -4877
rect -470 -4885 -468 -4877
rect -464 -4885 -462 -4877
rect -460 -4885 -459 -4877
rect -455 -4885 -454 -4877
rect -452 -4885 -447 -4877
rect -443 -4885 -438 -4877
rect -436 -4885 -435 -4877
rect -431 -4885 -430 -4877
rect -428 -4885 -426 -4877
rect -422 -4885 -420 -4877
rect -418 -4885 -417 -4877
rect -413 -4885 -412 -4877
rect -410 -4885 -405 -4877
rect -401 -4885 -396 -4877
rect -394 -4885 -393 -4877
rect -389 -4885 -388 -4877
rect -386 -4885 -385 -4877
rect -215 -4885 -214 -4877
rect -212 -4885 -210 -4877
rect -206 -4885 -204 -4877
rect -202 -4885 -201 -4877
rect -189 -4885 -188 -4877
rect -186 -4885 -185 -4877
rect -181 -4885 -180 -4877
rect -178 -4885 -173 -4877
rect -169 -4885 -164 -4877
rect -162 -4885 -161 -4877
rect -157 -4885 -156 -4877
rect -154 -4885 -152 -4877
rect -148 -4885 -146 -4877
rect -144 -4885 -143 -4877
rect -139 -4885 -138 -4877
rect -136 -4885 -131 -4877
rect -127 -4885 -122 -4877
rect -120 -4885 -119 -4877
rect -115 -4885 -114 -4877
rect -112 -4885 -110 -4877
rect -106 -4885 -104 -4877
rect -102 -4885 -101 -4877
rect -97 -4885 -96 -4877
rect -94 -4885 -89 -4877
rect -85 -4885 -80 -4877
rect -78 -4885 -77 -4877
rect -73 -4885 -72 -4877
rect -70 -4885 -68 -4877
rect -64 -4885 -62 -4877
rect -60 -4885 -59 -4877
rect -55 -4885 -54 -4877
rect -52 -4885 -47 -4877
rect -43 -4885 -38 -4877
rect -36 -4885 -35 -4877
rect -31 -4885 -30 -4877
rect -28 -4885 -27 -4877
rect 213 -4885 214 -4877
rect 216 -4885 218 -4877
rect 222 -4885 224 -4877
rect 226 -4885 227 -4877
rect 239 -4885 240 -4877
rect 242 -4885 243 -4877
rect 247 -4885 248 -4877
rect 250 -4885 255 -4877
rect 259 -4885 264 -4877
rect 266 -4885 267 -4877
rect 271 -4885 272 -4877
rect 274 -4885 276 -4877
rect 280 -4885 282 -4877
rect 284 -4885 285 -4877
rect 289 -4885 290 -4877
rect 292 -4885 297 -4877
rect 301 -4885 306 -4877
rect 308 -4885 309 -4877
rect 313 -4885 314 -4877
rect 316 -4885 318 -4877
rect 322 -4885 324 -4877
rect 326 -4885 327 -4877
rect 331 -4885 332 -4877
rect 334 -4885 339 -4877
rect 343 -4885 348 -4877
rect 350 -4885 351 -4877
rect 355 -4885 356 -4877
rect 358 -4885 360 -4877
rect 364 -4885 366 -4877
rect 368 -4885 369 -4877
rect 373 -4885 374 -4877
rect 376 -4885 381 -4877
rect 385 -4885 390 -4877
rect 392 -4885 393 -4877
rect 397 -4885 398 -4877
rect 400 -4885 401 -4877
rect -1335 -5002 -1334 -4994
rect -1332 -5002 -1331 -4994
rect -1327 -5002 -1326 -4994
rect -1324 -5002 -1322 -4994
rect -1318 -5002 -1316 -4994
rect -1314 -5002 -1313 -4994
rect -931 -5002 -930 -4994
rect -928 -5002 -927 -4994
rect -923 -5002 -922 -4994
rect -920 -5002 -918 -4994
rect -914 -5002 -912 -4994
rect -910 -5002 -909 -4994
rect -573 -5002 -572 -4994
rect -570 -5002 -569 -4994
rect -565 -5002 -564 -4994
rect -562 -5002 -560 -4994
rect -556 -5002 -554 -4994
rect -552 -5002 -551 -4994
rect -215 -5002 -214 -4994
rect -212 -5002 -211 -4994
rect -207 -5002 -206 -4994
rect -204 -5002 -202 -4994
rect -198 -5002 -196 -4994
rect -194 -5002 -193 -4994
rect 213 -5002 214 -4994
rect 216 -5002 217 -4994
rect 221 -5002 222 -4994
rect 224 -5002 226 -4994
rect 230 -5002 232 -4994
rect 234 -5002 235 -4994
rect 569 -5002 570 -4994
rect 572 -5002 573 -4994
rect 577 -5002 578 -4994
rect 580 -5002 582 -4994
rect 586 -5002 588 -4994
rect 590 -5002 591 -4994
rect 967 -5002 968 -4994
rect 970 -5002 971 -4994
rect 975 -5002 976 -4994
rect 978 -5002 980 -4994
rect 984 -5002 986 -4994
rect 988 -5002 989 -4994
rect 1325 -5002 1326 -4994
rect 1328 -5002 1329 -4994
rect 1333 -5002 1334 -4994
rect 1336 -5002 1338 -4994
rect 1342 -5002 1344 -4994
rect 1346 -5002 1347 -4994
rect -1260 -5121 -1259 -5113
rect -1257 -5121 -1255 -5113
rect -1251 -5121 -1249 -5113
rect -1247 -5121 -1246 -5113
rect -1234 -5121 -1233 -5113
rect -1231 -5121 -1223 -5113
rect -1221 -5121 -1220 -5113
rect -1216 -5121 -1215 -5113
rect -1213 -5121 -1205 -5113
rect -1203 -5121 -1198 -5113
rect -1194 -5121 -1189 -5113
rect -1187 -5121 -1186 -5113
rect -1182 -5121 -1181 -5113
rect -1179 -5121 -1177 -5113
rect -1173 -5121 -1171 -5113
rect -1169 -5121 -1168 -5113
rect -931 -5121 -930 -5113
rect -928 -5121 -926 -5113
rect -922 -5121 -920 -5113
rect -918 -5121 -917 -5113
rect -905 -5121 -904 -5113
rect -902 -5121 -900 -5113
rect -896 -5121 -894 -5113
rect -892 -5121 -891 -5113
rect -879 -5121 -878 -5113
rect -876 -5121 -868 -5113
rect -866 -5121 -865 -5113
rect -861 -5121 -860 -5113
rect -858 -5121 -850 -5113
rect -848 -5121 -843 -5113
rect -839 -5121 -834 -5113
rect -832 -5121 -831 -5113
rect -827 -5121 -826 -5113
rect -824 -5121 -822 -5113
rect -818 -5121 -816 -5113
rect -814 -5121 -813 -5113
rect -801 -5121 -800 -5113
rect -798 -5121 -790 -5113
rect -788 -5121 -787 -5113
rect -783 -5121 -782 -5113
rect -780 -5121 -772 -5113
rect -770 -5121 -765 -5113
rect -761 -5121 -756 -5113
rect -754 -5121 -753 -5113
rect -749 -5121 -748 -5113
rect -746 -5121 -741 -5113
rect -737 -5121 -732 -5113
rect -730 -5121 -729 -5113
rect -717 -5121 -716 -5113
rect -714 -5121 -708 -5113
rect -706 -5121 -704 -5113
rect -700 -5121 -698 -5113
rect -696 -5121 -695 -5113
rect -573 -5121 -572 -5113
rect -570 -5121 -568 -5113
rect -564 -5121 -562 -5113
rect -560 -5121 -559 -5113
rect -547 -5121 -546 -5113
rect -544 -5121 -542 -5113
rect -538 -5121 -536 -5113
rect -534 -5121 -533 -5113
rect -521 -5121 -520 -5113
rect -518 -5121 -510 -5113
rect -508 -5121 -507 -5113
rect -503 -5121 -502 -5113
rect -500 -5121 -492 -5113
rect -490 -5121 -485 -5113
rect -481 -5121 -476 -5113
rect -474 -5121 -473 -5113
rect -469 -5121 -468 -5113
rect -466 -5121 -464 -5113
rect -460 -5121 -458 -5113
rect -456 -5121 -455 -5113
rect -443 -5121 -442 -5113
rect -440 -5121 -432 -5113
rect -430 -5121 -429 -5113
rect -425 -5121 -424 -5113
rect -422 -5121 -414 -5113
rect -412 -5121 -407 -5113
rect -403 -5121 -398 -5113
rect -396 -5121 -395 -5113
rect -391 -5121 -390 -5113
rect -388 -5121 -383 -5113
rect -379 -5121 -374 -5113
rect -372 -5121 -371 -5113
rect -359 -5121 -358 -5113
rect -356 -5121 -350 -5113
rect -348 -5121 -346 -5113
rect -342 -5121 -340 -5113
rect -338 -5121 -337 -5113
rect -215 -5121 -214 -5113
rect -212 -5121 -210 -5113
rect -206 -5121 -204 -5113
rect -202 -5121 -201 -5113
rect -189 -5121 -188 -5113
rect -186 -5121 -184 -5113
rect -180 -5121 -178 -5113
rect -176 -5121 -175 -5113
rect -163 -5121 -162 -5113
rect -160 -5121 -152 -5113
rect -150 -5121 -149 -5113
rect -145 -5121 -144 -5113
rect -142 -5121 -134 -5113
rect -132 -5121 -127 -5113
rect -123 -5121 -118 -5113
rect -116 -5121 -115 -5113
rect -111 -5121 -110 -5113
rect -108 -5121 -106 -5113
rect -102 -5121 -100 -5113
rect -98 -5121 -97 -5113
rect -85 -5121 -84 -5113
rect -82 -5121 -74 -5113
rect -72 -5121 -71 -5113
rect -67 -5121 -66 -5113
rect -64 -5121 -56 -5113
rect -54 -5121 -49 -5113
rect -45 -5121 -40 -5113
rect -38 -5121 -37 -5113
rect -33 -5121 -32 -5113
rect -30 -5121 -25 -5113
rect -21 -5121 -16 -5113
rect -14 -5121 -13 -5113
rect -1 -5121 0 -5113
rect 2 -5121 8 -5113
rect 10 -5121 12 -5113
rect 16 -5121 18 -5113
rect 20 -5121 21 -5113
rect 213 -5121 214 -5113
rect 216 -5121 218 -5113
rect 222 -5121 224 -5113
rect 226 -5121 227 -5113
rect 239 -5121 240 -5113
rect 242 -5121 244 -5113
rect 248 -5121 250 -5113
rect 252 -5121 253 -5113
rect 265 -5121 266 -5113
rect 268 -5121 276 -5113
rect 278 -5121 279 -5113
rect 283 -5121 284 -5113
rect 286 -5121 294 -5113
rect 296 -5121 301 -5113
rect 305 -5121 310 -5113
rect 312 -5121 313 -5113
rect 317 -5121 318 -5113
rect 320 -5121 322 -5113
rect 326 -5121 328 -5113
rect 330 -5121 331 -5113
rect 343 -5121 344 -5113
rect 346 -5121 354 -5113
rect 356 -5121 357 -5113
rect 361 -5121 362 -5113
rect 364 -5121 372 -5113
rect 374 -5121 379 -5113
rect 383 -5121 388 -5113
rect 390 -5121 391 -5113
rect 395 -5121 396 -5113
rect 398 -5121 403 -5113
rect 407 -5121 412 -5113
rect 414 -5121 415 -5113
rect 427 -5121 428 -5113
rect 430 -5121 436 -5113
rect 438 -5121 440 -5113
rect 444 -5121 446 -5113
rect 448 -5121 449 -5113
rect 569 -5121 570 -5113
rect 572 -5121 574 -5113
rect 578 -5121 580 -5113
rect 582 -5121 583 -5113
rect 595 -5121 596 -5113
rect 598 -5121 600 -5113
rect 604 -5121 606 -5113
rect 608 -5121 609 -5113
rect 621 -5121 622 -5113
rect 624 -5121 632 -5113
rect 634 -5121 635 -5113
rect 639 -5121 640 -5113
rect 642 -5121 650 -5113
rect 652 -5121 657 -5113
rect 661 -5121 666 -5113
rect 668 -5121 669 -5113
rect 673 -5121 674 -5113
rect 676 -5121 678 -5113
rect 682 -5121 684 -5113
rect 686 -5121 687 -5113
rect 699 -5121 700 -5113
rect 702 -5121 710 -5113
rect 712 -5121 713 -5113
rect 717 -5121 718 -5113
rect 720 -5121 728 -5113
rect 730 -5121 735 -5113
rect 739 -5121 744 -5113
rect 746 -5121 747 -5113
rect 751 -5121 752 -5113
rect 754 -5121 759 -5113
rect 763 -5121 768 -5113
rect 770 -5121 771 -5113
rect 783 -5121 784 -5113
rect 786 -5121 792 -5113
rect 794 -5121 796 -5113
rect 800 -5121 802 -5113
rect 804 -5121 805 -5113
rect 967 -5121 968 -5113
rect 970 -5121 972 -5113
rect 976 -5121 978 -5113
rect 980 -5121 981 -5113
rect 993 -5121 994 -5113
rect 996 -5121 998 -5113
rect 1002 -5121 1004 -5113
rect 1006 -5121 1007 -5113
rect 1019 -5121 1020 -5113
rect 1022 -5121 1030 -5113
rect 1032 -5121 1033 -5113
rect 1037 -5121 1038 -5113
rect 1040 -5121 1048 -5113
rect 1050 -5121 1055 -5113
rect 1059 -5121 1064 -5113
rect 1066 -5121 1067 -5113
rect 1071 -5121 1072 -5113
rect 1074 -5121 1076 -5113
rect 1080 -5121 1082 -5113
rect 1084 -5121 1085 -5113
rect 1097 -5121 1098 -5113
rect 1100 -5121 1108 -5113
rect 1110 -5121 1111 -5113
rect 1115 -5121 1116 -5113
rect 1118 -5121 1126 -5113
rect 1128 -5121 1133 -5113
rect 1137 -5121 1142 -5113
rect 1144 -5121 1145 -5113
rect 1149 -5121 1150 -5113
rect 1152 -5121 1157 -5113
rect 1161 -5121 1166 -5113
rect 1168 -5121 1169 -5113
rect 1181 -5121 1182 -5113
rect 1184 -5121 1190 -5113
rect 1192 -5121 1194 -5113
rect 1198 -5121 1200 -5113
rect 1202 -5121 1203 -5113
rect 1325 -5121 1326 -5113
rect 1328 -5121 1330 -5113
rect 1334 -5121 1336 -5113
rect 1338 -5121 1339 -5113
rect 1351 -5121 1352 -5113
rect 1354 -5121 1356 -5113
rect 1360 -5121 1362 -5113
rect 1364 -5121 1365 -5113
rect 1377 -5121 1378 -5113
rect 1380 -5121 1388 -5113
rect 1390 -5121 1391 -5113
rect 1395 -5121 1396 -5113
rect 1398 -5121 1406 -5113
rect 1408 -5121 1413 -5113
rect 1417 -5121 1422 -5113
rect 1424 -5121 1425 -5113
rect 1429 -5121 1430 -5113
rect 1432 -5121 1434 -5113
rect 1438 -5121 1440 -5113
rect 1442 -5121 1443 -5113
rect 1455 -5121 1456 -5113
rect 1458 -5121 1466 -5113
rect 1468 -5121 1469 -5113
rect 1473 -5121 1474 -5113
rect 1476 -5121 1484 -5113
rect 1486 -5121 1491 -5113
rect 1495 -5121 1500 -5113
rect 1502 -5121 1503 -5113
rect 1507 -5121 1508 -5113
rect 1510 -5121 1515 -5113
rect 1519 -5121 1524 -5113
rect 1526 -5121 1527 -5113
rect 1539 -5121 1540 -5113
rect 1542 -5121 1548 -5113
rect 1550 -5121 1552 -5113
rect 1556 -5121 1558 -5113
rect 1560 -5121 1561 -5113
rect -1260 -5240 -1259 -5232
rect -1257 -5240 -1255 -5232
rect -1251 -5240 -1249 -5232
rect -1247 -5240 -1246 -5232
rect -1234 -5240 -1233 -5232
rect -1231 -5240 -1230 -5232
rect -1226 -5240 -1225 -5232
rect -1223 -5240 -1218 -5232
rect -1214 -5240 -1209 -5232
rect -1207 -5240 -1206 -5232
rect -1202 -5240 -1201 -5232
rect -1199 -5240 -1197 -5232
rect -1193 -5240 -1191 -5232
rect -1189 -5240 -1188 -5232
rect -1184 -5240 -1183 -5232
rect -1181 -5240 -1176 -5232
rect -1172 -5240 -1167 -5232
rect -1165 -5240 -1164 -5232
rect -1160 -5240 -1159 -5232
rect -1157 -5240 -1155 -5232
rect -1151 -5240 -1149 -5232
rect -1147 -5240 -1146 -5232
rect -1142 -5240 -1141 -5232
rect -1139 -5240 -1134 -5232
rect -1130 -5240 -1125 -5232
rect -1123 -5240 -1122 -5232
rect -1118 -5240 -1117 -5232
rect -1115 -5240 -1113 -5232
rect -1109 -5240 -1107 -5232
rect -1105 -5240 -1104 -5232
rect -1100 -5240 -1099 -5232
rect -1097 -5240 -1092 -5232
rect -1088 -5240 -1083 -5232
rect -1081 -5240 -1080 -5232
rect -1076 -5240 -1075 -5232
rect -1073 -5240 -1072 -5232
rect -931 -5240 -930 -5232
rect -928 -5240 -926 -5232
rect -922 -5240 -920 -5232
rect -918 -5240 -917 -5232
rect -905 -5240 -904 -5232
rect -902 -5240 -901 -5232
rect -897 -5240 -896 -5232
rect -894 -5240 -889 -5232
rect -885 -5240 -880 -5232
rect -878 -5240 -877 -5232
rect -873 -5240 -872 -5232
rect -870 -5240 -868 -5232
rect -864 -5240 -862 -5232
rect -860 -5240 -859 -5232
rect -855 -5240 -854 -5232
rect -852 -5240 -847 -5232
rect -843 -5240 -838 -5232
rect -836 -5240 -835 -5232
rect -831 -5240 -830 -5232
rect -828 -5240 -826 -5232
rect -822 -5240 -820 -5232
rect -818 -5240 -817 -5232
rect -813 -5240 -812 -5232
rect -810 -5240 -805 -5232
rect -801 -5240 -796 -5232
rect -794 -5240 -793 -5232
rect -789 -5240 -788 -5232
rect -786 -5240 -784 -5232
rect -780 -5240 -778 -5232
rect -776 -5240 -775 -5232
rect -771 -5240 -770 -5232
rect -768 -5240 -763 -5232
rect -759 -5240 -754 -5232
rect -752 -5240 -751 -5232
rect -747 -5240 -746 -5232
rect -744 -5240 -743 -5232
rect -1260 -5361 -1259 -5353
rect -1257 -5361 -1255 -5353
rect -1251 -5361 -1249 -5353
rect -1247 -5361 -1246 -5353
rect -1234 -5361 -1233 -5353
rect -1231 -5361 -1230 -5353
rect -1226 -5361 -1225 -5353
rect -1223 -5361 -1218 -5353
rect -1214 -5361 -1209 -5353
rect -1207 -5361 -1206 -5353
rect -1202 -5361 -1201 -5353
rect -1199 -5361 -1197 -5353
rect -1193 -5361 -1191 -5353
rect -1189 -5361 -1188 -5353
rect -1184 -5361 -1183 -5353
rect -1181 -5361 -1176 -5353
rect -1172 -5361 -1167 -5353
rect -1165 -5361 -1164 -5353
rect -1160 -5361 -1159 -5353
rect -1157 -5361 -1155 -5353
rect -1151 -5361 -1149 -5353
rect -1147 -5361 -1146 -5353
rect -1142 -5361 -1141 -5353
rect -1139 -5361 -1134 -5353
rect -1130 -5361 -1125 -5353
rect -1123 -5361 -1122 -5353
rect -1118 -5361 -1117 -5353
rect -1115 -5361 -1113 -5353
rect -1109 -5361 -1107 -5353
rect -1105 -5361 -1104 -5353
rect -1100 -5361 -1099 -5353
rect -1097 -5361 -1092 -5353
rect -1088 -5361 -1083 -5353
rect -1081 -5361 -1080 -5353
rect -1076 -5361 -1075 -5353
rect -1073 -5361 -1072 -5353
rect -1022 -5361 -1021 -5353
rect -1019 -5361 -1018 -5353
rect -931 -5361 -930 -5353
rect -928 -5361 -926 -5353
rect -922 -5361 -920 -5353
rect -918 -5361 -917 -5353
rect -905 -5361 -904 -5353
rect -902 -5361 -901 -5353
rect -897 -5361 -896 -5353
rect -894 -5361 -889 -5353
rect -885 -5361 -880 -5353
rect -878 -5361 -877 -5353
rect -873 -5361 -872 -5353
rect -870 -5361 -868 -5353
rect -864 -5361 -862 -5353
rect -860 -5361 -859 -5353
rect -855 -5361 -854 -5353
rect -852 -5361 -847 -5353
rect -843 -5361 -838 -5353
rect -836 -5361 -835 -5353
rect -831 -5361 -830 -5353
rect -828 -5361 -826 -5353
rect -822 -5361 -820 -5353
rect -818 -5361 -817 -5353
rect -813 -5361 -812 -5353
rect -810 -5361 -805 -5353
rect -801 -5361 -796 -5353
rect -794 -5361 -793 -5353
rect -789 -5361 -788 -5353
rect -786 -5361 -784 -5353
rect -780 -5361 -778 -5353
rect -776 -5361 -775 -5353
rect -771 -5361 -770 -5353
rect -768 -5361 -763 -5353
rect -759 -5361 -754 -5353
rect -752 -5361 -751 -5353
rect -747 -5361 -746 -5353
rect -744 -5361 -743 -5353
rect -669 -5369 -668 -5353
rect -666 -5369 -665 -5353
rect -573 -5361 -572 -5353
rect -570 -5361 -568 -5353
rect -564 -5361 -562 -5353
rect -560 -5361 -559 -5353
rect -547 -5361 -546 -5353
rect -544 -5361 -543 -5353
rect -539 -5361 -538 -5353
rect -536 -5361 -531 -5353
rect -527 -5361 -522 -5353
rect -520 -5361 -519 -5353
rect -515 -5361 -514 -5353
rect -512 -5361 -510 -5353
rect -506 -5361 -504 -5353
rect -502 -5361 -501 -5353
rect -497 -5361 -496 -5353
rect -494 -5361 -489 -5353
rect -485 -5361 -480 -5353
rect -478 -5361 -477 -5353
rect -473 -5361 -472 -5353
rect -470 -5361 -468 -5353
rect -464 -5361 -462 -5353
rect -460 -5361 -459 -5353
rect -455 -5361 -454 -5353
rect -452 -5361 -447 -5353
rect -443 -5361 -438 -5353
rect -436 -5361 -435 -5353
rect -431 -5361 -430 -5353
rect -428 -5361 -426 -5353
rect -422 -5361 -420 -5353
rect -418 -5361 -417 -5353
rect -413 -5361 -412 -5353
rect -410 -5361 -405 -5353
rect -401 -5361 -396 -5353
rect -394 -5361 -393 -5353
rect -389 -5361 -388 -5353
rect -386 -5361 -385 -5353
rect -323 -5361 -322 -5353
rect -320 -5361 -319 -5353
rect -215 -5361 -214 -5353
rect -212 -5361 -210 -5353
rect -206 -5361 -204 -5353
rect -202 -5361 -201 -5353
rect -189 -5361 -188 -5353
rect -186 -5361 -185 -5353
rect -181 -5361 -180 -5353
rect -178 -5361 -173 -5353
rect -169 -5361 -164 -5353
rect -162 -5361 -161 -5353
rect -157 -5361 -156 -5353
rect -154 -5361 -152 -5353
rect -148 -5361 -146 -5353
rect -144 -5361 -143 -5353
rect -139 -5361 -138 -5353
rect -136 -5361 -131 -5353
rect -127 -5361 -122 -5353
rect -120 -5361 -119 -5353
rect -115 -5361 -114 -5353
rect -112 -5361 -110 -5353
rect -106 -5361 -104 -5353
rect -102 -5361 -101 -5353
rect -97 -5361 -96 -5353
rect -94 -5361 -89 -5353
rect -85 -5361 -80 -5353
rect -78 -5361 -77 -5353
rect -73 -5361 -72 -5353
rect -70 -5361 -68 -5353
rect -64 -5361 -62 -5353
rect -60 -5361 -59 -5353
rect -55 -5361 -54 -5353
rect -52 -5361 -47 -5353
rect -43 -5361 -38 -5353
rect -36 -5361 -35 -5353
rect -31 -5361 -30 -5353
rect -28 -5361 -27 -5353
rect 213 -5361 214 -5353
rect 216 -5361 218 -5353
rect 222 -5361 224 -5353
rect 226 -5361 227 -5353
rect 239 -5361 240 -5353
rect 242 -5361 243 -5353
rect 247 -5361 248 -5353
rect 250 -5361 255 -5353
rect 259 -5361 264 -5353
rect 266 -5361 267 -5353
rect 271 -5361 272 -5353
rect 274 -5361 276 -5353
rect 280 -5361 282 -5353
rect 284 -5361 285 -5353
rect 289 -5361 290 -5353
rect 292 -5361 297 -5353
rect 301 -5361 306 -5353
rect 308 -5361 309 -5353
rect 313 -5361 314 -5353
rect 316 -5361 318 -5353
rect 322 -5361 324 -5353
rect 326 -5361 327 -5353
rect 331 -5361 332 -5353
rect 334 -5361 339 -5353
rect 343 -5361 348 -5353
rect 350 -5361 351 -5353
rect 355 -5361 356 -5353
rect 358 -5361 360 -5353
rect 364 -5361 366 -5353
rect 368 -5361 369 -5353
rect 373 -5361 374 -5353
rect 376 -5361 381 -5353
rect 385 -5361 390 -5353
rect 392 -5361 393 -5353
rect 397 -5361 398 -5353
rect 400 -5361 401 -5353
rect 470 -5361 471 -5353
rect 473 -5361 474 -5353
rect 569 -5361 570 -5353
rect 572 -5361 574 -5353
rect 578 -5361 580 -5353
rect 582 -5361 583 -5353
rect 595 -5361 596 -5353
rect 598 -5361 599 -5353
rect 603 -5361 604 -5353
rect 606 -5361 611 -5353
rect 615 -5361 620 -5353
rect 622 -5361 623 -5353
rect 627 -5361 628 -5353
rect 630 -5361 632 -5353
rect 636 -5361 638 -5353
rect 640 -5361 641 -5353
rect 645 -5361 646 -5353
rect 648 -5361 653 -5353
rect 657 -5361 662 -5353
rect 664 -5361 665 -5353
rect 669 -5361 670 -5353
rect 672 -5361 674 -5353
rect 678 -5361 680 -5353
rect 682 -5361 683 -5353
rect 687 -5361 688 -5353
rect 690 -5361 695 -5353
rect 699 -5361 704 -5353
rect 706 -5361 707 -5353
rect 711 -5361 712 -5353
rect 714 -5361 716 -5353
rect 720 -5361 722 -5353
rect 724 -5361 725 -5353
rect 729 -5361 730 -5353
rect 732 -5361 737 -5353
rect 741 -5361 746 -5353
rect 748 -5361 749 -5353
rect 753 -5361 754 -5353
rect 756 -5361 757 -5353
rect 871 -5369 872 -5353
rect 874 -5369 875 -5353
rect 967 -5361 968 -5353
rect 970 -5361 972 -5353
rect 976 -5361 978 -5353
rect 980 -5361 981 -5353
rect 993 -5361 994 -5353
rect 996 -5361 997 -5353
rect 1001 -5361 1002 -5353
rect 1004 -5361 1009 -5353
rect 1013 -5361 1018 -5353
rect 1020 -5361 1021 -5353
rect 1025 -5361 1026 -5353
rect 1028 -5361 1030 -5353
rect 1034 -5361 1036 -5353
rect 1038 -5361 1039 -5353
rect 1043 -5361 1044 -5353
rect 1046 -5361 1051 -5353
rect 1055 -5361 1060 -5353
rect 1062 -5361 1063 -5353
rect 1067 -5361 1068 -5353
rect 1070 -5361 1072 -5353
rect 1076 -5361 1078 -5353
rect 1080 -5361 1081 -5353
rect 1085 -5361 1086 -5353
rect 1088 -5361 1093 -5353
rect 1097 -5361 1102 -5353
rect 1104 -5361 1105 -5353
rect 1109 -5361 1110 -5353
rect 1112 -5361 1114 -5353
rect 1118 -5361 1120 -5353
rect 1122 -5361 1123 -5353
rect 1127 -5361 1128 -5353
rect 1130 -5361 1135 -5353
rect 1139 -5361 1144 -5353
rect 1146 -5361 1147 -5353
rect 1151 -5361 1152 -5353
rect 1154 -5361 1155 -5353
rect 1214 -5361 1215 -5353
rect 1217 -5361 1218 -5353
rect 1325 -5361 1326 -5353
rect 1328 -5361 1330 -5353
rect 1334 -5361 1336 -5353
rect 1338 -5361 1339 -5353
rect 1351 -5361 1352 -5353
rect 1354 -5361 1355 -5353
rect 1359 -5361 1360 -5353
rect 1362 -5361 1367 -5353
rect 1371 -5361 1376 -5353
rect 1378 -5361 1379 -5353
rect 1383 -5361 1384 -5353
rect 1386 -5361 1388 -5353
rect 1392 -5361 1394 -5353
rect 1396 -5361 1397 -5353
rect 1401 -5361 1402 -5353
rect 1404 -5361 1409 -5353
rect 1413 -5361 1418 -5353
rect 1420 -5361 1421 -5353
rect 1425 -5361 1426 -5353
rect 1428 -5361 1430 -5353
rect 1434 -5361 1436 -5353
rect 1438 -5361 1439 -5353
rect 1443 -5361 1444 -5353
rect 1446 -5361 1451 -5353
rect 1455 -5361 1460 -5353
rect 1462 -5361 1463 -5353
rect 1467 -5361 1468 -5353
rect 1470 -5361 1472 -5353
rect 1476 -5361 1478 -5353
rect 1480 -5361 1481 -5353
rect 1485 -5361 1486 -5353
rect 1488 -5361 1493 -5353
rect 1497 -5361 1502 -5353
rect 1504 -5361 1505 -5353
rect 1509 -5361 1510 -5353
rect 1512 -5361 1513 -5353
rect -1260 -5481 -1259 -5473
rect -1257 -5481 -1255 -5473
rect -1251 -5481 -1249 -5473
rect -1247 -5481 -1246 -5473
rect -1234 -5481 -1233 -5473
rect -1231 -5481 -1230 -5473
rect -1226 -5481 -1225 -5473
rect -1223 -5481 -1218 -5473
rect -1214 -5481 -1209 -5473
rect -1207 -5481 -1206 -5473
rect -1202 -5481 -1201 -5473
rect -1199 -5481 -1197 -5473
rect -1193 -5481 -1191 -5473
rect -1189 -5481 -1188 -5473
rect -1184 -5481 -1183 -5473
rect -1181 -5481 -1176 -5473
rect -1172 -5481 -1167 -5473
rect -1165 -5481 -1164 -5473
rect -1160 -5481 -1159 -5473
rect -1157 -5481 -1155 -5473
rect -1151 -5481 -1149 -5473
rect -1147 -5481 -1146 -5473
rect -1142 -5481 -1141 -5473
rect -1139 -5481 -1134 -5473
rect -1130 -5481 -1125 -5473
rect -1123 -5481 -1122 -5473
rect -1118 -5481 -1117 -5473
rect -1115 -5481 -1113 -5473
rect -1109 -5481 -1107 -5473
rect -1105 -5481 -1104 -5473
rect -1100 -5481 -1099 -5473
rect -1097 -5481 -1092 -5473
rect -1088 -5481 -1083 -5473
rect -1081 -5481 -1080 -5473
rect -1076 -5481 -1075 -5473
rect -1073 -5481 -1072 -5473
rect -1022 -5481 -1021 -5473
rect -1019 -5481 -1018 -5473
rect -931 -5481 -930 -5473
rect -928 -5481 -926 -5473
rect -922 -5481 -920 -5473
rect -918 -5481 -917 -5473
rect -905 -5481 -904 -5473
rect -902 -5481 -901 -5473
rect -897 -5481 -896 -5473
rect -894 -5481 -889 -5473
rect -885 -5481 -880 -5473
rect -878 -5481 -877 -5473
rect -873 -5481 -872 -5473
rect -870 -5481 -868 -5473
rect -864 -5481 -862 -5473
rect -860 -5481 -859 -5473
rect -855 -5481 -854 -5473
rect -852 -5481 -847 -5473
rect -843 -5481 -838 -5473
rect -836 -5481 -835 -5473
rect -831 -5481 -830 -5473
rect -828 -5481 -826 -5473
rect -822 -5481 -820 -5473
rect -818 -5481 -817 -5473
rect -813 -5481 -812 -5473
rect -810 -5481 -805 -5473
rect -801 -5481 -796 -5473
rect -794 -5481 -793 -5473
rect -789 -5481 -788 -5473
rect -786 -5481 -784 -5473
rect -780 -5481 -778 -5473
rect -776 -5481 -775 -5473
rect -771 -5481 -770 -5473
rect -768 -5481 -763 -5473
rect -759 -5481 -754 -5473
rect -752 -5481 -751 -5473
rect -747 -5481 -746 -5473
rect -744 -5481 -743 -5473
rect -573 -5481 -572 -5473
rect -570 -5481 -568 -5473
rect -564 -5481 -562 -5473
rect -560 -5481 -559 -5473
rect -547 -5481 -546 -5473
rect -544 -5481 -543 -5473
rect -539 -5481 -538 -5473
rect -536 -5481 -531 -5473
rect -527 -5481 -522 -5473
rect -520 -5481 -519 -5473
rect -515 -5481 -514 -5473
rect -512 -5481 -510 -5473
rect -506 -5481 -504 -5473
rect -502 -5481 -501 -5473
rect -497 -5481 -496 -5473
rect -494 -5481 -489 -5473
rect -485 -5481 -480 -5473
rect -478 -5481 -477 -5473
rect -473 -5481 -472 -5473
rect -470 -5481 -468 -5473
rect -464 -5481 -462 -5473
rect -460 -5481 -459 -5473
rect -455 -5481 -454 -5473
rect -452 -5481 -447 -5473
rect -443 -5481 -438 -5473
rect -436 -5481 -435 -5473
rect -431 -5481 -430 -5473
rect -428 -5481 -426 -5473
rect -422 -5481 -420 -5473
rect -418 -5481 -417 -5473
rect -413 -5481 -412 -5473
rect -410 -5481 -405 -5473
rect -401 -5481 -396 -5473
rect -394 -5481 -393 -5473
rect -389 -5481 -388 -5473
rect -386 -5481 -385 -5473
rect -323 -5481 -322 -5473
rect -320 -5481 -319 -5473
rect -215 -5481 -214 -5473
rect -212 -5481 -210 -5473
rect -206 -5481 -204 -5473
rect -202 -5481 -201 -5473
rect -189 -5481 -188 -5473
rect -186 -5481 -185 -5473
rect -181 -5481 -180 -5473
rect -178 -5481 -173 -5473
rect -169 -5481 -164 -5473
rect -162 -5481 -161 -5473
rect -157 -5481 -156 -5473
rect -154 -5481 -152 -5473
rect -148 -5481 -146 -5473
rect -144 -5481 -143 -5473
rect -139 -5481 -138 -5473
rect -136 -5481 -131 -5473
rect -127 -5481 -122 -5473
rect -120 -5481 -119 -5473
rect -115 -5481 -114 -5473
rect -112 -5481 -110 -5473
rect -106 -5481 -104 -5473
rect -102 -5481 -101 -5473
rect -97 -5481 -96 -5473
rect -94 -5481 -89 -5473
rect -85 -5481 -80 -5473
rect -78 -5481 -77 -5473
rect -73 -5481 -72 -5473
rect -70 -5481 -68 -5473
rect -64 -5481 -62 -5473
rect -60 -5481 -59 -5473
rect -55 -5481 -54 -5473
rect -52 -5481 -47 -5473
rect -43 -5481 -38 -5473
rect -36 -5481 -35 -5473
rect -31 -5481 -30 -5473
rect -28 -5481 -27 -5473
rect 213 -5481 214 -5473
rect 216 -5481 218 -5473
rect 222 -5481 224 -5473
rect 226 -5481 227 -5473
rect 239 -5481 240 -5473
rect 242 -5481 243 -5473
rect 247 -5481 248 -5473
rect 250 -5481 255 -5473
rect 259 -5481 264 -5473
rect 266 -5481 267 -5473
rect 271 -5481 272 -5473
rect 274 -5481 276 -5473
rect 280 -5481 282 -5473
rect 284 -5481 285 -5473
rect 289 -5481 290 -5473
rect 292 -5481 297 -5473
rect 301 -5481 306 -5473
rect 308 -5481 309 -5473
rect 313 -5481 314 -5473
rect 316 -5481 318 -5473
rect 322 -5481 324 -5473
rect 326 -5481 327 -5473
rect 331 -5481 332 -5473
rect 334 -5481 339 -5473
rect 343 -5481 348 -5473
rect 350 -5481 351 -5473
rect 355 -5481 356 -5473
rect 358 -5481 360 -5473
rect 364 -5481 366 -5473
rect 368 -5481 369 -5473
rect 373 -5481 374 -5473
rect 376 -5481 381 -5473
rect 385 -5481 390 -5473
rect 392 -5481 393 -5473
rect 397 -5481 398 -5473
rect 400 -5481 401 -5473
rect 470 -5481 471 -5473
rect 473 -5481 474 -5473
rect 569 -5481 570 -5473
rect 572 -5481 574 -5473
rect 578 -5481 580 -5473
rect 582 -5481 583 -5473
rect 595 -5481 596 -5473
rect 598 -5481 599 -5473
rect 603 -5481 604 -5473
rect 606 -5481 611 -5473
rect 615 -5481 620 -5473
rect 622 -5481 623 -5473
rect 627 -5481 628 -5473
rect 630 -5481 632 -5473
rect 636 -5481 638 -5473
rect 640 -5481 641 -5473
rect 645 -5481 646 -5473
rect 648 -5481 653 -5473
rect 657 -5481 662 -5473
rect 664 -5481 665 -5473
rect 669 -5481 670 -5473
rect 672 -5481 674 -5473
rect 678 -5481 680 -5473
rect 682 -5481 683 -5473
rect 687 -5481 688 -5473
rect 690 -5481 695 -5473
rect 699 -5481 704 -5473
rect 706 -5481 707 -5473
rect 711 -5481 712 -5473
rect 714 -5481 716 -5473
rect 720 -5481 722 -5473
rect 724 -5481 725 -5473
rect 729 -5481 730 -5473
rect 732 -5481 737 -5473
rect 741 -5481 746 -5473
rect 748 -5481 749 -5473
rect 753 -5481 754 -5473
rect 756 -5481 757 -5473
rect 967 -5481 968 -5473
rect 970 -5481 972 -5473
rect 976 -5481 978 -5473
rect 980 -5481 981 -5473
rect 993 -5481 994 -5473
rect 996 -5481 997 -5473
rect 1001 -5481 1002 -5473
rect 1004 -5481 1009 -5473
rect 1013 -5481 1018 -5473
rect 1020 -5481 1021 -5473
rect 1025 -5481 1026 -5473
rect 1028 -5481 1030 -5473
rect 1034 -5481 1036 -5473
rect 1038 -5481 1039 -5473
rect 1043 -5481 1044 -5473
rect 1046 -5481 1051 -5473
rect 1055 -5481 1060 -5473
rect 1062 -5481 1063 -5473
rect 1067 -5481 1068 -5473
rect 1070 -5481 1072 -5473
rect 1076 -5481 1078 -5473
rect 1080 -5481 1081 -5473
rect 1085 -5481 1086 -5473
rect 1088 -5481 1093 -5473
rect 1097 -5481 1102 -5473
rect 1104 -5481 1105 -5473
rect 1109 -5481 1110 -5473
rect 1112 -5481 1114 -5473
rect 1118 -5481 1120 -5473
rect 1122 -5481 1123 -5473
rect 1127 -5481 1128 -5473
rect 1130 -5481 1135 -5473
rect 1139 -5481 1144 -5473
rect 1146 -5481 1147 -5473
rect 1151 -5481 1152 -5473
rect 1154 -5481 1155 -5473
rect 1214 -5481 1215 -5473
rect 1217 -5481 1218 -5473
rect 1325 -5481 1326 -5473
rect 1328 -5481 1330 -5473
rect 1334 -5481 1336 -5473
rect 1338 -5481 1339 -5473
rect 1351 -5481 1352 -5473
rect 1354 -5481 1355 -5473
rect 1359 -5481 1360 -5473
rect 1362 -5481 1367 -5473
rect 1371 -5481 1376 -5473
rect 1378 -5481 1379 -5473
rect 1383 -5481 1384 -5473
rect 1386 -5481 1388 -5473
rect 1392 -5481 1394 -5473
rect 1396 -5481 1397 -5473
rect 1401 -5481 1402 -5473
rect 1404 -5481 1409 -5473
rect 1413 -5481 1418 -5473
rect 1420 -5481 1421 -5473
rect 1425 -5481 1426 -5473
rect 1428 -5481 1430 -5473
rect 1434 -5481 1436 -5473
rect 1438 -5481 1439 -5473
rect 1443 -5481 1444 -5473
rect 1446 -5481 1451 -5473
rect 1455 -5481 1460 -5473
rect 1462 -5481 1463 -5473
rect 1467 -5481 1468 -5473
rect 1470 -5481 1472 -5473
rect 1476 -5481 1478 -5473
rect 1480 -5481 1481 -5473
rect 1485 -5481 1486 -5473
rect 1488 -5481 1493 -5473
rect 1497 -5481 1502 -5473
rect 1504 -5481 1505 -5473
rect 1509 -5481 1510 -5473
rect 1512 -5481 1513 -5473
rect -1260 -5598 -1259 -5590
rect -1257 -5598 -1255 -5590
rect -1251 -5598 -1249 -5590
rect -1247 -5598 -1246 -5590
rect -1234 -5598 -1233 -5590
rect -1231 -5598 -1230 -5590
rect -1226 -5598 -1225 -5590
rect -1223 -5598 -1218 -5590
rect -1214 -5598 -1209 -5590
rect -1207 -5598 -1206 -5590
rect -1202 -5598 -1201 -5590
rect -1199 -5598 -1197 -5590
rect -1193 -5598 -1191 -5590
rect -1189 -5598 -1188 -5590
rect -1184 -5598 -1183 -5590
rect -1181 -5598 -1176 -5590
rect -1172 -5598 -1167 -5590
rect -1165 -5598 -1164 -5590
rect -1160 -5598 -1159 -5590
rect -1157 -5598 -1155 -5590
rect -1151 -5598 -1149 -5590
rect -1147 -5598 -1146 -5590
rect -1142 -5598 -1141 -5590
rect -1139 -5598 -1134 -5590
rect -1130 -5598 -1125 -5590
rect -1123 -5598 -1122 -5590
rect -1118 -5598 -1117 -5590
rect -1115 -5598 -1113 -5590
rect -1109 -5598 -1107 -5590
rect -1105 -5598 -1104 -5590
rect -1100 -5598 -1099 -5590
rect -1097 -5598 -1092 -5590
rect -1088 -5598 -1083 -5590
rect -1081 -5598 -1080 -5590
rect -1076 -5598 -1075 -5590
rect -1073 -5598 -1072 -5590
rect -931 -5598 -930 -5590
rect -928 -5598 -926 -5590
rect -922 -5598 -920 -5590
rect -918 -5598 -917 -5590
rect -905 -5598 -904 -5590
rect -902 -5598 -901 -5590
rect -897 -5598 -896 -5590
rect -894 -5598 -889 -5590
rect -885 -5598 -880 -5590
rect -878 -5598 -877 -5590
rect -873 -5598 -872 -5590
rect -870 -5598 -868 -5590
rect -864 -5598 -862 -5590
rect -860 -5598 -859 -5590
rect -855 -5598 -854 -5590
rect -852 -5598 -847 -5590
rect -843 -5598 -838 -5590
rect -836 -5598 -835 -5590
rect -831 -5598 -830 -5590
rect -828 -5598 -826 -5590
rect -822 -5598 -820 -5590
rect -818 -5598 -817 -5590
rect -813 -5598 -812 -5590
rect -810 -5598 -805 -5590
rect -801 -5598 -796 -5590
rect -794 -5598 -793 -5590
rect -789 -5598 -788 -5590
rect -786 -5598 -784 -5590
rect -780 -5598 -778 -5590
rect -776 -5598 -775 -5590
rect -771 -5598 -770 -5590
rect -768 -5598 -763 -5590
rect -759 -5598 -754 -5590
rect -752 -5598 -751 -5590
rect -747 -5598 -746 -5590
rect -744 -5598 -743 -5590
rect -573 -5598 -572 -5590
rect -570 -5598 -568 -5590
rect -564 -5598 -562 -5590
rect -560 -5598 -559 -5590
rect -547 -5598 -546 -5590
rect -544 -5598 -543 -5590
rect -539 -5598 -538 -5590
rect -536 -5598 -531 -5590
rect -527 -5598 -522 -5590
rect -520 -5598 -519 -5590
rect -515 -5598 -514 -5590
rect -512 -5598 -510 -5590
rect -506 -5598 -504 -5590
rect -502 -5598 -501 -5590
rect -497 -5598 -496 -5590
rect -494 -5598 -489 -5590
rect -485 -5598 -480 -5590
rect -478 -5598 -477 -5590
rect -473 -5598 -472 -5590
rect -470 -5598 -468 -5590
rect -464 -5598 -462 -5590
rect -460 -5598 -459 -5590
rect -455 -5598 -454 -5590
rect -452 -5598 -447 -5590
rect -443 -5598 -438 -5590
rect -436 -5598 -435 -5590
rect -431 -5598 -430 -5590
rect -428 -5598 -426 -5590
rect -422 -5598 -420 -5590
rect -418 -5598 -417 -5590
rect -413 -5598 -412 -5590
rect -410 -5598 -405 -5590
rect -401 -5598 -396 -5590
rect -394 -5598 -393 -5590
rect -389 -5598 -388 -5590
rect -386 -5598 -385 -5590
rect -215 -5598 -214 -5590
rect -212 -5598 -210 -5590
rect -206 -5598 -204 -5590
rect -202 -5598 -201 -5590
rect -189 -5598 -188 -5590
rect -186 -5598 -185 -5590
rect -181 -5598 -180 -5590
rect -178 -5598 -173 -5590
rect -169 -5598 -164 -5590
rect -162 -5598 -161 -5590
rect -157 -5598 -156 -5590
rect -154 -5598 -152 -5590
rect -148 -5598 -146 -5590
rect -144 -5598 -143 -5590
rect -139 -5598 -138 -5590
rect -136 -5598 -131 -5590
rect -127 -5598 -122 -5590
rect -120 -5598 -119 -5590
rect -115 -5598 -114 -5590
rect -112 -5598 -110 -5590
rect -106 -5598 -104 -5590
rect -102 -5598 -101 -5590
rect -97 -5598 -96 -5590
rect -94 -5598 -89 -5590
rect -85 -5598 -80 -5590
rect -78 -5598 -77 -5590
rect -73 -5598 -72 -5590
rect -70 -5598 -68 -5590
rect -64 -5598 -62 -5590
rect -60 -5598 -59 -5590
rect -55 -5598 -54 -5590
rect -52 -5598 -47 -5590
rect -43 -5598 -38 -5590
rect -36 -5598 -35 -5590
rect -31 -5598 -30 -5590
rect -28 -5598 -27 -5590
rect 213 -5598 214 -5590
rect 216 -5598 218 -5590
rect 222 -5598 224 -5590
rect 226 -5598 227 -5590
rect 239 -5598 240 -5590
rect 242 -5598 243 -5590
rect 247 -5598 248 -5590
rect 250 -5598 255 -5590
rect 259 -5598 264 -5590
rect 266 -5598 267 -5590
rect 271 -5598 272 -5590
rect 274 -5598 276 -5590
rect 280 -5598 282 -5590
rect 284 -5598 285 -5590
rect 289 -5598 290 -5590
rect 292 -5598 297 -5590
rect 301 -5598 306 -5590
rect 308 -5598 309 -5590
rect 313 -5598 314 -5590
rect 316 -5598 318 -5590
rect 322 -5598 324 -5590
rect 326 -5598 327 -5590
rect 331 -5598 332 -5590
rect 334 -5598 339 -5590
rect 343 -5598 348 -5590
rect 350 -5598 351 -5590
rect 355 -5598 356 -5590
rect 358 -5598 360 -5590
rect 364 -5598 366 -5590
rect 368 -5598 369 -5590
rect 373 -5598 374 -5590
rect 376 -5598 381 -5590
rect 385 -5598 390 -5590
rect 392 -5598 393 -5590
rect 397 -5598 398 -5590
rect 400 -5598 401 -5590
rect 569 -5598 570 -5590
rect 572 -5598 574 -5590
rect 578 -5598 580 -5590
rect 582 -5598 583 -5590
rect 595 -5598 596 -5590
rect 598 -5598 599 -5590
rect 603 -5598 604 -5590
rect 606 -5598 611 -5590
rect 615 -5598 620 -5590
rect 622 -5598 623 -5590
rect 627 -5598 628 -5590
rect 630 -5598 632 -5590
rect 636 -5598 638 -5590
rect 640 -5598 641 -5590
rect 645 -5598 646 -5590
rect 648 -5598 653 -5590
rect 657 -5598 662 -5590
rect 664 -5598 665 -5590
rect 669 -5598 670 -5590
rect 672 -5598 674 -5590
rect 678 -5598 680 -5590
rect 682 -5598 683 -5590
rect 687 -5598 688 -5590
rect 690 -5598 695 -5590
rect 699 -5598 704 -5590
rect 706 -5598 707 -5590
rect 711 -5598 712 -5590
rect 714 -5598 716 -5590
rect 720 -5598 722 -5590
rect 724 -5598 725 -5590
rect 729 -5598 730 -5590
rect 732 -5598 737 -5590
rect 741 -5598 746 -5590
rect 748 -5598 749 -5590
rect 753 -5598 754 -5590
rect 756 -5598 757 -5590
rect -1335 -5715 -1334 -5707
rect -1332 -5715 -1331 -5707
rect -1327 -5715 -1326 -5707
rect -1324 -5715 -1322 -5707
rect -1318 -5715 -1316 -5707
rect -1314 -5715 -1313 -5707
rect -931 -5715 -930 -5707
rect -928 -5715 -927 -5707
rect -923 -5715 -922 -5707
rect -920 -5715 -918 -5707
rect -914 -5715 -912 -5707
rect -910 -5715 -909 -5707
rect -573 -5715 -572 -5707
rect -570 -5715 -569 -5707
rect -565 -5715 -564 -5707
rect -562 -5715 -560 -5707
rect -556 -5715 -554 -5707
rect -552 -5715 -551 -5707
rect -215 -5715 -214 -5707
rect -212 -5715 -211 -5707
rect -207 -5715 -206 -5707
rect -204 -5715 -202 -5707
rect -198 -5715 -196 -5707
rect -194 -5715 -193 -5707
rect 213 -5715 214 -5707
rect 216 -5715 217 -5707
rect 221 -5715 222 -5707
rect 224 -5715 226 -5707
rect 230 -5715 232 -5707
rect 234 -5715 235 -5707
rect 569 -5715 570 -5707
rect 572 -5715 573 -5707
rect 577 -5715 578 -5707
rect 580 -5715 582 -5707
rect 586 -5715 588 -5707
rect 590 -5715 591 -5707
rect 967 -5715 968 -5707
rect 970 -5715 971 -5707
rect 975 -5715 976 -5707
rect 978 -5715 980 -5707
rect 984 -5715 986 -5707
rect 988 -5715 989 -5707
rect 1325 -5715 1326 -5707
rect 1328 -5715 1329 -5707
rect 1333 -5715 1334 -5707
rect 1336 -5715 1338 -5707
rect 1342 -5715 1344 -5707
rect 1346 -5715 1347 -5707
rect -1260 -5834 -1259 -5826
rect -1257 -5834 -1255 -5826
rect -1251 -5834 -1249 -5826
rect -1247 -5834 -1246 -5826
rect -1234 -5834 -1233 -5826
rect -1231 -5834 -1223 -5826
rect -1221 -5834 -1220 -5826
rect -1216 -5834 -1215 -5826
rect -1213 -5834 -1205 -5826
rect -1203 -5834 -1198 -5826
rect -1194 -5834 -1189 -5826
rect -1187 -5834 -1186 -5826
rect -1182 -5834 -1181 -5826
rect -1179 -5834 -1177 -5826
rect -1173 -5834 -1171 -5826
rect -1169 -5834 -1168 -5826
rect -931 -5834 -930 -5826
rect -928 -5834 -926 -5826
rect -922 -5834 -920 -5826
rect -918 -5834 -917 -5826
rect -905 -5834 -904 -5826
rect -902 -5834 -900 -5826
rect -896 -5834 -894 -5826
rect -892 -5834 -891 -5826
rect -879 -5834 -878 -5826
rect -876 -5834 -868 -5826
rect -866 -5834 -865 -5826
rect -861 -5834 -860 -5826
rect -858 -5834 -850 -5826
rect -848 -5834 -843 -5826
rect -839 -5834 -834 -5826
rect -832 -5834 -831 -5826
rect -827 -5834 -826 -5826
rect -824 -5834 -822 -5826
rect -818 -5834 -816 -5826
rect -814 -5834 -813 -5826
rect -801 -5834 -800 -5826
rect -798 -5834 -790 -5826
rect -788 -5834 -787 -5826
rect -783 -5834 -782 -5826
rect -780 -5834 -772 -5826
rect -770 -5834 -765 -5826
rect -761 -5834 -756 -5826
rect -754 -5834 -753 -5826
rect -749 -5834 -748 -5826
rect -746 -5834 -741 -5826
rect -737 -5834 -732 -5826
rect -730 -5834 -729 -5826
rect -717 -5834 -716 -5826
rect -714 -5834 -708 -5826
rect -706 -5834 -704 -5826
rect -700 -5834 -698 -5826
rect -696 -5834 -695 -5826
rect -573 -5834 -572 -5826
rect -570 -5834 -568 -5826
rect -564 -5834 -562 -5826
rect -560 -5834 -559 -5826
rect -547 -5834 -546 -5826
rect -544 -5834 -542 -5826
rect -538 -5834 -536 -5826
rect -534 -5834 -533 -5826
rect -521 -5834 -520 -5826
rect -518 -5834 -510 -5826
rect -508 -5834 -507 -5826
rect -503 -5834 -502 -5826
rect -500 -5834 -492 -5826
rect -490 -5834 -485 -5826
rect -481 -5834 -476 -5826
rect -474 -5834 -473 -5826
rect -469 -5834 -468 -5826
rect -466 -5834 -464 -5826
rect -460 -5834 -458 -5826
rect -456 -5834 -455 -5826
rect -443 -5834 -442 -5826
rect -440 -5834 -432 -5826
rect -430 -5834 -429 -5826
rect -425 -5834 -424 -5826
rect -422 -5834 -414 -5826
rect -412 -5834 -407 -5826
rect -403 -5834 -398 -5826
rect -396 -5834 -395 -5826
rect -391 -5834 -390 -5826
rect -388 -5834 -383 -5826
rect -379 -5834 -374 -5826
rect -372 -5834 -371 -5826
rect -359 -5834 -358 -5826
rect -356 -5834 -350 -5826
rect -348 -5834 -346 -5826
rect -342 -5834 -340 -5826
rect -338 -5834 -337 -5826
rect -215 -5834 -214 -5826
rect -212 -5834 -210 -5826
rect -206 -5834 -204 -5826
rect -202 -5834 -201 -5826
rect -189 -5834 -188 -5826
rect -186 -5834 -184 -5826
rect -180 -5834 -178 -5826
rect -176 -5834 -175 -5826
rect -163 -5834 -162 -5826
rect -160 -5834 -152 -5826
rect -150 -5834 -149 -5826
rect -145 -5834 -144 -5826
rect -142 -5834 -134 -5826
rect -132 -5834 -127 -5826
rect -123 -5834 -118 -5826
rect -116 -5834 -115 -5826
rect -111 -5834 -110 -5826
rect -108 -5834 -106 -5826
rect -102 -5834 -100 -5826
rect -98 -5834 -97 -5826
rect -85 -5834 -84 -5826
rect -82 -5834 -74 -5826
rect -72 -5834 -71 -5826
rect -67 -5834 -66 -5826
rect -64 -5834 -56 -5826
rect -54 -5834 -49 -5826
rect -45 -5834 -40 -5826
rect -38 -5834 -37 -5826
rect -33 -5834 -32 -5826
rect -30 -5834 -25 -5826
rect -21 -5834 -16 -5826
rect -14 -5834 -13 -5826
rect -1 -5834 0 -5826
rect 2 -5834 8 -5826
rect 10 -5834 12 -5826
rect 16 -5834 18 -5826
rect 20 -5834 21 -5826
rect 213 -5834 214 -5826
rect 216 -5834 218 -5826
rect 222 -5834 224 -5826
rect 226 -5834 227 -5826
rect 239 -5834 240 -5826
rect 242 -5834 244 -5826
rect 248 -5834 250 -5826
rect 252 -5834 253 -5826
rect 265 -5834 266 -5826
rect 268 -5834 276 -5826
rect 278 -5834 279 -5826
rect 283 -5834 284 -5826
rect 286 -5834 294 -5826
rect 296 -5834 301 -5826
rect 305 -5834 310 -5826
rect 312 -5834 313 -5826
rect 317 -5834 318 -5826
rect 320 -5834 322 -5826
rect 326 -5834 328 -5826
rect 330 -5834 331 -5826
rect 343 -5834 344 -5826
rect 346 -5834 354 -5826
rect 356 -5834 357 -5826
rect 361 -5834 362 -5826
rect 364 -5834 372 -5826
rect 374 -5834 379 -5826
rect 383 -5834 388 -5826
rect 390 -5834 391 -5826
rect 395 -5834 396 -5826
rect 398 -5834 403 -5826
rect 407 -5834 412 -5826
rect 414 -5834 415 -5826
rect 427 -5834 428 -5826
rect 430 -5834 436 -5826
rect 438 -5834 440 -5826
rect 444 -5834 446 -5826
rect 448 -5834 449 -5826
rect 569 -5834 570 -5826
rect 572 -5834 574 -5826
rect 578 -5834 580 -5826
rect 582 -5834 583 -5826
rect 595 -5834 596 -5826
rect 598 -5834 600 -5826
rect 604 -5834 606 -5826
rect 608 -5834 609 -5826
rect 621 -5834 622 -5826
rect 624 -5834 632 -5826
rect 634 -5834 635 -5826
rect 639 -5834 640 -5826
rect 642 -5834 650 -5826
rect 652 -5834 657 -5826
rect 661 -5834 666 -5826
rect 668 -5834 669 -5826
rect 673 -5834 674 -5826
rect 676 -5834 678 -5826
rect 682 -5834 684 -5826
rect 686 -5834 687 -5826
rect 699 -5834 700 -5826
rect 702 -5834 710 -5826
rect 712 -5834 713 -5826
rect 717 -5834 718 -5826
rect 720 -5834 728 -5826
rect 730 -5834 735 -5826
rect 739 -5834 744 -5826
rect 746 -5834 747 -5826
rect 751 -5834 752 -5826
rect 754 -5834 759 -5826
rect 763 -5834 768 -5826
rect 770 -5834 771 -5826
rect 783 -5834 784 -5826
rect 786 -5834 792 -5826
rect 794 -5834 796 -5826
rect 800 -5834 802 -5826
rect 804 -5834 805 -5826
rect 967 -5834 968 -5826
rect 970 -5834 972 -5826
rect 976 -5834 978 -5826
rect 980 -5834 981 -5826
rect 993 -5834 994 -5826
rect 996 -5834 998 -5826
rect 1002 -5834 1004 -5826
rect 1006 -5834 1007 -5826
rect 1019 -5834 1020 -5826
rect 1022 -5834 1030 -5826
rect 1032 -5834 1033 -5826
rect 1037 -5834 1038 -5826
rect 1040 -5834 1048 -5826
rect 1050 -5834 1055 -5826
rect 1059 -5834 1064 -5826
rect 1066 -5834 1067 -5826
rect 1071 -5834 1072 -5826
rect 1074 -5834 1076 -5826
rect 1080 -5834 1082 -5826
rect 1084 -5834 1085 -5826
rect 1097 -5834 1098 -5826
rect 1100 -5834 1108 -5826
rect 1110 -5834 1111 -5826
rect 1115 -5834 1116 -5826
rect 1118 -5834 1126 -5826
rect 1128 -5834 1133 -5826
rect 1137 -5834 1142 -5826
rect 1144 -5834 1145 -5826
rect 1149 -5834 1150 -5826
rect 1152 -5834 1157 -5826
rect 1161 -5834 1166 -5826
rect 1168 -5834 1169 -5826
rect 1181 -5834 1182 -5826
rect 1184 -5834 1190 -5826
rect 1192 -5834 1194 -5826
rect 1198 -5834 1200 -5826
rect 1202 -5834 1203 -5826
rect 1325 -5834 1326 -5826
rect 1328 -5834 1330 -5826
rect 1334 -5834 1336 -5826
rect 1338 -5834 1339 -5826
rect 1351 -5834 1352 -5826
rect 1354 -5834 1356 -5826
rect 1360 -5834 1362 -5826
rect 1364 -5834 1365 -5826
rect 1377 -5834 1378 -5826
rect 1380 -5834 1388 -5826
rect 1390 -5834 1391 -5826
rect 1395 -5834 1396 -5826
rect 1398 -5834 1406 -5826
rect 1408 -5834 1413 -5826
rect 1417 -5834 1422 -5826
rect 1424 -5834 1425 -5826
rect 1429 -5834 1430 -5826
rect 1432 -5834 1434 -5826
rect 1438 -5834 1440 -5826
rect 1442 -5834 1443 -5826
rect 1455 -5834 1456 -5826
rect 1458 -5834 1466 -5826
rect 1468 -5834 1469 -5826
rect 1473 -5834 1474 -5826
rect 1476 -5834 1484 -5826
rect 1486 -5834 1491 -5826
rect 1495 -5834 1500 -5826
rect 1502 -5834 1503 -5826
rect 1507 -5834 1508 -5826
rect 1510 -5834 1515 -5826
rect 1519 -5834 1524 -5826
rect 1526 -5834 1527 -5826
rect 1539 -5834 1540 -5826
rect 1542 -5834 1548 -5826
rect 1550 -5834 1552 -5826
rect 1556 -5834 1558 -5826
rect 1560 -5834 1561 -5826
rect -1260 -5957 -1259 -5949
rect -1257 -5957 -1255 -5949
rect -1251 -5957 -1249 -5949
rect -1247 -5957 -1246 -5949
rect -1234 -5957 -1233 -5949
rect -1231 -5957 -1230 -5949
rect -1226 -5957 -1225 -5949
rect -1223 -5957 -1218 -5949
rect -1214 -5957 -1209 -5949
rect -1207 -5957 -1206 -5949
rect -1202 -5957 -1201 -5949
rect -1199 -5957 -1197 -5949
rect -1193 -5957 -1191 -5949
rect -1189 -5957 -1188 -5949
rect -1184 -5957 -1183 -5949
rect -1181 -5957 -1176 -5949
rect -1172 -5957 -1167 -5949
rect -1165 -5957 -1164 -5949
rect -1160 -5957 -1159 -5949
rect -1157 -5957 -1155 -5949
rect -1151 -5957 -1149 -5949
rect -1147 -5957 -1146 -5949
rect -1142 -5957 -1141 -5949
rect -1139 -5957 -1134 -5949
rect -1130 -5957 -1125 -5949
rect -1123 -5957 -1122 -5949
rect -1118 -5957 -1117 -5949
rect -1115 -5957 -1113 -5949
rect -1109 -5957 -1107 -5949
rect -1105 -5957 -1104 -5949
rect -1100 -5957 -1099 -5949
rect -1097 -5957 -1092 -5949
rect -1088 -5957 -1083 -5949
rect -1081 -5957 -1080 -5949
rect -1076 -5957 -1075 -5949
rect -1073 -5957 -1072 -5949
rect -931 -5957 -930 -5949
rect -928 -5957 -926 -5949
rect -922 -5957 -920 -5949
rect -918 -5957 -917 -5949
rect -905 -5957 -904 -5949
rect -902 -5957 -901 -5949
rect -897 -5957 -896 -5949
rect -894 -5957 -889 -5949
rect -885 -5957 -880 -5949
rect -878 -5957 -877 -5949
rect -873 -5957 -872 -5949
rect -870 -5957 -868 -5949
rect -864 -5957 -862 -5949
rect -860 -5957 -859 -5949
rect -855 -5957 -854 -5949
rect -852 -5957 -847 -5949
rect -843 -5957 -838 -5949
rect -836 -5957 -835 -5949
rect -831 -5957 -830 -5949
rect -828 -5957 -826 -5949
rect -822 -5957 -820 -5949
rect -818 -5957 -817 -5949
rect -813 -5957 -812 -5949
rect -810 -5957 -805 -5949
rect -801 -5957 -796 -5949
rect -794 -5957 -793 -5949
rect -789 -5957 -788 -5949
rect -786 -5957 -784 -5949
rect -780 -5957 -778 -5949
rect -776 -5957 -775 -5949
rect -771 -5957 -770 -5949
rect -768 -5957 -763 -5949
rect -759 -5957 -754 -5949
rect -752 -5957 -751 -5949
rect -747 -5957 -746 -5949
rect -744 -5957 -743 -5949
rect -573 -5957 -572 -5949
rect -570 -5957 -568 -5949
rect -564 -5957 -562 -5949
rect -560 -5957 -559 -5949
rect -547 -5957 -546 -5949
rect -544 -5957 -543 -5949
rect -539 -5957 -538 -5949
rect -536 -5957 -531 -5949
rect -527 -5957 -522 -5949
rect -520 -5957 -519 -5949
rect -515 -5957 -514 -5949
rect -512 -5957 -510 -5949
rect -506 -5957 -504 -5949
rect -502 -5957 -501 -5949
rect -497 -5957 -496 -5949
rect -494 -5957 -489 -5949
rect -485 -5957 -480 -5949
rect -478 -5957 -477 -5949
rect -473 -5957 -472 -5949
rect -470 -5957 -468 -5949
rect -464 -5957 -462 -5949
rect -460 -5957 -459 -5949
rect -455 -5957 -454 -5949
rect -452 -5957 -447 -5949
rect -443 -5957 -438 -5949
rect -436 -5957 -435 -5949
rect -431 -5957 -430 -5949
rect -428 -5957 -426 -5949
rect -422 -5957 -420 -5949
rect -418 -5957 -417 -5949
rect -413 -5957 -412 -5949
rect -410 -5957 -405 -5949
rect -401 -5957 -396 -5949
rect -394 -5957 -393 -5949
rect -389 -5957 -388 -5949
rect -386 -5957 -385 -5949
rect -215 -5957 -214 -5949
rect -212 -5957 -210 -5949
rect -206 -5957 -204 -5949
rect -202 -5957 -201 -5949
rect -189 -5957 -188 -5949
rect -186 -5957 -185 -5949
rect -181 -5957 -180 -5949
rect -178 -5957 -173 -5949
rect -169 -5957 -164 -5949
rect -162 -5957 -161 -5949
rect -157 -5957 -156 -5949
rect -154 -5957 -152 -5949
rect -148 -5957 -146 -5949
rect -144 -5957 -143 -5949
rect -139 -5957 -138 -5949
rect -136 -5957 -131 -5949
rect -127 -5957 -122 -5949
rect -120 -5957 -119 -5949
rect -115 -5957 -114 -5949
rect -112 -5957 -110 -5949
rect -106 -5957 -104 -5949
rect -102 -5957 -101 -5949
rect -97 -5957 -96 -5949
rect -94 -5957 -89 -5949
rect -85 -5957 -80 -5949
rect -78 -5957 -77 -5949
rect -73 -5957 -72 -5949
rect -70 -5957 -68 -5949
rect -64 -5957 -62 -5949
rect -60 -5957 -59 -5949
rect -55 -5957 -54 -5949
rect -52 -5957 -47 -5949
rect -43 -5957 -38 -5949
rect -36 -5957 -35 -5949
rect -31 -5957 -30 -5949
rect -28 -5957 -27 -5949
rect 213 -5957 214 -5949
rect 216 -5957 218 -5949
rect 222 -5957 224 -5949
rect 226 -5957 227 -5949
rect 239 -5957 240 -5949
rect 242 -5957 243 -5949
rect 247 -5957 248 -5949
rect 250 -5957 255 -5949
rect 259 -5957 264 -5949
rect 266 -5957 267 -5949
rect 271 -5957 272 -5949
rect 274 -5957 276 -5949
rect 280 -5957 282 -5949
rect 284 -5957 285 -5949
rect 289 -5957 290 -5949
rect 292 -5957 297 -5949
rect 301 -5957 306 -5949
rect 308 -5957 309 -5949
rect 313 -5957 314 -5949
rect 316 -5957 318 -5949
rect 322 -5957 324 -5949
rect 326 -5957 327 -5949
rect 331 -5957 332 -5949
rect 334 -5957 339 -5949
rect 343 -5957 348 -5949
rect 350 -5957 351 -5949
rect 355 -5957 356 -5949
rect 358 -5957 360 -5949
rect 364 -5957 366 -5949
rect 368 -5957 369 -5949
rect 373 -5957 374 -5949
rect 376 -5957 381 -5949
rect 385 -5957 390 -5949
rect 392 -5957 393 -5949
rect 397 -5957 398 -5949
rect 400 -5957 401 -5949
rect 569 -5957 570 -5949
rect 572 -5957 574 -5949
rect 578 -5957 580 -5949
rect 582 -5957 583 -5949
rect 595 -5957 596 -5949
rect 598 -5957 599 -5949
rect 603 -5957 604 -5949
rect 606 -5957 611 -5949
rect 615 -5957 620 -5949
rect 622 -5957 623 -5949
rect 627 -5957 628 -5949
rect 630 -5957 632 -5949
rect 636 -5957 638 -5949
rect 640 -5957 641 -5949
rect 645 -5957 646 -5949
rect 648 -5957 653 -5949
rect 657 -5957 662 -5949
rect 664 -5957 665 -5949
rect 669 -5957 670 -5949
rect 672 -5957 674 -5949
rect 678 -5957 680 -5949
rect 682 -5957 683 -5949
rect 687 -5957 688 -5949
rect 690 -5957 695 -5949
rect 699 -5957 704 -5949
rect 706 -5957 707 -5949
rect 711 -5957 712 -5949
rect 714 -5957 716 -5949
rect 720 -5957 722 -5949
rect 724 -5957 725 -5949
rect 729 -5957 730 -5949
rect 732 -5957 737 -5949
rect 741 -5957 746 -5949
rect 748 -5957 749 -5949
rect 753 -5957 754 -5949
rect 756 -5957 757 -5949
rect 967 -5957 968 -5949
rect 970 -5957 972 -5949
rect 976 -5957 978 -5949
rect 980 -5957 981 -5949
rect 993 -5957 994 -5949
rect 996 -5957 997 -5949
rect 1001 -5957 1002 -5949
rect 1004 -5957 1009 -5949
rect 1013 -5957 1018 -5949
rect 1020 -5957 1021 -5949
rect 1025 -5957 1026 -5949
rect 1028 -5957 1030 -5949
rect 1034 -5957 1036 -5949
rect 1038 -5957 1039 -5949
rect 1043 -5957 1044 -5949
rect 1046 -5957 1051 -5949
rect 1055 -5957 1060 -5949
rect 1062 -5957 1063 -5949
rect 1067 -5957 1068 -5949
rect 1070 -5957 1072 -5949
rect 1076 -5957 1078 -5949
rect 1080 -5957 1081 -5949
rect 1085 -5957 1086 -5949
rect 1088 -5957 1093 -5949
rect 1097 -5957 1102 -5949
rect 1104 -5957 1105 -5949
rect 1109 -5957 1110 -5949
rect 1112 -5957 1114 -5949
rect 1118 -5957 1120 -5949
rect 1122 -5957 1123 -5949
rect 1127 -5957 1128 -5949
rect 1130 -5957 1135 -5949
rect 1139 -5957 1144 -5949
rect 1146 -5957 1147 -5949
rect 1151 -5957 1152 -5949
rect 1154 -5957 1155 -5949
rect 1325 -5957 1326 -5949
rect 1328 -5957 1330 -5949
rect 1334 -5957 1336 -5949
rect 1338 -5957 1339 -5949
rect 1351 -5957 1352 -5949
rect 1354 -5957 1355 -5949
rect 1359 -5957 1360 -5949
rect 1362 -5957 1367 -5949
rect 1371 -5957 1376 -5949
rect 1378 -5957 1379 -5949
rect 1383 -5957 1384 -5949
rect 1386 -5957 1388 -5949
rect 1392 -5957 1394 -5949
rect 1396 -5957 1397 -5949
rect 1401 -5957 1402 -5949
rect 1404 -5957 1409 -5949
rect 1413 -5957 1418 -5949
rect 1420 -5957 1421 -5949
rect 1425 -5957 1426 -5949
rect 1428 -5957 1430 -5949
rect 1434 -5957 1436 -5949
rect 1438 -5957 1439 -5949
rect 1443 -5957 1444 -5949
rect 1446 -5957 1451 -5949
rect 1455 -5957 1460 -5949
rect 1462 -5957 1463 -5949
rect 1467 -5957 1468 -5949
rect 1470 -5957 1472 -5949
rect 1476 -5957 1478 -5949
rect 1480 -5957 1481 -5949
rect 1485 -5957 1486 -5949
rect 1488 -5957 1493 -5949
rect 1497 -5957 1502 -5949
rect 1504 -5957 1505 -5949
rect 1509 -5957 1510 -5949
rect 1512 -5957 1513 -5949
rect 1325 -6075 1326 -6067
rect 1328 -6075 1330 -6067
rect 1334 -6075 1336 -6067
rect 1338 -6075 1339 -6067
rect 1351 -6075 1352 -6067
rect 1354 -6075 1355 -6067
rect 1359 -6075 1360 -6067
rect 1362 -6075 1367 -6067
rect 1371 -6075 1376 -6067
rect 1378 -6075 1379 -6067
rect 1383 -6075 1384 -6067
rect 1386 -6075 1388 -6067
rect 1392 -6075 1394 -6067
rect 1396 -6075 1397 -6067
rect 1401 -6075 1402 -6067
rect 1404 -6075 1409 -6067
rect 1413 -6075 1418 -6067
rect 1420 -6075 1421 -6067
rect 1425 -6075 1426 -6067
rect 1428 -6075 1430 -6067
rect 1434 -6075 1436 -6067
rect 1438 -6075 1439 -6067
rect 1443 -6075 1444 -6067
rect 1446 -6075 1451 -6067
rect 1455 -6075 1460 -6067
rect 1462 -6075 1463 -6067
rect 1467 -6075 1468 -6067
rect 1470 -6075 1472 -6067
rect 1476 -6075 1478 -6067
rect 1480 -6075 1481 -6067
rect 1485 -6075 1486 -6067
rect 1488 -6075 1493 -6067
rect 1497 -6075 1502 -6067
rect 1504 -6075 1505 -6067
rect 1509 -6075 1510 -6067
rect 1512 -6075 1513 -6067
<< metal1 >>
rect -1349 -1062 -1345 -998
rect -1337 -1038 -1333 -1034
rect -1320 -1038 -1316 -1034
rect -1329 -1049 -1325 -1046
rect -1329 -1053 -1314 -1049
rect -1349 -1066 -1336 -1062
rect -1349 -1292 -1345 -1066
rect -1318 -1092 -1314 -1053
rect -1318 -1107 -1314 -1096
rect -1337 -1111 -1314 -1107
rect -1337 -1114 -1333 -1111
rect -1311 -1114 -1307 -1046
rect -942 -1062 -938 -998
rect -936 -1038 -932 -1034
rect -919 -1038 -915 -1034
rect -928 -1049 -924 -1046
rect -928 -1053 -913 -1049
rect -942 -1066 -935 -1062
rect -1320 -1122 -1316 -1118
rect -1311 -1200 -1307 -1118
rect -1339 -1268 -1335 -1264
rect -1322 -1268 -1318 -1264
rect -1331 -1279 -1327 -1276
rect -1331 -1283 -1316 -1279
rect -1349 -1296 -1338 -1292
rect -1349 -1795 -1345 -1296
rect -1320 -1322 -1316 -1283
rect -1320 -1337 -1316 -1326
rect -1339 -1341 -1316 -1337
rect -1339 -1344 -1335 -1341
rect -1313 -1344 -1309 -1276
rect -1322 -1352 -1318 -1348
rect -1313 -1437 -1309 -1348
rect -1266 -1430 -1262 -1090
rect -1251 -1152 -1247 -1148
rect -1234 -1152 -1230 -1148
rect -1214 -1152 -1210 -1148
rect -1193 -1152 -1189 -1148
rect -1172 -1152 -1168 -1148
rect -1151 -1152 -1147 -1148
rect -1130 -1152 -1126 -1148
rect -1109 -1152 -1105 -1148
rect -1088 -1152 -1084 -1148
rect -1068 -1152 -1064 -1148
rect -1260 -1207 -1256 -1160
rect -1260 -1228 -1256 -1211
rect -1242 -1221 -1238 -1160
rect -1226 -1221 -1222 -1160
rect -1202 -1200 -1198 -1160
rect -1202 -1221 -1198 -1204
rect -1184 -1221 -1180 -1160
rect -1160 -1207 -1156 -1160
rect -1160 -1221 -1156 -1211
rect -1142 -1200 -1138 -1160
rect -1142 -1221 -1138 -1204
rect -1118 -1214 -1114 -1160
rect -1100 -1192 -1096 -1160
rect -1100 -1200 -1096 -1196
rect -1118 -1221 -1114 -1218
rect -1242 -1225 -1233 -1221
rect -1226 -1225 -1218 -1221
rect -1242 -1228 -1238 -1225
rect -1218 -1228 -1214 -1225
rect -1210 -1225 -1198 -1221
rect -1184 -1225 -1176 -1221
rect -1210 -1228 -1206 -1225
rect -1176 -1228 -1172 -1225
rect -1168 -1225 -1156 -1221
rect -1142 -1225 -1130 -1221
rect -1168 -1228 -1164 -1225
rect -1134 -1228 -1130 -1225
rect -1126 -1225 -1114 -1221
rect -1100 -1221 -1096 -1204
rect -1076 -1207 -1072 -1160
rect -1076 -1221 -1072 -1211
rect -1100 -1225 -1088 -1221
rect -1126 -1228 -1122 -1225
rect -1092 -1228 -1088 -1225
rect -1084 -1225 -1072 -1221
rect -1084 -1228 -1080 -1225
rect -1251 -1236 -1247 -1232
rect -1234 -1236 -1230 -1232
rect -1193 -1236 -1189 -1232
rect -1151 -1236 -1147 -1232
rect -1109 -1236 -1105 -1232
rect -1068 -1236 -1064 -1232
rect -1251 -1382 -1247 -1378
rect -1234 -1382 -1230 -1378
rect -1194 -1382 -1190 -1378
rect -1173 -1382 -1169 -1378
rect -1260 -1423 -1256 -1390
rect -1260 -1458 -1256 -1427
rect -1242 -1417 -1238 -1390
rect -1242 -1421 -1233 -1417
rect -1242 -1458 -1238 -1421
rect -1216 -1444 -1212 -1390
rect -1216 -1451 -1212 -1448
rect -1182 -1451 -1178 -1390
rect -1164 -1422 -1160 -1390
rect -1234 -1458 -1230 -1455
rect -1225 -1455 -1212 -1451
rect -1225 -1458 -1221 -1455
rect -1198 -1458 -1194 -1455
rect -1190 -1455 -1171 -1451
rect -1190 -1458 -1186 -1455
rect -1164 -1458 -1160 -1426
rect -954 -1429 -950 -1317
rect -948 -1414 -944 -1082
rect -942 -1292 -938 -1066
rect -917 -1094 -913 -1053
rect -917 -1107 -913 -1098
rect -936 -1111 -913 -1107
rect -910 -1086 -906 -1046
rect -583 -1062 -579 -999
rect -577 -1038 -573 -1034
rect -560 -1038 -556 -1034
rect -569 -1049 -565 -1046
rect -569 -1053 -554 -1049
rect -583 -1066 -576 -1062
rect -936 -1114 -932 -1111
rect -910 -1114 -906 -1090
rect -919 -1122 -915 -1118
rect -926 -1152 -922 -1148
rect -909 -1152 -905 -1148
rect -889 -1152 -885 -1148
rect -868 -1152 -864 -1148
rect -847 -1152 -843 -1148
rect -826 -1152 -822 -1148
rect -805 -1152 -801 -1148
rect -784 -1152 -780 -1148
rect -763 -1152 -759 -1148
rect -743 -1152 -739 -1148
rect -935 -1207 -931 -1160
rect -935 -1228 -931 -1211
rect -917 -1221 -913 -1160
rect -901 -1221 -897 -1160
rect -877 -1200 -873 -1160
rect -877 -1221 -873 -1204
rect -859 -1221 -855 -1160
rect -835 -1207 -831 -1160
rect -835 -1221 -831 -1211
rect -817 -1200 -813 -1160
rect -817 -1221 -813 -1204
rect -793 -1214 -789 -1160
rect -775 -1192 -771 -1160
rect -775 -1200 -771 -1196
rect -793 -1221 -789 -1218
rect -917 -1225 -908 -1221
rect -901 -1225 -893 -1221
rect -917 -1228 -913 -1225
rect -893 -1228 -889 -1225
rect -885 -1225 -873 -1221
rect -859 -1225 -851 -1221
rect -885 -1228 -881 -1225
rect -851 -1228 -847 -1225
rect -843 -1225 -831 -1221
rect -817 -1225 -805 -1221
rect -843 -1228 -839 -1225
rect -809 -1228 -805 -1225
rect -801 -1225 -789 -1221
rect -775 -1221 -771 -1204
rect -751 -1207 -747 -1160
rect -751 -1221 -747 -1211
rect -775 -1225 -763 -1221
rect -801 -1228 -797 -1225
rect -767 -1228 -763 -1225
rect -759 -1225 -747 -1221
rect -759 -1228 -755 -1225
rect -926 -1236 -922 -1232
rect -909 -1236 -905 -1232
rect -868 -1236 -864 -1232
rect -826 -1236 -822 -1232
rect -784 -1236 -780 -1232
rect -743 -1236 -739 -1232
rect -935 -1268 -931 -1264
rect -918 -1268 -914 -1264
rect -927 -1279 -923 -1276
rect -927 -1283 -912 -1279
rect -942 -1296 -934 -1292
rect -1251 -1466 -1247 -1462
rect -1207 -1466 -1203 -1462
rect -1173 -1466 -1169 -1462
rect -1272 -1674 -1268 -1477
rect -1158 -1480 -1154 -1448
rect -1266 -1553 -1262 -1484
rect -1251 -1505 -1247 -1501
rect -1234 -1505 -1230 -1501
rect -1214 -1505 -1210 -1501
rect -1193 -1505 -1189 -1501
rect -1172 -1505 -1168 -1501
rect -1151 -1505 -1147 -1501
rect -1130 -1505 -1126 -1501
rect -1109 -1505 -1105 -1501
rect -1088 -1505 -1084 -1501
rect -1068 -1505 -1064 -1501
rect -1260 -1560 -1256 -1513
rect -1260 -1581 -1256 -1564
rect -1242 -1574 -1238 -1513
rect -1226 -1574 -1222 -1513
rect -1202 -1553 -1198 -1513
rect -1202 -1574 -1198 -1557
rect -1184 -1574 -1180 -1513
rect -1160 -1560 -1156 -1513
rect -1160 -1574 -1156 -1564
rect -1142 -1553 -1138 -1513
rect -1142 -1574 -1138 -1557
rect -1118 -1567 -1114 -1513
rect -1100 -1545 -1096 -1513
rect -1100 -1553 -1096 -1549
rect -1118 -1574 -1114 -1571
rect -1242 -1578 -1233 -1574
rect -1226 -1578 -1218 -1574
rect -1242 -1581 -1238 -1578
rect -1218 -1581 -1214 -1578
rect -1210 -1578 -1198 -1574
rect -1184 -1578 -1176 -1574
rect -1210 -1581 -1206 -1578
rect -1176 -1581 -1172 -1578
rect -1168 -1578 -1156 -1574
rect -1142 -1578 -1130 -1574
rect -1168 -1581 -1164 -1578
rect -1134 -1581 -1130 -1578
rect -1126 -1578 -1114 -1574
rect -1100 -1574 -1096 -1557
rect -1076 -1560 -1072 -1513
rect -1076 -1574 -1072 -1564
rect -1100 -1578 -1088 -1574
rect -1126 -1581 -1122 -1578
rect -1092 -1581 -1088 -1578
rect -1084 -1578 -1072 -1574
rect -1084 -1581 -1080 -1578
rect -1251 -1589 -1247 -1585
rect -1234 -1589 -1230 -1585
rect -1193 -1589 -1189 -1585
rect -1151 -1589 -1147 -1585
rect -1109 -1589 -1105 -1585
rect -1068 -1589 -1064 -1585
rect -1251 -1626 -1247 -1622
rect -1234 -1626 -1230 -1622
rect -1214 -1626 -1210 -1622
rect -1193 -1626 -1189 -1622
rect -1172 -1626 -1168 -1622
rect -1151 -1626 -1147 -1622
rect -1130 -1626 -1126 -1622
rect -1109 -1626 -1105 -1622
rect -1088 -1626 -1084 -1622
rect -1068 -1626 -1064 -1622
rect -1260 -1681 -1256 -1634
rect -1260 -1702 -1256 -1685
rect -1242 -1695 -1238 -1634
rect -1226 -1695 -1222 -1634
rect -1202 -1674 -1198 -1634
rect -1202 -1695 -1198 -1678
rect -1184 -1695 -1180 -1634
rect -1160 -1681 -1156 -1634
rect -1160 -1695 -1156 -1685
rect -1142 -1674 -1138 -1634
rect -1142 -1695 -1138 -1678
rect -1118 -1688 -1114 -1634
rect -1100 -1666 -1096 -1634
rect -1100 -1674 -1096 -1670
rect -1118 -1695 -1114 -1692
rect -1242 -1699 -1233 -1695
rect -1226 -1699 -1218 -1695
rect -1242 -1702 -1238 -1699
rect -1218 -1702 -1214 -1699
rect -1210 -1699 -1198 -1695
rect -1184 -1699 -1176 -1695
rect -1210 -1702 -1206 -1699
rect -1176 -1702 -1172 -1699
rect -1168 -1699 -1156 -1695
rect -1142 -1699 -1130 -1695
rect -1168 -1702 -1164 -1699
rect -1134 -1702 -1130 -1699
rect -1126 -1699 -1114 -1695
rect -1100 -1695 -1096 -1678
rect -1076 -1681 -1072 -1634
rect -1076 -1695 -1072 -1685
rect -1100 -1699 -1088 -1695
rect -1126 -1702 -1122 -1699
rect -1092 -1702 -1088 -1699
rect -1084 -1699 -1072 -1695
rect -1084 -1702 -1080 -1699
rect -1251 -1710 -1247 -1706
rect -1234 -1710 -1230 -1706
rect -1193 -1710 -1189 -1706
rect -1151 -1710 -1147 -1706
rect -1109 -1710 -1105 -1706
rect -1068 -1710 -1064 -1706
rect -1062 -1717 -1058 -1670
rect -948 -1674 -944 -1484
rect -1339 -1974 -1335 -1970
rect -1322 -1974 -1318 -1970
rect -1331 -1985 -1327 -1982
rect -1331 -1989 -1316 -1985
rect -1349 -2002 -1338 -1998
rect -1349 -2547 -1345 -2002
rect -1320 -2028 -1316 -1989
rect -1320 -2043 -1316 -2032
rect -1339 -2047 -1316 -2043
rect -1339 -2050 -1335 -2047
rect -1313 -2050 -1309 -1982
rect -1322 -2058 -1318 -2054
rect -1313 -2148 -1309 -2054
rect -1266 -2141 -1262 -1721
rect -1251 -1747 -1247 -1743
rect -1234 -1747 -1230 -1743
rect -1214 -1747 -1210 -1743
rect -1193 -1747 -1189 -1743
rect -1172 -1747 -1168 -1743
rect -1151 -1747 -1147 -1743
rect -1130 -1747 -1126 -1743
rect -1109 -1747 -1105 -1743
rect -1088 -1747 -1084 -1743
rect -1068 -1747 -1064 -1743
rect -1029 -1747 -1025 -1743
rect -1260 -1802 -1256 -1755
rect -1260 -1823 -1256 -1806
rect -1242 -1816 -1238 -1755
rect -1226 -1816 -1222 -1755
rect -1202 -1795 -1198 -1755
rect -1202 -1816 -1198 -1799
rect -1184 -1816 -1180 -1755
rect -1160 -1802 -1156 -1755
rect -1160 -1816 -1156 -1806
rect -1142 -1795 -1138 -1755
rect -1142 -1816 -1138 -1799
rect -1118 -1809 -1114 -1755
rect -1100 -1787 -1096 -1755
rect -1100 -1795 -1096 -1791
rect -1118 -1816 -1114 -1813
rect -1242 -1820 -1233 -1816
rect -1226 -1820 -1218 -1816
rect -1242 -1823 -1238 -1820
rect -1218 -1823 -1214 -1820
rect -1210 -1820 -1198 -1816
rect -1184 -1820 -1176 -1816
rect -1210 -1823 -1206 -1820
rect -1176 -1823 -1172 -1820
rect -1168 -1820 -1156 -1816
rect -1142 -1820 -1130 -1816
rect -1168 -1823 -1164 -1820
rect -1134 -1823 -1130 -1820
rect -1126 -1820 -1114 -1816
rect -1100 -1816 -1096 -1799
rect -1076 -1802 -1072 -1755
rect -1076 -1816 -1072 -1806
rect -1100 -1820 -1088 -1816
rect -1126 -1823 -1122 -1820
rect -1092 -1823 -1088 -1820
rect -1084 -1820 -1072 -1816
rect -1084 -1823 -1080 -1820
rect -1251 -1831 -1247 -1827
rect -1234 -1831 -1230 -1827
rect -1193 -1831 -1189 -1827
rect -1151 -1831 -1147 -1827
rect -1109 -1831 -1105 -1827
rect -1068 -1831 -1064 -1827
rect -1251 -1862 -1247 -1858
rect -1234 -1862 -1230 -1858
rect -1214 -1862 -1210 -1858
rect -1193 -1862 -1189 -1858
rect -1172 -1862 -1168 -1858
rect -1151 -1862 -1147 -1858
rect -1130 -1862 -1126 -1858
rect -1109 -1862 -1105 -1858
rect -1088 -1862 -1084 -1858
rect -1068 -1862 -1064 -1858
rect -1260 -1917 -1256 -1870
rect -1260 -1938 -1256 -1921
rect -1242 -1931 -1238 -1870
rect -1226 -1931 -1222 -1870
rect -1202 -1910 -1198 -1870
rect -1202 -1931 -1198 -1914
rect -1184 -1931 -1180 -1870
rect -1160 -1917 -1156 -1870
rect -1160 -1931 -1156 -1921
rect -1142 -1910 -1138 -1870
rect -1142 -1931 -1138 -1914
rect -1118 -1924 -1114 -1870
rect -1100 -1894 -1096 -1870
rect -1100 -1910 -1096 -1898
rect -1118 -1931 -1114 -1928
rect -1242 -1935 -1233 -1931
rect -1226 -1935 -1218 -1931
rect -1242 -1938 -1238 -1935
rect -1218 -1938 -1214 -1935
rect -1210 -1935 -1198 -1931
rect -1184 -1935 -1176 -1931
rect -1210 -1938 -1206 -1935
rect -1176 -1938 -1172 -1935
rect -1168 -1935 -1156 -1931
rect -1142 -1935 -1130 -1931
rect -1168 -1938 -1164 -1935
rect -1134 -1938 -1130 -1935
rect -1126 -1935 -1114 -1931
rect -1100 -1931 -1096 -1914
rect -1076 -1917 -1072 -1870
rect -1076 -1931 -1072 -1921
rect -1100 -1935 -1088 -1931
rect -1126 -1938 -1122 -1935
rect -1092 -1938 -1088 -1935
rect -1084 -1935 -1072 -1931
rect -1084 -1938 -1080 -1935
rect -1251 -1946 -1247 -1942
rect -1234 -1946 -1230 -1942
rect -1193 -1946 -1189 -1942
rect -1151 -1946 -1147 -1942
rect -1109 -1946 -1105 -1942
rect -1068 -1946 -1064 -1942
rect -1062 -2006 -1058 -1898
rect -1056 -1998 -1052 -1791
rect -1021 -1788 -1017 -1755
rect -1021 -1823 -1017 -1792
rect -1029 -1831 -1025 -1827
rect -1029 -1862 -1025 -1858
rect -1021 -1903 -1017 -1870
rect -1021 -1938 -1017 -1907
rect -1029 -1946 -1025 -1942
rect -1251 -2093 -1247 -2089
rect -1234 -2093 -1230 -2089
rect -1194 -2093 -1190 -2089
rect -1173 -2093 -1169 -2089
rect -1260 -2134 -1256 -2101
rect -1260 -2169 -1256 -2138
rect -1242 -2128 -1238 -2101
rect -1242 -2132 -1233 -2128
rect -1242 -2169 -1238 -2132
rect -1216 -2155 -1212 -2101
rect -1216 -2162 -1212 -2159
rect -1182 -2162 -1178 -2101
rect -1164 -2133 -1160 -2101
rect -953 -2125 -949 -1722
rect -942 -1795 -938 -1296
rect -916 -1322 -912 -1283
rect -916 -1337 -912 -1326
rect -935 -1341 -912 -1337
rect -909 -1313 -905 -1276
rect -935 -1344 -931 -1341
rect -909 -1344 -905 -1317
rect -918 -1352 -914 -1348
rect -926 -1382 -922 -1378
rect -900 -1382 -896 -1378
rect -883 -1382 -879 -1378
rect -843 -1382 -839 -1378
rect -822 -1382 -818 -1378
rect -805 -1382 -801 -1378
rect -765 -1382 -761 -1378
rect -741 -1382 -737 -1378
rect -704 -1382 -700 -1378
rect -935 -1407 -931 -1390
rect -935 -1458 -931 -1411
rect -917 -1400 -913 -1390
rect -917 -1458 -913 -1404
rect -909 -1429 -905 -1390
rect -891 -1422 -887 -1390
rect -909 -1458 -905 -1433
rect -891 -1458 -887 -1426
rect -865 -1414 -861 -1390
rect -865 -1451 -861 -1418
rect -831 -1451 -827 -1390
rect -813 -1407 -809 -1390
rect -883 -1458 -879 -1455
rect -875 -1455 -861 -1451
rect -875 -1458 -871 -1455
rect -847 -1458 -843 -1455
rect -839 -1455 -820 -1451
rect -839 -1458 -835 -1455
rect -813 -1458 -809 -1411
rect -787 -1422 -783 -1390
rect -787 -1451 -783 -1426
rect -753 -1444 -749 -1390
rect -753 -1448 -736 -1444
rect -805 -1458 -801 -1455
rect -796 -1455 -783 -1451
rect -796 -1458 -792 -1455
rect -769 -1458 -765 -1455
rect -745 -1458 -741 -1448
rect -729 -1451 -725 -1390
rect -721 -1444 -717 -1390
rect -695 -1414 -691 -1390
rect -721 -1448 -702 -1444
rect -737 -1455 -720 -1451
rect -737 -1458 -733 -1455
rect -713 -1458 -709 -1448
rect -695 -1458 -691 -1418
rect -926 -1466 -922 -1462
rect -900 -1466 -896 -1462
rect -857 -1466 -853 -1462
rect -822 -1466 -818 -1462
rect -778 -1466 -774 -1462
rect -761 -1466 -757 -1462
rect -725 -1466 -721 -1462
rect -704 -1466 -700 -1462
rect -689 -1473 -685 -1426
rect -595 -1429 -591 -1317
rect -589 -1414 -585 -1090
rect -583 -1292 -579 -1066
rect -558 -1094 -554 -1053
rect -558 -1107 -554 -1098
rect -577 -1111 -554 -1107
rect -551 -1078 -547 -1046
rect -225 -1062 -221 -998
rect -219 -1038 -215 -1034
rect -202 -1038 -198 -1034
rect -211 -1049 -207 -1046
rect -211 -1053 -196 -1049
rect -225 -1066 -218 -1062
rect -577 -1114 -573 -1111
rect -551 -1114 -547 -1082
rect -560 -1122 -556 -1118
rect -568 -1152 -564 -1148
rect -551 -1152 -547 -1148
rect -531 -1152 -527 -1148
rect -510 -1152 -506 -1148
rect -489 -1152 -485 -1148
rect -468 -1152 -464 -1148
rect -447 -1152 -443 -1148
rect -426 -1152 -422 -1148
rect -405 -1152 -401 -1148
rect -385 -1152 -381 -1148
rect -577 -1207 -573 -1160
rect -577 -1228 -573 -1211
rect -559 -1221 -555 -1160
rect -543 -1221 -539 -1160
rect -519 -1200 -515 -1160
rect -519 -1221 -515 -1204
rect -501 -1221 -497 -1160
rect -477 -1207 -473 -1160
rect -477 -1221 -473 -1211
rect -459 -1200 -455 -1160
rect -459 -1221 -455 -1204
rect -435 -1214 -431 -1160
rect -417 -1192 -413 -1160
rect -417 -1200 -413 -1196
rect -435 -1221 -431 -1218
rect -559 -1225 -550 -1221
rect -543 -1225 -535 -1221
rect -559 -1228 -555 -1225
rect -535 -1228 -531 -1225
rect -527 -1225 -515 -1221
rect -501 -1225 -493 -1221
rect -527 -1228 -523 -1225
rect -493 -1228 -489 -1225
rect -485 -1225 -473 -1221
rect -459 -1225 -447 -1221
rect -485 -1228 -481 -1225
rect -451 -1228 -447 -1225
rect -443 -1225 -431 -1221
rect -417 -1221 -413 -1204
rect -393 -1207 -389 -1160
rect -393 -1221 -389 -1211
rect -417 -1225 -405 -1221
rect -443 -1228 -439 -1225
rect -409 -1228 -405 -1225
rect -401 -1225 -389 -1221
rect -401 -1228 -397 -1225
rect -568 -1236 -564 -1232
rect -551 -1236 -547 -1232
rect -510 -1236 -506 -1232
rect -468 -1236 -464 -1232
rect -426 -1236 -422 -1232
rect -385 -1236 -381 -1232
rect -577 -1268 -573 -1264
rect -560 -1268 -556 -1264
rect -569 -1279 -565 -1276
rect -569 -1283 -554 -1279
rect -583 -1296 -576 -1292
rect -926 -1505 -922 -1501
rect -909 -1505 -905 -1501
rect -889 -1505 -885 -1501
rect -868 -1505 -864 -1501
rect -847 -1505 -843 -1501
rect -826 -1505 -822 -1501
rect -805 -1505 -801 -1501
rect -784 -1505 -780 -1501
rect -763 -1505 -759 -1501
rect -743 -1505 -739 -1501
rect -935 -1560 -931 -1513
rect -935 -1581 -931 -1564
rect -917 -1574 -913 -1513
rect -901 -1574 -897 -1513
rect -877 -1553 -873 -1513
rect -877 -1574 -873 -1557
rect -859 -1574 -855 -1513
rect -835 -1560 -831 -1513
rect -835 -1574 -831 -1564
rect -817 -1553 -813 -1513
rect -817 -1574 -813 -1557
rect -793 -1567 -789 -1513
rect -775 -1545 -771 -1513
rect -775 -1553 -771 -1549
rect -793 -1574 -789 -1571
rect -917 -1578 -908 -1574
rect -901 -1578 -893 -1574
rect -917 -1581 -913 -1578
rect -893 -1581 -889 -1578
rect -885 -1578 -873 -1574
rect -859 -1578 -851 -1574
rect -885 -1581 -881 -1578
rect -851 -1581 -847 -1578
rect -843 -1578 -831 -1574
rect -817 -1578 -805 -1574
rect -843 -1581 -839 -1578
rect -809 -1581 -805 -1578
rect -801 -1578 -789 -1574
rect -775 -1574 -771 -1557
rect -751 -1560 -747 -1513
rect -751 -1574 -747 -1564
rect -775 -1578 -763 -1574
rect -801 -1581 -797 -1578
rect -767 -1581 -763 -1578
rect -759 -1578 -747 -1574
rect -759 -1581 -755 -1578
rect -926 -1589 -922 -1585
rect -909 -1589 -905 -1585
rect -868 -1589 -864 -1585
rect -826 -1589 -822 -1585
rect -784 -1589 -780 -1585
rect -743 -1589 -739 -1585
rect -926 -1626 -922 -1622
rect -909 -1626 -905 -1622
rect -889 -1626 -885 -1622
rect -868 -1626 -864 -1622
rect -847 -1626 -843 -1622
rect -826 -1626 -822 -1622
rect -805 -1626 -801 -1622
rect -784 -1626 -780 -1622
rect -763 -1626 -759 -1622
rect -743 -1626 -739 -1622
rect -935 -1681 -931 -1634
rect -935 -1702 -931 -1685
rect -917 -1695 -913 -1634
rect -901 -1695 -897 -1634
rect -877 -1674 -873 -1634
rect -877 -1695 -873 -1678
rect -859 -1695 -855 -1634
rect -835 -1681 -831 -1634
rect -835 -1695 -831 -1685
rect -817 -1674 -813 -1634
rect -817 -1695 -813 -1678
rect -793 -1688 -789 -1634
rect -775 -1666 -771 -1634
rect -775 -1674 -771 -1670
rect -793 -1695 -789 -1692
rect -917 -1699 -908 -1695
rect -901 -1699 -893 -1695
rect -917 -1702 -913 -1699
rect -893 -1702 -889 -1699
rect -885 -1699 -873 -1695
rect -859 -1699 -851 -1695
rect -885 -1702 -881 -1699
rect -851 -1702 -847 -1699
rect -843 -1699 -831 -1695
rect -817 -1699 -805 -1695
rect -843 -1702 -839 -1699
rect -809 -1702 -805 -1699
rect -801 -1699 -789 -1695
rect -775 -1695 -771 -1678
rect -751 -1681 -747 -1634
rect -751 -1695 -747 -1685
rect -775 -1699 -763 -1695
rect -801 -1702 -797 -1699
rect -767 -1702 -763 -1699
rect -759 -1699 -747 -1695
rect -759 -1702 -755 -1699
rect -926 -1710 -922 -1706
rect -909 -1710 -905 -1706
rect -868 -1710 -864 -1706
rect -826 -1710 -822 -1706
rect -784 -1710 -780 -1706
rect -743 -1710 -739 -1706
rect -737 -1718 -733 -1670
rect -589 -1674 -585 -1491
rect -926 -1747 -922 -1743
rect -909 -1747 -905 -1743
rect -889 -1747 -885 -1743
rect -868 -1747 -864 -1743
rect -847 -1747 -843 -1743
rect -826 -1747 -822 -1743
rect -805 -1747 -801 -1743
rect -784 -1747 -780 -1743
rect -763 -1747 -759 -1743
rect -743 -1747 -739 -1743
rect -935 -1802 -931 -1755
rect -935 -1823 -931 -1806
rect -917 -1816 -913 -1755
rect -901 -1816 -897 -1755
rect -877 -1795 -873 -1755
rect -877 -1816 -873 -1799
rect -859 -1816 -855 -1755
rect -835 -1802 -831 -1755
rect -835 -1816 -831 -1806
rect -817 -1795 -813 -1755
rect -817 -1816 -813 -1799
rect -793 -1809 -789 -1755
rect -775 -1787 -771 -1755
rect -775 -1795 -771 -1791
rect -793 -1816 -789 -1813
rect -917 -1820 -908 -1816
rect -901 -1820 -893 -1816
rect -917 -1823 -913 -1820
rect -893 -1823 -889 -1820
rect -885 -1820 -873 -1816
rect -859 -1820 -851 -1816
rect -885 -1823 -881 -1820
rect -851 -1823 -847 -1820
rect -843 -1820 -831 -1816
rect -817 -1820 -805 -1816
rect -843 -1823 -839 -1820
rect -809 -1823 -805 -1820
rect -801 -1820 -789 -1816
rect -775 -1816 -771 -1799
rect -751 -1802 -747 -1755
rect -751 -1816 -747 -1806
rect -775 -1820 -763 -1816
rect -801 -1823 -797 -1820
rect -767 -1823 -763 -1820
rect -759 -1820 -747 -1816
rect -759 -1823 -755 -1820
rect -926 -1831 -922 -1827
rect -909 -1831 -905 -1827
rect -868 -1831 -864 -1827
rect -826 -1831 -822 -1827
rect -784 -1831 -780 -1827
rect -743 -1831 -739 -1827
rect -935 -1974 -931 -1970
rect -918 -1974 -914 -1970
rect -927 -1985 -923 -1982
rect -927 -1989 -912 -1985
rect -941 -2002 -934 -1998
rect -1234 -2169 -1230 -2166
rect -1225 -2166 -1212 -2162
rect -1225 -2169 -1221 -2166
rect -1198 -2169 -1194 -2166
rect -1190 -2166 -1171 -2162
rect -1190 -2169 -1186 -2166
rect -1164 -2169 -1160 -2137
rect -947 -2140 -943 -2023
rect -1251 -2177 -1247 -2173
rect -1207 -2177 -1203 -2173
rect -1173 -2177 -1169 -2173
rect -1276 -2416 -1272 -2188
rect -1158 -2191 -1154 -2159
rect -1270 -2285 -1266 -2195
rect -1255 -2237 -1251 -2233
rect -1238 -2237 -1234 -2233
rect -1218 -2237 -1214 -2233
rect -1197 -2237 -1193 -2233
rect -1176 -2237 -1172 -2233
rect -1155 -2237 -1151 -2233
rect -1134 -2237 -1130 -2233
rect -1113 -2237 -1109 -2233
rect -1092 -2237 -1088 -2233
rect -1072 -2237 -1068 -2233
rect -1264 -2292 -1260 -2245
rect -1264 -2313 -1260 -2296
rect -1246 -2306 -1242 -2245
rect -1230 -2306 -1226 -2245
rect -1206 -2285 -1202 -2245
rect -1206 -2306 -1202 -2289
rect -1188 -2306 -1184 -2245
rect -1164 -2292 -1160 -2245
rect -1164 -2306 -1160 -2296
rect -1146 -2285 -1142 -2245
rect -1146 -2306 -1142 -2289
rect -1122 -2299 -1118 -2245
rect -1104 -2277 -1100 -2245
rect -1104 -2285 -1100 -2281
rect -1122 -2306 -1118 -2303
rect -1246 -2310 -1237 -2306
rect -1230 -2310 -1222 -2306
rect -1246 -2313 -1242 -2310
rect -1222 -2313 -1218 -2310
rect -1214 -2310 -1202 -2306
rect -1188 -2310 -1180 -2306
rect -1214 -2313 -1210 -2310
rect -1180 -2313 -1176 -2310
rect -1172 -2310 -1160 -2306
rect -1146 -2310 -1134 -2306
rect -1172 -2313 -1168 -2310
rect -1138 -2313 -1134 -2310
rect -1130 -2310 -1118 -2306
rect -1104 -2306 -1100 -2289
rect -1080 -2292 -1076 -2245
rect -1080 -2306 -1076 -2296
rect -1104 -2310 -1092 -2306
rect -1130 -2313 -1126 -2310
rect -1096 -2313 -1092 -2310
rect -1088 -2310 -1076 -2306
rect -1088 -2313 -1084 -2310
rect -1255 -2321 -1251 -2317
rect -1238 -2321 -1234 -2317
rect -1197 -2321 -1193 -2317
rect -1155 -2321 -1151 -2317
rect -1113 -2321 -1109 -2317
rect -1072 -2321 -1068 -2317
rect -1255 -2368 -1251 -2364
rect -1238 -2368 -1234 -2364
rect -1218 -2368 -1214 -2364
rect -1197 -2368 -1193 -2364
rect -1176 -2368 -1172 -2364
rect -1155 -2368 -1151 -2364
rect -1134 -2368 -1130 -2364
rect -1113 -2368 -1109 -2364
rect -1092 -2368 -1088 -2364
rect -1072 -2368 -1068 -2364
rect -1264 -2423 -1260 -2376
rect -1264 -2444 -1260 -2427
rect -1246 -2437 -1242 -2376
rect -1230 -2437 -1226 -2376
rect -1206 -2416 -1202 -2376
rect -1206 -2437 -1202 -2420
rect -1188 -2437 -1184 -2376
rect -1164 -2423 -1160 -2376
rect -1164 -2437 -1160 -2427
rect -1146 -2416 -1142 -2376
rect -1146 -2437 -1142 -2420
rect -1122 -2430 -1118 -2376
rect -1104 -2408 -1100 -2376
rect -1104 -2416 -1100 -2412
rect -1122 -2437 -1118 -2434
rect -1246 -2441 -1237 -2437
rect -1230 -2441 -1222 -2437
rect -1246 -2444 -1242 -2441
rect -1222 -2444 -1218 -2441
rect -1214 -2441 -1202 -2437
rect -1188 -2441 -1180 -2437
rect -1214 -2444 -1210 -2441
rect -1180 -2444 -1176 -2441
rect -1172 -2441 -1160 -2437
rect -1146 -2441 -1134 -2437
rect -1172 -2444 -1168 -2441
rect -1138 -2444 -1134 -2441
rect -1130 -2441 -1118 -2437
rect -1104 -2437 -1100 -2420
rect -1080 -2423 -1076 -2376
rect -1080 -2437 -1076 -2427
rect -1104 -2441 -1092 -2437
rect -1130 -2444 -1126 -2441
rect -1096 -2444 -1092 -2441
rect -1088 -2441 -1076 -2437
rect -1088 -2444 -1084 -2441
rect -1255 -2452 -1251 -2448
rect -1238 -2452 -1234 -2448
rect -1197 -2452 -1193 -2448
rect -1155 -2452 -1151 -2448
rect -1113 -2452 -1109 -2448
rect -1072 -2452 -1068 -2448
rect -1066 -2460 -1062 -2412
rect -947 -2416 -943 -2195
rect -1339 -2724 -1335 -2720
rect -1322 -2724 -1318 -2720
rect -1331 -2735 -1327 -2732
rect -1331 -2739 -1316 -2735
rect -1349 -2752 -1338 -2748
rect -1349 -3247 -1345 -2752
rect -1320 -2778 -1316 -2739
rect -1320 -2793 -1316 -2782
rect -1339 -2797 -1316 -2793
rect -1339 -2800 -1335 -2797
rect -1313 -2800 -1309 -2732
rect -1322 -2808 -1318 -2804
rect -1313 -2898 -1309 -2804
rect -1270 -2891 -1266 -2464
rect -1255 -2499 -1251 -2495
rect -1238 -2499 -1234 -2495
rect -1218 -2499 -1214 -2495
rect -1197 -2499 -1193 -2495
rect -1176 -2499 -1172 -2495
rect -1155 -2499 -1151 -2495
rect -1134 -2499 -1130 -2495
rect -1113 -2499 -1109 -2495
rect -1092 -2499 -1088 -2495
rect -1072 -2499 -1068 -2495
rect -1264 -2554 -1260 -2507
rect -1264 -2575 -1260 -2558
rect -1246 -2568 -1242 -2507
rect -1230 -2568 -1226 -2507
rect -1206 -2547 -1202 -2507
rect -1206 -2568 -1202 -2551
rect -1188 -2568 -1184 -2507
rect -1164 -2554 -1160 -2507
rect -1164 -2568 -1160 -2558
rect -1146 -2547 -1142 -2507
rect -1146 -2568 -1142 -2551
rect -1122 -2561 -1118 -2507
rect -1104 -2539 -1100 -2507
rect -1104 -2547 -1100 -2543
rect -1122 -2568 -1118 -2565
rect -1246 -2572 -1237 -2568
rect -1230 -2572 -1222 -2568
rect -1246 -2575 -1242 -2572
rect -1222 -2575 -1218 -2572
rect -1214 -2572 -1202 -2568
rect -1188 -2572 -1180 -2568
rect -1214 -2575 -1210 -2572
rect -1180 -2575 -1176 -2572
rect -1172 -2572 -1160 -2568
rect -1146 -2572 -1134 -2568
rect -1172 -2575 -1168 -2572
rect -1138 -2575 -1134 -2572
rect -1130 -2572 -1118 -2568
rect -1104 -2568 -1100 -2551
rect -1080 -2554 -1076 -2507
rect -1080 -2568 -1076 -2558
rect -1104 -2572 -1092 -2568
rect -1130 -2575 -1126 -2572
rect -1096 -2575 -1092 -2572
rect -1088 -2572 -1076 -2568
rect -1088 -2575 -1084 -2572
rect -1255 -2583 -1251 -2579
rect -1238 -2583 -1234 -2579
rect -1197 -2583 -1193 -2579
rect -1155 -2583 -1151 -2579
rect -1113 -2583 -1109 -2579
rect -1072 -2583 -1068 -2579
rect -1255 -2611 -1251 -2607
rect -1238 -2611 -1234 -2607
rect -1218 -2611 -1214 -2607
rect -1197 -2611 -1193 -2607
rect -1176 -2611 -1172 -2607
rect -1155 -2611 -1151 -2607
rect -1134 -2611 -1130 -2607
rect -1113 -2611 -1109 -2607
rect -1092 -2611 -1088 -2607
rect -1072 -2611 -1068 -2607
rect -1264 -2666 -1260 -2619
rect -1264 -2687 -1260 -2670
rect -1246 -2680 -1242 -2619
rect -1230 -2680 -1226 -2619
rect -1206 -2659 -1202 -2619
rect -1206 -2680 -1202 -2663
rect -1188 -2680 -1184 -2619
rect -1164 -2666 -1160 -2619
rect -1164 -2680 -1160 -2670
rect -1146 -2659 -1142 -2619
rect -1146 -2680 -1142 -2663
rect -1122 -2673 -1118 -2619
rect -1104 -2651 -1100 -2619
rect -1104 -2659 -1100 -2655
rect -1122 -2680 -1118 -2677
rect -1246 -2684 -1237 -2680
rect -1230 -2684 -1222 -2680
rect -1246 -2687 -1242 -2684
rect -1222 -2687 -1218 -2684
rect -1214 -2684 -1202 -2680
rect -1188 -2684 -1180 -2680
rect -1214 -2687 -1210 -2684
rect -1180 -2687 -1176 -2684
rect -1172 -2684 -1160 -2680
rect -1146 -2684 -1134 -2680
rect -1172 -2687 -1168 -2684
rect -1138 -2687 -1134 -2684
rect -1130 -2684 -1118 -2680
rect -1104 -2680 -1100 -2663
rect -1080 -2666 -1076 -2619
rect -1080 -2680 -1076 -2670
rect -1104 -2684 -1092 -2680
rect -1130 -2687 -1126 -2684
rect -1096 -2687 -1092 -2684
rect -1088 -2684 -1076 -2680
rect -1088 -2687 -1084 -2684
rect -1255 -2695 -1251 -2691
rect -1238 -2695 -1234 -2691
rect -1197 -2695 -1193 -2691
rect -1155 -2695 -1151 -2691
rect -1113 -2695 -1109 -2691
rect -1072 -2695 -1068 -2691
rect -1066 -2748 -1062 -2543
rect -1255 -2843 -1251 -2839
rect -1238 -2843 -1234 -2839
rect -1198 -2843 -1194 -2839
rect -1177 -2843 -1173 -2839
rect -1264 -2884 -1260 -2851
rect -1264 -2919 -1260 -2888
rect -1246 -2878 -1242 -2851
rect -1246 -2882 -1237 -2878
rect -1246 -2919 -1242 -2882
rect -1220 -2905 -1216 -2851
rect -1220 -2912 -1216 -2909
rect -1186 -2912 -1182 -2851
rect -1168 -2883 -1164 -2851
rect -953 -2875 -949 -2773
rect -1238 -2919 -1234 -2916
rect -1229 -2916 -1216 -2912
rect -1229 -2919 -1225 -2916
rect -1202 -2919 -1198 -2916
rect -1194 -2916 -1175 -2912
rect -1194 -2919 -1190 -2916
rect -1168 -2919 -1164 -2887
rect -947 -2890 -943 -2463
rect -941 -2547 -937 -2002
rect -916 -2028 -912 -1989
rect -916 -2043 -912 -2032
rect -935 -2047 -912 -2043
rect -909 -2019 -905 -1982
rect -737 -1998 -733 -1791
rect -673 -1862 -669 -1858
rect -665 -1903 -661 -1878
rect -665 -1934 -661 -1907
rect -673 -1946 -669 -1942
rect -935 -2050 -931 -2047
rect -909 -2050 -905 -2023
rect -918 -2058 -914 -2054
rect -926 -2093 -922 -2089
rect -900 -2093 -896 -2089
rect -883 -2093 -879 -2089
rect -843 -2093 -839 -2089
rect -822 -2093 -818 -2089
rect -805 -2093 -801 -2089
rect -765 -2093 -761 -2089
rect -741 -2093 -737 -2089
rect -704 -2093 -700 -2089
rect -935 -2118 -931 -2101
rect -935 -2169 -931 -2122
rect -917 -2111 -913 -2101
rect -917 -2169 -913 -2115
rect -909 -2140 -905 -2101
rect -891 -2133 -887 -2101
rect -909 -2169 -905 -2144
rect -891 -2169 -887 -2137
rect -865 -2125 -861 -2101
rect -865 -2162 -861 -2129
rect -831 -2162 -827 -2101
rect -813 -2118 -809 -2101
rect -883 -2169 -879 -2166
rect -875 -2166 -861 -2162
rect -875 -2169 -871 -2166
rect -847 -2169 -843 -2166
rect -839 -2166 -820 -2162
rect -839 -2169 -835 -2166
rect -813 -2169 -809 -2122
rect -787 -2133 -783 -2101
rect -787 -2162 -783 -2137
rect -753 -2155 -749 -2101
rect -753 -2159 -736 -2155
rect -805 -2169 -801 -2166
rect -796 -2166 -783 -2162
rect -796 -2169 -792 -2166
rect -769 -2169 -765 -2166
rect -745 -2169 -741 -2159
rect -729 -2162 -725 -2101
rect -721 -2155 -717 -2101
rect -695 -2125 -691 -2101
rect -721 -2159 -702 -2155
rect -737 -2166 -720 -2162
rect -737 -2169 -733 -2166
rect -713 -2169 -709 -2159
rect -695 -2169 -691 -2129
rect -926 -2177 -922 -2173
rect -900 -2177 -896 -2173
rect -857 -2177 -853 -2173
rect -822 -2177 -818 -2173
rect -778 -2177 -774 -2173
rect -761 -2177 -757 -2173
rect -725 -2177 -721 -2173
rect -704 -2177 -700 -2173
rect -689 -2184 -685 -2137
rect -595 -2140 -591 -2023
rect -589 -2125 -585 -1722
rect -583 -1795 -579 -1296
rect -558 -1322 -554 -1283
rect -558 -1337 -554 -1326
rect -577 -1341 -554 -1337
rect -551 -1313 -547 -1276
rect -577 -1344 -573 -1341
rect -551 -1344 -547 -1317
rect -560 -1352 -556 -1348
rect -568 -1382 -564 -1378
rect -542 -1382 -538 -1378
rect -525 -1382 -521 -1378
rect -485 -1382 -481 -1378
rect -464 -1382 -460 -1378
rect -447 -1382 -443 -1378
rect -407 -1382 -403 -1378
rect -383 -1382 -379 -1378
rect -346 -1382 -342 -1378
rect -577 -1407 -573 -1390
rect -577 -1458 -573 -1411
rect -559 -1400 -555 -1390
rect -559 -1458 -555 -1404
rect -551 -1429 -547 -1390
rect -533 -1422 -529 -1390
rect -551 -1458 -547 -1433
rect -533 -1458 -529 -1426
rect -507 -1414 -503 -1390
rect -507 -1451 -503 -1418
rect -473 -1451 -469 -1390
rect -455 -1407 -451 -1390
rect -525 -1458 -521 -1455
rect -517 -1455 -503 -1451
rect -517 -1458 -513 -1455
rect -489 -1458 -485 -1455
rect -481 -1455 -462 -1451
rect -481 -1458 -477 -1455
rect -455 -1458 -451 -1411
rect -429 -1422 -425 -1390
rect -429 -1451 -425 -1426
rect -395 -1444 -391 -1390
rect -395 -1448 -378 -1444
rect -447 -1458 -443 -1455
rect -438 -1455 -425 -1451
rect -438 -1458 -434 -1455
rect -411 -1458 -407 -1455
rect -387 -1458 -383 -1448
rect -371 -1451 -367 -1390
rect -363 -1444 -359 -1390
rect -337 -1414 -333 -1390
rect -363 -1448 -344 -1444
rect -379 -1455 -362 -1451
rect -379 -1458 -375 -1455
rect -355 -1458 -351 -1448
rect -337 -1458 -333 -1418
rect -568 -1466 -564 -1462
rect -542 -1466 -538 -1462
rect -499 -1466 -495 -1462
rect -464 -1466 -460 -1462
rect -420 -1466 -416 -1462
rect -403 -1466 -399 -1462
rect -367 -1466 -363 -1462
rect -346 -1466 -342 -1462
rect -331 -1480 -327 -1426
rect -237 -1429 -233 -1317
rect -231 -1414 -227 -1082
rect -225 -1292 -221 -1066
rect -200 -1094 -196 -1053
rect -200 -1107 -196 -1098
rect -219 -1111 -196 -1107
rect -193 -1086 -189 -1046
rect 203 -1062 207 -998
rect 209 -1038 213 -1034
rect 226 -1038 230 -1034
rect 217 -1049 221 -1046
rect 217 -1053 232 -1049
rect 203 -1066 210 -1062
rect -219 -1114 -215 -1111
rect -193 -1114 -189 -1090
rect -202 -1122 -198 -1118
rect -210 -1152 -206 -1148
rect -193 -1152 -189 -1148
rect -173 -1152 -169 -1148
rect -152 -1152 -148 -1148
rect -131 -1152 -127 -1148
rect -110 -1152 -106 -1148
rect -89 -1152 -85 -1148
rect -68 -1152 -64 -1148
rect -47 -1152 -43 -1148
rect -27 -1152 -23 -1148
rect -219 -1207 -215 -1160
rect -219 -1228 -215 -1211
rect -201 -1221 -197 -1160
rect -185 -1221 -181 -1160
rect -161 -1200 -157 -1160
rect -161 -1221 -157 -1204
rect -143 -1221 -139 -1160
rect -119 -1207 -115 -1160
rect -119 -1221 -115 -1211
rect -101 -1200 -97 -1160
rect -101 -1221 -97 -1204
rect -77 -1214 -73 -1160
rect -59 -1192 -55 -1160
rect -59 -1200 -55 -1196
rect -77 -1221 -73 -1218
rect -201 -1225 -192 -1221
rect -185 -1225 -177 -1221
rect -201 -1228 -197 -1225
rect -177 -1228 -173 -1225
rect -169 -1225 -157 -1221
rect -143 -1225 -135 -1221
rect -169 -1228 -165 -1225
rect -135 -1228 -131 -1225
rect -127 -1225 -115 -1221
rect -101 -1225 -89 -1221
rect -127 -1228 -123 -1225
rect -93 -1228 -89 -1225
rect -85 -1225 -73 -1221
rect -59 -1221 -55 -1204
rect -35 -1207 -31 -1160
rect -35 -1221 -31 -1211
rect -59 -1225 -47 -1221
rect -85 -1228 -81 -1225
rect -51 -1228 -47 -1225
rect -43 -1225 -31 -1221
rect -43 -1228 -39 -1225
rect -210 -1236 -206 -1232
rect -193 -1236 -189 -1232
rect -152 -1236 -148 -1232
rect -110 -1236 -106 -1232
rect -68 -1236 -64 -1232
rect -27 -1236 -23 -1232
rect -219 -1268 -215 -1264
rect -202 -1268 -198 -1264
rect -211 -1279 -207 -1276
rect -211 -1283 -196 -1279
rect -225 -1296 -218 -1292
rect -568 -1505 -564 -1501
rect -551 -1505 -547 -1501
rect -531 -1505 -527 -1501
rect -510 -1505 -506 -1501
rect -489 -1505 -485 -1501
rect -468 -1505 -464 -1501
rect -447 -1505 -443 -1501
rect -426 -1505 -422 -1501
rect -405 -1505 -401 -1501
rect -385 -1505 -381 -1501
rect -577 -1560 -573 -1513
rect -577 -1581 -573 -1564
rect -559 -1574 -555 -1513
rect -543 -1574 -539 -1513
rect -519 -1553 -515 -1513
rect -519 -1574 -515 -1557
rect -501 -1574 -497 -1513
rect -477 -1560 -473 -1513
rect -477 -1574 -473 -1564
rect -459 -1553 -455 -1513
rect -459 -1574 -455 -1557
rect -435 -1567 -431 -1513
rect -417 -1545 -413 -1513
rect -417 -1553 -413 -1549
rect -435 -1574 -431 -1571
rect -559 -1578 -550 -1574
rect -543 -1578 -535 -1574
rect -559 -1581 -555 -1578
rect -535 -1581 -531 -1578
rect -527 -1578 -515 -1574
rect -501 -1578 -493 -1574
rect -527 -1581 -523 -1578
rect -493 -1581 -489 -1578
rect -485 -1578 -473 -1574
rect -459 -1578 -447 -1574
rect -485 -1581 -481 -1578
rect -451 -1581 -447 -1578
rect -443 -1578 -431 -1574
rect -417 -1574 -413 -1557
rect -393 -1560 -389 -1513
rect -393 -1574 -389 -1564
rect -417 -1578 -405 -1574
rect -443 -1581 -439 -1578
rect -409 -1581 -405 -1578
rect -401 -1578 -389 -1574
rect -401 -1581 -397 -1578
rect -568 -1589 -564 -1585
rect -551 -1589 -547 -1585
rect -510 -1589 -506 -1585
rect -468 -1589 -464 -1585
rect -426 -1589 -422 -1585
rect -385 -1589 -381 -1585
rect -568 -1626 -564 -1622
rect -551 -1626 -547 -1622
rect -531 -1626 -527 -1622
rect -510 -1626 -506 -1622
rect -489 -1626 -485 -1622
rect -468 -1626 -464 -1622
rect -447 -1626 -443 -1622
rect -426 -1626 -422 -1622
rect -405 -1626 -401 -1622
rect -385 -1626 -381 -1622
rect -577 -1681 -573 -1634
rect -577 -1702 -573 -1685
rect -559 -1695 -555 -1634
rect -543 -1695 -539 -1634
rect -519 -1674 -515 -1634
rect -519 -1695 -515 -1678
rect -501 -1695 -497 -1634
rect -477 -1681 -473 -1634
rect -477 -1695 -473 -1685
rect -459 -1674 -455 -1634
rect -459 -1695 -455 -1678
rect -435 -1688 -431 -1634
rect -417 -1666 -413 -1634
rect -417 -1674 -413 -1670
rect -435 -1695 -431 -1692
rect -559 -1699 -550 -1695
rect -543 -1699 -535 -1695
rect -559 -1702 -555 -1699
rect -535 -1702 -531 -1699
rect -527 -1699 -515 -1695
rect -501 -1699 -493 -1695
rect -527 -1702 -523 -1699
rect -493 -1702 -489 -1699
rect -485 -1699 -473 -1695
rect -459 -1699 -447 -1695
rect -485 -1702 -481 -1699
rect -451 -1702 -447 -1699
rect -443 -1699 -431 -1695
rect -417 -1695 -413 -1678
rect -393 -1681 -389 -1634
rect -393 -1695 -389 -1685
rect -417 -1699 -405 -1695
rect -443 -1702 -439 -1699
rect -409 -1702 -405 -1699
rect -401 -1699 -389 -1695
rect -401 -1702 -397 -1699
rect -568 -1710 -564 -1706
rect -551 -1710 -547 -1706
rect -510 -1710 -506 -1706
rect -468 -1710 -464 -1706
rect -426 -1710 -422 -1706
rect -385 -1710 -381 -1706
rect -379 -1718 -375 -1670
rect -231 -1674 -227 -1484
rect -568 -1747 -564 -1743
rect -551 -1747 -547 -1743
rect -531 -1747 -527 -1743
rect -510 -1747 -506 -1743
rect -489 -1747 -485 -1743
rect -468 -1747 -464 -1743
rect -447 -1747 -443 -1743
rect -426 -1747 -422 -1743
rect -405 -1747 -401 -1743
rect -385 -1747 -381 -1743
rect -332 -1747 -328 -1743
rect -577 -1802 -573 -1755
rect -577 -1823 -573 -1806
rect -559 -1816 -555 -1755
rect -543 -1816 -539 -1755
rect -519 -1795 -515 -1755
rect -519 -1816 -515 -1799
rect -501 -1816 -497 -1755
rect -477 -1802 -473 -1755
rect -477 -1816 -473 -1806
rect -459 -1795 -455 -1755
rect -459 -1816 -455 -1799
rect -435 -1809 -431 -1755
rect -417 -1787 -413 -1755
rect -417 -1795 -413 -1791
rect -435 -1816 -431 -1813
rect -559 -1820 -550 -1816
rect -543 -1820 -535 -1816
rect -559 -1823 -555 -1820
rect -535 -1823 -531 -1820
rect -527 -1820 -515 -1816
rect -501 -1820 -493 -1816
rect -527 -1823 -523 -1820
rect -493 -1823 -489 -1820
rect -485 -1820 -473 -1816
rect -459 -1820 -447 -1816
rect -485 -1823 -481 -1820
rect -451 -1823 -447 -1820
rect -443 -1820 -431 -1816
rect -417 -1816 -413 -1799
rect -393 -1802 -389 -1755
rect -393 -1816 -389 -1806
rect -417 -1820 -405 -1816
rect -443 -1823 -439 -1820
rect -409 -1823 -405 -1820
rect -401 -1820 -389 -1816
rect -401 -1823 -397 -1820
rect -568 -1831 -564 -1827
rect -551 -1831 -547 -1827
rect -510 -1831 -506 -1827
rect -468 -1831 -464 -1827
rect -426 -1831 -422 -1827
rect -385 -1831 -381 -1827
rect -577 -1974 -573 -1970
rect -560 -1974 -556 -1970
rect -569 -1985 -565 -1982
rect -569 -1989 -554 -1985
rect -583 -2002 -576 -1998
rect -926 -2237 -922 -2233
rect -909 -2237 -905 -2233
rect -889 -2237 -885 -2233
rect -868 -2237 -864 -2233
rect -847 -2237 -843 -2233
rect -826 -2237 -822 -2233
rect -805 -2237 -801 -2233
rect -784 -2237 -780 -2233
rect -763 -2237 -759 -2233
rect -743 -2237 -739 -2233
rect -935 -2292 -931 -2245
rect -935 -2313 -931 -2296
rect -917 -2306 -913 -2245
rect -901 -2306 -897 -2245
rect -877 -2285 -873 -2245
rect -877 -2306 -873 -2289
rect -859 -2306 -855 -2245
rect -835 -2292 -831 -2245
rect -835 -2306 -831 -2296
rect -817 -2285 -813 -2245
rect -817 -2306 -813 -2289
rect -793 -2299 -789 -2245
rect -775 -2277 -771 -2245
rect -775 -2285 -771 -2281
rect -793 -2306 -789 -2303
rect -917 -2310 -908 -2306
rect -901 -2310 -893 -2306
rect -917 -2313 -913 -2310
rect -893 -2313 -889 -2310
rect -885 -2310 -873 -2306
rect -859 -2310 -851 -2306
rect -885 -2313 -881 -2310
rect -851 -2313 -847 -2310
rect -843 -2310 -831 -2306
rect -817 -2310 -805 -2306
rect -843 -2313 -839 -2310
rect -809 -2313 -805 -2310
rect -801 -2310 -789 -2306
rect -775 -2306 -771 -2289
rect -751 -2292 -747 -2245
rect -751 -2306 -747 -2296
rect -775 -2310 -763 -2306
rect -801 -2313 -797 -2310
rect -767 -2313 -763 -2310
rect -759 -2310 -747 -2306
rect -759 -2313 -755 -2310
rect -926 -2321 -922 -2317
rect -909 -2321 -905 -2317
rect -868 -2321 -864 -2317
rect -826 -2321 -822 -2317
rect -784 -2321 -780 -2317
rect -743 -2321 -739 -2317
rect -926 -2368 -922 -2364
rect -909 -2368 -905 -2364
rect -889 -2368 -885 -2364
rect -868 -2368 -864 -2364
rect -847 -2368 -843 -2364
rect -826 -2368 -822 -2364
rect -805 -2368 -801 -2364
rect -784 -2368 -780 -2364
rect -763 -2368 -759 -2364
rect -743 -2368 -739 -2364
rect -935 -2423 -931 -2376
rect -935 -2444 -931 -2427
rect -917 -2437 -913 -2376
rect -901 -2437 -897 -2376
rect -877 -2416 -873 -2376
rect -877 -2437 -873 -2420
rect -859 -2437 -855 -2376
rect -835 -2423 -831 -2376
rect -835 -2437 -831 -2427
rect -817 -2416 -813 -2376
rect -817 -2437 -813 -2420
rect -793 -2430 -789 -2376
rect -775 -2408 -771 -2376
rect -775 -2416 -771 -2412
rect -793 -2437 -789 -2434
rect -917 -2441 -908 -2437
rect -901 -2441 -893 -2437
rect -917 -2444 -913 -2441
rect -893 -2444 -889 -2441
rect -885 -2441 -873 -2437
rect -859 -2441 -851 -2437
rect -885 -2444 -881 -2441
rect -851 -2444 -847 -2441
rect -843 -2441 -831 -2437
rect -817 -2441 -805 -2437
rect -843 -2444 -839 -2441
rect -809 -2444 -805 -2441
rect -801 -2441 -789 -2437
rect -775 -2437 -771 -2420
rect -751 -2423 -747 -2376
rect -751 -2437 -747 -2427
rect -775 -2441 -763 -2437
rect -801 -2444 -797 -2441
rect -767 -2444 -763 -2441
rect -759 -2441 -747 -2437
rect -759 -2444 -755 -2441
rect -926 -2452 -922 -2448
rect -909 -2452 -905 -2448
rect -868 -2452 -864 -2448
rect -826 -2452 -822 -2448
rect -784 -2452 -780 -2448
rect -743 -2452 -739 -2448
rect -737 -2459 -733 -2412
rect -589 -2416 -585 -2188
rect -926 -2499 -922 -2495
rect -909 -2499 -905 -2495
rect -889 -2499 -885 -2495
rect -868 -2499 -864 -2495
rect -847 -2499 -843 -2495
rect -826 -2499 -822 -2495
rect -805 -2499 -801 -2495
rect -784 -2499 -780 -2495
rect -763 -2499 -759 -2495
rect -743 -2499 -739 -2495
rect -935 -2554 -931 -2507
rect -935 -2575 -931 -2558
rect -917 -2568 -913 -2507
rect -901 -2568 -897 -2507
rect -877 -2547 -873 -2507
rect -877 -2568 -873 -2551
rect -859 -2568 -855 -2507
rect -835 -2554 -831 -2507
rect -835 -2568 -831 -2558
rect -817 -2547 -813 -2507
rect -817 -2568 -813 -2551
rect -793 -2561 -789 -2507
rect -775 -2539 -771 -2507
rect -775 -2547 -771 -2543
rect -793 -2568 -789 -2565
rect -917 -2572 -908 -2568
rect -901 -2572 -893 -2568
rect -917 -2575 -913 -2572
rect -893 -2575 -889 -2572
rect -885 -2572 -873 -2568
rect -859 -2572 -851 -2568
rect -885 -2575 -881 -2572
rect -851 -2575 -847 -2572
rect -843 -2572 -831 -2568
rect -817 -2572 -805 -2568
rect -843 -2575 -839 -2572
rect -809 -2575 -805 -2572
rect -801 -2572 -789 -2568
rect -775 -2568 -771 -2551
rect -751 -2554 -747 -2507
rect -751 -2568 -747 -2558
rect -775 -2572 -763 -2568
rect -801 -2575 -797 -2572
rect -767 -2575 -763 -2572
rect -759 -2572 -747 -2568
rect -759 -2575 -755 -2572
rect -926 -2583 -922 -2579
rect -909 -2583 -905 -2579
rect -868 -2583 -864 -2579
rect -826 -2583 -822 -2579
rect -784 -2583 -780 -2579
rect -743 -2583 -739 -2579
rect -926 -2611 -922 -2607
rect -909 -2611 -905 -2607
rect -889 -2611 -885 -2607
rect -868 -2611 -864 -2607
rect -847 -2611 -843 -2607
rect -826 -2611 -822 -2607
rect -805 -2611 -801 -2607
rect -784 -2611 -780 -2607
rect -763 -2611 -759 -2607
rect -743 -2611 -739 -2607
rect -935 -2666 -931 -2619
rect -935 -2687 -931 -2670
rect -917 -2680 -913 -2619
rect -901 -2680 -897 -2619
rect -877 -2659 -873 -2619
rect -877 -2680 -873 -2663
rect -859 -2680 -855 -2619
rect -835 -2666 -831 -2619
rect -835 -2680 -831 -2670
rect -817 -2659 -813 -2619
rect -817 -2680 -813 -2663
rect -793 -2673 -789 -2619
rect -775 -2651 -771 -2619
rect -775 -2659 -771 -2655
rect -793 -2680 -789 -2677
rect -917 -2684 -908 -2680
rect -901 -2684 -893 -2680
rect -917 -2687 -913 -2684
rect -893 -2687 -889 -2684
rect -885 -2684 -873 -2680
rect -859 -2684 -851 -2680
rect -885 -2687 -881 -2684
rect -851 -2687 -847 -2684
rect -843 -2684 -831 -2680
rect -817 -2684 -805 -2680
rect -843 -2687 -839 -2684
rect -809 -2687 -805 -2684
rect -801 -2684 -789 -2680
rect -775 -2680 -771 -2663
rect -751 -2666 -747 -2619
rect -751 -2680 -747 -2670
rect -775 -2684 -763 -2680
rect -801 -2687 -797 -2684
rect -767 -2687 -763 -2684
rect -759 -2684 -747 -2680
rect -759 -2687 -755 -2684
rect -926 -2695 -922 -2691
rect -909 -2695 -905 -2691
rect -868 -2695 -864 -2691
rect -826 -2695 -822 -2691
rect -784 -2695 -780 -2691
rect -743 -2695 -739 -2691
rect -935 -2724 -931 -2720
rect -918 -2724 -914 -2720
rect -927 -2735 -923 -2732
rect -927 -2739 -912 -2735
rect -941 -2752 -934 -2748
rect -1255 -2927 -1251 -2923
rect -1211 -2927 -1207 -2923
rect -1177 -2927 -1173 -2923
rect -1276 -3126 -1272 -2938
rect -1162 -2942 -1158 -2909
rect -1270 -3010 -1266 -2946
rect -1255 -2962 -1251 -2958
rect -1238 -2962 -1234 -2958
rect -1218 -2962 -1214 -2958
rect -1197 -2962 -1193 -2958
rect -1176 -2962 -1172 -2958
rect -1155 -2962 -1151 -2958
rect -1134 -2962 -1130 -2958
rect -1113 -2962 -1109 -2958
rect -1092 -2962 -1088 -2958
rect -1072 -2962 -1068 -2958
rect -1026 -2962 -1022 -2958
rect -1264 -3017 -1260 -2970
rect -1264 -3038 -1260 -3021
rect -1246 -3031 -1242 -2970
rect -1230 -3031 -1226 -2970
rect -1206 -3010 -1202 -2970
rect -1206 -3031 -1202 -3014
rect -1188 -3031 -1184 -2970
rect -1164 -3017 -1160 -2970
rect -1164 -3031 -1160 -3021
rect -1146 -3010 -1142 -2970
rect -1146 -3031 -1142 -3014
rect -1122 -3024 -1118 -2970
rect -1104 -2975 -1100 -2970
rect -1104 -3010 -1100 -2979
rect -1122 -3031 -1118 -3028
rect -1246 -3035 -1237 -3031
rect -1230 -3035 -1222 -3031
rect -1246 -3038 -1242 -3035
rect -1222 -3038 -1218 -3035
rect -1214 -3035 -1202 -3031
rect -1188 -3035 -1180 -3031
rect -1214 -3038 -1210 -3035
rect -1180 -3038 -1176 -3035
rect -1172 -3035 -1160 -3031
rect -1146 -3035 -1134 -3031
rect -1172 -3038 -1168 -3035
rect -1138 -3038 -1134 -3035
rect -1130 -3035 -1118 -3031
rect -1104 -3031 -1100 -3014
rect -1080 -3017 -1076 -2970
rect -1018 -3004 -1014 -2970
rect -1080 -3031 -1076 -3021
rect -1104 -3035 -1092 -3031
rect -1130 -3038 -1126 -3035
rect -1096 -3038 -1092 -3035
rect -1088 -3035 -1076 -3031
rect -1088 -3038 -1084 -3035
rect -1018 -3038 -1014 -3008
rect -1255 -3046 -1251 -3042
rect -1238 -3046 -1234 -3042
rect -1197 -3046 -1193 -3042
rect -1155 -3046 -1151 -3042
rect -1113 -3046 -1109 -3042
rect -1072 -3046 -1068 -3042
rect -1026 -3046 -1022 -3042
rect -1255 -3078 -1251 -3074
rect -1238 -3078 -1234 -3074
rect -1218 -3078 -1214 -3074
rect -1197 -3078 -1193 -3074
rect -1176 -3078 -1172 -3074
rect -1155 -3078 -1151 -3074
rect -1134 -3078 -1130 -3074
rect -1113 -3078 -1109 -3074
rect -1092 -3078 -1088 -3074
rect -1072 -3078 -1068 -3074
rect -1026 -3078 -1022 -3074
rect -1264 -3133 -1260 -3086
rect -1264 -3154 -1260 -3137
rect -1246 -3147 -1242 -3086
rect -1230 -3147 -1226 -3086
rect -1206 -3126 -1202 -3086
rect -1206 -3147 -1202 -3130
rect -1188 -3147 -1184 -3086
rect -1164 -3133 -1160 -3086
rect -1164 -3147 -1160 -3137
rect -1146 -3126 -1142 -3086
rect -1146 -3147 -1142 -3130
rect -1122 -3140 -1118 -3086
rect -1104 -3118 -1100 -3086
rect -1104 -3126 -1100 -3122
rect -1122 -3147 -1118 -3144
rect -1246 -3151 -1237 -3147
rect -1230 -3151 -1222 -3147
rect -1246 -3154 -1242 -3151
rect -1222 -3154 -1218 -3151
rect -1214 -3151 -1202 -3147
rect -1188 -3151 -1180 -3147
rect -1214 -3154 -1210 -3151
rect -1180 -3154 -1176 -3151
rect -1172 -3151 -1160 -3147
rect -1146 -3151 -1134 -3147
rect -1172 -3154 -1168 -3151
rect -1138 -3154 -1134 -3151
rect -1130 -3151 -1118 -3147
rect -1104 -3147 -1100 -3130
rect -1080 -3133 -1076 -3086
rect -1080 -3147 -1076 -3137
rect -1104 -3151 -1092 -3147
rect -1130 -3154 -1126 -3151
rect -1096 -3154 -1092 -3151
rect -1088 -3151 -1076 -3147
rect -1088 -3154 -1084 -3151
rect -1255 -3162 -1251 -3158
rect -1238 -3162 -1234 -3158
rect -1197 -3162 -1193 -3158
rect -1155 -3162 -1151 -3158
rect -1113 -3162 -1109 -3158
rect -1072 -3162 -1068 -3158
rect -1066 -3170 -1062 -3122
rect -1018 -3119 -1014 -3086
rect -1018 -3154 -1014 -3123
rect -947 -3126 -943 -2945
rect -1026 -3162 -1022 -3158
rect -1339 -3430 -1335 -3426
rect -1322 -3430 -1318 -3426
rect -1331 -3441 -1327 -3438
rect -1331 -3445 -1316 -3441
rect -1349 -3458 -1338 -3454
rect -1629 -3851 -1621 -3837
rect -1349 -4088 -1345 -3458
rect -1320 -3484 -1316 -3445
rect -1320 -3499 -1316 -3488
rect -1339 -3503 -1316 -3499
rect -1339 -3506 -1335 -3503
rect -1313 -3506 -1309 -3438
rect -1322 -3514 -1318 -3510
rect -1313 -3609 -1309 -3510
rect -1270 -3602 -1266 -3174
rect -1255 -3199 -1251 -3195
rect -1238 -3199 -1234 -3195
rect -1218 -3199 -1214 -3195
rect -1197 -3199 -1193 -3195
rect -1176 -3199 -1172 -3195
rect -1155 -3199 -1151 -3195
rect -1134 -3199 -1130 -3195
rect -1113 -3199 -1109 -3195
rect -1092 -3199 -1088 -3195
rect -1072 -3199 -1068 -3195
rect -1264 -3254 -1260 -3207
rect -1264 -3275 -1260 -3258
rect -1246 -3268 -1242 -3207
rect -1230 -3268 -1226 -3207
rect -1206 -3247 -1202 -3207
rect -1206 -3268 -1202 -3251
rect -1188 -3268 -1184 -3207
rect -1164 -3254 -1160 -3207
rect -1164 -3268 -1160 -3258
rect -1146 -3247 -1142 -3207
rect -1146 -3268 -1142 -3251
rect -1122 -3261 -1118 -3207
rect -1104 -3239 -1100 -3207
rect -1104 -3247 -1100 -3243
rect -1122 -3268 -1118 -3265
rect -1246 -3272 -1237 -3268
rect -1230 -3272 -1222 -3268
rect -1246 -3275 -1242 -3272
rect -1222 -3275 -1218 -3272
rect -1214 -3272 -1202 -3268
rect -1188 -3272 -1180 -3268
rect -1214 -3275 -1210 -3272
rect -1180 -3275 -1176 -3272
rect -1172 -3272 -1160 -3268
rect -1146 -3272 -1134 -3268
rect -1172 -3275 -1168 -3272
rect -1138 -3275 -1134 -3272
rect -1130 -3272 -1118 -3268
rect -1104 -3268 -1100 -3251
rect -1080 -3254 -1076 -3207
rect -1080 -3268 -1076 -3258
rect -1104 -3272 -1092 -3268
rect -1130 -3275 -1126 -3272
rect -1096 -3275 -1092 -3272
rect -1088 -3272 -1076 -3268
rect -1088 -3275 -1084 -3272
rect -1255 -3283 -1251 -3279
rect -1238 -3283 -1234 -3279
rect -1197 -3283 -1193 -3279
rect -1155 -3283 -1151 -3279
rect -1113 -3283 -1109 -3279
rect -1072 -3283 -1068 -3279
rect -1255 -3313 -1251 -3309
rect -1238 -3313 -1234 -3309
rect -1218 -3313 -1214 -3309
rect -1197 -3313 -1193 -3309
rect -1176 -3313 -1172 -3309
rect -1155 -3313 -1151 -3309
rect -1134 -3313 -1130 -3309
rect -1113 -3313 -1109 -3309
rect -1092 -3313 -1088 -3309
rect -1072 -3313 -1068 -3309
rect -1264 -3368 -1260 -3321
rect -1264 -3389 -1260 -3372
rect -1246 -3382 -1242 -3321
rect -1230 -3382 -1226 -3321
rect -1206 -3361 -1202 -3321
rect -1206 -3382 -1202 -3365
rect -1188 -3382 -1184 -3321
rect -1164 -3368 -1160 -3321
rect -1164 -3382 -1160 -3372
rect -1146 -3361 -1142 -3321
rect -1146 -3382 -1142 -3365
rect -1122 -3375 -1118 -3321
rect -1104 -3353 -1100 -3321
rect -1104 -3361 -1100 -3357
rect -1122 -3382 -1118 -3379
rect -1246 -3386 -1237 -3382
rect -1230 -3386 -1222 -3382
rect -1246 -3389 -1242 -3386
rect -1222 -3389 -1218 -3386
rect -1214 -3386 -1202 -3382
rect -1188 -3386 -1180 -3382
rect -1214 -3389 -1210 -3386
rect -1180 -3389 -1176 -3386
rect -1172 -3386 -1160 -3382
rect -1146 -3386 -1134 -3382
rect -1172 -3389 -1168 -3386
rect -1138 -3389 -1134 -3386
rect -1130 -3386 -1118 -3382
rect -1104 -3382 -1100 -3365
rect -1080 -3368 -1076 -3321
rect -1080 -3382 -1076 -3372
rect -1104 -3386 -1092 -3382
rect -1130 -3389 -1126 -3386
rect -1096 -3389 -1092 -3386
rect -1088 -3386 -1076 -3382
rect -1088 -3389 -1084 -3386
rect -1255 -3397 -1251 -3393
rect -1238 -3397 -1234 -3393
rect -1197 -3397 -1193 -3393
rect -1155 -3397 -1151 -3393
rect -1113 -3397 -1109 -3393
rect -1072 -3397 -1068 -3393
rect -1066 -3454 -1062 -3243
rect -1255 -3554 -1251 -3550
rect -1238 -3554 -1234 -3550
rect -1198 -3554 -1194 -3550
rect -1177 -3554 -1173 -3550
rect -1264 -3595 -1260 -3562
rect -1264 -3630 -1260 -3599
rect -1246 -3589 -1242 -3562
rect -1246 -3593 -1237 -3589
rect -1246 -3630 -1242 -3593
rect -1220 -3616 -1216 -3562
rect -1220 -3623 -1216 -3620
rect -1186 -3623 -1182 -3562
rect -1168 -3594 -1164 -3562
rect -953 -3586 -949 -3479
rect -1238 -3630 -1234 -3627
rect -1229 -3627 -1216 -3623
rect -1229 -3630 -1225 -3627
rect -1202 -3630 -1198 -3627
rect -1194 -3627 -1175 -3623
rect -1194 -3630 -1190 -3627
rect -1168 -3630 -1164 -3598
rect -947 -3601 -943 -3174
rect -941 -3247 -937 -2752
rect -916 -2778 -912 -2739
rect -916 -2793 -912 -2782
rect -935 -2797 -912 -2793
rect -909 -2769 -905 -2732
rect -737 -2756 -733 -2655
rect -731 -2748 -727 -2543
rect -935 -2800 -931 -2797
rect -909 -2800 -905 -2773
rect -918 -2808 -914 -2804
rect -926 -2843 -922 -2839
rect -900 -2843 -896 -2839
rect -883 -2843 -879 -2839
rect -843 -2843 -839 -2839
rect -822 -2843 -818 -2839
rect -805 -2843 -801 -2839
rect -765 -2843 -761 -2839
rect -741 -2843 -737 -2839
rect -704 -2843 -700 -2839
rect -935 -2868 -931 -2851
rect -935 -2919 -931 -2872
rect -917 -2861 -913 -2851
rect -917 -2919 -913 -2865
rect -909 -2890 -905 -2851
rect -891 -2883 -887 -2851
rect -909 -2919 -905 -2894
rect -891 -2919 -887 -2887
rect -865 -2875 -861 -2851
rect -865 -2912 -861 -2879
rect -831 -2912 -827 -2851
rect -813 -2868 -809 -2851
rect -883 -2919 -879 -2916
rect -875 -2916 -861 -2912
rect -875 -2919 -871 -2916
rect -847 -2919 -843 -2916
rect -839 -2916 -820 -2912
rect -839 -2919 -835 -2916
rect -813 -2919 -809 -2872
rect -787 -2883 -783 -2851
rect -787 -2912 -783 -2887
rect -753 -2905 -749 -2851
rect -753 -2909 -736 -2905
rect -805 -2919 -801 -2916
rect -796 -2916 -783 -2912
rect -796 -2919 -792 -2916
rect -769 -2919 -765 -2916
rect -745 -2919 -741 -2909
rect -729 -2912 -725 -2851
rect -721 -2905 -717 -2851
rect -695 -2875 -691 -2851
rect -721 -2909 -702 -2905
rect -737 -2916 -720 -2912
rect -737 -2919 -733 -2916
rect -713 -2919 -709 -2909
rect -695 -2919 -691 -2879
rect -926 -2927 -922 -2923
rect -900 -2927 -896 -2923
rect -857 -2927 -853 -2923
rect -822 -2927 -818 -2923
rect -778 -2927 -774 -2923
rect -761 -2927 -757 -2923
rect -725 -2927 -721 -2923
rect -704 -2927 -700 -2923
rect -689 -2934 -685 -2887
rect -595 -2890 -591 -2773
rect -589 -2875 -585 -2464
rect -583 -2547 -579 -2002
rect -558 -2028 -554 -1989
rect -558 -2043 -554 -2032
rect -577 -2047 -554 -2043
rect -551 -2019 -547 -1982
rect -379 -1998 -375 -1791
rect -324 -1788 -320 -1755
rect -324 -1823 -320 -1792
rect -332 -1831 -328 -1827
rect -332 -1862 -328 -1858
rect -324 -1903 -320 -1870
rect -324 -1938 -320 -1907
rect -332 -1946 -328 -1942
rect -577 -2050 -573 -2047
rect -551 -2050 -547 -2023
rect -560 -2058 -556 -2054
rect -568 -2093 -564 -2089
rect -542 -2093 -538 -2089
rect -525 -2093 -521 -2089
rect -485 -2093 -481 -2089
rect -464 -2093 -460 -2089
rect -447 -2093 -443 -2089
rect -407 -2093 -403 -2089
rect -383 -2093 -379 -2089
rect -346 -2093 -342 -2089
rect -577 -2118 -573 -2101
rect -577 -2169 -573 -2122
rect -559 -2111 -555 -2101
rect -559 -2169 -555 -2115
rect -551 -2140 -547 -2101
rect -533 -2133 -529 -2101
rect -551 -2169 -547 -2144
rect -533 -2169 -529 -2137
rect -507 -2125 -503 -2101
rect -507 -2162 -503 -2129
rect -473 -2162 -469 -2101
rect -455 -2118 -451 -2101
rect -525 -2169 -521 -2166
rect -517 -2166 -503 -2162
rect -517 -2169 -513 -2166
rect -489 -2169 -485 -2166
rect -481 -2166 -462 -2162
rect -481 -2169 -477 -2166
rect -455 -2169 -451 -2122
rect -429 -2133 -425 -2101
rect -429 -2162 -425 -2137
rect -395 -2155 -391 -2101
rect -395 -2159 -378 -2155
rect -447 -2169 -443 -2166
rect -438 -2166 -425 -2162
rect -438 -2169 -434 -2166
rect -411 -2169 -407 -2166
rect -387 -2169 -383 -2159
rect -371 -2162 -367 -2101
rect -363 -2155 -359 -2101
rect -337 -2122 -333 -2101
rect -363 -2159 -344 -2155
rect -379 -2166 -362 -2162
rect -379 -2169 -375 -2166
rect -355 -2169 -351 -2159
rect -337 -2169 -333 -2126
rect -568 -2177 -564 -2173
rect -542 -2177 -538 -2173
rect -499 -2177 -495 -2173
rect -464 -2177 -460 -2173
rect -420 -2177 -416 -2173
rect -403 -2177 -399 -2173
rect -367 -2177 -363 -2173
rect -346 -2177 -342 -2173
rect -331 -2191 -327 -2137
rect -237 -2140 -233 -2023
rect -231 -2125 -227 -1721
rect -225 -1795 -221 -1296
rect -200 -1322 -196 -1283
rect -200 -1337 -196 -1326
rect -219 -1341 -196 -1337
rect -193 -1313 -189 -1276
rect -219 -1344 -215 -1341
rect -193 -1344 -189 -1317
rect -202 -1352 -198 -1348
rect -210 -1382 -206 -1378
rect -184 -1382 -180 -1378
rect -167 -1382 -163 -1378
rect -127 -1382 -123 -1378
rect -106 -1382 -102 -1378
rect -89 -1382 -85 -1378
rect -49 -1382 -45 -1378
rect -25 -1382 -21 -1378
rect 12 -1382 16 -1378
rect -219 -1407 -215 -1390
rect -219 -1458 -215 -1411
rect -201 -1400 -197 -1390
rect -201 -1458 -197 -1404
rect -193 -1429 -189 -1390
rect -175 -1422 -171 -1390
rect -193 -1458 -189 -1433
rect -175 -1458 -171 -1426
rect -149 -1414 -145 -1390
rect -149 -1451 -145 -1418
rect -115 -1451 -111 -1390
rect -97 -1407 -93 -1390
rect -167 -1458 -163 -1455
rect -159 -1455 -145 -1451
rect -159 -1458 -155 -1455
rect -131 -1458 -127 -1455
rect -123 -1455 -104 -1451
rect -123 -1458 -119 -1455
rect -97 -1458 -93 -1411
rect -71 -1422 -67 -1390
rect -71 -1451 -67 -1426
rect -37 -1444 -33 -1390
rect -37 -1448 -20 -1444
rect -89 -1458 -85 -1455
rect -80 -1455 -67 -1451
rect -80 -1458 -76 -1455
rect -53 -1458 -49 -1455
rect -29 -1458 -25 -1448
rect -13 -1451 -9 -1390
rect -5 -1444 -1 -1390
rect 21 -1414 25 -1390
rect -5 -1448 14 -1444
rect -21 -1455 -4 -1451
rect -21 -1458 -17 -1455
rect 3 -1458 7 -1448
rect 21 -1458 25 -1418
rect -210 -1466 -206 -1462
rect -184 -1466 -180 -1462
rect -141 -1466 -137 -1462
rect -106 -1466 -102 -1462
rect -62 -1466 -58 -1462
rect -45 -1466 -41 -1462
rect -9 -1466 -5 -1462
rect 12 -1466 16 -1462
rect 27 -1487 31 -1426
rect 191 -1429 195 -1317
rect 197 -1414 201 -1090
rect 203 -1292 207 -1066
rect 228 -1107 232 -1053
rect 209 -1111 228 -1107
rect 235 -1078 239 -1046
rect 559 -1062 563 -998
rect 565 -1038 569 -1034
rect 582 -1038 586 -1034
rect 573 -1049 577 -1046
rect 573 -1053 588 -1049
rect 559 -1066 566 -1062
rect 209 -1114 213 -1111
rect 235 -1114 239 -1082
rect 226 -1122 230 -1118
rect 218 -1152 222 -1148
rect 235 -1152 239 -1148
rect 255 -1152 259 -1148
rect 276 -1152 280 -1148
rect 297 -1152 301 -1148
rect 318 -1152 322 -1148
rect 339 -1152 343 -1148
rect 360 -1152 364 -1148
rect 381 -1152 385 -1148
rect 401 -1152 405 -1148
rect 209 -1207 213 -1160
rect 209 -1228 213 -1211
rect 227 -1221 231 -1160
rect 243 -1221 247 -1160
rect 267 -1200 271 -1160
rect 267 -1221 271 -1204
rect 285 -1221 289 -1160
rect 309 -1207 313 -1160
rect 309 -1221 313 -1211
rect 327 -1200 331 -1160
rect 327 -1221 331 -1204
rect 351 -1214 355 -1160
rect 369 -1192 373 -1160
rect 369 -1200 373 -1196
rect 351 -1221 355 -1218
rect 227 -1225 236 -1221
rect 243 -1225 251 -1221
rect 227 -1228 231 -1225
rect 251 -1228 255 -1225
rect 259 -1225 271 -1221
rect 285 -1225 293 -1221
rect 259 -1228 263 -1225
rect 293 -1228 297 -1225
rect 301 -1225 313 -1221
rect 327 -1225 339 -1221
rect 301 -1228 305 -1225
rect 335 -1228 339 -1225
rect 343 -1225 355 -1221
rect 369 -1221 373 -1204
rect 393 -1207 397 -1160
rect 393 -1221 397 -1211
rect 369 -1225 381 -1221
rect 343 -1228 347 -1225
rect 377 -1228 381 -1225
rect 385 -1225 397 -1221
rect 385 -1228 389 -1225
rect 218 -1236 222 -1232
rect 235 -1236 239 -1232
rect 276 -1236 280 -1232
rect 318 -1236 322 -1232
rect 360 -1236 364 -1232
rect 401 -1236 405 -1232
rect 209 -1268 213 -1264
rect 226 -1268 230 -1264
rect 217 -1279 221 -1276
rect 217 -1283 232 -1279
rect 203 -1296 210 -1292
rect -210 -1505 -206 -1501
rect -193 -1505 -189 -1501
rect -173 -1505 -169 -1501
rect -152 -1505 -148 -1501
rect -131 -1505 -127 -1501
rect -110 -1505 -106 -1501
rect -89 -1505 -85 -1501
rect -68 -1505 -64 -1501
rect -47 -1505 -43 -1501
rect -27 -1505 -23 -1501
rect -219 -1560 -215 -1513
rect -219 -1581 -215 -1564
rect -201 -1574 -197 -1513
rect -185 -1574 -181 -1513
rect -161 -1553 -157 -1513
rect -161 -1574 -157 -1557
rect -143 -1574 -139 -1513
rect -119 -1560 -115 -1513
rect -119 -1574 -115 -1564
rect -101 -1553 -97 -1513
rect -101 -1574 -97 -1557
rect -77 -1567 -73 -1513
rect -59 -1545 -55 -1513
rect -59 -1553 -55 -1549
rect -77 -1574 -73 -1571
rect -201 -1578 -192 -1574
rect -185 -1578 -177 -1574
rect -201 -1581 -197 -1578
rect -177 -1581 -173 -1578
rect -169 -1578 -157 -1574
rect -143 -1578 -135 -1574
rect -169 -1581 -165 -1578
rect -135 -1581 -131 -1578
rect -127 -1578 -115 -1574
rect -101 -1578 -89 -1574
rect -127 -1581 -123 -1578
rect -93 -1581 -89 -1578
rect -85 -1578 -73 -1574
rect -59 -1574 -55 -1557
rect -35 -1560 -31 -1513
rect -35 -1574 -31 -1564
rect -59 -1578 -47 -1574
rect -85 -1581 -81 -1578
rect -51 -1581 -47 -1578
rect -43 -1578 -31 -1574
rect -43 -1581 -39 -1578
rect -210 -1589 -206 -1585
rect -193 -1589 -189 -1585
rect -152 -1589 -148 -1585
rect -110 -1589 -106 -1585
rect -68 -1589 -64 -1585
rect -27 -1589 -23 -1585
rect -210 -1626 -206 -1622
rect -193 -1626 -189 -1622
rect -173 -1626 -169 -1622
rect -152 -1626 -148 -1622
rect -131 -1626 -127 -1622
rect -110 -1626 -106 -1622
rect -89 -1626 -85 -1622
rect -68 -1626 -64 -1622
rect -47 -1626 -43 -1622
rect -27 -1626 -23 -1622
rect -219 -1681 -215 -1634
rect -219 -1702 -215 -1685
rect -201 -1695 -197 -1634
rect -185 -1695 -181 -1634
rect -161 -1674 -157 -1634
rect -161 -1695 -157 -1678
rect -143 -1695 -139 -1634
rect -119 -1681 -115 -1634
rect -119 -1695 -115 -1685
rect -101 -1674 -97 -1634
rect -101 -1695 -97 -1678
rect -77 -1688 -73 -1634
rect -59 -1666 -55 -1634
rect -59 -1674 -55 -1670
rect -77 -1695 -73 -1692
rect -201 -1699 -192 -1695
rect -185 -1699 -177 -1695
rect -201 -1702 -197 -1699
rect -177 -1702 -173 -1699
rect -169 -1699 -157 -1695
rect -143 -1699 -135 -1695
rect -169 -1702 -165 -1699
rect -135 -1702 -131 -1699
rect -127 -1699 -115 -1695
rect -101 -1699 -89 -1695
rect -127 -1702 -123 -1699
rect -93 -1702 -89 -1699
rect -85 -1699 -73 -1695
rect -59 -1695 -55 -1678
rect -35 -1681 -31 -1634
rect -35 -1695 -31 -1685
rect -59 -1699 -47 -1695
rect -85 -1702 -81 -1699
rect -51 -1702 -47 -1699
rect -43 -1699 -31 -1695
rect -43 -1702 -39 -1699
rect -210 -1710 -206 -1706
rect -193 -1710 -189 -1706
rect -152 -1710 -148 -1706
rect -110 -1710 -106 -1706
rect -68 -1710 -64 -1706
rect -27 -1710 -23 -1706
rect -21 -1717 -17 -1670
rect 197 -1674 201 -1491
rect -210 -1747 -206 -1743
rect -193 -1747 -189 -1743
rect -173 -1747 -169 -1743
rect -152 -1747 -148 -1743
rect -131 -1747 -127 -1743
rect -110 -1747 -106 -1743
rect -89 -1747 -85 -1743
rect -68 -1747 -64 -1743
rect -47 -1747 -43 -1743
rect -27 -1747 -23 -1743
rect -219 -1802 -215 -1755
rect -219 -1823 -215 -1806
rect -201 -1816 -197 -1755
rect -185 -1816 -181 -1755
rect -161 -1795 -157 -1755
rect -161 -1816 -157 -1799
rect -143 -1816 -139 -1755
rect -119 -1802 -115 -1755
rect -119 -1816 -115 -1806
rect -101 -1795 -97 -1755
rect -101 -1816 -97 -1799
rect -77 -1809 -73 -1755
rect -59 -1787 -55 -1755
rect -59 -1795 -55 -1791
rect -77 -1816 -73 -1813
rect -201 -1820 -192 -1816
rect -185 -1820 -177 -1816
rect -201 -1823 -197 -1820
rect -177 -1823 -173 -1820
rect -169 -1820 -157 -1816
rect -143 -1820 -135 -1816
rect -169 -1823 -165 -1820
rect -135 -1823 -131 -1820
rect -127 -1820 -115 -1816
rect -101 -1820 -89 -1816
rect -127 -1823 -123 -1820
rect -93 -1823 -89 -1820
rect -85 -1820 -73 -1816
rect -59 -1816 -55 -1799
rect -35 -1802 -31 -1755
rect -35 -1816 -31 -1806
rect -59 -1820 -47 -1816
rect -85 -1823 -81 -1820
rect -51 -1823 -47 -1820
rect -43 -1820 -31 -1816
rect -43 -1823 -39 -1820
rect -210 -1831 -206 -1827
rect -193 -1831 -189 -1827
rect -152 -1831 -148 -1827
rect -110 -1831 -106 -1827
rect -68 -1831 -64 -1827
rect -27 -1831 -23 -1827
rect -219 -1974 -215 -1970
rect -202 -1974 -198 -1970
rect -211 -1985 -207 -1982
rect -211 -1989 -196 -1985
rect -225 -2002 -218 -1998
rect -568 -2237 -564 -2233
rect -551 -2237 -547 -2233
rect -531 -2237 -527 -2233
rect -510 -2237 -506 -2233
rect -489 -2237 -485 -2233
rect -468 -2237 -464 -2233
rect -447 -2237 -443 -2233
rect -426 -2237 -422 -2233
rect -405 -2237 -401 -2233
rect -385 -2237 -381 -2233
rect -577 -2292 -573 -2245
rect -577 -2313 -573 -2296
rect -559 -2306 -555 -2245
rect -543 -2306 -539 -2245
rect -519 -2285 -515 -2245
rect -519 -2306 -515 -2289
rect -501 -2306 -497 -2245
rect -477 -2292 -473 -2245
rect -477 -2306 -473 -2296
rect -459 -2285 -455 -2245
rect -459 -2306 -455 -2289
rect -435 -2299 -431 -2245
rect -417 -2277 -413 -2245
rect -417 -2285 -413 -2281
rect -435 -2306 -431 -2303
rect -559 -2310 -550 -2306
rect -543 -2310 -535 -2306
rect -559 -2313 -555 -2310
rect -535 -2313 -531 -2310
rect -527 -2310 -515 -2306
rect -501 -2310 -493 -2306
rect -527 -2313 -523 -2310
rect -493 -2313 -489 -2310
rect -485 -2310 -473 -2306
rect -459 -2310 -447 -2306
rect -485 -2313 -481 -2310
rect -451 -2313 -447 -2310
rect -443 -2310 -431 -2306
rect -417 -2306 -413 -2289
rect -393 -2292 -389 -2245
rect -393 -2306 -389 -2296
rect -417 -2310 -405 -2306
rect -443 -2313 -439 -2310
rect -409 -2313 -405 -2310
rect -401 -2310 -389 -2306
rect -401 -2313 -397 -2310
rect -568 -2321 -564 -2317
rect -551 -2321 -547 -2317
rect -510 -2321 -506 -2317
rect -468 -2321 -464 -2317
rect -426 -2321 -422 -2317
rect -385 -2321 -381 -2317
rect -568 -2368 -564 -2364
rect -551 -2368 -547 -2364
rect -531 -2368 -527 -2364
rect -510 -2368 -506 -2364
rect -489 -2368 -485 -2364
rect -468 -2368 -464 -2364
rect -447 -2368 -443 -2364
rect -426 -2368 -422 -2364
rect -405 -2368 -401 -2364
rect -385 -2368 -381 -2364
rect -577 -2423 -573 -2376
rect -577 -2444 -573 -2427
rect -559 -2437 -555 -2376
rect -543 -2437 -539 -2376
rect -519 -2416 -515 -2376
rect -519 -2437 -515 -2420
rect -501 -2437 -497 -2376
rect -477 -2423 -473 -2376
rect -477 -2437 -473 -2427
rect -459 -2416 -455 -2376
rect -459 -2437 -455 -2420
rect -435 -2430 -431 -2376
rect -417 -2408 -413 -2376
rect -417 -2416 -413 -2412
rect -435 -2437 -431 -2434
rect -559 -2441 -550 -2437
rect -543 -2441 -535 -2437
rect -559 -2444 -555 -2441
rect -535 -2444 -531 -2441
rect -527 -2441 -515 -2437
rect -501 -2441 -493 -2437
rect -527 -2444 -523 -2441
rect -493 -2444 -489 -2441
rect -485 -2441 -473 -2437
rect -459 -2441 -447 -2437
rect -485 -2444 -481 -2441
rect -451 -2444 -447 -2441
rect -443 -2441 -431 -2437
rect -417 -2437 -413 -2420
rect -393 -2423 -389 -2376
rect -393 -2437 -389 -2427
rect -417 -2441 -405 -2437
rect -443 -2444 -439 -2441
rect -409 -2444 -405 -2441
rect -401 -2441 -389 -2437
rect -401 -2444 -397 -2441
rect -568 -2452 -564 -2448
rect -551 -2452 -547 -2448
rect -510 -2452 -506 -2448
rect -468 -2452 -464 -2448
rect -426 -2452 -422 -2448
rect -385 -2452 -381 -2448
rect -379 -2460 -375 -2412
rect -231 -2416 -227 -2195
rect -568 -2499 -564 -2495
rect -551 -2499 -547 -2495
rect -531 -2499 -527 -2495
rect -510 -2499 -506 -2495
rect -489 -2499 -485 -2495
rect -468 -2499 -464 -2495
rect -447 -2499 -443 -2495
rect -426 -2499 -422 -2495
rect -405 -2499 -401 -2495
rect -385 -2499 -381 -2495
rect -577 -2554 -573 -2507
rect -577 -2575 -573 -2558
rect -559 -2568 -555 -2507
rect -543 -2568 -539 -2507
rect -519 -2547 -515 -2507
rect -519 -2568 -515 -2551
rect -501 -2568 -497 -2507
rect -477 -2554 -473 -2507
rect -477 -2568 -473 -2558
rect -459 -2547 -455 -2507
rect -459 -2568 -455 -2551
rect -435 -2561 -431 -2507
rect -417 -2539 -413 -2507
rect -417 -2547 -413 -2543
rect -435 -2568 -431 -2565
rect -559 -2572 -550 -2568
rect -543 -2572 -535 -2568
rect -559 -2575 -555 -2572
rect -535 -2575 -531 -2572
rect -527 -2572 -515 -2568
rect -501 -2572 -493 -2568
rect -527 -2575 -523 -2572
rect -493 -2575 -489 -2572
rect -485 -2572 -473 -2568
rect -459 -2572 -447 -2568
rect -485 -2575 -481 -2572
rect -451 -2575 -447 -2572
rect -443 -2572 -431 -2568
rect -417 -2568 -413 -2551
rect -393 -2554 -389 -2507
rect -393 -2568 -389 -2558
rect -417 -2572 -405 -2568
rect -443 -2575 -439 -2572
rect -409 -2575 -405 -2572
rect -401 -2572 -389 -2568
rect -401 -2575 -397 -2572
rect -568 -2583 -564 -2579
rect -551 -2583 -547 -2579
rect -510 -2583 -506 -2579
rect -468 -2583 -464 -2579
rect -426 -2583 -422 -2579
rect -385 -2583 -381 -2579
rect -577 -2724 -573 -2720
rect -560 -2724 -556 -2720
rect -569 -2735 -565 -2732
rect -569 -2739 -554 -2735
rect -583 -2752 -576 -2748
rect -926 -2962 -922 -2958
rect -909 -2962 -905 -2958
rect -889 -2962 -885 -2958
rect -868 -2962 -864 -2958
rect -847 -2962 -843 -2958
rect -826 -2962 -822 -2958
rect -805 -2962 -801 -2958
rect -784 -2962 -780 -2958
rect -763 -2962 -759 -2958
rect -743 -2962 -739 -2958
rect -672 -2962 -668 -2958
rect -935 -3017 -931 -2970
rect -935 -3038 -931 -3021
rect -917 -3031 -913 -2970
rect -901 -3031 -897 -2970
rect -877 -3010 -873 -2970
rect -877 -3031 -873 -3014
rect -859 -3031 -855 -2970
rect -835 -3017 -831 -2970
rect -835 -3031 -831 -3021
rect -817 -3010 -813 -2970
rect -817 -3031 -813 -3014
rect -793 -3024 -789 -2970
rect -775 -2992 -771 -2970
rect -775 -3010 -771 -2996
rect -793 -3031 -789 -3028
rect -917 -3035 -908 -3031
rect -901 -3035 -893 -3031
rect -917 -3038 -913 -3035
rect -893 -3038 -889 -3035
rect -885 -3035 -873 -3031
rect -859 -3035 -851 -3031
rect -885 -3038 -881 -3035
rect -851 -3038 -847 -3035
rect -843 -3035 -831 -3031
rect -817 -3035 -805 -3031
rect -843 -3038 -839 -3035
rect -809 -3038 -805 -3035
rect -801 -3035 -789 -3031
rect -775 -3031 -771 -3014
rect -751 -3017 -747 -2970
rect -664 -3003 -660 -2978
rect -751 -3031 -747 -3021
rect -775 -3035 -763 -3031
rect -801 -3038 -797 -3035
rect -767 -3038 -763 -3035
rect -759 -3035 -747 -3031
rect -664 -3034 -660 -3007
rect -759 -3038 -755 -3035
rect -926 -3046 -922 -3042
rect -909 -3046 -905 -3042
rect -868 -3046 -864 -3042
rect -826 -3046 -822 -3042
rect -784 -3046 -780 -3042
rect -743 -3046 -739 -3042
rect -672 -3046 -668 -3042
rect -926 -3078 -922 -3074
rect -909 -3078 -905 -3074
rect -889 -3078 -885 -3074
rect -868 -3078 -864 -3074
rect -847 -3078 -843 -3074
rect -826 -3078 -822 -3074
rect -805 -3078 -801 -3074
rect -784 -3078 -780 -3074
rect -763 -3078 -759 -3074
rect -743 -3078 -739 -3074
rect -935 -3133 -931 -3086
rect -935 -3154 -931 -3137
rect -917 -3147 -913 -3086
rect -901 -3147 -897 -3086
rect -877 -3126 -873 -3086
rect -877 -3147 -873 -3130
rect -859 -3147 -855 -3086
rect -835 -3133 -831 -3086
rect -835 -3147 -831 -3137
rect -817 -3126 -813 -3086
rect -817 -3147 -813 -3130
rect -793 -3140 -789 -3086
rect -775 -3118 -771 -3086
rect -775 -3126 -771 -3122
rect -793 -3147 -789 -3144
rect -917 -3151 -908 -3147
rect -901 -3151 -893 -3147
rect -917 -3154 -913 -3151
rect -893 -3154 -889 -3151
rect -885 -3151 -873 -3147
rect -859 -3151 -851 -3147
rect -885 -3154 -881 -3151
rect -851 -3154 -847 -3151
rect -843 -3151 -831 -3147
rect -817 -3151 -805 -3147
rect -843 -3154 -839 -3151
rect -809 -3154 -805 -3151
rect -801 -3151 -789 -3147
rect -775 -3147 -771 -3130
rect -751 -3133 -747 -3086
rect -751 -3147 -747 -3137
rect -775 -3151 -763 -3147
rect -801 -3154 -797 -3151
rect -767 -3154 -763 -3151
rect -759 -3151 -747 -3147
rect -759 -3154 -755 -3151
rect -926 -3162 -922 -3158
rect -909 -3162 -905 -3158
rect -868 -3162 -864 -3158
rect -826 -3162 -822 -3158
rect -784 -3162 -780 -3158
rect -743 -3162 -739 -3158
rect -737 -3170 -733 -3122
rect -589 -3126 -585 -2938
rect -926 -3199 -922 -3195
rect -909 -3199 -905 -3195
rect -889 -3199 -885 -3195
rect -868 -3199 -864 -3195
rect -847 -3199 -843 -3195
rect -826 -3199 -822 -3195
rect -805 -3199 -801 -3195
rect -784 -3199 -780 -3195
rect -763 -3199 -759 -3195
rect -743 -3199 -739 -3195
rect -935 -3254 -931 -3207
rect -935 -3275 -931 -3258
rect -917 -3268 -913 -3207
rect -901 -3268 -897 -3207
rect -877 -3247 -873 -3207
rect -877 -3268 -873 -3251
rect -859 -3268 -855 -3207
rect -835 -3254 -831 -3207
rect -835 -3268 -831 -3258
rect -817 -3247 -813 -3207
rect -817 -3268 -813 -3251
rect -793 -3261 -789 -3207
rect -775 -3239 -771 -3207
rect -775 -3247 -771 -3243
rect -793 -3268 -789 -3265
rect -917 -3272 -908 -3268
rect -901 -3272 -893 -3268
rect -917 -3275 -913 -3272
rect -893 -3275 -889 -3272
rect -885 -3272 -873 -3268
rect -859 -3272 -851 -3268
rect -885 -3275 -881 -3272
rect -851 -3275 -847 -3272
rect -843 -3272 -831 -3268
rect -817 -3272 -805 -3268
rect -843 -3275 -839 -3272
rect -809 -3275 -805 -3272
rect -801 -3272 -789 -3268
rect -775 -3268 -771 -3251
rect -751 -3254 -747 -3207
rect -751 -3268 -747 -3258
rect -775 -3272 -763 -3268
rect -801 -3275 -797 -3272
rect -767 -3275 -763 -3272
rect -759 -3272 -747 -3268
rect -759 -3275 -755 -3272
rect -926 -3283 -922 -3279
rect -909 -3283 -905 -3279
rect -868 -3283 -864 -3279
rect -826 -3283 -822 -3279
rect -784 -3283 -780 -3279
rect -743 -3283 -739 -3279
rect -926 -3313 -922 -3309
rect -909 -3313 -905 -3309
rect -889 -3313 -885 -3309
rect -868 -3313 -864 -3309
rect -847 -3313 -843 -3309
rect -826 -3313 -822 -3309
rect -805 -3313 -801 -3309
rect -784 -3313 -780 -3309
rect -763 -3313 -759 -3309
rect -743 -3313 -739 -3309
rect -935 -3368 -931 -3321
rect -935 -3389 -931 -3372
rect -917 -3382 -913 -3321
rect -901 -3382 -897 -3321
rect -877 -3361 -873 -3321
rect -877 -3382 -873 -3365
rect -859 -3382 -855 -3321
rect -835 -3368 -831 -3321
rect -835 -3382 -831 -3372
rect -817 -3361 -813 -3321
rect -817 -3382 -813 -3365
rect -793 -3375 -789 -3321
rect -775 -3353 -771 -3321
rect -775 -3361 -771 -3357
rect -793 -3382 -789 -3379
rect -917 -3386 -908 -3382
rect -901 -3386 -893 -3382
rect -917 -3389 -913 -3386
rect -893 -3389 -889 -3386
rect -885 -3386 -873 -3382
rect -859 -3386 -851 -3382
rect -885 -3389 -881 -3386
rect -851 -3389 -847 -3386
rect -843 -3386 -831 -3382
rect -817 -3386 -805 -3382
rect -843 -3389 -839 -3386
rect -809 -3389 -805 -3386
rect -801 -3386 -789 -3382
rect -775 -3382 -771 -3365
rect -751 -3368 -747 -3321
rect -751 -3382 -747 -3372
rect -775 -3386 -763 -3382
rect -801 -3389 -797 -3386
rect -767 -3389 -763 -3386
rect -759 -3386 -747 -3382
rect -759 -3389 -755 -3386
rect -926 -3397 -922 -3393
rect -909 -3397 -905 -3393
rect -868 -3397 -864 -3393
rect -826 -3397 -822 -3393
rect -784 -3397 -780 -3393
rect -743 -3397 -739 -3393
rect -935 -3430 -931 -3426
rect -918 -3430 -914 -3426
rect -927 -3441 -923 -3438
rect -927 -3445 -912 -3441
rect -941 -3458 -934 -3454
rect -1255 -3638 -1251 -3634
rect -1211 -3638 -1207 -3634
rect -1177 -3638 -1173 -3634
rect -1276 -3963 -1272 -3649
rect -1162 -3652 -1158 -3620
rect -1270 -3732 -1266 -3656
rect -1255 -3684 -1251 -3680
rect -1238 -3684 -1234 -3680
rect -1218 -3684 -1214 -3680
rect -1197 -3684 -1193 -3680
rect -1176 -3684 -1172 -3680
rect -1155 -3684 -1151 -3680
rect -1134 -3684 -1130 -3680
rect -1113 -3684 -1109 -3680
rect -1092 -3684 -1088 -3680
rect -1072 -3684 -1068 -3680
rect -1264 -3739 -1260 -3692
rect -1264 -3760 -1260 -3743
rect -1246 -3753 -1242 -3692
rect -1230 -3753 -1226 -3692
rect -1206 -3732 -1202 -3692
rect -1206 -3753 -1202 -3736
rect -1188 -3753 -1184 -3692
rect -1164 -3739 -1160 -3692
rect -1164 -3753 -1160 -3743
rect -1146 -3732 -1142 -3692
rect -1146 -3753 -1142 -3736
rect -1122 -3746 -1118 -3692
rect -1104 -3724 -1100 -3692
rect -1104 -3732 -1100 -3728
rect -1122 -3753 -1118 -3750
rect -1246 -3757 -1237 -3753
rect -1230 -3757 -1222 -3753
rect -1246 -3760 -1242 -3757
rect -1222 -3760 -1218 -3757
rect -1214 -3757 -1202 -3753
rect -1188 -3757 -1180 -3753
rect -1214 -3760 -1210 -3757
rect -1180 -3760 -1176 -3757
rect -1172 -3757 -1160 -3753
rect -1146 -3757 -1134 -3753
rect -1172 -3760 -1168 -3757
rect -1138 -3760 -1134 -3757
rect -1130 -3757 -1118 -3753
rect -1104 -3753 -1100 -3736
rect -1080 -3739 -1076 -3692
rect -1080 -3753 -1076 -3743
rect -1104 -3757 -1092 -3753
rect -1130 -3760 -1126 -3757
rect -1096 -3760 -1092 -3757
rect -1088 -3757 -1076 -3753
rect -1088 -3760 -1084 -3757
rect -1255 -3768 -1251 -3764
rect -1238 -3768 -1234 -3764
rect -1197 -3768 -1193 -3764
rect -1155 -3768 -1151 -3764
rect -1113 -3768 -1109 -3764
rect -1072 -3768 -1068 -3764
rect -1255 -3915 -1251 -3911
rect -1238 -3915 -1234 -3911
rect -1218 -3915 -1214 -3911
rect -1197 -3915 -1193 -3911
rect -1176 -3915 -1172 -3911
rect -1155 -3915 -1151 -3911
rect -1134 -3915 -1130 -3911
rect -1113 -3915 -1109 -3911
rect -1092 -3915 -1088 -3911
rect -1072 -3915 -1068 -3911
rect -1264 -3970 -1260 -3923
rect -1264 -3991 -1260 -3974
rect -1246 -3984 -1242 -3923
rect -1230 -3984 -1226 -3923
rect -1206 -3963 -1202 -3923
rect -1206 -3984 -1202 -3967
rect -1188 -3984 -1184 -3923
rect -1164 -3970 -1160 -3923
rect -1164 -3984 -1160 -3974
rect -1146 -3963 -1142 -3923
rect -1146 -3984 -1142 -3967
rect -1122 -3977 -1118 -3923
rect -1104 -3955 -1100 -3923
rect -1104 -3963 -1100 -3959
rect -1122 -3984 -1118 -3981
rect -1246 -3988 -1237 -3984
rect -1230 -3988 -1222 -3984
rect -1246 -3991 -1242 -3988
rect -1222 -3991 -1218 -3988
rect -1214 -3988 -1202 -3984
rect -1188 -3988 -1180 -3984
rect -1214 -3991 -1210 -3988
rect -1180 -3991 -1176 -3988
rect -1172 -3988 -1160 -3984
rect -1146 -3988 -1134 -3984
rect -1172 -3991 -1168 -3988
rect -1138 -3991 -1134 -3988
rect -1130 -3988 -1118 -3984
rect -1104 -3984 -1100 -3967
rect -1080 -3970 -1076 -3923
rect -1080 -3984 -1076 -3974
rect -1104 -3988 -1092 -3984
rect -1130 -3991 -1126 -3988
rect -1096 -3991 -1092 -3988
rect -1088 -3988 -1076 -3984
rect -1088 -3991 -1084 -3988
rect -1255 -3999 -1251 -3995
rect -1238 -3999 -1234 -3995
rect -1197 -3999 -1193 -3995
rect -1155 -3999 -1151 -3995
rect -1113 -3999 -1109 -3995
rect -1072 -3999 -1068 -3995
rect -1066 -4006 -1062 -3959
rect -947 -3963 -943 -3656
rect -1339 -4275 -1335 -4271
rect -1322 -4275 -1318 -4271
rect -1331 -4286 -1327 -4283
rect -1331 -4290 -1316 -4286
rect -1349 -4303 -1338 -4299
rect -1349 -4807 -1345 -4303
rect -1320 -4329 -1316 -4290
rect -1320 -4344 -1316 -4333
rect -1339 -4348 -1316 -4344
rect -1339 -4351 -1335 -4348
rect -1313 -4351 -1309 -4283
rect -1322 -4359 -1318 -4355
rect -1313 -4449 -1309 -4355
rect -1270 -4442 -1266 -4010
rect -1255 -4040 -1251 -4036
rect -1238 -4040 -1234 -4036
rect -1218 -4040 -1214 -4036
rect -1197 -4040 -1193 -4036
rect -1176 -4040 -1172 -4036
rect -1155 -4040 -1151 -4036
rect -1134 -4040 -1130 -4036
rect -1113 -4040 -1109 -4036
rect -1092 -4040 -1088 -4036
rect -1072 -4040 -1068 -4036
rect -1264 -4095 -1260 -4048
rect -1264 -4116 -1260 -4099
rect -1246 -4109 -1242 -4048
rect -1230 -4109 -1226 -4048
rect -1206 -4088 -1202 -4048
rect -1206 -4109 -1202 -4092
rect -1188 -4109 -1184 -4048
rect -1164 -4095 -1160 -4048
rect -1164 -4109 -1160 -4099
rect -1146 -4088 -1142 -4048
rect -1146 -4109 -1142 -4092
rect -1122 -4102 -1118 -4048
rect -1104 -4080 -1100 -4048
rect -1104 -4088 -1100 -4084
rect -1122 -4109 -1118 -4106
rect -1246 -4113 -1237 -4109
rect -1230 -4113 -1222 -4109
rect -1246 -4116 -1242 -4113
rect -1222 -4116 -1218 -4113
rect -1214 -4113 -1202 -4109
rect -1188 -4113 -1180 -4109
rect -1214 -4116 -1210 -4113
rect -1180 -4116 -1176 -4113
rect -1172 -4113 -1160 -4109
rect -1146 -4113 -1134 -4109
rect -1172 -4116 -1168 -4113
rect -1138 -4116 -1134 -4113
rect -1130 -4113 -1118 -4109
rect -1104 -4109 -1100 -4092
rect -1080 -4095 -1076 -4048
rect -1080 -4109 -1076 -4099
rect -1104 -4113 -1092 -4109
rect -1130 -4116 -1126 -4113
rect -1096 -4116 -1092 -4113
rect -1088 -4113 -1076 -4109
rect -1088 -4116 -1084 -4113
rect -1255 -4124 -1251 -4120
rect -1238 -4124 -1234 -4120
rect -1197 -4124 -1193 -4120
rect -1155 -4124 -1151 -4120
rect -1113 -4124 -1109 -4120
rect -1072 -4124 -1068 -4120
rect -1255 -4164 -1251 -4160
rect -1238 -4164 -1234 -4160
rect -1218 -4164 -1214 -4160
rect -1197 -4164 -1193 -4160
rect -1176 -4164 -1172 -4160
rect -1155 -4164 -1151 -4160
rect -1134 -4164 -1130 -4160
rect -1113 -4164 -1109 -4160
rect -1092 -4164 -1088 -4160
rect -1072 -4164 -1068 -4160
rect -1264 -4219 -1260 -4172
rect -1264 -4240 -1260 -4223
rect -1246 -4233 -1242 -4172
rect -1230 -4233 -1226 -4172
rect -1206 -4212 -1202 -4172
rect -1206 -4233 -1202 -4216
rect -1188 -4233 -1184 -4172
rect -1164 -4219 -1160 -4172
rect -1164 -4233 -1160 -4223
rect -1146 -4212 -1142 -4172
rect -1146 -4233 -1142 -4216
rect -1122 -4226 -1118 -4172
rect -1104 -4179 -1100 -4172
rect -1104 -4212 -1100 -4183
rect -1122 -4233 -1118 -4230
rect -1246 -4237 -1237 -4233
rect -1230 -4237 -1222 -4233
rect -1246 -4240 -1242 -4237
rect -1222 -4240 -1218 -4237
rect -1214 -4237 -1202 -4233
rect -1188 -4237 -1180 -4233
rect -1214 -4240 -1210 -4237
rect -1180 -4240 -1176 -4237
rect -1172 -4237 -1160 -4233
rect -1146 -4237 -1134 -4233
rect -1172 -4240 -1168 -4237
rect -1138 -4240 -1134 -4237
rect -1130 -4237 -1118 -4233
rect -1104 -4233 -1100 -4216
rect -1080 -4219 -1076 -4172
rect -1080 -4233 -1076 -4223
rect -1104 -4237 -1092 -4233
rect -1130 -4240 -1126 -4237
rect -1096 -4240 -1092 -4237
rect -1088 -4237 -1076 -4233
rect -1088 -4240 -1084 -4237
rect -1255 -4248 -1251 -4244
rect -1238 -4248 -1234 -4244
rect -1197 -4248 -1193 -4244
rect -1155 -4248 -1151 -4244
rect -1113 -4248 -1109 -4244
rect -1072 -4248 -1068 -4244
rect -1066 -4299 -1062 -4084
rect -1029 -4164 -1025 -4160
rect -1021 -4201 -1017 -4172
rect -1021 -4240 -1017 -4205
rect -1029 -4248 -1025 -4244
rect -1029 -4275 -1025 -4271
rect -1021 -4316 -1017 -4283
rect -1021 -4351 -1017 -4320
rect -1029 -4359 -1025 -4355
rect -1255 -4394 -1251 -4390
rect -1238 -4394 -1234 -4390
rect -1198 -4394 -1194 -4390
rect -1177 -4394 -1173 -4390
rect -1264 -4435 -1260 -4402
rect -1264 -4470 -1260 -4439
rect -1246 -4429 -1242 -4402
rect -1246 -4433 -1237 -4429
rect -1246 -4470 -1242 -4433
rect -1220 -4456 -1216 -4402
rect -1220 -4463 -1216 -4460
rect -1186 -4463 -1182 -4402
rect -1168 -4434 -1164 -4402
rect -953 -4426 -949 -4324
rect -1238 -4470 -1234 -4467
rect -1229 -4467 -1216 -4463
rect -1229 -4470 -1225 -4467
rect -1202 -4470 -1198 -4467
rect -1194 -4467 -1175 -4463
rect -1194 -4470 -1190 -4467
rect -1168 -4470 -1164 -4438
rect -947 -4441 -943 -4011
rect -941 -4088 -937 -3458
rect -916 -3484 -912 -3445
rect -916 -3499 -912 -3488
rect -935 -3503 -912 -3499
rect -909 -3475 -905 -3438
rect -737 -3454 -733 -3243
rect -935 -3506 -931 -3503
rect -909 -3506 -905 -3479
rect -918 -3514 -914 -3510
rect -926 -3554 -922 -3550
rect -900 -3554 -896 -3550
rect -883 -3554 -879 -3550
rect -843 -3554 -839 -3550
rect -822 -3554 -818 -3550
rect -805 -3554 -801 -3550
rect -765 -3554 -761 -3550
rect -741 -3554 -737 -3550
rect -704 -3554 -700 -3550
rect -935 -3579 -931 -3562
rect -935 -3630 -931 -3583
rect -917 -3572 -913 -3562
rect -917 -3630 -913 -3576
rect -909 -3601 -905 -3562
rect -891 -3594 -887 -3562
rect -909 -3630 -905 -3605
rect -891 -3630 -887 -3598
rect -865 -3586 -861 -3562
rect -865 -3623 -861 -3590
rect -831 -3623 -827 -3562
rect -813 -3579 -809 -3562
rect -883 -3630 -879 -3627
rect -875 -3627 -861 -3623
rect -875 -3630 -871 -3627
rect -847 -3630 -843 -3627
rect -839 -3627 -820 -3623
rect -839 -3630 -835 -3627
rect -813 -3630 -809 -3583
rect -787 -3594 -783 -3562
rect -787 -3623 -783 -3598
rect -753 -3616 -749 -3562
rect -753 -3620 -736 -3616
rect -805 -3630 -801 -3627
rect -796 -3627 -783 -3623
rect -796 -3630 -792 -3627
rect -769 -3630 -765 -3627
rect -745 -3630 -741 -3620
rect -729 -3623 -725 -3562
rect -721 -3616 -717 -3562
rect -695 -3586 -691 -3562
rect -721 -3620 -702 -3616
rect -737 -3627 -720 -3623
rect -737 -3630 -733 -3627
rect -713 -3630 -709 -3620
rect -695 -3630 -691 -3590
rect -926 -3638 -922 -3634
rect -900 -3638 -896 -3634
rect -857 -3638 -853 -3634
rect -822 -3638 -818 -3634
rect -778 -3638 -774 -3634
rect -761 -3638 -757 -3634
rect -725 -3638 -721 -3634
rect -704 -3638 -700 -3634
rect -689 -3645 -685 -3598
rect -595 -3601 -591 -3479
rect -589 -3586 -585 -3173
rect -583 -3247 -579 -2752
rect -558 -2778 -554 -2739
rect -558 -2793 -554 -2782
rect -577 -2797 -554 -2793
rect -551 -2769 -547 -2732
rect -379 -2748 -375 -2543
rect -577 -2800 -573 -2797
rect -551 -2800 -547 -2773
rect -560 -2808 -556 -2804
rect -568 -2843 -564 -2839
rect -542 -2843 -538 -2839
rect -525 -2843 -521 -2839
rect -485 -2843 -481 -2839
rect -464 -2843 -460 -2839
rect -447 -2843 -443 -2839
rect -407 -2843 -403 -2839
rect -383 -2843 -379 -2839
rect -346 -2843 -342 -2839
rect -577 -2868 -573 -2851
rect -577 -2919 -573 -2872
rect -559 -2861 -555 -2851
rect -559 -2919 -555 -2865
rect -551 -2890 -547 -2851
rect -533 -2883 -529 -2851
rect -551 -2919 -547 -2894
rect -533 -2919 -529 -2887
rect -507 -2875 -503 -2851
rect -507 -2912 -503 -2879
rect -473 -2912 -469 -2851
rect -455 -2868 -451 -2851
rect -525 -2919 -521 -2916
rect -517 -2916 -503 -2912
rect -517 -2919 -513 -2916
rect -489 -2919 -485 -2916
rect -481 -2916 -462 -2912
rect -481 -2919 -477 -2916
rect -455 -2919 -451 -2872
rect -429 -2883 -425 -2851
rect -429 -2912 -425 -2887
rect -395 -2905 -391 -2851
rect -395 -2909 -378 -2905
rect -447 -2919 -443 -2916
rect -438 -2916 -425 -2912
rect -438 -2919 -434 -2916
rect -411 -2919 -407 -2916
rect -387 -2919 -383 -2909
rect -371 -2912 -367 -2851
rect -363 -2905 -359 -2851
rect -337 -2874 -333 -2851
rect -363 -2909 -344 -2905
rect -379 -2916 -362 -2912
rect -379 -2919 -375 -2916
rect -355 -2919 -351 -2909
rect -337 -2919 -333 -2878
rect -568 -2927 -564 -2923
rect -542 -2927 -538 -2923
rect -499 -2927 -495 -2923
rect -464 -2927 -460 -2923
rect -420 -2927 -416 -2923
rect -403 -2927 -399 -2923
rect -367 -2927 -363 -2923
rect -346 -2927 -342 -2923
rect -331 -2941 -327 -2887
rect -237 -2890 -233 -2773
rect -231 -2875 -227 -2464
rect -225 -2547 -221 -2002
rect -200 -2028 -196 -1989
rect -200 -2043 -196 -2032
rect -219 -2047 -196 -2043
rect -193 -2019 -189 -1982
rect -21 -1998 -17 -1791
rect -219 -2050 -215 -2047
rect -193 -2050 -189 -2023
rect -202 -2058 -198 -2054
rect -210 -2093 -206 -2089
rect -184 -2093 -180 -2089
rect -167 -2093 -163 -2089
rect -127 -2093 -123 -2089
rect -106 -2093 -102 -2089
rect -89 -2093 -85 -2089
rect -49 -2093 -45 -2089
rect -25 -2093 -21 -2089
rect 12 -2093 16 -2089
rect -219 -2118 -215 -2101
rect -219 -2169 -215 -2122
rect -201 -2111 -197 -2101
rect -201 -2169 -197 -2115
rect -193 -2140 -189 -2101
rect -175 -2133 -171 -2101
rect -193 -2169 -189 -2144
rect -175 -2169 -171 -2137
rect -149 -2125 -145 -2101
rect -149 -2162 -145 -2129
rect -115 -2162 -111 -2101
rect -97 -2118 -93 -2101
rect -167 -2169 -163 -2166
rect -159 -2166 -145 -2162
rect -159 -2169 -155 -2166
rect -131 -2169 -127 -2166
rect -123 -2166 -104 -2162
rect -123 -2169 -119 -2166
rect -97 -2169 -93 -2122
rect -71 -2133 -67 -2101
rect -71 -2162 -67 -2137
rect -37 -2155 -33 -2101
rect -37 -2159 -20 -2155
rect -89 -2169 -85 -2166
rect -80 -2166 -67 -2162
rect -80 -2169 -76 -2166
rect -53 -2169 -49 -2166
rect -29 -2169 -25 -2159
rect -13 -2162 -9 -2101
rect -5 -2155 -1 -2101
rect 21 -2125 25 -2101
rect -5 -2159 14 -2155
rect -21 -2166 -4 -2162
rect -21 -2169 -17 -2166
rect 3 -2169 7 -2159
rect 21 -2169 25 -2129
rect -210 -2177 -206 -2173
rect -184 -2177 -180 -2173
rect -141 -2177 -137 -2173
rect -106 -2177 -102 -2173
rect -62 -2177 -58 -2173
rect -45 -2177 -41 -2173
rect -9 -2177 -5 -2173
rect 12 -2177 16 -2173
rect 27 -2184 31 -2137
rect 191 -2140 195 -2023
rect 197 -2125 201 -1722
rect 203 -1795 207 -1296
rect 228 -1322 232 -1283
rect 228 -1337 232 -1326
rect 209 -1341 232 -1337
rect 235 -1313 239 -1276
rect 209 -1344 213 -1341
rect 235 -1344 239 -1317
rect 226 -1352 230 -1348
rect 218 -1382 222 -1378
rect 244 -1382 248 -1378
rect 261 -1382 265 -1378
rect 301 -1382 305 -1378
rect 322 -1382 326 -1378
rect 339 -1382 343 -1378
rect 379 -1382 383 -1378
rect 403 -1382 407 -1378
rect 440 -1382 444 -1378
rect 209 -1407 213 -1390
rect 209 -1458 213 -1411
rect 227 -1400 231 -1390
rect 227 -1458 231 -1404
rect 235 -1429 239 -1390
rect 253 -1422 257 -1390
rect 235 -1458 239 -1433
rect 253 -1458 257 -1426
rect 279 -1414 283 -1390
rect 279 -1451 283 -1418
rect 313 -1451 317 -1390
rect 331 -1407 335 -1390
rect 261 -1458 265 -1455
rect 269 -1455 283 -1451
rect 269 -1458 273 -1455
rect 297 -1458 301 -1455
rect 305 -1455 324 -1451
rect 305 -1458 309 -1455
rect 331 -1458 335 -1411
rect 357 -1422 361 -1390
rect 357 -1451 361 -1426
rect 391 -1444 395 -1390
rect 391 -1448 408 -1444
rect 339 -1458 343 -1455
rect 348 -1455 361 -1451
rect 348 -1458 352 -1455
rect 375 -1458 379 -1455
rect 399 -1458 403 -1448
rect 415 -1451 419 -1390
rect 423 -1444 427 -1390
rect 449 -1414 453 -1390
rect 423 -1448 442 -1444
rect 407 -1455 424 -1451
rect 407 -1458 411 -1455
rect 431 -1458 435 -1448
rect 449 -1458 453 -1418
rect 218 -1466 222 -1462
rect 244 -1466 248 -1462
rect 287 -1466 291 -1462
rect 322 -1466 326 -1462
rect 366 -1466 370 -1462
rect 383 -1466 387 -1462
rect 419 -1466 423 -1462
rect 440 -1466 444 -1462
rect 455 -1480 459 -1426
rect 547 -1429 551 -1317
rect 553 -1414 557 -1082
rect 559 -1292 563 -1066
rect 584 -1107 588 -1053
rect 565 -1111 584 -1107
rect 591 -1086 595 -1046
rect 957 -1062 961 -998
rect 963 -1038 967 -1034
rect 980 -1038 984 -1034
rect 971 -1049 975 -1046
rect 971 -1053 986 -1049
rect 957 -1066 964 -1062
rect 565 -1114 569 -1111
rect 591 -1114 595 -1090
rect 582 -1122 586 -1118
rect 574 -1152 578 -1148
rect 591 -1152 595 -1148
rect 611 -1152 615 -1148
rect 632 -1152 636 -1148
rect 653 -1152 657 -1148
rect 674 -1152 678 -1148
rect 695 -1152 699 -1148
rect 716 -1152 720 -1148
rect 737 -1152 741 -1148
rect 757 -1152 761 -1148
rect 565 -1207 569 -1160
rect 565 -1228 569 -1211
rect 583 -1221 587 -1160
rect 599 -1221 603 -1160
rect 623 -1200 627 -1160
rect 623 -1221 627 -1204
rect 641 -1221 645 -1160
rect 665 -1207 669 -1160
rect 665 -1221 669 -1211
rect 683 -1200 687 -1160
rect 683 -1221 687 -1204
rect 707 -1214 711 -1160
rect 725 -1192 729 -1160
rect 725 -1200 729 -1196
rect 707 -1221 711 -1218
rect 583 -1225 592 -1221
rect 599 -1225 607 -1221
rect 583 -1228 587 -1225
rect 607 -1228 611 -1225
rect 615 -1225 627 -1221
rect 641 -1225 649 -1221
rect 615 -1228 619 -1225
rect 649 -1228 653 -1225
rect 657 -1225 669 -1221
rect 683 -1225 695 -1221
rect 657 -1228 661 -1225
rect 691 -1228 695 -1225
rect 699 -1225 711 -1221
rect 725 -1221 729 -1204
rect 749 -1207 753 -1160
rect 749 -1221 753 -1211
rect 725 -1225 737 -1221
rect 699 -1228 703 -1225
rect 733 -1228 737 -1225
rect 741 -1225 753 -1221
rect 741 -1228 745 -1225
rect 574 -1236 578 -1232
rect 591 -1236 595 -1232
rect 632 -1236 636 -1232
rect 674 -1236 678 -1232
rect 716 -1236 720 -1232
rect 757 -1236 761 -1232
rect 565 -1268 569 -1264
rect 582 -1268 586 -1264
rect 573 -1279 577 -1276
rect 573 -1283 588 -1279
rect 559 -1296 566 -1292
rect 218 -1505 222 -1501
rect 235 -1505 239 -1501
rect 255 -1505 259 -1501
rect 276 -1505 280 -1501
rect 297 -1505 301 -1501
rect 318 -1505 322 -1501
rect 339 -1505 343 -1501
rect 360 -1505 364 -1501
rect 381 -1505 385 -1501
rect 401 -1505 405 -1501
rect 209 -1560 213 -1513
rect 209 -1581 213 -1564
rect 227 -1574 231 -1513
rect 243 -1574 247 -1513
rect 267 -1553 271 -1513
rect 267 -1574 271 -1557
rect 285 -1574 289 -1513
rect 309 -1560 313 -1513
rect 309 -1574 313 -1564
rect 327 -1553 331 -1513
rect 327 -1574 331 -1557
rect 351 -1567 355 -1513
rect 369 -1545 373 -1513
rect 369 -1553 373 -1549
rect 351 -1574 355 -1571
rect 227 -1578 236 -1574
rect 243 -1578 251 -1574
rect 227 -1581 231 -1578
rect 251 -1581 255 -1578
rect 259 -1578 271 -1574
rect 285 -1578 293 -1574
rect 259 -1581 263 -1578
rect 293 -1581 297 -1578
rect 301 -1578 313 -1574
rect 327 -1578 339 -1574
rect 301 -1581 305 -1578
rect 335 -1581 339 -1578
rect 343 -1578 355 -1574
rect 369 -1574 373 -1557
rect 393 -1560 397 -1513
rect 393 -1574 397 -1564
rect 369 -1578 381 -1574
rect 343 -1581 347 -1578
rect 377 -1581 381 -1578
rect 385 -1578 397 -1574
rect 385 -1581 389 -1578
rect 218 -1589 222 -1585
rect 235 -1589 239 -1585
rect 276 -1589 280 -1585
rect 318 -1589 322 -1585
rect 360 -1589 364 -1585
rect 401 -1589 405 -1585
rect 218 -1626 222 -1622
rect 235 -1626 239 -1622
rect 255 -1626 259 -1622
rect 276 -1626 280 -1622
rect 297 -1626 301 -1622
rect 318 -1626 322 -1622
rect 339 -1626 343 -1622
rect 360 -1626 364 -1622
rect 381 -1626 385 -1622
rect 401 -1626 405 -1622
rect 209 -1681 213 -1634
rect 209 -1702 213 -1685
rect 227 -1695 231 -1634
rect 243 -1695 247 -1634
rect 267 -1674 271 -1634
rect 267 -1695 271 -1678
rect 285 -1695 289 -1634
rect 309 -1681 313 -1634
rect 309 -1695 313 -1685
rect 327 -1674 331 -1634
rect 327 -1695 331 -1678
rect 351 -1688 355 -1634
rect 369 -1666 373 -1634
rect 369 -1674 373 -1670
rect 351 -1695 355 -1692
rect 227 -1699 236 -1695
rect 243 -1699 251 -1695
rect 227 -1702 231 -1699
rect 251 -1702 255 -1699
rect 259 -1699 271 -1695
rect 285 -1699 293 -1695
rect 259 -1702 263 -1699
rect 293 -1702 297 -1699
rect 301 -1699 313 -1695
rect 327 -1699 339 -1695
rect 301 -1702 305 -1699
rect 335 -1702 339 -1699
rect 343 -1699 355 -1695
rect 369 -1695 373 -1678
rect 393 -1681 397 -1634
rect 393 -1695 397 -1685
rect 369 -1699 381 -1695
rect 343 -1702 347 -1699
rect 377 -1702 381 -1699
rect 385 -1699 397 -1695
rect 385 -1702 389 -1699
rect 218 -1710 222 -1706
rect 235 -1710 239 -1706
rect 276 -1710 280 -1706
rect 318 -1710 322 -1706
rect 360 -1710 364 -1706
rect 401 -1710 405 -1706
rect 407 -1718 411 -1670
rect 553 -1674 557 -1484
rect 218 -1747 222 -1743
rect 235 -1747 239 -1743
rect 255 -1747 259 -1743
rect 276 -1747 280 -1743
rect 297 -1747 301 -1743
rect 318 -1747 322 -1743
rect 339 -1747 343 -1743
rect 360 -1747 364 -1743
rect 381 -1747 385 -1743
rect 401 -1747 405 -1743
rect 464 -1747 468 -1743
rect 209 -1802 213 -1755
rect 209 -1823 213 -1806
rect 227 -1816 231 -1755
rect 243 -1816 247 -1755
rect 267 -1795 271 -1755
rect 267 -1816 271 -1799
rect 285 -1816 289 -1755
rect 309 -1802 313 -1755
rect 309 -1816 313 -1806
rect 327 -1795 331 -1755
rect 327 -1816 331 -1799
rect 351 -1809 355 -1755
rect 369 -1787 373 -1755
rect 369 -1795 373 -1791
rect 351 -1816 355 -1813
rect 227 -1820 236 -1816
rect 243 -1820 251 -1816
rect 227 -1823 231 -1820
rect 251 -1823 255 -1820
rect 259 -1820 271 -1816
rect 285 -1820 293 -1816
rect 259 -1823 263 -1820
rect 293 -1823 297 -1820
rect 301 -1820 313 -1816
rect 327 -1820 339 -1816
rect 301 -1823 305 -1820
rect 335 -1823 339 -1820
rect 343 -1820 355 -1816
rect 369 -1816 373 -1799
rect 393 -1802 397 -1755
rect 393 -1816 397 -1806
rect 369 -1820 381 -1816
rect 343 -1823 347 -1820
rect 377 -1823 381 -1820
rect 385 -1820 397 -1816
rect 385 -1823 389 -1820
rect 218 -1831 222 -1827
rect 235 -1831 239 -1827
rect 276 -1831 280 -1827
rect 318 -1831 322 -1827
rect 360 -1831 364 -1827
rect 401 -1831 405 -1827
rect 209 -1974 213 -1970
rect 226 -1974 230 -1970
rect 217 -1985 221 -1982
rect 217 -1989 232 -1985
rect 203 -2002 210 -1998
rect -210 -2237 -206 -2233
rect -193 -2237 -189 -2233
rect -173 -2237 -169 -2233
rect -152 -2237 -148 -2233
rect -131 -2237 -127 -2233
rect -110 -2237 -106 -2233
rect -89 -2237 -85 -2233
rect -68 -2237 -64 -2233
rect -47 -2237 -43 -2233
rect -27 -2237 -23 -2233
rect -219 -2292 -215 -2245
rect -219 -2313 -215 -2296
rect -201 -2306 -197 -2245
rect -185 -2306 -181 -2245
rect -161 -2285 -157 -2245
rect -161 -2306 -157 -2289
rect -143 -2306 -139 -2245
rect -119 -2292 -115 -2245
rect -119 -2306 -115 -2296
rect -101 -2285 -97 -2245
rect -101 -2306 -97 -2289
rect -77 -2299 -73 -2245
rect -59 -2277 -55 -2245
rect -59 -2285 -55 -2281
rect -77 -2306 -73 -2303
rect -201 -2310 -192 -2306
rect -185 -2310 -177 -2306
rect -201 -2313 -197 -2310
rect -177 -2313 -173 -2310
rect -169 -2310 -157 -2306
rect -143 -2310 -135 -2306
rect -169 -2313 -165 -2310
rect -135 -2313 -131 -2310
rect -127 -2310 -115 -2306
rect -101 -2310 -89 -2306
rect -127 -2313 -123 -2310
rect -93 -2313 -89 -2310
rect -85 -2310 -73 -2306
rect -59 -2306 -55 -2289
rect -35 -2292 -31 -2245
rect -35 -2306 -31 -2296
rect -59 -2310 -47 -2306
rect -85 -2313 -81 -2310
rect -51 -2313 -47 -2310
rect -43 -2310 -31 -2306
rect -43 -2313 -39 -2310
rect -210 -2321 -206 -2317
rect -193 -2321 -189 -2317
rect -152 -2321 -148 -2317
rect -110 -2321 -106 -2317
rect -68 -2321 -64 -2317
rect -27 -2321 -23 -2317
rect -210 -2368 -206 -2364
rect -193 -2368 -189 -2364
rect -173 -2368 -169 -2364
rect -152 -2368 -148 -2364
rect -131 -2368 -127 -2364
rect -110 -2368 -106 -2364
rect -89 -2368 -85 -2364
rect -68 -2368 -64 -2364
rect -47 -2368 -43 -2364
rect -27 -2368 -23 -2364
rect -219 -2423 -215 -2376
rect -219 -2444 -215 -2427
rect -201 -2437 -197 -2376
rect -185 -2437 -181 -2376
rect -161 -2416 -157 -2376
rect -161 -2437 -157 -2420
rect -143 -2437 -139 -2376
rect -119 -2423 -115 -2376
rect -119 -2437 -115 -2427
rect -101 -2416 -97 -2376
rect -101 -2437 -97 -2420
rect -77 -2430 -73 -2376
rect -59 -2408 -55 -2376
rect -59 -2416 -55 -2412
rect -77 -2437 -73 -2434
rect -201 -2441 -192 -2437
rect -185 -2441 -177 -2437
rect -201 -2444 -197 -2441
rect -177 -2444 -173 -2441
rect -169 -2441 -157 -2437
rect -143 -2441 -135 -2437
rect -169 -2444 -165 -2441
rect -135 -2444 -131 -2441
rect -127 -2441 -115 -2437
rect -101 -2441 -89 -2437
rect -127 -2444 -123 -2441
rect -93 -2444 -89 -2441
rect -85 -2441 -73 -2437
rect -59 -2437 -55 -2420
rect -35 -2423 -31 -2376
rect -35 -2437 -31 -2427
rect -59 -2441 -47 -2437
rect -85 -2444 -81 -2441
rect -51 -2444 -47 -2441
rect -43 -2441 -31 -2437
rect -43 -2444 -39 -2441
rect -210 -2452 -206 -2448
rect -193 -2452 -189 -2448
rect -152 -2452 -148 -2448
rect -110 -2452 -106 -2448
rect -68 -2452 -64 -2448
rect -27 -2452 -23 -2448
rect -21 -2460 -17 -2412
rect 197 -2416 201 -2188
rect -210 -2499 -206 -2495
rect -193 -2499 -189 -2495
rect -173 -2499 -169 -2495
rect -152 -2499 -148 -2495
rect -131 -2499 -127 -2495
rect -110 -2499 -106 -2495
rect -89 -2499 -85 -2495
rect -68 -2499 -64 -2495
rect -47 -2499 -43 -2495
rect -27 -2499 -23 -2495
rect 90 -2499 94 -2495
rect -219 -2554 -215 -2507
rect -219 -2575 -215 -2558
rect -201 -2568 -197 -2507
rect -185 -2568 -181 -2507
rect -161 -2547 -157 -2507
rect -161 -2568 -157 -2551
rect -143 -2568 -139 -2507
rect -119 -2554 -115 -2507
rect -119 -2568 -115 -2558
rect -101 -2547 -97 -2507
rect -101 -2568 -97 -2551
rect -77 -2561 -73 -2507
rect -59 -2539 -55 -2507
rect -59 -2547 -55 -2543
rect -77 -2568 -73 -2565
rect -201 -2572 -192 -2568
rect -185 -2572 -177 -2568
rect -201 -2575 -197 -2572
rect -177 -2575 -173 -2572
rect -169 -2572 -157 -2568
rect -143 -2572 -135 -2568
rect -169 -2575 -165 -2572
rect -135 -2575 -131 -2572
rect -127 -2572 -115 -2568
rect -101 -2572 -89 -2568
rect -127 -2575 -123 -2572
rect -93 -2575 -89 -2572
rect -85 -2572 -73 -2568
rect -59 -2568 -55 -2551
rect -35 -2554 -31 -2507
rect -35 -2568 -31 -2558
rect -59 -2572 -47 -2568
rect -85 -2575 -81 -2572
rect -51 -2575 -47 -2572
rect -43 -2572 -31 -2568
rect -43 -2575 -39 -2572
rect -210 -2583 -206 -2579
rect -193 -2583 -189 -2579
rect -152 -2583 -148 -2579
rect -110 -2583 -106 -2579
rect -68 -2583 -64 -2579
rect -27 -2583 -23 -2579
rect -219 -2724 -215 -2720
rect -202 -2724 -198 -2720
rect -211 -2735 -207 -2732
rect -211 -2739 -196 -2735
rect -225 -2752 -218 -2748
rect -568 -2962 -564 -2958
rect -551 -2962 -547 -2958
rect -531 -2962 -527 -2958
rect -510 -2962 -506 -2958
rect -489 -2962 -485 -2958
rect -468 -2962 -464 -2958
rect -447 -2962 -443 -2958
rect -426 -2962 -422 -2958
rect -405 -2962 -401 -2958
rect -385 -2962 -381 -2958
rect -329 -2962 -325 -2958
rect -577 -3017 -573 -2970
rect -577 -3038 -573 -3021
rect -559 -3031 -555 -2970
rect -543 -3031 -539 -2970
rect -519 -3010 -515 -2970
rect -519 -3031 -515 -3014
rect -501 -3031 -497 -2970
rect -477 -3017 -473 -2970
rect -477 -3031 -473 -3021
rect -459 -3010 -455 -2970
rect -459 -3031 -455 -3014
rect -435 -3024 -431 -2970
rect -417 -2976 -413 -2970
rect -417 -3010 -413 -2980
rect -435 -3031 -431 -3028
rect -559 -3035 -550 -3031
rect -543 -3035 -535 -3031
rect -559 -3038 -555 -3035
rect -535 -3038 -531 -3035
rect -527 -3035 -515 -3031
rect -501 -3035 -493 -3031
rect -527 -3038 -523 -3035
rect -493 -3038 -489 -3035
rect -485 -3035 -473 -3031
rect -459 -3035 -447 -3031
rect -485 -3038 -481 -3035
rect -451 -3038 -447 -3035
rect -443 -3035 -431 -3031
rect -417 -3031 -413 -3014
rect -393 -3017 -389 -2970
rect -321 -3005 -317 -2970
rect -393 -3031 -389 -3021
rect -417 -3035 -405 -3031
rect -443 -3038 -439 -3035
rect -409 -3038 -405 -3035
rect -401 -3035 -389 -3031
rect -401 -3038 -397 -3035
rect -321 -3038 -317 -3009
rect -568 -3046 -564 -3042
rect -551 -3046 -547 -3042
rect -510 -3046 -506 -3042
rect -468 -3046 -464 -3042
rect -426 -3046 -422 -3042
rect -385 -3046 -381 -3042
rect -329 -3046 -325 -3042
rect -568 -3078 -564 -3074
rect -551 -3078 -547 -3074
rect -531 -3078 -527 -3074
rect -510 -3078 -506 -3074
rect -489 -3078 -485 -3074
rect -468 -3078 -464 -3074
rect -447 -3078 -443 -3074
rect -426 -3078 -422 -3074
rect -405 -3078 -401 -3074
rect -385 -3078 -381 -3074
rect -329 -3078 -325 -3074
rect -577 -3133 -573 -3086
rect -577 -3154 -573 -3137
rect -559 -3147 -555 -3086
rect -543 -3147 -539 -3086
rect -519 -3126 -515 -3086
rect -519 -3147 -515 -3130
rect -501 -3147 -497 -3086
rect -477 -3133 -473 -3086
rect -477 -3147 -473 -3137
rect -459 -3126 -455 -3086
rect -459 -3147 -455 -3130
rect -435 -3140 -431 -3086
rect -417 -3118 -413 -3086
rect -417 -3126 -413 -3122
rect -435 -3147 -431 -3144
rect -559 -3151 -550 -3147
rect -543 -3151 -535 -3147
rect -559 -3154 -555 -3151
rect -535 -3154 -531 -3151
rect -527 -3151 -515 -3147
rect -501 -3151 -493 -3147
rect -527 -3154 -523 -3151
rect -493 -3154 -489 -3151
rect -485 -3151 -473 -3147
rect -459 -3151 -447 -3147
rect -485 -3154 -481 -3151
rect -451 -3154 -447 -3151
rect -443 -3151 -431 -3147
rect -417 -3147 -413 -3130
rect -393 -3133 -389 -3086
rect -393 -3147 -389 -3137
rect -417 -3151 -405 -3147
rect -443 -3154 -439 -3151
rect -409 -3154 -405 -3151
rect -401 -3151 -389 -3147
rect -401 -3154 -397 -3151
rect -568 -3162 -564 -3158
rect -551 -3162 -547 -3158
rect -510 -3162 -506 -3158
rect -468 -3162 -464 -3158
rect -426 -3162 -422 -3158
rect -385 -3162 -381 -3158
rect -379 -3169 -375 -3122
rect -321 -3120 -317 -3086
rect -321 -3154 -317 -3124
rect -231 -3126 -227 -2945
rect -329 -3162 -325 -3158
rect -568 -3199 -564 -3195
rect -551 -3199 -547 -3195
rect -531 -3199 -527 -3195
rect -510 -3199 -506 -3195
rect -489 -3199 -485 -3195
rect -468 -3199 -464 -3195
rect -447 -3199 -443 -3195
rect -426 -3199 -422 -3195
rect -405 -3199 -401 -3195
rect -385 -3199 -381 -3195
rect -577 -3254 -573 -3207
rect -577 -3275 -573 -3258
rect -559 -3268 -555 -3207
rect -543 -3268 -539 -3207
rect -519 -3247 -515 -3207
rect -519 -3268 -515 -3251
rect -501 -3268 -497 -3207
rect -477 -3254 -473 -3207
rect -477 -3268 -473 -3258
rect -459 -3247 -455 -3207
rect -459 -3268 -455 -3251
rect -435 -3261 -431 -3207
rect -417 -3239 -413 -3207
rect -417 -3247 -413 -3243
rect -435 -3268 -431 -3265
rect -559 -3272 -550 -3268
rect -543 -3272 -535 -3268
rect -559 -3275 -555 -3272
rect -535 -3275 -531 -3272
rect -527 -3272 -515 -3268
rect -501 -3272 -493 -3268
rect -527 -3275 -523 -3272
rect -493 -3275 -489 -3272
rect -485 -3272 -473 -3268
rect -459 -3272 -447 -3268
rect -485 -3275 -481 -3272
rect -451 -3275 -447 -3272
rect -443 -3272 -431 -3268
rect -417 -3268 -413 -3251
rect -393 -3254 -389 -3207
rect -393 -3268 -389 -3258
rect -417 -3272 -405 -3268
rect -443 -3275 -439 -3272
rect -409 -3275 -405 -3272
rect -401 -3272 -389 -3268
rect -401 -3275 -397 -3272
rect -568 -3283 -564 -3279
rect -551 -3283 -547 -3279
rect -510 -3283 -506 -3279
rect -468 -3283 -464 -3279
rect -426 -3283 -422 -3279
rect -385 -3283 -381 -3279
rect -568 -3313 -564 -3309
rect -551 -3313 -547 -3309
rect -531 -3313 -527 -3309
rect -510 -3313 -506 -3309
rect -489 -3313 -485 -3309
rect -468 -3313 -464 -3309
rect -447 -3313 -443 -3309
rect -426 -3313 -422 -3309
rect -405 -3313 -401 -3309
rect -385 -3313 -381 -3309
rect -577 -3368 -573 -3321
rect -577 -3389 -573 -3372
rect -559 -3382 -555 -3321
rect -543 -3382 -539 -3321
rect -519 -3361 -515 -3321
rect -519 -3382 -515 -3365
rect -501 -3382 -497 -3321
rect -477 -3368 -473 -3321
rect -477 -3382 -473 -3372
rect -459 -3361 -455 -3321
rect -459 -3382 -455 -3365
rect -435 -3375 -431 -3321
rect -417 -3353 -413 -3321
rect -417 -3361 -413 -3357
rect -435 -3382 -431 -3379
rect -559 -3386 -550 -3382
rect -543 -3386 -535 -3382
rect -559 -3389 -555 -3386
rect -535 -3389 -531 -3386
rect -527 -3386 -515 -3382
rect -501 -3386 -493 -3382
rect -527 -3389 -523 -3386
rect -493 -3389 -489 -3386
rect -485 -3386 -473 -3382
rect -459 -3386 -447 -3382
rect -485 -3389 -481 -3386
rect -451 -3389 -447 -3386
rect -443 -3386 -431 -3382
rect -417 -3382 -413 -3365
rect -393 -3368 -389 -3321
rect -393 -3382 -389 -3372
rect -417 -3386 -405 -3382
rect -443 -3389 -439 -3386
rect -409 -3389 -405 -3386
rect -401 -3386 -389 -3382
rect -401 -3389 -397 -3386
rect -568 -3397 -564 -3393
rect -551 -3397 -547 -3393
rect -510 -3397 -506 -3393
rect -468 -3397 -464 -3393
rect -426 -3397 -422 -3393
rect -385 -3397 -381 -3393
rect -577 -3430 -573 -3426
rect -560 -3430 -556 -3426
rect -569 -3441 -565 -3438
rect -569 -3445 -554 -3441
rect -583 -3458 -576 -3454
rect -926 -3684 -922 -3680
rect -909 -3684 -905 -3680
rect -889 -3684 -885 -3680
rect -868 -3684 -864 -3680
rect -847 -3684 -843 -3680
rect -826 -3684 -822 -3680
rect -805 -3684 -801 -3680
rect -784 -3684 -780 -3680
rect -763 -3684 -759 -3680
rect -743 -3684 -739 -3680
rect -935 -3739 -931 -3692
rect -935 -3760 -931 -3743
rect -917 -3753 -913 -3692
rect -901 -3753 -897 -3692
rect -877 -3732 -873 -3692
rect -877 -3753 -873 -3736
rect -859 -3753 -855 -3692
rect -835 -3739 -831 -3692
rect -835 -3753 -831 -3743
rect -817 -3732 -813 -3692
rect -817 -3753 -813 -3736
rect -793 -3746 -789 -3692
rect -775 -3724 -771 -3692
rect -775 -3732 -771 -3728
rect -793 -3753 -789 -3750
rect -917 -3757 -908 -3753
rect -901 -3757 -893 -3753
rect -917 -3760 -913 -3757
rect -893 -3760 -889 -3757
rect -885 -3757 -873 -3753
rect -859 -3757 -851 -3753
rect -885 -3760 -881 -3757
rect -851 -3760 -847 -3757
rect -843 -3757 -831 -3753
rect -817 -3757 -805 -3753
rect -843 -3760 -839 -3757
rect -809 -3760 -805 -3757
rect -801 -3757 -789 -3753
rect -775 -3753 -771 -3736
rect -751 -3739 -747 -3692
rect -751 -3753 -747 -3743
rect -775 -3757 -763 -3753
rect -801 -3760 -797 -3757
rect -767 -3760 -763 -3757
rect -759 -3757 -747 -3753
rect -759 -3760 -755 -3757
rect -926 -3768 -922 -3764
rect -909 -3768 -905 -3764
rect -868 -3768 -864 -3764
rect -826 -3768 -822 -3764
rect -784 -3768 -780 -3764
rect -743 -3768 -739 -3764
rect -926 -3915 -922 -3911
rect -909 -3915 -905 -3911
rect -889 -3915 -885 -3911
rect -868 -3915 -864 -3911
rect -847 -3915 -843 -3911
rect -826 -3915 -822 -3911
rect -805 -3915 -801 -3911
rect -784 -3915 -780 -3911
rect -763 -3915 -759 -3911
rect -743 -3915 -739 -3911
rect -935 -3970 -931 -3923
rect -935 -3991 -931 -3974
rect -917 -3984 -913 -3923
rect -901 -3984 -897 -3923
rect -877 -3963 -873 -3923
rect -877 -3984 -873 -3967
rect -859 -3984 -855 -3923
rect -835 -3970 -831 -3923
rect -835 -3984 -831 -3974
rect -817 -3963 -813 -3923
rect -817 -3984 -813 -3967
rect -793 -3977 -789 -3923
rect -775 -3955 -771 -3923
rect -775 -3963 -771 -3959
rect -793 -3984 -789 -3981
rect -917 -3988 -908 -3984
rect -901 -3988 -893 -3984
rect -917 -3991 -913 -3988
rect -893 -3991 -889 -3988
rect -885 -3988 -873 -3984
rect -859 -3988 -851 -3984
rect -885 -3991 -881 -3988
rect -851 -3991 -847 -3988
rect -843 -3988 -831 -3984
rect -817 -3988 -805 -3984
rect -843 -3991 -839 -3988
rect -809 -3991 -805 -3988
rect -801 -3988 -789 -3984
rect -775 -3984 -771 -3967
rect -751 -3970 -747 -3923
rect -751 -3984 -747 -3974
rect -775 -3988 -763 -3984
rect -801 -3991 -797 -3988
rect -767 -3991 -763 -3988
rect -759 -3988 -747 -3984
rect -759 -3991 -755 -3988
rect -926 -3999 -922 -3995
rect -909 -3999 -905 -3995
rect -868 -3999 -864 -3995
rect -826 -3999 -822 -3995
rect -784 -3999 -780 -3995
rect -743 -3999 -739 -3995
rect -737 -4007 -733 -3959
rect -589 -3963 -585 -3649
rect -926 -4040 -922 -4036
rect -909 -4040 -905 -4036
rect -889 -4040 -885 -4036
rect -868 -4040 -864 -4036
rect -847 -4040 -843 -4036
rect -826 -4040 -822 -4036
rect -805 -4040 -801 -4036
rect -784 -4040 -780 -4036
rect -763 -4040 -759 -4036
rect -743 -4040 -739 -4036
rect -935 -4088 -931 -4048
rect -937 -4092 -931 -4088
rect -935 -4095 -931 -4092
rect -935 -4116 -931 -4099
rect -917 -4109 -913 -4048
rect -901 -4109 -897 -4048
rect -877 -4088 -873 -4048
rect -877 -4109 -873 -4092
rect -859 -4109 -855 -4048
rect -835 -4095 -831 -4048
rect -835 -4109 -831 -4099
rect -817 -4088 -813 -4048
rect -817 -4109 -813 -4092
rect -793 -4102 -789 -4048
rect -775 -4080 -771 -4048
rect -775 -4088 -771 -4084
rect -793 -4109 -789 -4106
rect -917 -4113 -908 -4109
rect -901 -4113 -893 -4109
rect -917 -4116 -913 -4113
rect -893 -4116 -889 -4113
rect -885 -4113 -873 -4109
rect -859 -4113 -851 -4109
rect -885 -4116 -881 -4113
rect -851 -4116 -847 -4113
rect -843 -4113 -831 -4109
rect -817 -4113 -805 -4109
rect -843 -4116 -839 -4113
rect -809 -4116 -805 -4113
rect -801 -4113 -789 -4109
rect -775 -4109 -771 -4092
rect -751 -4095 -747 -4048
rect -751 -4109 -747 -4099
rect -775 -4113 -763 -4109
rect -801 -4116 -797 -4113
rect -767 -4116 -763 -4113
rect -759 -4113 -747 -4109
rect -759 -4116 -755 -4113
rect -926 -4124 -922 -4120
rect -909 -4124 -905 -4120
rect -868 -4124 -864 -4120
rect -826 -4124 -822 -4120
rect -784 -4124 -780 -4120
rect -743 -4124 -739 -4120
rect -926 -4164 -922 -4160
rect -909 -4164 -905 -4160
rect -889 -4164 -885 -4160
rect -868 -4164 -864 -4160
rect -847 -4164 -843 -4160
rect -826 -4164 -822 -4160
rect -805 -4164 -801 -4160
rect -784 -4164 -780 -4160
rect -763 -4164 -759 -4160
rect -743 -4164 -739 -4160
rect -935 -4219 -931 -4172
rect -935 -4240 -931 -4223
rect -917 -4233 -913 -4172
rect -901 -4233 -897 -4172
rect -877 -4212 -873 -4172
rect -877 -4233 -873 -4216
rect -859 -4233 -855 -4172
rect -835 -4219 -831 -4172
rect -835 -4233 -831 -4223
rect -817 -4212 -813 -4172
rect -817 -4233 -813 -4216
rect -793 -4226 -789 -4172
rect -775 -4204 -771 -4172
rect -775 -4212 -771 -4208
rect -793 -4233 -789 -4230
rect -917 -4237 -908 -4233
rect -901 -4237 -893 -4233
rect -917 -4240 -913 -4237
rect -893 -4240 -889 -4237
rect -885 -4237 -873 -4233
rect -859 -4237 -851 -4233
rect -885 -4240 -881 -4237
rect -851 -4240 -847 -4237
rect -843 -4237 -831 -4233
rect -817 -4237 -805 -4233
rect -843 -4240 -839 -4237
rect -809 -4240 -805 -4237
rect -801 -4237 -789 -4233
rect -775 -4233 -771 -4216
rect -751 -4219 -747 -4172
rect -751 -4233 -747 -4223
rect -775 -4237 -763 -4233
rect -801 -4240 -797 -4237
rect -767 -4240 -763 -4237
rect -759 -4237 -747 -4233
rect -759 -4240 -755 -4237
rect -926 -4248 -922 -4244
rect -909 -4248 -905 -4244
rect -868 -4248 -864 -4244
rect -826 -4248 -822 -4244
rect -784 -4248 -780 -4244
rect -743 -4248 -739 -4244
rect -935 -4275 -931 -4271
rect -918 -4275 -914 -4271
rect -927 -4286 -923 -4283
rect -927 -4290 -912 -4286
rect -941 -4303 -934 -4299
rect -1255 -4478 -1251 -4474
rect -1211 -4478 -1207 -4474
rect -1177 -4478 -1173 -4474
rect -1276 -4686 -1272 -4489
rect -1162 -4492 -1158 -4460
rect -1270 -4565 -1266 -4496
rect -1255 -4517 -1251 -4513
rect -1238 -4517 -1234 -4513
rect -1218 -4517 -1214 -4513
rect -1197 -4517 -1193 -4513
rect -1176 -4517 -1172 -4513
rect -1155 -4517 -1151 -4513
rect -1134 -4517 -1130 -4513
rect -1113 -4517 -1109 -4513
rect -1092 -4517 -1088 -4513
rect -1072 -4517 -1068 -4513
rect -1264 -4572 -1260 -4525
rect -1264 -4593 -1260 -4576
rect -1246 -4586 -1242 -4525
rect -1230 -4586 -1226 -4525
rect -1206 -4565 -1202 -4525
rect -1206 -4586 -1202 -4569
rect -1188 -4586 -1184 -4525
rect -1164 -4572 -1160 -4525
rect -1164 -4586 -1160 -4576
rect -1146 -4565 -1142 -4525
rect -1146 -4586 -1142 -4569
rect -1122 -4579 -1118 -4525
rect -1104 -4557 -1100 -4525
rect -1104 -4565 -1100 -4561
rect -1122 -4586 -1118 -4583
rect -1246 -4590 -1237 -4586
rect -1230 -4590 -1222 -4586
rect -1246 -4593 -1242 -4590
rect -1222 -4593 -1218 -4590
rect -1214 -4590 -1202 -4586
rect -1188 -4590 -1180 -4586
rect -1214 -4593 -1210 -4590
rect -1180 -4593 -1176 -4590
rect -1172 -4590 -1160 -4586
rect -1146 -4590 -1134 -4586
rect -1172 -4593 -1168 -4590
rect -1138 -4593 -1134 -4590
rect -1130 -4590 -1118 -4586
rect -1104 -4586 -1100 -4569
rect -1080 -4572 -1076 -4525
rect -1080 -4586 -1076 -4576
rect -1104 -4590 -1092 -4586
rect -1130 -4593 -1126 -4590
rect -1096 -4593 -1092 -4590
rect -1088 -4590 -1076 -4586
rect -1088 -4593 -1084 -4590
rect -1255 -4601 -1251 -4597
rect -1238 -4601 -1234 -4597
rect -1197 -4601 -1193 -4597
rect -1155 -4601 -1151 -4597
rect -1113 -4601 -1109 -4597
rect -1072 -4601 -1068 -4597
rect -1255 -4638 -1251 -4634
rect -1238 -4638 -1234 -4634
rect -1218 -4638 -1214 -4634
rect -1197 -4638 -1193 -4634
rect -1176 -4638 -1172 -4634
rect -1155 -4638 -1151 -4634
rect -1134 -4638 -1130 -4634
rect -1113 -4638 -1109 -4634
rect -1092 -4638 -1088 -4634
rect -1072 -4638 -1068 -4634
rect -1264 -4693 -1260 -4646
rect -1264 -4714 -1260 -4697
rect -1246 -4707 -1242 -4646
rect -1230 -4707 -1226 -4646
rect -1206 -4686 -1202 -4646
rect -1206 -4707 -1202 -4690
rect -1188 -4707 -1184 -4646
rect -1164 -4693 -1160 -4646
rect -1164 -4707 -1160 -4697
rect -1146 -4686 -1142 -4646
rect -1146 -4707 -1142 -4690
rect -1122 -4700 -1118 -4646
rect -1104 -4678 -1100 -4646
rect -1104 -4686 -1100 -4682
rect -1122 -4707 -1118 -4704
rect -1246 -4711 -1237 -4707
rect -1230 -4711 -1222 -4707
rect -1246 -4714 -1242 -4711
rect -1222 -4714 -1218 -4711
rect -1214 -4711 -1202 -4707
rect -1188 -4711 -1180 -4707
rect -1214 -4714 -1210 -4711
rect -1180 -4714 -1176 -4711
rect -1172 -4711 -1160 -4707
rect -1146 -4711 -1134 -4707
rect -1172 -4714 -1168 -4711
rect -1138 -4714 -1134 -4711
rect -1130 -4711 -1118 -4707
rect -1104 -4707 -1100 -4690
rect -1080 -4693 -1076 -4646
rect -1080 -4707 -1076 -4697
rect -1104 -4711 -1092 -4707
rect -1130 -4714 -1126 -4711
rect -1096 -4714 -1092 -4711
rect -1088 -4711 -1076 -4707
rect -1088 -4714 -1084 -4711
rect -1255 -4722 -1251 -4718
rect -1238 -4722 -1234 -4718
rect -1197 -4722 -1193 -4718
rect -1155 -4722 -1151 -4718
rect -1113 -4722 -1109 -4718
rect -1072 -4722 -1068 -4718
rect -1066 -4730 -1062 -4682
rect -947 -4686 -943 -4496
rect -1339 -4994 -1335 -4990
rect -1322 -4994 -1318 -4990
rect -1331 -5005 -1327 -5002
rect -1331 -5009 -1316 -5005
rect -1349 -5022 -1338 -5018
rect -1349 -5521 -1345 -5022
rect -1320 -5048 -1316 -5009
rect -1320 -5063 -1316 -5052
rect -1339 -5067 -1316 -5063
rect -1339 -5070 -1335 -5067
rect -1313 -5070 -1309 -5002
rect -1322 -5078 -1318 -5074
rect -1313 -5168 -1309 -5074
rect -1270 -5161 -1266 -4734
rect -1255 -4759 -1251 -4755
rect -1238 -4759 -1234 -4755
rect -1218 -4759 -1214 -4755
rect -1197 -4759 -1193 -4755
rect -1176 -4759 -1172 -4755
rect -1155 -4759 -1151 -4755
rect -1134 -4759 -1130 -4755
rect -1113 -4759 -1109 -4755
rect -1092 -4759 -1088 -4755
rect -1072 -4759 -1068 -4755
rect -1264 -4814 -1260 -4767
rect -1264 -4835 -1260 -4818
rect -1246 -4828 -1242 -4767
rect -1230 -4828 -1226 -4767
rect -1206 -4807 -1202 -4767
rect -1206 -4828 -1202 -4811
rect -1188 -4828 -1184 -4767
rect -1164 -4814 -1160 -4767
rect -1164 -4828 -1160 -4818
rect -1146 -4807 -1142 -4767
rect -1146 -4828 -1142 -4811
rect -1122 -4821 -1118 -4767
rect -1104 -4799 -1100 -4767
rect -1104 -4807 -1100 -4803
rect -1122 -4828 -1118 -4825
rect -1246 -4832 -1237 -4828
rect -1230 -4832 -1222 -4828
rect -1246 -4835 -1242 -4832
rect -1222 -4835 -1218 -4832
rect -1214 -4832 -1202 -4828
rect -1188 -4832 -1180 -4828
rect -1214 -4835 -1210 -4832
rect -1180 -4835 -1176 -4832
rect -1172 -4832 -1160 -4828
rect -1146 -4832 -1134 -4828
rect -1172 -4835 -1168 -4832
rect -1138 -4835 -1134 -4832
rect -1130 -4832 -1118 -4828
rect -1104 -4828 -1100 -4811
rect -1080 -4814 -1076 -4767
rect -1080 -4828 -1076 -4818
rect -1104 -4832 -1092 -4828
rect -1130 -4835 -1126 -4832
rect -1096 -4835 -1092 -4832
rect -1088 -4832 -1076 -4828
rect -1088 -4835 -1084 -4832
rect -1255 -4843 -1251 -4839
rect -1238 -4843 -1234 -4839
rect -1197 -4843 -1193 -4839
rect -1155 -4843 -1151 -4839
rect -1113 -4843 -1109 -4839
rect -1072 -4843 -1068 -4839
rect -1255 -4877 -1251 -4873
rect -1238 -4877 -1234 -4873
rect -1218 -4877 -1214 -4873
rect -1197 -4877 -1193 -4873
rect -1176 -4877 -1172 -4873
rect -1155 -4877 -1151 -4873
rect -1134 -4877 -1130 -4873
rect -1113 -4877 -1109 -4873
rect -1092 -4877 -1088 -4873
rect -1072 -4877 -1068 -4873
rect -1264 -4932 -1260 -4885
rect -1264 -4953 -1260 -4936
rect -1246 -4946 -1242 -4885
rect -1230 -4946 -1226 -4885
rect -1206 -4925 -1202 -4885
rect -1206 -4946 -1202 -4929
rect -1188 -4946 -1184 -4885
rect -1164 -4932 -1160 -4885
rect -1164 -4946 -1160 -4936
rect -1146 -4925 -1142 -4885
rect -1146 -4946 -1142 -4929
rect -1122 -4939 -1118 -4885
rect -1104 -4917 -1100 -4885
rect -1104 -4925 -1100 -4921
rect -1122 -4946 -1118 -4943
rect -1246 -4950 -1237 -4946
rect -1230 -4950 -1222 -4946
rect -1246 -4953 -1242 -4950
rect -1222 -4953 -1218 -4950
rect -1214 -4950 -1202 -4946
rect -1188 -4950 -1180 -4946
rect -1214 -4953 -1210 -4950
rect -1180 -4953 -1176 -4950
rect -1172 -4950 -1160 -4946
rect -1146 -4950 -1134 -4946
rect -1172 -4953 -1168 -4950
rect -1138 -4953 -1134 -4950
rect -1130 -4950 -1118 -4946
rect -1104 -4946 -1100 -4929
rect -1080 -4932 -1076 -4885
rect -1080 -4946 -1076 -4936
rect -1104 -4950 -1092 -4946
rect -1130 -4953 -1126 -4950
rect -1096 -4953 -1092 -4950
rect -1088 -4950 -1076 -4946
rect -1088 -4953 -1084 -4950
rect -1255 -4961 -1251 -4957
rect -1238 -4961 -1234 -4957
rect -1197 -4961 -1193 -4957
rect -1155 -4961 -1151 -4957
rect -1113 -4961 -1109 -4957
rect -1072 -4961 -1068 -4957
rect -1066 -5018 -1062 -4803
rect -1255 -5113 -1251 -5109
rect -1238 -5113 -1234 -5109
rect -1198 -5113 -1194 -5109
rect -1177 -5113 -1173 -5109
rect -1264 -5154 -1260 -5121
rect -1264 -5189 -1260 -5158
rect -1246 -5148 -1242 -5121
rect -1246 -5152 -1237 -5148
rect -1246 -5189 -1242 -5152
rect -1220 -5175 -1216 -5121
rect -1220 -5182 -1216 -5179
rect -1186 -5182 -1182 -5121
rect -1168 -5153 -1164 -5121
rect -953 -5145 -949 -5043
rect -1238 -5189 -1234 -5186
rect -1229 -5186 -1216 -5182
rect -1229 -5189 -1225 -5186
rect -1202 -5189 -1198 -5186
rect -1194 -5186 -1175 -5182
rect -1194 -5189 -1190 -5186
rect -1168 -5189 -1164 -5157
rect -947 -5160 -943 -4733
rect -941 -4807 -937 -4303
rect -916 -4329 -912 -4290
rect -916 -4344 -912 -4333
rect -935 -4348 -912 -4344
rect -909 -4320 -905 -4283
rect -737 -4299 -733 -4084
rect -673 -4275 -669 -4271
rect -665 -4317 -661 -4291
rect -935 -4351 -931 -4348
rect -909 -4351 -905 -4324
rect -665 -4347 -661 -4321
rect -918 -4359 -914 -4355
rect -673 -4359 -669 -4355
rect -926 -4394 -922 -4390
rect -900 -4394 -896 -4390
rect -883 -4394 -879 -4390
rect -843 -4394 -839 -4390
rect -822 -4394 -818 -4390
rect -805 -4394 -801 -4390
rect -765 -4394 -761 -4390
rect -741 -4394 -737 -4390
rect -704 -4394 -700 -4390
rect -935 -4419 -931 -4402
rect -935 -4470 -931 -4423
rect -917 -4412 -913 -4402
rect -917 -4470 -913 -4416
rect -909 -4441 -905 -4402
rect -891 -4434 -887 -4402
rect -909 -4470 -905 -4445
rect -891 -4470 -887 -4438
rect -865 -4426 -861 -4402
rect -865 -4463 -861 -4430
rect -831 -4463 -827 -4402
rect -813 -4419 -809 -4402
rect -883 -4470 -879 -4467
rect -875 -4467 -861 -4463
rect -875 -4470 -871 -4467
rect -847 -4470 -843 -4467
rect -839 -4467 -820 -4463
rect -839 -4470 -835 -4467
rect -813 -4470 -809 -4423
rect -787 -4434 -783 -4402
rect -787 -4463 -783 -4438
rect -753 -4456 -749 -4402
rect -753 -4460 -736 -4456
rect -805 -4470 -801 -4467
rect -796 -4467 -783 -4463
rect -796 -4470 -792 -4467
rect -769 -4470 -765 -4467
rect -745 -4470 -741 -4460
rect -729 -4463 -725 -4402
rect -721 -4456 -717 -4402
rect -695 -4426 -691 -4402
rect -721 -4460 -702 -4456
rect -737 -4467 -720 -4463
rect -737 -4470 -733 -4467
rect -713 -4470 -709 -4460
rect -695 -4470 -691 -4430
rect -926 -4478 -922 -4474
rect -900 -4478 -896 -4474
rect -857 -4478 -853 -4474
rect -822 -4478 -818 -4474
rect -778 -4478 -774 -4474
rect -761 -4478 -757 -4474
rect -725 -4478 -721 -4474
rect -704 -4478 -700 -4474
rect -689 -4485 -685 -4438
rect -595 -4441 -591 -4324
rect -589 -4426 -585 -4010
rect -583 -4088 -579 -3458
rect -558 -3484 -554 -3445
rect -558 -3499 -554 -3488
rect -577 -3503 -554 -3499
rect -551 -3475 -547 -3438
rect -379 -3462 -375 -3357
rect -373 -3454 -369 -3243
rect -577 -3506 -573 -3503
rect -551 -3506 -547 -3479
rect -560 -3514 -556 -3510
rect -568 -3554 -564 -3550
rect -542 -3554 -538 -3550
rect -525 -3554 -521 -3550
rect -485 -3554 -481 -3550
rect -464 -3554 -460 -3550
rect -447 -3554 -443 -3550
rect -407 -3554 -403 -3550
rect -383 -3554 -379 -3550
rect -346 -3554 -342 -3550
rect -577 -3579 -573 -3562
rect -577 -3630 -573 -3583
rect -559 -3572 -555 -3562
rect -559 -3630 -555 -3576
rect -551 -3601 -547 -3562
rect -533 -3594 -529 -3562
rect -551 -3630 -547 -3605
rect -533 -3630 -529 -3598
rect -507 -3586 -503 -3562
rect -507 -3623 -503 -3590
rect -473 -3623 -469 -3562
rect -455 -3579 -451 -3562
rect -525 -3630 -521 -3627
rect -517 -3627 -503 -3623
rect -517 -3630 -513 -3627
rect -489 -3630 -485 -3627
rect -481 -3627 -462 -3623
rect -481 -3630 -477 -3627
rect -455 -3630 -451 -3583
rect -429 -3594 -425 -3562
rect -429 -3623 -425 -3598
rect -395 -3616 -391 -3562
rect -395 -3620 -378 -3616
rect -447 -3630 -443 -3627
rect -438 -3627 -425 -3623
rect -438 -3630 -434 -3627
rect -411 -3630 -407 -3627
rect -387 -3630 -383 -3620
rect -371 -3623 -367 -3562
rect -363 -3616 -359 -3562
rect -337 -3585 -333 -3562
rect -363 -3620 -344 -3616
rect -379 -3627 -362 -3623
rect -379 -3630 -375 -3627
rect -355 -3630 -351 -3620
rect -337 -3630 -333 -3589
rect -568 -3638 -564 -3634
rect -542 -3638 -538 -3634
rect -499 -3638 -495 -3634
rect -464 -3638 -460 -3634
rect -420 -3638 -416 -3634
rect -403 -3638 -399 -3634
rect -367 -3638 -363 -3634
rect -346 -3638 -342 -3634
rect -331 -3652 -327 -3598
rect -237 -3601 -233 -3479
rect -231 -3586 -227 -3174
rect -225 -3247 -221 -2752
rect -200 -2778 -196 -2739
rect -200 -2793 -196 -2782
rect -219 -2797 -196 -2793
rect -193 -2769 -189 -2732
rect -21 -2748 -17 -2543
rect 98 -2542 102 -2531
rect 98 -2563 102 -2546
rect 90 -2583 94 -2579
rect -219 -2800 -215 -2797
rect -193 -2800 -189 -2773
rect -202 -2808 -198 -2804
rect -210 -2843 -206 -2839
rect -184 -2843 -180 -2839
rect -167 -2843 -163 -2839
rect -127 -2843 -123 -2839
rect -106 -2843 -102 -2839
rect -89 -2843 -85 -2839
rect -49 -2843 -45 -2839
rect -25 -2843 -21 -2839
rect 12 -2843 16 -2839
rect -219 -2868 -215 -2851
rect -219 -2919 -215 -2872
rect -201 -2861 -197 -2851
rect -201 -2919 -197 -2865
rect -193 -2890 -189 -2851
rect -175 -2883 -171 -2851
rect -193 -2919 -189 -2894
rect -175 -2919 -171 -2887
rect -149 -2875 -145 -2851
rect -149 -2912 -145 -2879
rect -115 -2912 -111 -2851
rect -97 -2868 -93 -2851
rect -167 -2919 -163 -2916
rect -159 -2916 -145 -2912
rect -159 -2919 -155 -2916
rect -131 -2919 -127 -2916
rect -123 -2916 -104 -2912
rect -123 -2919 -119 -2916
rect -97 -2919 -93 -2872
rect -71 -2883 -67 -2851
rect -71 -2912 -67 -2887
rect -37 -2905 -33 -2851
rect -37 -2909 -20 -2905
rect -89 -2919 -85 -2916
rect -80 -2916 -67 -2912
rect -80 -2919 -76 -2916
rect -53 -2919 -49 -2916
rect -29 -2919 -25 -2909
rect -13 -2912 -9 -2851
rect -5 -2905 -1 -2851
rect 21 -2875 25 -2851
rect -5 -2909 14 -2905
rect -21 -2916 -4 -2912
rect -21 -2919 -17 -2916
rect 3 -2919 7 -2909
rect 21 -2919 25 -2879
rect -210 -2927 -206 -2923
rect -184 -2927 -180 -2923
rect -141 -2927 -137 -2923
rect -106 -2927 -102 -2923
rect -62 -2927 -58 -2923
rect -45 -2927 -41 -2923
rect -9 -2927 -5 -2923
rect 12 -2927 16 -2923
rect 27 -2934 31 -2887
rect 191 -2890 195 -2773
rect 197 -2875 201 -2463
rect 203 -2547 207 -2002
rect 228 -2028 232 -1989
rect 228 -2043 232 -2032
rect 209 -2047 232 -2043
rect 235 -2019 239 -1982
rect 407 -1998 411 -1791
rect 472 -1788 476 -1755
rect 472 -1823 476 -1792
rect 464 -1831 468 -1827
rect 464 -1862 468 -1858
rect 472 -1903 476 -1870
rect 472 -1938 476 -1907
rect 464 -1946 468 -1942
rect 209 -2050 213 -2047
rect 235 -2050 239 -2023
rect 226 -2058 230 -2054
rect 218 -2093 222 -2089
rect 244 -2093 248 -2089
rect 261 -2093 265 -2089
rect 301 -2093 305 -2089
rect 322 -2093 326 -2089
rect 339 -2093 343 -2089
rect 379 -2093 383 -2089
rect 403 -2093 407 -2089
rect 440 -2093 444 -2089
rect 209 -2118 213 -2101
rect 209 -2169 213 -2122
rect 227 -2111 231 -2101
rect 227 -2169 231 -2115
rect 235 -2140 239 -2101
rect 253 -2133 257 -2101
rect 235 -2169 239 -2144
rect 253 -2169 257 -2137
rect 279 -2125 283 -2101
rect 279 -2162 283 -2129
rect 313 -2162 317 -2101
rect 331 -2118 335 -2101
rect 261 -2169 265 -2166
rect 269 -2166 283 -2162
rect 269 -2169 273 -2166
rect 297 -2169 301 -2166
rect 305 -2166 324 -2162
rect 305 -2169 309 -2166
rect 331 -2169 335 -2122
rect 357 -2133 361 -2101
rect 357 -2162 361 -2137
rect 391 -2155 395 -2101
rect 391 -2159 408 -2155
rect 339 -2169 343 -2166
rect 348 -2166 361 -2162
rect 348 -2169 352 -2166
rect 375 -2169 379 -2166
rect 399 -2169 403 -2159
rect 415 -2162 419 -2101
rect 423 -2155 427 -2101
rect 449 -2125 453 -2101
rect 423 -2159 442 -2155
rect 407 -2166 424 -2162
rect 407 -2169 411 -2166
rect 431 -2169 435 -2159
rect 449 -2169 453 -2129
rect 218 -2177 222 -2173
rect 244 -2177 248 -2173
rect 287 -2177 291 -2173
rect 322 -2177 326 -2173
rect 366 -2177 370 -2173
rect 383 -2177 387 -2173
rect 419 -2177 423 -2173
rect 440 -2177 444 -2173
rect 455 -2191 459 -2137
rect 547 -2140 551 -2023
rect 553 -2125 557 -1721
rect 559 -1795 563 -1296
rect 584 -1322 588 -1283
rect 584 -1337 588 -1326
rect 565 -1341 588 -1337
rect 591 -1313 595 -1276
rect 565 -1344 569 -1341
rect 591 -1344 595 -1317
rect 582 -1352 586 -1348
rect 574 -1382 578 -1378
rect 600 -1382 604 -1378
rect 617 -1382 621 -1378
rect 657 -1382 661 -1378
rect 678 -1382 682 -1378
rect 695 -1382 699 -1378
rect 735 -1382 739 -1378
rect 759 -1382 763 -1378
rect 796 -1382 800 -1378
rect 565 -1407 569 -1390
rect 565 -1458 569 -1411
rect 583 -1400 587 -1390
rect 583 -1458 587 -1404
rect 591 -1429 595 -1390
rect 609 -1422 613 -1390
rect 591 -1458 595 -1433
rect 609 -1458 613 -1426
rect 635 -1414 639 -1390
rect 635 -1451 639 -1418
rect 669 -1451 673 -1390
rect 687 -1407 691 -1390
rect 617 -1458 621 -1455
rect 625 -1455 639 -1451
rect 625 -1458 629 -1455
rect 653 -1458 657 -1455
rect 661 -1455 680 -1451
rect 661 -1458 665 -1455
rect 687 -1458 691 -1411
rect 713 -1422 717 -1390
rect 713 -1451 717 -1426
rect 747 -1444 751 -1390
rect 747 -1448 764 -1444
rect 695 -1458 699 -1455
rect 704 -1455 717 -1451
rect 704 -1458 708 -1455
rect 731 -1458 735 -1455
rect 755 -1458 759 -1448
rect 771 -1451 775 -1390
rect 779 -1444 783 -1390
rect 805 -1414 809 -1390
rect 779 -1448 798 -1444
rect 763 -1455 780 -1451
rect 763 -1458 767 -1455
rect 787 -1458 791 -1448
rect 805 -1458 809 -1418
rect 574 -1466 578 -1462
rect 600 -1466 604 -1462
rect 643 -1466 647 -1462
rect 678 -1466 682 -1462
rect 722 -1466 726 -1462
rect 739 -1466 743 -1462
rect 775 -1466 779 -1462
rect 796 -1466 800 -1462
rect 811 -1487 815 -1426
rect 945 -1429 949 -1317
rect 951 -1414 955 -1090
rect 957 -1292 961 -1066
rect 982 -1107 986 -1053
rect 963 -1111 982 -1107
rect 989 -1078 993 -1046
rect 963 -1114 967 -1111
rect 989 -1114 993 -1082
rect 1315 -1062 1319 -998
rect 1321 -1038 1325 -1034
rect 1338 -1038 1342 -1034
rect 1329 -1049 1333 -1046
rect 1329 -1053 1344 -1049
rect 1315 -1066 1322 -1062
rect 980 -1122 984 -1118
rect 972 -1152 976 -1148
rect 989 -1152 993 -1148
rect 1009 -1152 1013 -1148
rect 1030 -1152 1034 -1148
rect 1051 -1152 1055 -1148
rect 1072 -1152 1076 -1148
rect 1093 -1152 1097 -1148
rect 1114 -1152 1118 -1148
rect 1135 -1152 1139 -1148
rect 1155 -1152 1159 -1148
rect 963 -1207 967 -1160
rect 963 -1228 967 -1211
rect 981 -1221 985 -1160
rect 997 -1221 1001 -1160
rect 1021 -1200 1025 -1160
rect 1021 -1221 1025 -1204
rect 1039 -1221 1043 -1160
rect 1063 -1207 1067 -1160
rect 1063 -1221 1067 -1211
rect 1081 -1200 1085 -1160
rect 1081 -1221 1085 -1204
rect 1105 -1214 1109 -1160
rect 1123 -1192 1127 -1160
rect 1123 -1200 1127 -1196
rect 1105 -1221 1109 -1218
rect 981 -1225 990 -1221
rect 997 -1225 1005 -1221
rect 981 -1228 985 -1225
rect 1005 -1228 1009 -1225
rect 1013 -1225 1025 -1221
rect 1039 -1225 1047 -1221
rect 1013 -1228 1017 -1225
rect 1047 -1228 1051 -1225
rect 1055 -1225 1067 -1221
rect 1081 -1225 1093 -1221
rect 1055 -1228 1059 -1225
rect 1089 -1228 1093 -1225
rect 1097 -1225 1109 -1221
rect 1123 -1221 1127 -1204
rect 1147 -1207 1151 -1160
rect 1147 -1221 1151 -1211
rect 1123 -1225 1135 -1221
rect 1097 -1228 1101 -1225
rect 1131 -1228 1135 -1225
rect 1139 -1225 1151 -1221
rect 1139 -1228 1143 -1225
rect 972 -1236 976 -1232
rect 989 -1236 993 -1232
rect 1030 -1236 1034 -1232
rect 1072 -1236 1076 -1232
rect 1114 -1236 1118 -1232
rect 1155 -1236 1159 -1232
rect 963 -1268 967 -1264
rect 980 -1268 984 -1264
rect 971 -1279 975 -1276
rect 971 -1283 986 -1279
rect 957 -1296 964 -1292
rect 574 -1505 578 -1501
rect 591 -1505 595 -1501
rect 611 -1505 615 -1501
rect 632 -1505 636 -1501
rect 653 -1505 657 -1501
rect 674 -1505 678 -1501
rect 695 -1505 699 -1501
rect 716 -1505 720 -1501
rect 737 -1505 741 -1501
rect 757 -1505 761 -1501
rect 565 -1560 569 -1513
rect 565 -1581 569 -1564
rect 583 -1574 587 -1513
rect 599 -1574 603 -1513
rect 623 -1553 627 -1513
rect 623 -1574 627 -1557
rect 641 -1574 645 -1513
rect 665 -1560 669 -1513
rect 665 -1574 669 -1564
rect 683 -1553 687 -1513
rect 683 -1574 687 -1557
rect 707 -1567 711 -1513
rect 725 -1545 729 -1513
rect 725 -1553 729 -1549
rect 707 -1574 711 -1571
rect 583 -1578 592 -1574
rect 599 -1578 607 -1574
rect 583 -1581 587 -1578
rect 607 -1581 611 -1578
rect 615 -1578 627 -1574
rect 641 -1578 649 -1574
rect 615 -1581 619 -1578
rect 649 -1581 653 -1578
rect 657 -1578 669 -1574
rect 683 -1578 695 -1574
rect 657 -1581 661 -1578
rect 691 -1581 695 -1578
rect 699 -1578 711 -1574
rect 725 -1574 729 -1557
rect 749 -1560 753 -1513
rect 749 -1574 753 -1564
rect 725 -1578 737 -1574
rect 699 -1581 703 -1578
rect 733 -1581 737 -1578
rect 741 -1578 753 -1574
rect 741 -1581 745 -1578
rect 574 -1589 578 -1585
rect 591 -1589 595 -1585
rect 632 -1589 636 -1585
rect 674 -1589 678 -1585
rect 716 -1589 720 -1585
rect 757 -1589 761 -1585
rect 574 -1626 578 -1622
rect 591 -1626 595 -1622
rect 611 -1626 615 -1622
rect 632 -1626 636 -1622
rect 653 -1626 657 -1622
rect 674 -1626 678 -1622
rect 695 -1626 699 -1622
rect 716 -1626 720 -1622
rect 737 -1626 741 -1622
rect 757 -1626 761 -1622
rect 565 -1681 569 -1634
rect 565 -1702 569 -1685
rect 583 -1695 587 -1634
rect 599 -1695 603 -1634
rect 623 -1674 627 -1634
rect 623 -1695 627 -1678
rect 641 -1695 645 -1634
rect 665 -1681 669 -1634
rect 665 -1695 669 -1685
rect 683 -1674 687 -1634
rect 683 -1695 687 -1678
rect 707 -1688 711 -1634
rect 725 -1666 729 -1634
rect 725 -1674 729 -1670
rect 707 -1695 711 -1692
rect 583 -1699 592 -1695
rect 599 -1699 607 -1695
rect 583 -1702 587 -1699
rect 607 -1702 611 -1699
rect 615 -1699 627 -1695
rect 641 -1699 649 -1695
rect 615 -1702 619 -1699
rect 649 -1702 653 -1699
rect 657 -1699 669 -1695
rect 683 -1699 695 -1695
rect 657 -1702 661 -1699
rect 691 -1702 695 -1699
rect 699 -1699 711 -1695
rect 725 -1695 729 -1678
rect 749 -1681 753 -1634
rect 749 -1695 753 -1685
rect 725 -1699 737 -1695
rect 699 -1702 703 -1699
rect 733 -1702 737 -1699
rect 741 -1699 753 -1695
rect 741 -1702 745 -1699
rect 574 -1710 578 -1706
rect 591 -1710 595 -1706
rect 632 -1710 636 -1706
rect 674 -1710 678 -1706
rect 716 -1710 720 -1706
rect 757 -1710 761 -1706
rect 763 -1717 767 -1670
rect 951 -1674 955 -1491
rect 574 -1747 578 -1743
rect 591 -1747 595 -1743
rect 611 -1747 615 -1743
rect 632 -1747 636 -1743
rect 653 -1747 657 -1743
rect 674 -1747 678 -1743
rect 695 -1747 699 -1743
rect 716 -1747 720 -1743
rect 737 -1747 741 -1743
rect 757 -1747 761 -1743
rect 565 -1802 569 -1755
rect 565 -1823 569 -1806
rect 583 -1816 587 -1755
rect 599 -1816 603 -1755
rect 623 -1795 627 -1755
rect 623 -1816 627 -1799
rect 641 -1816 645 -1755
rect 665 -1802 669 -1755
rect 665 -1816 669 -1806
rect 683 -1795 687 -1755
rect 683 -1816 687 -1799
rect 707 -1809 711 -1755
rect 725 -1787 729 -1755
rect 725 -1795 729 -1791
rect 707 -1816 711 -1813
rect 583 -1820 592 -1816
rect 599 -1820 607 -1816
rect 583 -1823 587 -1820
rect 607 -1823 611 -1820
rect 615 -1820 627 -1816
rect 641 -1820 649 -1816
rect 615 -1823 619 -1820
rect 649 -1823 653 -1820
rect 657 -1820 669 -1816
rect 683 -1820 695 -1816
rect 657 -1823 661 -1820
rect 691 -1823 695 -1820
rect 699 -1820 711 -1816
rect 725 -1816 729 -1799
rect 749 -1802 753 -1755
rect 749 -1816 753 -1806
rect 725 -1820 737 -1816
rect 699 -1823 703 -1820
rect 733 -1823 737 -1820
rect 741 -1820 753 -1816
rect 741 -1823 745 -1820
rect 574 -1831 578 -1827
rect 591 -1831 595 -1827
rect 632 -1831 636 -1827
rect 674 -1831 678 -1827
rect 716 -1831 720 -1827
rect 757 -1831 761 -1827
rect 565 -1974 569 -1970
rect 582 -1974 586 -1970
rect 573 -1985 577 -1982
rect 573 -1989 588 -1985
rect 559 -2002 566 -1998
rect 218 -2237 222 -2233
rect 235 -2237 239 -2233
rect 255 -2237 259 -2233
rect 276 -2237 280 -2233
rect 297 -2237 301 -2233
rect 318 -2237 322 -2233
rect 339 -2237 343 -2233
rect 360 -2237 364 -2233
rect 381 -2237 385 -2233
rect 401 -2237 405 -2233
rect 209 -2292 213 -2245
rect 209 -2313 213 -2296
rect 227 -2306 231 -2245
rect 243 -2306 247 -2245
rect 267 -2285 271 -2245
rect 267 -2306 271 -2289
rect 285 -2306 289 -2245
rect 309 -2292 313 -2245
rect 309 -2306 313 -2296
rect 327 -2285 331 -2245
rect 327 -2306 331 -2289
rect 351 -2299 355 -2245
rect 369 -2277 373 -2245
rect 369 -2285 373 -2281
rect 351 -2306 355 -2303
rect 227 -2310 236 -2306
rect 243 -2310 251 -2306
rect 227 -2313 231 -2310
rect 251 -2313 255 -2310
rect 259 -2310 271 -2306
rect 285 -2310 293 -2306
rect 259 -2313 263 -2310
rect 293 -2313 297 -2310
rect 301 -2310 313 -2306
rect 327 -2310 339 -2306
rect 301 -2313 305 -2310
rect 335 -2313 339 -2310
rect 343 -2310 355 -2306
rect 369 -2306 373 -2289
rect 393 -2292 397 -2245
rect 393 -2306 397 -2296
rect 369 -2310 381 -2306
rect 343 -2313 347 -2310
rect 377 -2313 381 -2310
rect 385 -2310 397 -2306
rect 385 -2313 389 -2310
rect 218 -2321 222 -2317
rect 235 -2321 239 -2317
rect 276 -2321 280 -2317
rect 318 -2321 322 -2317
rect 360 -2321 364 -2317
rect 401 -2321 405 -2317
rect 218 -2368 222 -2364
rect 235 -2368 239 -2364
rect 255 -2368 259 -2364
rect 276 -2368 280 -2364
rect 297 -2368 301 -2364
rect 318 -2368 322 -2364
rect 339 -2368 343 -2364
rect 360 -2368 364 -2364
rect 381 -2368 385 -2364
rect 401 -2368 405 -2364
rect 209 -2423 213 -2376
rect 209 -2444 213 -2427
rect 227 -2437 231 -2376
rect 243 -2437 247 -2376
rect 267 -2416 271 -2376
rect 267 -2437 271 -2420
rect 285 -2437 289 -2376
rect 309 -2423 313 -2376
rect 309 -2437 313 -2427
rect 327 -2416 331 -2376
rect 327 -2437 331 -2420
rect 351 -2430 355 -2376
rect 369 -2408 373 -2376
rect 369 -2416 373 -2412
rect 351 -2437 355 -2434
rect 227 -2441 236 -2437
rect 243 -2441 251 -2437
rect 227 -2444 231 -2441
rect 251 -2444 255 -2441
rect 259 -2441 271 -2437
rect 285 -2441 293 -2437
rect 259 -2444 263 -2441
rect 293 -2444 297 -2441
rect 301 -2441 313 -2437
rect 327 -2441 339 -2437
rect 301 -2444 305 -2441
rect 335 -2444 339 -2441
rect 343 -2441 355 -2437
rect 369 -2437 373 -2420
rect 393 -2423 397 -2376
rect 393 -2437 397 -2427
rect 369 -2441 381 -2437
rect 343 -2444 347 -2441
rect 377 -2444 381 -2441
rect 385 -2441 397 -2437
rect 385 -2444 389 -2441
rect 218 -2452 222 -2448
rect 235 -2452 239 -2448
rect 276 -2452 280 -2448
rect 318 -2452 322 -2448
rect 360 -2452 364 -2448
rect 401 -2452 405 -2448
rect 407 -2459 411 -2412
rect 553 -2416 557 -2195
rect 218 -2499 222 -2495
rect 235 -2499 239 -2495
rect 255 -2499 259 -2495
rect 276 -2499 280 -2495
rect 297 -2499 301 -2495
rect 318 -2499 322 -2495
rect 339 -2499 343 -2495
rect 360 -2499 364 -2495
rect 381 -2499 385 -2495
rect 401 -2499 405 -2495
rect 209 -2554 213 -2507
rect 209 -2575 213 -2558
rect 227 -2568 231 -2507
rect 243 -2568 247 -2507
rect 267 -2547 271 -2507
rect 267 -2568 271 -2551
rect 285 -2568 289 -2507
rect 309 -2554 313 -2507
rect 309 -2568 313 -2558
rect 327 -2547 331 -2507
rect 327 -2568 331 -2551
rect 351 -2561 355 -2507
rect 369 -2539 373 -2507
rect 369 -2547 373 -2543
rect 351 -2568 355 -2565
rect 227 -2572 236 -2568
rect 243 -2572 251 -2568
rect 227 -2575 231 -2572
rect 251 -2575 255 -2572
rect 259 -2572 271 -2568
rect 285 -2572 293 -2568
rect 259 -2575 263 -2572
rect 293 -2575 297 -2572
rect 301 -2572 313 -2568
rect 327 -2572 339 -2568
rect 301 -2575 305 -2572
rect 335 -2575 339 -2572
rect 343 -2572 355 -2568
rect 369 -2568 373 -2551
rect 393 -2554 397 -2507
rect 393 -2568 397 -2558
rect 369 -2572 381 -2568
rect 343 -2575 347 -2572
rect 377 -2575 381 -2572
rect 385 -2572 397 -2568
rect 385 -2575 389 -2572
rect 218 -2583 222 -2579
rect 235 -2583 239 -2579
rect 276 -2583 280 -2579
rect 318 -2583 322 -2579
rect 360 -2583 364 -2579
rect 401 -2583 405 -2579
rect 209 -2724 213 -2720
rect 226 -2724 230 -2720
rect 217 -2735 221 -2732
rect 217 -2739 232 -2735
rect 203 -2752 210 -2748
rect -210 -2962 -206 -2958
rect -193 -2962 -189 -2958
rect -173 -2962 -169 -2958
rect -152 -2962 -148 -2958
rect -131 -2962 -127 -2958
rect -110 -2962 -106 -2958
rect -89 -2962 -85 -2958
rect -68 -2962 -64 -2958
rect -47 -2962 -43 -2958
rect -27 -2962 -23 -2958
rect -219 -3017 -215 -2970
rect -219 -3038 -215 -3021
rect -201 -3031 -197 -2970
rect -185 -3031 -181 -2970
rect -161 -3010 -157 -2970
rect -161 -3031 -157 -3014
rect -143 -3031 -139 -2970
rect -119 -3017 -115 -2970
rect -119 -3031 -115 -3021
rect -101 -3010 -97 -2970
rect -101 -3031 -97 -3014
rect -77 -3024 -73 -2970
rect -59 -3002 -55 -2970
rect -59 -3010 -55 -3006
rect -77 -3031 -73 -3028
rect -201 -3035 -192 -3031
rect -185 -3035 -177 -3031
rect -201 -3038 -197 -3035
rect -177 -3038 -173 -3035
rect -169 -3035 -157 -3031
rect -143 -3035 -135 -3031
rect -169 -3038 -165 -3035
rect -135 -3038 -131 -3035
rect -127 -3035 -115 -3031
rect -101 -3035 -89 -3031
rect -127 -3038 -123 -3035
rect -93 -3038 -89 -3035
rect -85 -3035 -73 -3031
rect -59 -3031 -55 -3014
rect -35 -3017 -31 -2970
rect -35 -3031 -31 -3021
rect -59 -3035 -47 -3031
rect -85 -3038 -81 -3035
rect -51 -3038 -47 -3035
rect -43 -3035 -31 -3031
rect -43 -3038 -39 -3035
rect -210 -3046 -206 -3042
rect -193 -3046 -189 -3042
rect -152 -3046 -148 -3042
rect -110 -3046 -106 -3042
rect -68 -3046 -64 -3042
rect -27 -3046 -23 -3042
rect -210 -3078 -206 -3074
rect -193 -3078 -189 -3074
rect -173 -3078 -169 -3074
rect -152 -3078 -148 -3074
rect -131 -3078 -127 -3074
rect -110 -3078 -106 -3074
rect -89 -3078 -85 -3074
rect -68 -3078 -64 -3074
rect -47 -3078 -43 -3074
rect -27 -3078 -23 -3074
rect -219 -3133 -215 -3086
rect -219 -3154 -215 -3137
rect -201 -3147 -197 -3086
rect -185 -3147 -181 -3086
rect -161 -3126 -157 -3086
rect -161 -3147 -157 -3130
rect -143 -3147 -139 -3086
rect -119 -3133 -115 -3086
rect -119 -3147 -115 -3137
rect -101 -3126 -97 -3086
rect -101 -3147 -97 -3130
rect -77 -3140 -73 -3086
rect -59 -3118 -55 -3086
rect -59 -3126 -55 -3122
rect -77 -3147 -73 -3144
rect -201 -3151 -192 -3147
rect -185 -3151 -177 -3147
rect -201 -3154 -197 -3151
rect -177 -3154 -173 -3151
rect -169 -3151 -157 -3147
rect -143 -3151 -135 -3147
rect -169 -3154 -165 -3151
rect -135 -3154 -131 -3151
rect -127 -3151 -115 -3147
rect -101 -3151 -89 -3147
rect -127 -3154 -123 -3151
rect -93 -3154 -89 -3151
rect -85 -3151 -73 -3147
rect -59 -3147 -55 -3130
rect -35 -3133 -31 -3086
rect -35 -3147 -31 -3137
rect -59 -3151 -47 -3147
rect -85 -3154 -81 -3151
rect -51 -3154 -47 -3151
rect -43 -3151 -31 -3147
rect -43 -3154 -39 -3151
rect -210 -3162 -206 -3158
rect -193 -3162 -189 -3158
rect -152 -3162 -148 -3158
rect -110 -3162 -106 -3158
rect -68 -3162 -64 -3158
rect -27 -3162 -23 -3158
rect -21 -3170 -17 -3122
rect 197 -3126 201 -2938
rect -210 -3199 -206 -3195
rect -193 -3199 -189 -3195
rect -173 -3199 -169 -3195
rect -152 -3199 -148 -3195
rect -131 -3199 -127 -3195
rect -110 -3199 -106 -3195
rect -89 -3199 -85 -3195
rect -68 -3199 -64 -3195
rect -47 -3199 -43 -3195
rect -27 -3199 -23 -3195
rect -219 -3254 -215 -3207
rect -219 -3275 -215 -3258
rect -201 -3268 -197 -3207
rect -185 -3268 -181 -3207
rect -161 -3247 -157 -3207
rect -161 -3268 -157 -3251
rect -143 -3268 -139 -3207
rect -119 -3254 -115 -3207
rect -119 -3268 -115 -3258
rect -101 -3247 -97 -3207
rect -101 -3268 -97 -3251
rect -77 -3261 -73 -3207
rect -59 -3239 -55 -3207
rect -59 -3247 -55 -3243
rect -77 -3268 -73 -3265
rect -201 -3272 -192 -3268
rect -185 -3272 -177 -3268
rect -201 -3275 -197 -3272
rect -177 -3275 -173 -3272
rect -169 -3272 -157 -3268
rect -143 -3272 -135 -3268
rect -169 -3275 -165 -3272
rect -135 -3275 -131 -3272
rect -127 -3272 -115 -3268
rect -101 -3272 -89 -3268
rect -127 -3275 -123 -3272
rect -93 -3275 -89 -3272
rect -85 -3272 -73 -3268
rect -59 -3268 -55 -3251
rect -35 -3254 -31 -3207
rect -35 -3268 -31 -3258
rect -59 -3272 -47 -3268
rect -85 -3275 -81 -3272
rect -51 -3275 -47 -3272
rect -43 -3272 -31 -3268
rect -43 -3275 -39 -3272
rect -210 -3283 -206 -3279
rect -193 -3283 -189 -3279
rect -152 -3283 -148 -3279
rect -110 -3283 -106 -3279
rect -68 -3283 -64 -3279
rect -27 -3283 -23 -3279
rect -219 -3430 -215 -3426
rect -202 -3430 -198 -3426
rect -211 -3441 -207 -3438
rect -211 -3445 -196 -3441
rect -225 -3458 -218 -3454
rect -568 -3684 -564 -3680
rect -551 -3684 -547 -3680
rect -531 -3684 -527 -3680
rect -510 -3684 -506 -3680
rect -489 -3684 -485 -3680
rect -468 -3684 -464 -3680
rect -447 -3684 -443 -3680
rect -426 -3684 -422 -3680
rect -405 -3684 -401 -3680
rect -385 -3684 -381 -3680
rect -577 -3739 -573 -3692
rect -577 -3760 -573 -3743
rect -559 -3753 -555 -3692
rect -543 -3753 -539 -3692
rect -519 -3732 -515 -3692
rect -519 -3753 -515 -3736
rect -501 -3753 -497 -3692
rect -477 -3739 -473 -3692
rect -477 -3753 -473 -3743
rect -459 -3732 -455 -3692
rect -459 -3753 -455 -3736
rect -435 -3746 -431 -3692
rect -417 -3724 -413 -3692
rect -417 -3732 -413 -3728
rect -435 -3753 -431 -3750
rect -559 -3757 -550 -3753
rect -543 -3757 -535 -3753
rect -559 -3760 -555 -3757
rect -535 -3760 -531 -3757
rect -527 -3757 -515 -3753
rect -501 -3757 -493 -3753
rect -527 -3760 -523 -3757
rect -493 -3760 -489 -3757
rect -485 -3757 -473 -3753
rect -459 -3757 -447 -3753
rect -485 -3760 -481 -3757
rect -451 -3760 -447 -3757
rect -443 -3757 -431 -3753
rect -417 -3753 -413 -3736
rect -393 -3739 -389 -3692
rect -393 -3753 -389 -3743
rect -417 -3757 -405 -3753
rect -443 -3760 -439 -3757
rect -409 -3760 -405 -3757
rect -401 -3757 -389 -3753
rect -401 -3760 -397 -3757
rect -568 -3768 -564 -3764
rect -551 -3768 -547 -3764
rect -510 -3768 -506 -3764
rect -468 -3768 -464 -3764
rect -426 -3768 -422 -3764
rect -385 -3768 -381 -3764
rect -568 -3915 -564 -3911
rect -551 -3915 -547 -3911
rect -531 -3915 -527 -3911
rect -510 -3915 -506 -3911
rect -489 -3915 -485 -3911
rect -468 -3915 -464 -3911
rect -447 -3915 -443 -3911
rect -426 -3915 -422 -3911
rect -405 -3915 -401 -3911
rect -385 -3915 -381 -3911
rect -577 -3970 -573 -3923
rect -577 -3991 -573 -3974
rect -559 -3984 -555 -3923
rect -543 -3984 -539 -3923
rect -519 -3963 -515 -3923
rect -519 -3984 -515 -3967
rect -501 -3984 -497 -3923
rect -477 -3970 -473 -3923
rect -477 -3984 -473 -3974
rect -459 -3963 -455 -3923
rect -459 -3984 -455 -3967
rect -435 -3977 -431 -3923
rect -417 -3955 -413 -3923
rect -417 -3963 -413 -3959
rect -435 -3984 -431 -3981
rect -559 -3988 -550 -3984
rect -543 -3988 -535 -3984
rect -559 -3991 -555 -3988
rect -535 -3991 -531 -3988
rect -527 -3988 -515 -3984
rect -501 -3988 -493 -3984
rect -527 -3991 -523 -3988
rect -493 -3991 -489 -3988
rect -485 -3988 -473 -3984
rect -459 -3988 -447 -3984
rect -485 -3991 -481 -3988
rect -451 -3991 -447 -3988
rect -443 -3988 -431 -3984
rect -417 -3984 -413 -3967
rect -393 -3970 -389 -3923
rect -393 -3984 -389 -3974
rect -417 -3988 -405 -3984
rect -443 -3991 -439 -3988
rect -409 -3991 -405 -3988
rect -401 -3988 -389 -3984
rect -401 -3991 -397 -3988
rect -568 -3999 -564 -3995
rect -551 -3999 -547 -3995
rect -510 -3999 -506 -3995
rect -468 -3999 -464 -3995
rect -426 -3999 -422 -3995
rect -385 -3999 -381 -3995
rect -379 -4006 -375 -3959
rect -231 -3963 -227 -3656
rect -568 -4040 -564 -4036
rect -551 -4040 -547 -4036
rect -531 -4040 -527 -4036
rect -510 -4040 -506 -4036
rect -489 -4040 -485 -4036
rect -468 -4040 -464 -4036
rect -447 -4040 -443 -4036
rect -426 -4040 -422 -4036
rect -405 -4040 -401 -4036
rect -385 -4040 -381 -4036
rect -577 -4095 -573 -4048
rect -577 -4116 -573 -4099
rect -559 -4109 -555 -4048
rect -543 -4109 -539 -4048
rect -519 -4088 -515 -4048
rect -519 -4109 -515 -4092
rect -501 -4109 -497 -4048
rect -477 -4095 -473 -4048
rect -477 -4109 -473 -4099
rect -459 -4088 -455 -4048
rect -459 -4109 -455 -4092
rect -435 -4102 -431 -4048
rect -417 -4080 -413 -4048
rect -417 -4088 -413 -4084
rect -435 -4109 -431 -4106
rect -559 -4113 -550 -4109
rect -543 -4113 -535 -4109
rect -559 -4116 -555 -4113
rect -535 -4116 -531 -4113
rect -527 -4113 -515 -4109
rect -501 -4113 -493 -4109
rect -527 -4116 -523 -4113
rect -493 -4116 -489 -4113
rect -485 -4113 -473 -4109
rect -459 -4113 -447 -4109
rect -485 -4116 -481 -4113
rect -451 -4116 -447 -4113
rect -443 -4113 -431 -4109
rect -417 -4109 -413 -4092
rect -393 -4095 -389 -4048
rect -393 -4109 -389 -4099
rect -417 -4113 -405 -4109
rect -443 -4116 -439 -4113
rect -409 -4116 -405 -4113
rect -401 -4113 -389 -4109
rect -401 -4116 -397 -4113
rect -568 -4124 -564 -4120
rect -551 -4124 -547 -4120
rect -510 -4124 -506 -4120
rect -468 -4124 -464 -4120
rect -426 -4124 -422 -4120
rect -385 -4124 -381 -4120
rect -568 -4164 -564 -4160
rect -551 -4164 -547 -4160
rect -531 -4164 -527 -4160
rect -510 -4164 -506 -4160
rect -489 -4164 -485 -4160
rect -468 -4164 -464 -4160
rect -447 -4164 -443 -4160
rect -426 -4164 -422 -4160
rect -405 -4164 -401 -4160
rect -385 -4164 -381 -4160
rect -577 -4219 -573 -4172
rect -577 -4240 -573 -4223
rect -559 -4233 -555 -4172
rect -543 -4233 -539 -4172
rect -519 -4212 -515 -4172
rect -519 -4233 -515 -4216
rect -501 -4233 -497 -4172
rect -477 -4219 -473 -4172
rect -477 -4233 -473 -4223
rect -459 -4212 -455 -4172
rect -459 -4233 -455 -4216
rect -435 -4226 -431 -4172
rect -417 -4182 -413 -4172
rect -417 -4212 -413 -4186
rect -435 -4233 -431 -4230
rect -559 -4237 -550 -4233
rect -543 -4237 -535 -4233
rect -559 -4240 -555 -4237
rect -535 -4240 -531 -4237
rect -527 -4237 -515 -4233
rect -501 -4237 -493 -4233
rect -527 -4240 -523 -4237
rect -493 -4240 -489 -4237
rect -485 -4237 -473 -4233
rect -459 -4237 -447 -4233
rect -485 -4240 -481 -4237
rect -451 -4240 -447 -4237
rect -443 -4237 -431 -4233
rect -417 -4233 -413 -4216
rect -393 -4219 -389 -4172
rect -393 -4233 -389 -4223
rect -417 -4237 -405 -4233
rect -443 -4240 -439 -4237
rect -409 -4240 -405 -4237
rect -401 -4237 -389 -4233
rect -401 -4240 -397 -4237
rect -568 -4248 -564 -4244
rect -551 -4248 -547 -4244
rect -510 -4248 -506 -4244
rect -468 -4248 -464 -4244
rect -426 -4248 -422 -4244
rect -385 -4248 -381 -4244
rect -577 -4275 -573 -4271
rect -560 -4275 -556 -4271
rect -569 -4286 -565 -4283
rect -569 -4290 -554 -4286
rect -583 -4303 -576 -4299
rect -926 -4517 -922 -4513
rect -909 -4517 -905 -4513
rect -889 -4517 -885 -4513
rect -868 -4517 -864 -4513
rect -847 -4517 -843 -4513
rect -826 -4517 -822 -4513
rect -805 -4517 -801 -4513
rect -784 -4517 -780 -4513
rect -763 -4517 -759 -4513
rect -743 -4517 -739 -4513
rect -935 -4572 -931 -4525
rect -935 -4593 -931 -4576
rect -917 -4586 -913 -4525
rect -901 -4586 -897 -4525
rect -877 -4565 -873 -4525
rect -877 -4586 -873 -4569
rect -859 -4586 -855 -4525
rect -835 -4572 -831 -4525
rect -835 -4586 -831 -4576
rect -817 -4565 -813 -4525
rect -817 -4586 -813 -4569
rect -793 -4579 -789 -4525
rect -775 -4557 -771 -4525
rect -775 -4565 -771 -4561
rect -793 -4586 -789 -4583
rect -917 -4590 -908 -4586
rect -901 -4590 -893 -4586
rect -917 -4593 -913 -4590
rect -893 -4593 -889 -4590
rect -885 -4590 -873 -4586
rect -859 -4590 -851 -4586
rect -885 -4593 -881 -4590
rect -851 -4593 -847 -4590
rect -843 -4590 -831 -4586
rect -817 -4590 -805 -4586
rect -843 -4593 -839 -4590
rect -809 -4593 -805 -4590
rect -801 -4590 -789 -4586
rect -775 -4586 -771 -4569
rect -751 -4572 -747 -4525
rect -751 -4586 -747 -4576
rect -775 -4590 -763 -4586
rect -801 -4593 -797 -4590
rect -767 -4593 -763 -4590
rect -759 -4590 -747 -4586
rect -759 -4593 -755 -4590
rect -926 -4601 -922 -4597
rect -909 -4601 -905 -4597
rect -868 -4601 -864 -4597
rect -826 -4601 -822 -4597
rect -784 -4601 -780 -4597
rect -743 -4601 -739 -4597
rect -926 -4638 -922 -4634
rect -909 -4638 -905 -4634
rect -889 -4638 -885 -4634
rect -868 -4638 -864 -4634
rect -847 -4638 -843 -4634
rect -826 -4638 -822 -4634
rect -805 -4638 -801 -4634
rect -784 -4638 -780 -4634
rect -763 -4638 -759 -4634
rect -743 -4638 -739 -4634
rect -935 -4693 -931 -4646
rect -935 -4714 -931 -4697
rect -917 -4707 -913 -4646
rect -901 -4707 -897 -4646
rect -877 -4686 -873 -4646
rect -877 -4707 -873 -4690
rect -859 -4707 -855 -4646
rect -835 -4693 -831 -4646
rect -835 -4707 -831 -4697
rect -817 -4686 -813 -4646
rect -817 -4707 -813 -4690
rect -793 -4700 -789 -4646
rect -775 -4678 -771 -4646
rect -775 -4686 -771 -4682
rect -793 -4707 -789 -4704
rect -917 -4711 -908 -4707
rect -901 -4711 -893 -4707
rect -917 -4714 -913 -4711
rect -893 -4714 -889 -4711
rect -885 -4711 -873 -4707
rect -859 -4711 -851 -4707
rect -885 -4714 -881 -4711
rect -851 -4714 -847 -4711
rect -843 -4711 -831 -4707
rect -817 -4711 -805 -4707
rect -843 -4714 -839 -4711
rect -809 -4714 -805 -4711
rect -801 -4711 -789 -4707
rect -775 -4707 -771 -4690
rect -751 -4693 -747 -4646
rect -751 -4707 -747 -4697
rect -775 -4711 -763 -4707
rect -801 -4714 -797 -4711
rect -767 -4714 -763 -4711
rect -759 -4711 -747 -4707
rect -759 -4714 -755 -4711
rect -926 -4722 -922 -4718
rect -909 -4722 -905 -4718
rect -868 -4722 -864 -4718
rect -826 -4722 -822 -4718
rect -784 -4722 -780 -4718
rect -743 -4722 -739 -4718
rect -737 -4729 -733 -4682
rect -589 -4686 -585 -4489
rect -926 -4759 -922 -4755
rect -909 -4759 -905 -4755
rect -889 -4759 -885 -4755
rect -868 -4759 -864 -4755
rect -847 -4759 -843 -4755
rect -826 -4759 -822 -4755
rect -805 -4759 -801 -4755
rect -784 -4759 -780 -4755
rect -763 -4759 -759 -4755
rect -743 -4759 -739 -4755
rect -935 -4814 -931 -4767
rect -935 -4835 -931 -4818
rect -917 -4828 -913 -4767
rect -901 -4828 -897 -4767
rect -877 -4807 -873 -4767
rect -877 -4828 -873 -4811
rect -859 -4828 -855 -4767
rect -835 -4814 -831 -4767
rect -835 -4828 -831 -4818
rect -817 -4807 -813 -4767
rect -817 -4828 -813 -4811
rect -793 -4821 -789 -4767
rect -775 -4799 -771 -4767
rect -775 -4807 -771 -4803
rect -793 -4828 -789 -4825
rect -917 -4832 -908 -4828
rect -901 -4832 -893 -4828
rect -917 -4835 -913 -4832
rect -893 -4835 -889 -4832
rect -885 -4832 -873 -4828
rect -859 -4832 -851 -4828
rect -885 -4835 -881 -4832
rect -851 -4835 -847 -4832
rect -843 -4832 -831 -4828
rect -817 -4832 -805 -4828
rect -843 -4835 -839 -4832
rect -809 -4835 -805 -4832
rect -801 -4832 -789 -4828
rect -775 -4828 -771 -4811
rect -751 -4814 -747 -4767
rect -751 -4828 -747 -4818
rect -775 -4832 -763 -4828
rect -801 -4835 -797 -4832
rect -767 -4835 -763 -4832
rect -759 -4832 -747 -4828
rect -759 -4835 -755 -4832
rect -926 -4843 -922 -4839
rect -909 -4843 -905 -4839
rect -868 -4843 -864 -4839
rect -826 -4843 -822 -4839
rect -784 -4843 -780 -4839
rect -743 -4843 -739 -4839
rect -926 -4877 -922 -4873
rect -909 -4877 -905 -4873
rect -889 -4877 -885 -4873
rect -868 -4877 -864 -4873
rect -847 -4877 -843 -4873
rect -826 -4877 -822 -4873
rect -805 -4877 -801 -4873
rect -784 -4877 -780 -4873
rect -763 -4877 -759 -4873
rect -743 -4877 -739 -4873
rect -935 -4932 -931 -4885
rect -935 -4953 -931 -4936
rect -917 -4946 -913 -4885
rect -901 -4946 -897 -4885
rect -877 -4925 -873 -4885
rect -877 -4946 -873 -4929
rect -859 -4946 -855 -4885
rect -835 -4932 -831 -4885
rect -835 -4946 -831 -4936
rect -817 -4925 -813 -4885
rect -817 -4946 -813 -4929
rect -793 -4939 -789 -4885
rect -775 -4917 -771 -4885
rect -775 -4925 -771 -4921
rect -793 -4946 -789 -4943
rect -917 -4950 -908 -4946
rect -901 -4950 -893 -4946
rect -917 -4953 -913 -4950
rect -893 -4953 -889 -4950
rect -885 -4950 -873 -4946
rect -859 -4950 -851 -4946
rect -885 -4953 -881 -4950
rect -851 -4953 -847 -4950
rect -843 -4950 -831 -4946
rect -817 -4950 -805 -4946
rect -843 -4953 -839 -4950
rect -809 -4953 -805 -4950
rect -801 -4950 -789 -4946
rect -775 -4946 -771 -4929
rect -751 -4932 -747 -4885
rect -751 -4946 -747 -4936
rect -775 -4950 -763 -4946
rect -801 -4953 -797 -4950
rect -767 -4953 -763 -4950
rect -759 -4950 -747 -4946
rect -759 -4953 -755 -4950
rect -926 -4961 -922 -4957
rect -909 -4961 -905 -4957
rect -868 -4961 -864 -4957
rect -826 -4961 -822 -4957
rect -784 -4961 -780 -4957
rect -743 -4961 -739 -4957
rect -935 -4994 -931 -4990
rect -918 -4994 -914 -4990
rect -927 -5005 -923 -5002
rect -927 -5009 -912 -5005
rect -941 -5022 -934 -5018
rect -1255 -5197 -1251 -5193
rect -1211 -5197 -1207 -5193
rect -1177 -5197 -1173 -5193
rect -1276 -5401 -1272 -5208
rect -1162 -5212 -1158 -5179
rect -1270 -5280 -1266 -5216
rect -1255 -5232 -1251 -5228
rect -1238 -5232 -1234 -5228
rect -1218 -5232 -1214 -5228
rect -1197 -5232 -1193 -5228
rect -1176 -5232 -1172 -5228
rect -1155 -5232 -1151 -5228
rect -1134 -5232 -1130 -5228
rect -1113 -5232 -1109 -5228
rect -1092 -5232 -1088 -5228
rect -1072 -5232 -1068 -5228
rect -1264 -5287 -1260 -5240
rect -1264 -5308 -1260 -5291
rect -1246 -5301 -1242 -5240
rect -1230 -5301 -1226 -5240
rect -1206 -5280 -1202 -5240
rect -1206 -5301 -1202 -5284
rect -1188 -5301 -1184 -5240
rect -1164 -5287 -1160 -5240
rect -1164 -5301 -1160 -5291
rect -1146 -5280 -1142 -5240
rect -1146 -5301 -1142 -5284
rect -1122 -5294 -1118 -5240
rect -1104 -5272 -1100 -5240
rect -1104 -5280 -1100 -5276
rect -1122 -5301 -1118 -5298
rect -1246 -5305 -1237 -5301
rect -1230 -5305 -1222 -5301
rect -1246 -5308 -1242 -5305
rect -1222 -5308 -1218 -5305
rect -1214 -5305 -1202 -5301
rect -1188 -5305 -1180 -5301
rect -1214 -5308 -1210 -5305
rect -1180 -5308 -1176 -5305
rect -1172 -5305 -1160 -5301
rect -1146 -5305 -1134 -5301
rect -1172 -5308 -1168 -5305
rect -1138 -5308 -1134 -5305
rect -1130 -5305 -1118 -5301
rect -1104 -5301 -1100 -5284
rect -1080 -5287 -1076 -5240
rect -1080 -5301 -1076 -5291
rect -1104 -5305 -1092 -5301
rect -1130 -5308 -1126 -5305
rect -1096 -5308 -1092 -5305
rect -1088 -5305 -1076 -5301
rect -1088 -5308 -1084 -5305
rect -1255 -5316 -1251 -5312
rect -1238 -5316 -1234 -5312
rect -1197 -5316 -1193 -5312
rect -1155 -5316 -1151 -5312
rect -1113 -5316 -1109 -5312
rect -1072 -5316 -1068 -5312
rect -1255 -5353 -1251 -5349
rect -1238 -5353 -1234 -5349
rect -1218 -5353 -1214 -5349
rect -1197 -5353 -1193 -5349
rect -1176 -5353 -1172 -5349
rect -1155 -5353 -1151 -5349
rect -1134 -5353 -1130 -5349
rect -1113 -5353 -1109 -5349
rect -1092 -5353 -1088 -5349
rect -1072 -5353 -1068 -5349
rect -1026 -5353 -1022 -5349
rect -1264 -5408 -1260 -5361
rect -1264 -5429 -1260 -5412
rect -1246 -5422 -1242 -5361
rect -1230 -5422 -1226 -5361
rect -1206 -5401 -1202 -5361
rect -1206 -5422 -1202 -5405
rect -1188 -5422 -1184 -5361
rect -1164 -5408 -1160 -5361
rect -1164 -5422 -1160 -5412
rect -1146 -5401 -1142 -5361
rect -1146 -5422 -1142 -5405
rect -1122 -5415 -1118 -5361
rect -1104 -5393 -1100 -5361
rect -1104 -5401 -1100 -5397
rect -1122 -5422 -1118 -5419
rect -1246 -5426 -1237 -5422
rect -1230 -5426 -1222 -5422
rect -1246 -5429 -1242 -5426
rect -1222 -5429 -1218 -5426
rect -1214 -5426 -1202 -5422
rect -1188 -5426 -1180 -5422
rect -1214 -5429 -1210 -5426
rect -1180 -5429 -1176 -5426
rect -1172 -5426 -1160 -5422
rect -1146 -5426 -1134 -5422
rect -1172 -5429 -1168 -5426
rect -1138 -5429 -1134 -5426
rect -1130 -5426 -1118 -5422
rect -1104 -5422 -1100 -5405
rect -1080 -5408 -1076 -5361
rect -1018 -5390 -1014 -5361
rect -1080 -5422 -1076 -5412
rect -1104 -5426 -1092 -5422
rect -1130 -5429 -1126 -5426
rect -1096 -5429 -1092 -5426
rect -1088 -5426 -1076 -5422
rect -1088 -5429 -1084 -5426
rect -1255 -5437 -1251 -5433
rect -1238 -5437 -1234 -5433
rect -1197 -5437 -1193 -5433
rect -1155 -5437 -1151 -5433
rect -1113 -5437 -1109 -5433
rect -1072 -5437 -1068 -5433
rect -1066 -5444 -1062 -5397
rect -1018 -5429 -1014 -5394
rect -947 -5401 -943 -5215
rect -1026 -5437 -1022 -5433
rect -1339 -5707 -1335 -5703
rect -1322 -5707 -1318 -5703
rect -1331 -5718 -1327 -5715
rect -1331 -5722 -1316 -5718
rect -1320 -5761 -1316 -5722
rect -1320 -5776 -1316 -5765
rect -1339 -5780 -1316 -5776
rect -1339 -5783 -1335 -5780
rect -1313 -5783 -1309 -5715
rect -1322 -5791 -1318 -5787
rect -1313 -5881 -1309 -5787
rect -1270 -5874 -1266 -5448
rect -1255 -5473 -1251 -5469
rect -1238 -5473 -1234 -5469
rect -1218 -5473 -1214 -5469
rect -1197 -5473 -1193 -5469
rect -1176 -5473 -1172 -5469
rect -1155 -5473 -1151 -5469
rect -1134 -5473 -1130 -5469
rect -1113 -5473 -1109 -5469
rect -1092 -5473 -1088 -5469
rect -1072 -5473 -1068 -5469
rect -1026 -5473 -1022 -5469
rect -1264 -5528 -1260 -5481
rect -1264 -5549 -1260 -5532
rect -1246 -5542 -1242 -5481
rect -1230 -5542 -1226 -5481
rect -1206 -5521 -1202 -5481
rect -1206 -5542 -1202 -5525
rect -1188 -5542 -1184 -5481
rect -1164 -5528 -1160 -5481
rect -1164 -5542 -1160 -5532
rect -1146 -5521 -1142 -5481
rect -1146 -5542 -1142 -5525
rect -1122 -5535 -1118 -5481
rect -1104 -5513 -1100 -5481
rect -1104 -5521 -1100 -5517
rect -1122 -5542 -1118 -5539
rect -1246 -5546 -1237 -5542
rect -1230 -5546 -1222 -5542
rect -1246 -5549 -1242 -5546
rect -1222 -5549 -1218 -5546
rect -1214 -5546 -1202 -5542
rect -1188 -5546 -1180 -5542
rect -1214 -5549 -1210 -5546
rect -1180 -5549 -1176 -5546
rect -1172 -5546 -1160 -5542
rect -1146 -5546 -1134 -5542
rect -1172 -5549 -1168 -5546
rect -1138 -5549 -1134 -5546
rect -1130 -5546 -1118 -5542
rect -1104 -5542 -1100 -5525
rect -1080 -5528 -1076 -5481
rect -1080 -5542 -1076 -5532
rect -1104 -5546 -1092 -5542
rect -1130 -5549 -1126 -5546
rect -1096 -5549 -1092 -5546
rect -1088 -5546 -1076 -5542
rect -1088 -5549 -1084 -5546
rect -1255 -5557 -1251 -5553
rect -1238 -5557 -1234 -5553
rect -1197 -5557 -1193 -5553
rect -1155 -5557 -1151 -5553
rect -1113 -5557 -1109 -5553
rect -1072 -5557 -1068 -5553
rect -1255 -5590 -1251 -5586
rect -1238 -5590 -1234 -5586
rect -1218 -5590 -1214 -5586
rect -1197 -5590 -1193 -5586
rect -1176 -5590 -1172 -5586
rect -1155 -5590 -1151 -5586
rect -1134 -5590 -1130 -5586
rect -1113 -5590 -1109 -5586
rect -1092 -5590 -1088 -5586
rect -1072 -5590 -1068 -5586
rect -1264 -5645 -1260 -5598
rect -1264 -5666 -1260 -5649
rect -1246 -5659 -1242 -5598
rect -1230 -5659 -1226 -5598
rect -1206 -5638 -1202 -5598
rect -1206 -5659 -1202 -5642
rect -1188 -5659 -1184 -5598
rect -1164 -5645 -1160 -5598
rect -1164 -5659 -1160 -5649
rect -1146 -5638 -1142 -5598
rect -1146 -5659 -1142 -5642
rect -1122 -5652 -1118 -5598
rect -1104 -5630 -1100 -5598
rect -1104 -5638 -1100 -5634
rect -1122 -5659 -1118 -5656
rect -1246 -5663 -1237 -5659
rect -1230 -5663 -1222 -5659
rect -1246 -5666 -1242 -5663
rect -1222 -5666 -1218 -5663
rect -1214 -5663 -1202 -5659
rect -1188 -5663 -1180 -5659
rect -1214 -5666 -1210 -5663
rect -1180 -5666 -1176 -5663
rect -1172 -5663 -1160 -5659
rect -1146 -5663 -1134 -5659
rect -1172 -5666 -1168 -5663
rect -1138 -5666 -1134 -5663
rect -1130 -5663 -1118 -5659
rect -1104 -5659 -1100 -5642
rect -1080 -5645 -1076 -5598
rect -1080 -5659 -1076 -5649
rect -1104 -5663 -1092 -5659
rect -1130 -5666 -1126 -5663
rect -1096 -5666 -1092 -5663
rect -1088 -5663 -1076 -5659
rect -1088 -5666 -1084 -5663
rect -1255 -5674 -1251 -5670
rect -1238 -5674 -1234 -5670
rect -1197 -5674 -1193 -5670
rect -1155 -5674 -1151 -5670
rect -1113 -5674 -1109 -5670
rect -1072 -5674 -1068 -5670
rect -1066 -5731 -1062 -5517
rect -1018 -5514 -1014 -5481
rect -1018 -5549 -1014 -5518
rect -1026 -5557 -1022 -5553
rect -1255 -5826 -1251 -5822
rect -1238 -5826 -1234 -5822
rect -1198 -5826 -1194 -5822
rect -1177 -5826 -1173 -5822
rect -1264 -5867 -1260 -5834
rect -1264 -5902 -1260 -5871
rect -1246 -5861 -1242 -5834
rect -1246 -5865 -1237 -5861
rect -1246 -5902 -1242 -5865
rect -1220 -5888 -1216 -5834
rect -1220 -5895 -1216 -5892
rect -1186 -5895 -1182 -5834
rect -1168 -5866 -1164 -5834
rect -953 -5858 -949 -5756
rect -1238 -5902 -1234 -5899
rect -1229 -5899 -1216 -5895
rect -1229 -5902 -1225 -5899
rect -1202 -5902 -1198 -5899
rect -1194 -5899 -1175 -5895
rect -1194 -5902 -1190 -5899
rect -1168 -5902 -1164 -5870
rect -947 -5873 -943 -5448
rect -941 -5521 -937 -5022
rect -916 -5048 -912 -5009
rect -916 -5063 -912 -5052
rect -935 -5067 -912 -5063
rect -909 -5039 -905 -5002
rect -737 -5018 -733 -4803
rect -935 -5070 -931 -5067
rect -909 -5070 -905 -5043
rect -918 -5078 -914 -5074
rect -926 -5113 -922 -5109
rect -900 -5113 -896 -5109
rect -883 -5113 -879 -5109
rect -843 -5113 -839 -5109
rect -822 -5113 -818 -5109
rect -805 -5113 -801 -5109
rect -765 -5113 -761 -5109
rect -741 -5113 -737 -5109
rect -704 -5113 -700 -5109
rect -935 -5138 -931 -5121
rect -935 -5189 -931 -5142
rect -917 -5131 -913 -5121
rect -917 -5189 -913 -5135
rect -909 -5160 -905 -5121
rect -891 -5153 -887 -5121
rect -909 -5189 -905 -5164
rect -891 -5189 -887 -5157
rect -865 -5145 -861 -5121
rect -865 -5182 -861 -5149
rect -831 -5182 -827 -5121
rect -813 -5138 -809 -5121
rect -883 -5189 -879 -5186
rect -875 -5186 -861 -5182
rect -875 -5189 -871 -5186
rect -847 -5189 -843 -5186
rect -839 -5186 -820 -5182
rect -839 -5189 -835 -5186
rect -813 -5189 -809 -5142
rect -787 -5153 -783 -5121
rect -787 -5182 -783 -5157
rect -753 -5175 -749 -5121
rect -753 -5179 -736 -5175
rect -805 -5189 -801 -5186
rect -796 -5186 -783 -5182
rect -796 -5189 -792 -5186
rect -769 -5189 -765 -5186
rect -745 -5189 -741 -5179
rect -729 -5182 -725 -5121
rect -721 -5175 -717 -5121
rect -695 -5145 -691 -5121
rect -721 -5179 -702 -5175
rect -737 -5186 -720 -5182
rect -737 -5189 -733 -5186
rect -713 -5189 -709 -5179
rect -695 -5189 -691 -5149
rect -926 -5197 -922 -5193
rect -900 -5197 -896 -5193
rect -857 -5197 -853 -5193
rect -822 -5197 -818 -5193
rect -778 -5197 -774 -5193
rect -761 -5197 -757 -5193
rect -725 -5197 -721 -5193
rect -704 -5197 -700 -5193
rect -689 -5204 -685 -5157
rect -595 -5160 -591 -5043
rect -589 -5145 -585 -4733
rect -583 -4807 -579 -4303
rect -558 -4329 -554 -4290
rect -558 -4344 -554 -4333
rect -577 -4348 -554 -4344
rect -551 -4320 -547 -4283
rect -379 -4299 -375 -4084
rect -332 -4164 -328 -4160
rect -324 -4203 -320 -4172
rect -324 -4240 -320 -4207
rect -332 -4248 -328 -4244
rect -332 -4275 -328 -4271
rect -577 -4351 -573 -4348
rect -551 -4351 -547 -4324
rect -324 -4318 -320 -4283
rect -324 -4351 -320 -4322
rect -560 -4359 -556 -4355
rect -332 -4359 -328 -4355
rect -568 -4394 -564 -4390
rect -542 -4394 -538 -4390
rect -525 -4394 -521 -4390
rect -485 -4394 -481 -4390
rect -464 -4394 -460 -4390
rect -447 -4394 -443 -4390
rect -407 -4394 -403 -4390
rect -383 -4394 -379 -4390
rect -346 -4394 -342 -4390
rect -577 -4419 -573 -4402
rect -577 -4470 -573 -4423
rect -559 -4412 -555 -4402
rect -559 -4470 -555 -4416
rect -551 -4441 -547 -4402
rect -533 -4434 -529 -4402
rect -551 -4470 -547 -4445
rect -533 -4470 -529 -4438
rect -507 -4426 -503 -4402
rect -507 -4463 -503 -4430
rect -473 -4463 -469 -4402
rect -455 -4419 -451 -4402
rect -525 -4470 -521 -4467
rect -517 -4467 -503 -4463
rect -517 -4470 -513 -4467
rect -489 -4470 -485 -4467
rect -481 -4467 -462 -4463
rect -481 -4470 -477 -4467
rect -455 -4470 -451 -4423
rect -429 -4434 -425 -4402
rect -429 -4463 -425 -4438
rect -395 -4456 -391 -4402
rect -395 -4460 -378 -4456
rect -447 -4470 -443 -4467
rect -438 -4467 -425 -4463
rect -438 -4470 -434 -4467
rect -411 -4470 -407 -4467
rect -387 -4470 -383 -4460
rect -371 -4463 -367 -4402
rect -363 -4456 -359 -4402
rect -337 -4425 -333 -4402
rect -363 -4460 -344 -4456
rect -379 -4467 -362 -4463
rect -379 -4470 -375 -4467
rect -355 -4470 -351 -4460
rect -337 -4470 -333 -4429
rect -568 -4478 -564 -4474
rect -542 -4478 -538 -4474
rect -499 -4478 -495 -4474
rect -464 -4478 -460 -4474
rect -420 -4478 -416 -4474
rect -403 -4478 -399 -4474
rect -367 -4478 -363 -4474
rect -346 -4478 -342 -4474
rect -331 -4492 -327 -4438
rect -237 -4441 -233 -4324
rect -231 -4426 -227 -4010
rect -225 -4088 -221 -3458
rect -200 -3484 -196 -3445
rect -200 -3499 -196 -3488
rect -219 -3503 -196 -3499
rect -193 -3475 -189 -3438
rect -21 -3454 -17 -3243
rect -219 -3506 -215 -3503
rect -193 -3506 -189 -3479
rect -202 -3514 -198 -3510
rect -210 -3554 -206 -3550
rect -184 -3554 -180 -3550
rect -167 -3554 -163 -3550
rect -127 -3554 -123 -3550
rect -106 -3554 -102 -3550
rect -89 -3554 -85 -3550
rect -49 -3554 -45 -3550
rect -25 -3554 -21 -3550
rect 12 -3554 16 -3550
rect -219 -3579 -215 -3562
rect -219 -3630 -215 -3583
rect -201 -3572 -197 -3562
rect -201 -3630 -197 -3576
rect -193 -3601 -189 -3562
rect -175 -3594 -171 -3562
rect -193 -3630 -189 -3605
rect -175 -3630 -171 -3598
rect -149 -3586 -145 -3562
rect -149 -3623 -145 -3590
rect -115 -3623 -111 -3562
rect -97 -3579 -93 -3562
rect -167 -3630 -163 -3627
rect -159 -3627 -145 -3623
rect -159 -3630 -155 -3627
rect -131 -3630 -127 -3627
rect -123 -3627 -104 -3623
rect -123 -3630 -119 -3627
rect -97 -3630 -93 -3583
rect -71 -3594 -67 -3562
rect -71 -3623 -67 -3598
rect -37 -3616 -33 -3562
rect -37 -3620 -20 -3616
rect -89 -3630 -85 -3627
rect -80 -3627 -67 -3623
rect -80 -3630 -76 -3627
rect -53 -3630 -49 -3627
rect -29 -3630 -25 -3620
rect -13 -3623 -9 -3562
rect -5 -3616 -1 -3562
rect 21 -3586 25 -3562
rect -5 -3620 14 -3616
rect -21 -3627 -4 -3623
rect -21 -3630 -17 -3627
rect 3 -3630 7 -3620
rect 21 -3630 25 -3590
rect -210 -3638 -206 -3634
rect -184 -3638 -180 -3634
rect -141 -3638 -137 -3634
rect -106 -3638 -102 -3634
rect -62 -3638 -58 -3634
rect -45 -3638 -41 -3634
rect -9 -3638 -5 -3634
rect 12 -3638 16 -3634
rect 27 -3645 31 -3598
rect 191 -3601 195 -3479
rect 197 -3586 201 -3173
rect 203 -3247 207 -2752
rect 228 -2778 232 -2739
rect 228 -2793 232 -2782
rect 209 -2797 232 -2793
rect 235 -2769 239 -2732
rect 407 -2748 411 -2543
rect 209 -2800 213 -2797
rect 235 -2800 239 -2773
rect 226 -2808 230 -2804
rect 218 -2843 222 -2839
rect 244 -2843 248 -2839
rect 261 -2843 265 -2839
rect 301 -2843 305 -2839
rect 322 -2843 326 -2839
rect 339 -2843 343 -2839
rect 379 -2843 383 -2839
rect 403 -2843 407 -2839
rect 440 -2843 444 -2839
rect 209 -2868 213 -2851
rect 209 -2919 213 -2872
rect 227 -2861 231 -2851
rect 227 -2919 231 -2865
rect 235 -2890 239 -2851
rect 253 -2883 257 -2851
rect 235 -2919 239 -2894
rect 253 -2919 257 -2887
rect 279 -2875 283 -2851
rect 279 -2912 283 -2879
rect 313 -2912 317 -2851
rect 331 -2868 335 -2851
rect 261 -2919 265 -2916
rect 269 -2916 283 -2912
rect 269 -2919 273 -2916
rect 297 -2919 301 -2916
rect 305 -2916 324 -2912
rect 305 -2919 309 -2916
rect 331 -2919 335 -2872
rect 357 -2883 361 -2851
rect 357 -2912 361 -2887
rect 391 -2905 395 -2851
rect 391 -2909 408 -2905
rect 339 -2919 343 -2916
rect 348 -2916 361 -2912
rect 348 -2919 352 -2916
rect 375 -2919 379 -2916
rect 399 -2919 403 -2909
rect 415 -2912 419 -2851
rect 423 -2905 427 -2851
rect 449 -2875 453 -2851
rect 423 -2909 442 -2905
rect 407 -2916 424 -2912
rect 407 -2919 411 -2916
rect 431 -2919 435 -2909
rect 449 -2919 453 -2879
rect 218 -2927 222 -2923
rect 244 -2927 248 -2923
rect 287 -2927 291 -2923
rect 322 -2927 326 -2923
rect 366 -2927 370 -2923
rect 383 -2927 387 -2923
rect 419 -2927 423 -2923
rect 440 -2927 444 -2923
rect 455 -2941 459 -2887
rect 547 -2890 551 -2773
rect 553 -2875 557 -2463
rect 559 -2547 563 -2002
rect 584 -2028 588 -1989
rect 584 -2043 588 -2032
rect 565 -2047 588 -2043
rect 591 -2019 595 -1982
rect 763 -1998 767 -1791
rect 841 -1862 845 -1858
rect 849 -1903 853 -1878
rect 849 -1934 853 -1907
rect 841 -1946 845 -1942
rect 565 -2050 569 -2047
rect 591 -2050 595 -2023
rect 582 -2058 586 -2054
rect 574 -2093 578 -2089
rect 600 -2093 604 -2089
rect 617 -2093 621 -2089
rect 657 -2093 661 -2089
rect 678 -2093 682 -2089
rect 695 -2093 699 -2089
rect 735 -2093 739 -2089
rect 759 -2093 763 -2089
rect 796 -2093 800 -2089
rect 565 -2118 569 -2101
rect 565 -2169 569 -2122
rect 583 -2111 587 -2101
rect 583 -2169 587 -2115
rect 591 -2140 595 -2101
rect 609 -2133 613 -2101
rect 591 -2169 595 -2144
rect 609 -2169 613 -2137
rect 635 -2125 639 -2101
rect 635 -2162 639 -2129
rect 669 -2162 673 -2101
rect 687 -2118 691 -2101
rect 617 -2169 621 -2166
rect 625 -2166 639 -2162
rect 625 -2169 629 -2166
rect 653 -2169 657 -2166
rect 661 -2166 680 -2162
rect 661 -2169 665 -2166
rect 687 -2169 691 -2122
rect 713 -2133 717 -2101
rect 713 -2162 717 -2137
rect 747 -2155 751 -2101
rect 747 -2159 764 -2155
rect 695 -2169 699 -2166
rect 704 -2166 717 -2162
rect 704 -2169 708 -2166
rect 731 -2169 735 -2166
rect 755 -2169 759 -2159
rect 771 -2162 775 -2101
rect 779 -2155 783 -2101
rect 805 -2125 809 -2101
rect 779 -2159 798 -2155
rect 763 -2166 780 -2162
rect 763 -2169 767 -2166
rect 787 -2169 791 -2159
rect 805 -2169 809 -2129
rect 574 -2177 578 -2173
rect 600 -2177 604 -2173
rect 643 -2177 647 -2173
rect 678 -2177 682 -2173
rect 722 -2177 726 -2173
rect 739 -2177 743 -2173
rect 775 -2177 779 -2173
rect 796 -2177 800 -2173
rect 811 -2184 815 -2137
rect 945 -2140 949 -2023
rect 951 -2125 955 -1721
rect 957 -1795 961 -1296
rect 982 -1322 986 -1283
rect 982 -1337 986 -1326
rect 963 -1341 986 -1337
rect 989 -1313 993 -1276
rect 1315 -1292 1319 -1066
rect 1340 -1107 1344 -1053
rect 1321 -1111 1340 -1107
rect 1347 -1086 1351 -1046
rect 1321 -1114 1325 -1111
rect 1347 -1114 1351 -1090
rect 1338 -1122 1342 -1118
rect 1321 -1268 1325 -1264
rect 1338 -1268 1342 -1264
rect 1329 -1279 1333 -1276
rect 1329 -1283 1344 -1279
rect 1315 -1296 1322 -1292
rect 963 -1344 967 -1341
rect 989 -1344 993 -1317
rect 980 -1352 984 -1348
rect 972 -1382 976 -1378
rect 998 -1382 1002 -1378
rect 1015 -1382 1019 -1378
rect 1055 -1382 1059 -1378
rect 1076 -1382 1080 -1378
rect 1093 -1382 1097 -1378
rect 1133 -1382 1137 -1378
rect 1157 -1382 1161 -1378
rect 1194 -1382 1198 -1378
rect 963 -1407 967 -1390
rect 963 -1458 967 -1411
rect 981 -1400 985 -1390
rect 981 -1458 985 -1404
rect 989 -1429 993 -1390
rect 1007 -1422 1011 -1390
rect 989 -1458 993 -1433
rect 1007 -1458 1011 -1426
rect 1033 -1414 1037 -1390
rect 1033 -1451 1037 -1418
rect 1067 -1451 1071 -1390
rect 1085 -1407 1089 -1390
rect 1015 -1458 1019 -1455
rect 1023 -1455 1037 -1451
rect 1023 -1458 1027 -1455
rect 1051 -1458 1055 -1455
rect 1059 -1455 1078 -1451
rect 1059 -1458 1063 -1455
rect 1085 -1458 1089 -1411
rect 1111 -1422 1115 -1390
rect 1111 -1451 1115 -1426
rect 1145 -1444 1149 -1390
rect 1145 -1448 1162 -1444
rect 1093 -1458 1097 -1455
rect 1102 -1455 1115 -1451
rect 1102 -1458 1106 -1455
rect 1129 -1458 1133 -1455
rect 1153 -1458 1157 -1448
rect 1169 -1451 1173 -1390
rect 1177 -1444 1181 -1390
rect 1203 -1430 1207 -1390
rect 1177 -1448 1196 -1444
rect 1161 -1455 1178 -1451
rect 1161 -1458 1165 -1455
rect 1185 -1458 1189 -1448
rect 1203 -1458 1207 -1434
rect 972 -1466 976 -1462
rect 998 -1466 1002 -1462
rect 1041 -1466 1045 -1462
rect 1076 -1466 1080 -1462
rect 1120 -1466 1124 -1462
rect 1137 -1466 1141 -1462
rect 1173 -1466 1177 -1462
rect 1194 -1466 1198 -1462
rect 1209 -1480 1213 -1426
rect 1309 -1437 1313 -1317
rect 972 -1505 976 -1501
rect 989 -1505 993 -1501
rect 1009 -1505 1013 -1501
rect 1030 -1505 1034 -1501
rect 1051 -1505 1055 -1501
rect 1072 -1505 1076 -1501
rect 1093 -1505 1097 -1501
rect 1114 -1505 1118 -1501
rect 1135 -1505 1139 -1501
rect 1155 -1505 1159 -1501
rect 963 -1560 967 -1513
rect 963 -1581 967 -1564
rect 981 -1574 985 -1513
rect 997 -1574 1001 -1513
rect 1021 -1553 1025 -1513
rect 1021 -1574 1025 -1557
rect 1039 -1574 1043 -1513
rect 1063 -1560 1067 -1513
rect 1063 -1574 1067 -1564
rect 1081 -1553 1085 -1513
rect 1081 -1574 1085 -1557
rect 1105 -1567 1109 -1513
rect 1123 -1545 1127 -1513
rect 1123 -1553 1127 -1549
rect 1105 -1574 1109 -1571
rect 981 -1578 990 -1574
rect 997 -1578 1005 -1574
rect 981 -1581 985 -1578
rect 1005 -1581 1009 -1578
rect 1013 -1578 1025 -1574
rect 1039 -1578 1047 -1574
rect 1013 -1581 1017 -1578
rect 1047 -1581 1051 -1578
rect 1055 -1578 1067 -1574
rect 1081 -1578 1093 -1574
rect 1055 -1581 1059 -1578
rect 1089 -1581 1093 -1578
rect 1097 -1578 1109 -1574
rect 1123 -1574 1127 -1557
rect 1147 -1560 1151 -1513
rect 1147 -1574 1151 -1564
rect 1123 -1578 1135 -1574
rect 1097 -1581 1101 -1578
rect 1131 -1581 1135 -1578
rect 1139 -1578 1151 -1574
rect 1139 -1581 1143 -1578
rect 972 -1589 976 -1585
rect 989 -1589 993 -1585
rect 1030 -1589 1034 -1585
rect 1072 -1589 1076 -1585
rect 1114 -1589 1118 -1585
rect 1155 -1589 1159 -1585
rect 972 -1626 976 -1622
rect 989 -1626 993 -1622
rect 1009 -1626 1013 -1622
rect 1030 -1626 1034 -1622
rect 1051 -1626 1055 -1622
rect 1072 -1626 1076 -1622
rect 1093 -1626 1097 -1622
rect 1114 -1626 1118 -1622
rect 1135 -1626 1139 -1622
rect 1155 -1626 1159 -1622
rect 963 -1681 967 -1634
rect 963 -1702 967 -1685
rect 981 -1695 985 -1634
rect 997 -1695 1001 -1634
rect 1021 -1674 1025 -1634
rect 1021 -1695 1025 -1678
rect 1039 -1695 1043 -1634
rect 1063 -1681 1067 -1634
rect 1063 -1695 1067 -1685
rect 1081 -1674 1085 -1634
rect 1081 -1695 1085 -1678
rect 1105 -1688 1109 -1634
rect 1123 -1666 1127 -1634
rect 1123 -1674 1127 -1670
rect 1105 -1695 1109 -1692
rect 981 -1699 990 -1695
rect 997 -1699 1005 -1695
rect 981 -1702 985 -1699
rect 1005 -1702 1009 -1699
rect 1013 -1699 1025 -1695
rect 1039 -1699 1047 -1695
rect 1013 -1702 1017 -1699
rect 1047 -1702 1051 -1699
rect 1055 -1699 1067 -1695
rect 1081 -1699 1093 -1695
rect 1055 -1702 1059 -1699
rect 1089 -1702 1093 -1699
rect 1097 -1699 1109 -1695
rect 1123 -1695 1127 -1678
rect 1147 -1681 1151 -1634
rect 1147 -1695 1151 -1685
rect 1123 -1699 1135 -1695
rect 1097 -1702 1101 -1699
rect 1131 -1702 1135 -1699
rect 1139 -1699 1151 -1695
rect 1139 -1702 1143 -1699
rect 972 -1710 976 -1706
rect 989 -1710 993 -1706
rect 1030 -1710 1034 -1706
rect 1072 -1710 1076 -1706
rect 1114 -1710 1118 -1706
rect 1155 -1710 1159 -1706
rect 1161 -1717 1165 -1670
rect 1309 -1674 1313 -1484
rect 972 -1747 976 -1743
rect 989 -1747 993 -1743
rect 1009 -1747 1013 -1743
rect 1030 -1747 1034 -1743
rect 1051 -1747 1055 -1743
rect 1072 -1747 1076 -1743
rect 1093 -1747 1097 -1743
rect 1114 -1747 1118 -1743
rect 1135 -1747 1139 -1743
rect 1155 -1747 1159 -1743
rect 1203 -1747 1207 -1743
rect 963 -1802 967 -1755
rect 963 -1823 967 -1806
rect 981 -1816 985 -1755
rect 997 -1816 1001 -1755
rect 1021 -1795 1025 -1755
rect 1021 -1816 1025 -1799
rect 1039 -1816 1043 -1755
rect 1063 -1802 1067 -1755
rect 1063 -1816 1067 -1806
rect 1081 -1795 1085 -1755
rect 1081 -1816 1085 -1799
rect 1105 -1809 1109 -1755
rect 1123 -1787 1127 -1755
rect 1123 -1795 1127 -1791
rect 1105 -1816 1109 -1813
rect 981 -1820 990 -1816
rect 997 -1820 1005 -1816
rect 981 -1823 985 -1820
rect 1005 -1823 1009 -1820
rect 1013 -1820 1025 -1816
rect 1039 -1820 1047 -1816
rect 1013 -1823 1017 -1820
rect 1047 -1823 1051 -1820
rect 1055 -1820 1067 -1816
rect 1081 -1820 1093 -1816
rect 1055 -1823 1059 -1820
rect 1089 -1823 1093 -1820
rect 1097 -1820 1109 -1816
rect 1123 -1816 1127 -1799
rect 1147 -1802 1151 -1755
rect 1147 -1816 1151 -1806
rect 1123 -1820 1135 -1816
rect 1097 -1823 1101 -1820
rect 1131 -1823 1135 -1820
rect 1139 -1820 1151 -1816
rect 1139 -1823 1143 -1820
rect 972 -1831 976 -1827
rect 989 -1831 993 -1827
rect 1030 -1831 1034 -1827
rect 1072 -1831 1076 -1827
rect 1114 -1831 1118 -1827
rect 1155 -1831 1159 -1827
rect 963 -1974 967 -1970
rect 980 -1974 984 -1970
rect 971 -1985 975 -1982
rect 971 -1989 986 -1985
rect 957 -2002 964 -1998
rect 574 -2237 578 -2233
rect 591 -2237 595 -2233
rect 611 -2237 615 -2233
rect 632 -2237 636 -2233
rect 653 -2237 657 -2233
rect 674 -2237 678 -2233
rect 695 -2237 699 -2233
rect 716 -2237 720 -2233
rect 737 -2237 741 -2233
rect 757 -2237 761 -2233
rect 565 -2292 569 -2245
rect 565 -2313 569 -2296
rect 583 -2306 587 -2245
rect 599 -2306 603 -2245
rect 623 -2285 627 -2245
rect 623 -2306 627 -2289
rect 641 -2306 645 -2245
rect 665 -2292 669 -2245
rect 665 -2306 669 -2296
rect 683 -2285 687 -2245
rect 683 -2306 687 -2289
rect 707 -2299 711 -2245
rect 725 -2277 729 -2245
rect 725 -2285 729 -2281
rect 707 -2306 711 -2303
rect 583 -2310 592 -2306
rect 599 -2310 607 -2306
rect 583 -2313 587 -2310
rect 607 -2313 611 -2310
rect 615 -2310 627 -2306
rect 641 -2310 649 -2306
rect 615 -2313 619 -2310
rect 649 -2313 653 -2310
rect 657 -2310 669 -2306
rect 683 -2310 695 -2306
rect 657 -2313 661 -2310
rect 691 -2313 695 -2310
rect 699 -2310 711 -2306
rect 725 -2306 729 -2289
rect 749 -2292 753 -2245
rect 749 -2306 753 -2296
rect 725 -2310 737 -2306
rect 699 -2313 703 -2310
rect 733 -2313 737 -2310
rect 741 -2310 753 -2306
rect 741 -2313 745 -2310
rect 574 -2321 578 -2317
rect 591 -2321 595 -2317
rect 632 -2321 636 -2317
rect 674 -2321 678 -2317
rect 716 -2321 720 -2317
rect 757 -2321 761 -2317
rect 574 -2368 578 -2364
rect 591 -2368 595 -2364
rect 611 -2368 615 -2364
rect 632 -2368 636 -2364
rect 653 -2368 657 -2364
rect 674 -2368 678 -2364
rect 695 -2368 699 -2364
rect 716 -2368 720 -2364
rect 737 -2368 741 -2364
rect 757 -2368 761 -2364
rect 565 -2423 569 -2376
rect 565 -2444 569 -2427
rect 583 -2437 587 -2376
rect 599 -2437 603 -2376
rect 623 -2416 627 -2376
rect 623 -2437 627 -2420
rect 641 -2437 645 -2376
rect 665 -2423 669 -2376
rect 665 -2437 669 -2427
rect 683 -2416 687 -2376
rect 683 -2437 687 -2420
rect 707 -2430 711 -2376
rect 725 -2408 729 -2376
rect 725 -2416 729 -2412
rect 707 -2437 711 -2434
rect 583 -2441 592 -2437
rect 599 -2441 607 -2437
rect 583 -2444 587 -2441
rect 607 -2444 611 -2441
rect 615 -2441 627 -2437
rect 641 -2441 649 -2437
rect 615 -2444 619 -2441
rect 649 -2444 653 -2441
rect 657 -2441 669 -2437
rect 683 -2441 695 -2437
rect 657 -2444 661 -2441
rect 691 -2444 695 -2441
rect 699 -2441 711 -2437
rect 725 -2437 729 -2420
rect 749 -2423 753 -2376
rect 749 -2437 753 -2427
rect 725 -2441 737 -2437
rect 699 -2444 703 -2441
rect 733 -2444 737 -2441
rect 741 -2441 753 -2437
rect 741 -2444 745 -2441
rect 574 -2452 578 -2448
rect 591 -2452 595 -2448
rect 632 -2452 636 -2448
rect 674 -2452 678 -2448
rect 716 -2452 720 -2448
rect 757 -2452 761 -2448
rect 763 -2459 767 -2412
rect 951 -2416 955 -2188
rect 574 -2499 578 -2495
rect 591 -2499 595 -2495
rect 611 -2499 615 -2495
rect 632 -2499 636 -2495
rect 653 -2499 657 -2495
rect 674 -2499 678 -2495
rect 695 -2499 699 -2495
rect 716 -2499 720 -2495
rect 737 -2499 741 -2495
rect 757 -2499 761 -2495
rect 565 -2554 569 -2507
rect 565 -2575 569 -2558
rect 583 -2568 587 -2507
rect 599 -2568 603 -2507
rect 623 -2547 627 -2507
rect 623 -2568 627 -2551
rect 641 -2568 645 -2507
rect 665 -2554 669 -2507
rect 665 -2568 669 -2558
rect 683 -2547 687 -2507
rect 683 -2568 687 -2551
rect 707 -2561 711 -2507
rect 725 -2539 729 -2507
rect 725 -2547 729 -2543
rect 707 -2568 711 -2565
rect 583 -2572 592 -2568
rect 599 -2572 607 -2568
rect 583 -2575 587 -2572
rect 607 -2575 611 -2572
rect 615 -2572 627 -2568
rect 641 -2572 649 -2568
rect 615 -2575 619 -2572
rect 649 -2575 653 -2572
rect 657 -2572 669 -2568
rect 683 -2572 695 -2568
rect 657 -2575 661 -2572
rect 691 -2575 695 -2572
rect 699 -2572 711 -2568
rect 725 -2568 729 -2551
rect 749 -2554 753 -2507
rect 749 -2568 753 -2558
rect 725 -2572 737 -2568
rect 699 -2575 703 -2572
rect 733 -2575 737 -2572
rect 741 -2572 753 -2568
rect 741 -2575 745 -2572
rect 574 -2583 578 -2579
rect 591 -2583 595 -2579
rect 632 -2583 636 -2579
rect 674 -2583 678 -2579
rect 716 -2583 720 -2579
rect 757 -2583 761 -2579
rect 565 -2724 569 -2720
rect 582 -2724 586 -2720
rect 573 -2735 577 -2732
rect 573 -2739 588 -2735
rect 559 -2752 566 -2748
rect 218 -2962 222 -2958
rect 235 -2962 239 -2958
rect 255 -2962 259 -2958
rect 276 -2962 280 -2958
rect 297 -2962 301 -2958
rect 318 -2962 322 -2958
rect 339 -2962 343 -2958
rect 360 -2962 364 -2958
rect 381 -2962 385 -2958
rect 401 -2962 405 -2958
rect 472 -2962 476 -2958
rect 209 -3017 213 -2970
rect 209 -3038 213 -3021
rect 227 -3031 231 -2970
rect 243 -3031 247 -2970
rect 267 -3010 271 -2970
rect 267 -3031 271 -3014
rect 285 -3031 289 -2970
rect 309 -3017 313 -2970
rect 309 -3031 313 -3021
rect 327 -3010 331 -2970
rect 327 -3031 331 -3014
rect 351 -3024 355 -2970
rect 369 -3002 373 -2970
rect 369 -3010 373 -3006
rect 351 -3031 355 -3028
rect 227 -3035 236 -3031
rect 243 -3035 251 -3031
rect 227 -3038 231 -3035
rect 251 -3038 255 -3035
rect 259 -3035 271 -3031
rect 285 -3035 293 -3031
rect 259 -3038 263 -3035
rect 293 -3038 297 -3035
rect 301 -3035 313 -3031
rect 327 -3035 339 -3031
rect 301 -3038 305 -3035
rect 335 -3038 339 -3035
rect 343 -3035 355 -3031
rect 369 -3031 373 -3014
rect 393 -3017 397 -2970
rect 480 -3003 484 -2970
rect 393 -3031 397 -3021
rect 369 -3035 381 -3031
rect 343 -3038 347 -3035
rect 377 -3038 381 -3035
rect 385 -3035 397 -3031
rect 385 -3038 389 -3035
rect 480 -3038 484 -3007
rect 218 -3046 222 -3042
rect 235 -3046 239 -3042
rect 276 -3046 280 -3042
rect 318 -3046 322 -3042
rect 360 -3046 364 -3042
rect 401 -3046 405 -3042
rect 472 -3046 476 -3042
rect 218 -3078 222 -3074
rect 235 -3078 239 -3074
rect 255 -3078 259 -3074
rect 276 -3078 280 -3074
rect 297 -3078 301 -3074
rect 318 -3078 322 -3074
rect 339 -3078 343 -3074
rect 360 -3078 364 -3074
rect 381 -3078 385 -3074
rect 401 -3078 405 -3074
rect 472 -3078 476 -3074
rect 209 -3133 213 -3086
rect 209 -3154 213 -3137
rect 227 -3147 231 -3086
rect 243 -3147 247 -3086
rect 267 -3126 271 -3086
rect 267 -3147 271 -3130
rect 285 -3147 289 -3086
rect 309 -3133 313 -3086
rect 309 -3147 313 -3137
rect 327 -3126 331 -3086
rect 327 -3147 331 -3130
rect 351 -3140 355 -3086
rect 369 -3118 373 -3086
rect 369 -3126 373 -3122
rect 351 -3147 355 -3144
rect 227 -3151 236 -3147
rect 243 -3151 251 -3147
rect 227 -3154 231 -3151
rect 251 -3154 255 -3151
rect 259 -3151 271 -3147
rect 285 -3151 293 -3147
rect 259 -3154 263 -3151
rect 293 -3154 297 -3151
rect 301 -3151 313 -3147
rect 327 -3151 339 -3147
rect 301 -3154 305 -3151
rect 335 -3154 339 -3151
rect 343 -3151 355 -3147
rect 369 -3147 373 -3130
rect 393 -3133 397 -3086
rect 393 -3147 397 -3137
rect 369 -3151 381 -3147
rect 343 -3154 347 -3151
rect 377 -3154 381 -3151
rect 385 -3151 397 -3147
rect 385 -3154 389 -3151
rect 218 -3162 222 -3158
rect 235 -3162 239 -3158
rect 276 -3162 280 -3158
rect 318 -3162 322 -3158
rect 360 -3162 364 -3158
rect 401 -3162 405 -3158
rect 407 -3169 411 -3122
rect 480 -3119 484 -3086
rect 480 -3154 484 -3123
rect 553 -3126 557 -2945
rect 472 -3162 476 -3158
rect 218 -3199 222 -3195
rect 235 -3199 239 -3195
rect 255 -3199 259 -3195
rect 276 -3199 280 -3195
rect 297 -3199 301 -3195
rect 318 -3199 322 -3195
rect 339 -3199 343 -3195
rect 360 -3199 364 -3195
rect 381 -3199 385 -3195
rect 401 -3199 405 -3195
rect 209 -3254 213 -3207
rect 209 -3275 213 -3258
rect 227 -3268 231 -3207
rect 243 -3268 247 -3207
rect 267 -3247 271 -3207
rect 267 -3268 271 -3251
rect 285 -3268 289 -3207
rect 309 -3254 313 -3207
rect 309 -3268 313 -3258
rect 327 -3247 331 -3207
rect 327 -3268 331 -3251
rect 351 -3261 355 -3207
rect 369 -3239 373 -3207
rect 369 -3247 373 -3243
rect 351 -3268 355 -3265
rect 227 -3272 236 -3268
rect 243 -3272 251 -3268
rect 227 -3275 231 -3272
rect 251 -3275 255 -3272
rect 259 -3272 271 -3268
rect 285 -3272 293 -3268
rect 259 -3275 263 -3272
rect 293 -3275 297 -3272
rect 301 -3272 313 -3268
rect 327 -3272 339 -3268
rect 301 -3275 305 -3272
rect 335 -3275 339 -3272
rect 343 -3272 355 -3268
rect 369 -3268 373 -3251
rect 393 -3254 397 -3207
rect 393 -3268 397 -3258
rect 369 -3272 381 -3268
rect 343 -3275 347 -3272
rect 377 -3275 381 -3272
rect 385 -3272 397 -3268
rect 385 -3275 389 -3272
rect 218 -3283 222 -3279
rect 235 -3283 239 -3279
rect 276 -3283 280 -3279
rect 318 -3283 322 -3279
rect 360 -3283 364 -3279
rect 401 -3283 405 -3279
rect 209 -3430 213 -3426
rect 226 -3430 230 -3426
rect 217 -3441 221 -3438
rect 217 -3445 232 -3441
rect 203 -3458 210 -3454
rect -210 -3684 -206 -3680
rect -193 -3684 -189 -3680
rect -173 -3684 -169 -3680
rect -152 -3684 -148 -3680
rect -131 -3684 -127 -3680
rect -110 -3684 -106 -3680
rect -89 -3684 -85 -3680
rect -68 -3684 -64 -3680
rect -47 -3684 -43 -3680
rect -27 -3684 -23 -3680
rect -219 -3739 -215 -3692
rect -219 -3760 -215 -3743
rect -201 -3753 -197 -3692
rect -185 -3753 -181 -3692
rect -161 -3732 -157 -3692
rect -161 -3753 -157 -3736
rect -143 -3753 -139 -3692
rect -119 -3739 -115 -3692
rect -119 -3753 -115 -3743
rect -101 -3732 -97 -3692
rect -101 -3753 -97 -3736
rect -77 -3746 -73 -3692
rect -59 -3724 -55 -3692
rect -59 -3732 -55 -3728
rect -77 -3753 -73 -3750
rect -201 -3757 -192 -3753
rect -185 -3757 -177 -3753
rect -201 -3760 -197 -3757
rect -177 -3760 -173 -3757
rect -169 -3757 -157 -3753
rect -143 -3757 -135 -3753
rect -169 -3760 -165 -3757
rect -135 -3760 -131 -3757
rect -127 -3757 -115 -3753
rect -101 -3757 -89 -3753
rect -127 -3760 -123 -3757
rect -93 -3760 -89 -3757
rect -85 -3757 -73 -3753
rect -59 -3753 -55 -3736
rect -35 -3739 -31 -3692
rect -35 -3753 -31 -3743
rect -59 -3757 -47 -3753
rect -85 -3760 -81 -3757
rect -51 -3760 -47 -3757
rect -43 -3757 -31 -3753
rect -43 -3760 -39 -3757
rect -210 -3768 -206 -3764
rect -193 -3768 -189 -3764
rect -152 -3768 -148 -3764
rect -110 -3768 -106 -3764
rect -68 -3768 -64 -3764
rect -27 -3768 -23 -3764
rect 68 -3799 72 -3795
rect 76 -3842 80 -3831
rect 76 -3863 80 -3846
rect 68 -3883 72 -3879
rect -210 -3915 -206 -3911
rect -193 -3915 -189 -3911
rect -173 -3915 -169 -3911
rect -152 -3915 -148 -3911
rect -131 -3915 -127 -3911
rect -110 -3915 -106 -3911
rect -89 -3915 -85 -3911
rect -68 -3915 -64 -3911
rect -47 -3915 -43 -3911
rect -27 -3915 -23 -3911
rect -219 -3970 -215 -3923
rect -219 -3991 -215 -3974
rect -201 -3984 -197 -3923
rect -185 -3984 -181 -3923
rect -161 -3963 -157 -3923
rect -161 -3984 -157 -3967
rect -143 -3984 -139 -3923
rect -119 -3970 -115 -3923
rect -119 -3984 -115 -3974
rect -101 -3963 -97 -3923
rect -101 -3984 -97 -3967
rect -77 -3977 -73 -3923
rect -59 -3955 -55 -3923
rect -59 -3963 -55 -3959
rect -77 -3984 -73 -3981
rect -201 -3988 -192 -3984
rect -185 -3988 -177 -3984
rect -201 -3991 -197 -3988
rect -177 -3991 -173 -3988
rect -169 -3988 -157 -3984
rect -143 -3988 -135 -3984
rect -169 -3991 -165 -3988
rect -135 -3991 -131 -3988
rect -127 -3988 -115 -3984
rect -101 -3988 -89 -3984
rect -127 -3991 -123 -3988
rect -93 -3991 -89 -3988
rect -85 -3988 -73 -3984
rect -59 -3984 -55 -3967
rect -35 -3970 -31 -3923
rect -35 -3984 -31 -3974
rect -59 -3988 -47 -3984
rect -85 -3991 -81 -3988
rect -51 -3991 -47 -3988
rect -43 -3988 -31 -3984
rect -43 -3991 -39 -3988
rect -210 -3999 -206 -3995
rect -193 -3999 -189 -3995
rect -152 -3999 -148 -3995
rect -110 -3999 -106 -3995
rect -68 -3999 -64 -3995
rect -27 -3999 -23 -3995
rect -21 -4006 -17 -3959
rect 197 -3963 201 -3649
rect -210 -4040 -206 -4036
rect -193 -4040 -189 -4036
rect -173 -4040 -169 -4036
rect -152 -4040 -148 -4036
rect -131 -4040 -127 -4036
rect -110 -4040 -106 -4036
rect -89 -4040 -85 -4036
rect -68 -4040 -64 -4036
rect -47 -4040 -43 -4036
rect -27 -4040 -23 -4036
rect -219 -4095 -215 -4048
rect -219 -4116 -215 -4099
rect -201 -4109 -197 -4048
rect -185 -4109 -181 -4048
rect -161 -4088 -157 -4048
rect -161 -4109 -157 -4092
rect -143 -4109 -139 -4048
rect -119 -4095 -115 -4048
rect -119 -4109 -115 -4099
rect -101 -4088 -97 -4048
rect -101 -4109 -97 -4092
rect -77 -4102 -73 -4048
rect -59 -4080 -55 -4048
rect -59 -4088 -55 -4084
rect -77 -4109 -73 -4106
rect -201 -4113 -192 -4109
rect -185 -4113 -177 -4109
rect -201 -4116 -197 -4113
rect -177 -4116 -173 -4113
rect -169 -4113 -157 -4109
rect -143 -4113 -135 -4109
rect -169 -4116 -165 -4113
rect -135 -4116 -131 -4113
rect -127 -4113 -115 -4109
rect -101 -4113 -89 -4109
rect -127 -4116 -123 -4113
rect -93 -4116 -89 -4113
rect -85 -4113 -73 -4109
rect -59 -4109 -55 -4092
rect -35 -4095 -31 -4048
rect -35 -4109 -31 -4099
rect -59 -4113 -47 -4109
rect -85 -4116 -81 -4113
rect -51 -4116 -47 -4113
rect -43 -4113 -31 -4109
rect -43 -4116 -39 -4113
rect -210 -4124 -206 -4120
rect -193 -4124 -189 -4120
rect -152 -4124 -148 -4120
rect -110 -4124 -106 -4120
rect -68 -4124 -64 -4120
rect -27 -4124 -23 -4120
rect -210 -4164 -206 -4160
rect -193 -4164 -189 -4160
rect -173 -4164 -169 -4160
rect -152 -4164 -148 -4160
rect -131 -4164 -127 -4160
rect -110 -4164 -106 -4160
rect -89 -4164 -85 -4160
rect -68 -4164 -64 -4160
rect -47 -4164 -43 -4160
rect -27 -4164 -23 -4160
rect -219 -4219 -215 -4172
rect -219 -4240 -215 -4223
rect -201 -4233 -197 -4172
rect -185 -4233 -181 -4172
rect -161 -4212 -157 -4172
rect -161 -4233 -157 -4216
rect -143 -4233 -139 -4172
rect -119 -4219 -115 -4172
rect -119 -4233 -115 -4223
rect -101 -4212 -97 -4172
rect -101 -4233 -97 -4216
rect -77 -4226 -73 -4172
rect -59 -4204 -55 -4172
rect -59 -4212 -55 -4208
rect -77 -4233 -73 -4230
rect -201 -4237 -192 -4233
rect -185 -4237 -177 -4233
rect -201 -4240 -197 -4237
rect -177 -4240 -173 -4237
rect -169 -4237 -157 -4233
rect -143 -4237 -135 -4233
rect -169 -4240 -165 -4237
rect -135 -4240 -131 -4237
rect -127 -4237 -115 -4233
rect -101 -4237 -89 -4233
rect -127 -4240 -123 -4237
rect -93 -4240 -89 -4237
rect -85 -4237 -73 -4233
rect -59 -4233 -55 -4216
rect -35 -4219 -31 -4172
rect -35 -4233 -31 -4223
rect -59 -4237 -47 -4233
rect -85 -4240 -81 -4237
rect -51 -4240 -47 -4237
rect -43 -4237 -31 -4233
rect -43 -4240 -39 -4237
rect -210 -4248 -206 -4244
rect -193 -4248 -189 -4244
rect -152 -4248 -148 -4244
rect -110 -4248 -106 -4244
rect -68 -4248 -64 -4244
rect -27 -4248 -23 -4244
rect -219 -4275 -215 -4271
rect -202 -4275 -198 -4271
rect -211 -4286 -207 -4283
rect -211 -4290 -196 -4286
rect -225 -4303 -218 -4299
rect -568 -4517 -564 -4513
rect -551 -4517 -547 -4513
rect -531 -4517 -527 -4513
rect -510 -4517 -506 -4513
rect -489 -4517 -485 -4513
rect -468 -4517 -464 -4513
rect -447 -4517 -443 -4513
rect -426 -4517 -422 -4513
rect -405 -4517 -401 -4513
rect -385 -4517 -381 -4513
rect -577 -4572 -573 -4525
rect -577 -4593 -573 -4576
rect -559 -4586 -555 -4525
rect -543 -4586 -539 -4525
rect -519 -4565 -515 -4525
rect -519 -4586 -515 -4569
rect -501 -4586 -497 -4525
rect -477 -4572 -473 -4525
rect -477 -4586 -473 -4576
rect -459 -4565 -455 -4525
rect -459 -4586 -455 -4569
rect -435 -4579 -431 -4525
rect -417 -4557 -413 -4525
rect -417 -4565 -413 -4561
rect -435 -4586 -431 -4583
rect -559 -4590 -550 -4586
rect -543 -4590 -535 -4586
rect -559 -4593 -555 -4590
rect -535 -4593 -531 -4590
rect -527 -4590 -515 -4586
rect -501 -4590 -493 -4586
rect -527 -4593 -523 -4590
rect -493 -4593 -489 -4590
rect -485 -4590 -473 -4586
rect -459 -4590 -447 -4586
rect -485 -4593 -481 -4590
rect -451 -4593 -447 -4590
rect -443 -4590 -431 -4586
rect -417 -4586 -413 -4569
rect -393 -4572 -389 -4525
rect -393 -4586 -389 -4576
rect -417 -4590 -405 -4586
rect -443 -4593 -439 -4590
rect -409 -4593 -405 -4590
rect -401 -4590 -389 -4586
rect -401 -4593 -397 -4590
rect -568 -4601 -564 -4597
rect -551 -4601 -547 -4597
rect -510 -4601 -506 -4597
rect -468 -4601 -464 -4597
rect -426 -4601 -422 -4597
rect -385 -4601 -381 -4597
rect -568 -4638 -564 -4634
rect -551 -4638 -547 -4634
rect -531 -4638 -527 -4634
rect -510 -4638 -506 -4634
rect -489 -4638 -485 -4634
rect -468 -4638 -464 -4634
rect -447 -4638 -443 -4634
rect -426 -4638 -422 -4634
rect -405 -4638 -401 -4634
rect -385 -4638 -381 -4634
rect -577 -4693 -573 -4646
rect -577 -4714 -573 -4697
rect -559 -4707 -555 -4646
rect -543 -4707 -539 -4646
rect -519 -4686 -515 -4646
rect -519 -4707 -515 -4690
rect -501 -4707 -497 -4646
rect -477 -4693 -473 -4646
rect -477 -4707 -473 -4697
rect -459 -4686 -455 -4646
rect -459 -4707 -455 -4690
rect -435 -4700 -431 -4646
rect -417 -4678 -413 -4646
rect -417 -4686 -413 -4682
rect -435 -4707 -431 -4704
rect -559 -4711 -550 -4707
rect -543 -4711 -535 -4707
rect -559 -4714 -555 -4711
rect -535 -4714 -531 -4711
rect -527 -4711 -515 -4707
rect -501 -4711 -493 -4707
rect -527 -4714 -523 -4711
rect -493 -4714 -489 -4711
rect -485 -4711 -473 -4707
rect -459 -4711 -447 -4707
rect -485 -4714 -481 -4711
rect -451 -4714 -447 -4711
rect -443 -4711 -431 -4707
rect -417 -4707 -413 -4690
rect -393 -4693 -389 -4646
rect -393 -4707 -389 -4697
rect -417 -4711 -405 -4707
rect -443 -4714 -439 -4711
rect -409 -4714 -405 -4711
rect -401 -4711 -389 -4707
rect -401 -4714 -397 -4711
rect -568 -4722 -564 -4718
rect -551 -4722 -547 -4718
rect -510 -4722 -506 -4718
rect -468 -4722 -464 -4718
rect -426 -4722 -422 -4718
rect -385 -4722 -381 -4718
rect -379 -4729 -375 -4682
rect -231 -4686 -227 -4496
rect -568 -4759 -564 -4755
rect -551 -4759 -547 -4755
rect -531 -4759 -527 -4755
rect -510 -4759 -506 -4755
rect -489 -4759 -485 -4755
rect -468 -4759 -464 -4755
rect -447 -4759 -443 -4755
rect -426 -4759 -422 -4755
rect -405 -4759 -401 -4755
rect -385 -4759 -381 -4755
rect -577 -4814 -573 -4767
rect -577 -4835 -573 -4818
rect -559 -4828 -555 -4767
rect -543 -4828 -539 -4767
rect -519 -4807 -515 -4767
rect -519 -4828 -515 -4811
rect -501 -4828 -497 -4767
rect -477 -4814 -473 -4767
rect -477 -4828 -473 -4818
rect -459 -4807 -455 -4767
rect -459 -4828 -455 -4811
rect -435 -4821 -431 -4767
rect -417 -4799 -413 -4767
rect -417 -4807 -413 -4803
rect -435 -4828 -431 -4825
rect -559 -4832 -550 -4828
rect -543 -4832 -535 -4828
rect -559 -4835 -555 -4832
rect -535 -4835 -531 -4832
rect -527 -4832 -515 -4828
rect -501 -4832 -493 -4828
rect -527 -4835 -523 -4832
rect -493 -4835 -489 -4832
rect -485 -4832 -473 -4828
rect -459 -4832 -447 -4828
rect -485 -4835 -481 -4832
rect -451 -4835 -447 -4832
rect -443 -4832 -431 -4828
rect -417 -4828 -413 -4811
rect -393 -4814 -389 -4767
rect -393 -4828 -389 -4818
rect -417 -4832 -405 -4828
rect -443 -4835 -439 -4832
rect -409 -4835 -405 -4832
rect -401 -4832 -389 -4828
rect -401 -4835 -397 -4832
rect -568 -4843 -564 -4839
rect -551 -4843 -547 -4839
rect -510 -4843 -506 -4839
rect -468 -4843 -464 -4839
rect -426 -4843 -422 -4839
rect -385 -4843 -381 -4839
rect -568 -4877 -564 -4873
rect -551 -4877 -547 -4873
rect -531 -4877 -527 -4873
rect -510 -4877 -506 -4873
rect -489 -4877 -485 -4873
rect -468 -4877 -464 -4873
rect -447 -4877 -443 -4873
rect -426 -4877 -422 -4873
rect -405 -4877 -401 -4873
rect -385 -4877 -381 -4873
rect -577 -4932 -573 -4885
rect -577 -4953 -573 -4936
rect -559 -4946 -555 -4885
rect -543 -4946 -539 -4885
rect -519 -4925 -515 -4885
rect -519 -4946 -515 -4929
rect -501 -4946 -497 -4885
rect -477 -4932 -473 -4885
rect -477 -4946 -473 -4936
rect -459 -4925 -455 -4885
rect -459 -4946 -455 -4929
rect -435 -4939 -431 -4885
rect -417 -4917 -413 -4885
rect -417 -4925 -413 -4921
rect -435 -4946 -431 -4943
rect -559 -4950 -550 -4946
rect -543 -4950 -535 -4946
rect -559 -4953 -555 -4950
rect -535 -4953 -531 -4950
rect -527 -4950 -515 -4946
rect -501 -4950 -493 -4946
rect -527 -4953 -523 -4950
rect -493 -4953 -489 -4950
rect -485 -4950 -473 -4946
rect -459 -4950 -447 -4946
rect -485 -4953 -481 -4950
rect -451 -4953 -447 -4950
rect -443 -4950 -431 -4946
rect -417 -4946 -413 -4929
rect -393 -4932 -389 -4885
rect -393 -4946 -389 -4936
rect -417 -4950 -405 -4946
rect -443 -4953 -439 -4950
rect -409 -4953 -405 -4950
rect -401 -4950 -389 -4946
rect -401 -4953 -397 -4950
rect -568 -4961 -564 -4957
rect -551 -4961 -547 -4957
rect -510 -4961 -506 -4957
rect -468 -4961 -464 -4957
rect -426 -4961 -422 -4957
rect -385 -4961 -381 -4957
rect -577 -4994 -573 -4990
rect -560 -4994 -556 -4990
rect -569 -5005 -565 -5002
rect -569 -5009 -554 -5005
rect -583 -5022 -576 -5018
rect -926 -5232 -922 -5228
rect -909 -5232 -905 -5228
rect -889 -5232 -885 -5228
rect -868 -5232 -864 -5228
rect -847 -5232 -843 -5228
rect -826 -5232 -822 -5228
rect -805 -5232 -801 -5228
rect -784 -5232 -780 -5228
rect -763 -5232 -759 -5228
rect -743 -5232 -739 -5228
rect -935 -5287 -931 -5240
rect -935 -5308 -931 -5291
rect -917 -5301 -913 -5240
rect -901 -5301 -897 -5240
rect -877 -5280 -873 -5240
rect -877 -5301 -873 -5284
rect -859 -5301 -855 -5240
rect -835 -5287 -831 -5240
rect -835 -5301 -831 -5291
rect -817 -5280 -813 -5240
rect -817 -5301 -813 -5284
rect -793 -5294 -789 -5240
rect -775 -5272 -771 -5240
rect -775 -5280 -771 -5276
rect -793 -5301 -789 -5298
rect -917 -5305 -908 -5301
rect -901 -5305 -893 -5301
rect -917 -5308 -913 -5305
rect -893 -5308 -889 -5305
rect -885 -5305 -873 -5301
rect -859 -5305 -851 -5301
rect -885 -5308 -881 -5305
rect -851 -5308 -847 -5305
rect -843 -5305 -831 -5301
rect -817 -5305 -805 -5301
rect -843 -5308 -839 -5305
rect -809 -5308 -805 -5305
rect -801 -5305 -789 -5301
rect -775 -5301 -771 -5284
rect -751 -5287 -747 -5240
rect -751 -5301 -747 -5291
rect -775 -5305 -763 -5301
rect -801 -5308 -797 -5305
rect -767 -5308 -763 -5305
rect -759 -5305 -747 -5301
rect -759 -5308 -755 -5305
rect -926 -5316 -922 -5312
rect -909 -5316 -905 -5312
rect -868 -5316 -864 -5312
rect -826 -5316 -822 -5312
rect -784 -5316 -780 -5312
rect -743 -5316 -739 -5312
rect -926 -5353 -922 -5349
rect -909 -5353 -905 -5349
rect -889 -5353 -885 -5349
rect -868 -5353 -864 -5349
rect -847 -5353 -843 -5349
rect -826 -5353 -822 -5349
rect -805 -5353 -801 -5349
rect -784 -5353 -780 -5349
rect -763 -5353 -759 -5349
rect -743 -5353 -739 -5349
rect -673 -5353 -669 -5349
rect -935 -5408 -931 -5361
rect -935 -5429 -931 -5412
rect -917 -5422 -913 -5361
rect -901 -5422 -897 -5361
rect -877 -5401 -873 -5361
rect -877 -5422 -873 -5405
rect -859 -5422 -855 -5361
rect -835 -5408 -831 -5361
rect -835 -5422 -831 -5412
rect -817 -5401 -813 -5361
rect -817 -5422 -813 -5405
rect -793 -5415 -789 -5361
rect -775 -5393 -771 -5361
rect -775 -5401 -771 -5397
rect -793 -5422 -789 -5419
rect -917 -5426 -908 -5422
rect -901 -5426 -893 -5422
rect -917 -5429 -913 -5426
rect -893 -5429 -889 -5426
rect -885 -5426 -873 -5422
rect -859 -5426 -851 -5422
rect -885 -5429 -881 -5426
rect -851 -5429 -847 -5426
rect -843 -5426 -831 -5422
rect -817 -5426 -805 -5422
rect -843 -5429 -839 -5426
rect -809 -5429 -805 -5426
rect -801 -5426 -789 -5422
rect -775 -5422 -771 -5405
rect -751 -5408 -747 -5361
rect -751 -5422 -747 -5412
rect -775 -5426 -763 -5422
rect -801 -5429 -797 -5426
rect -767 -5429 -763 -5426
rect -759 -5426 -747 -5422
rect -759 -5429 -755 -5426
rect -926 -5437 -922 -5433
rect -909 -5437 -905 -5433
rect -868 -5437 -864 -5433
rect -826 -5437 -822 -5433
rect -784 -5437 -780 -5433
rect -743 -5437 -739 -5433
rect -737 -5444 -733 -5397
rect -665 -5395 -661 -5369
rect -665 -5425 -661 -5399
rect -589 -5401 -585 -5208
rect -673 -5437 -669 -5433
rect -926 -5473 -922 -5469
rect -909 -5473 -905 -5469
rect -889 -5473 -885 -5469
rect -868 -5473 -864 -5469
rect -847 -5473 -843 -5469
rect -826 -5473 -822 -5469
rect -805 -5473 -801 -5469
rect -784 -5473 -780 -5469
rect -763 -5473 -759 -5469
rect -743 -5473 -739 -5469
rect -935 -5528 -931 -5481
rect -935 -5549 -931 -5532
rect -917 -5542 -913 -5481
rect -901 -5542 -897 -5481
rect -877 -5521 -873 -5481
rect -877 -5542 -873 -5525
rect -859 -5542 -855 -5481
rect -835 -5528 -831 -5481
rect -835 -5542 -831 -5532
rect -817 -5521 -813 -5481
rect -817 -5542 -813 -5525
rect -793 -5535 -789 -5481
rect -775 -5513 -771 -5481
rect -775 -5521 -771 -5517
rect -793 -5542 -789 -5539
rect -917 -5546 -908 -5542
rect -901 -5546 -893 -5542
rect -917 -5549 -913 -5546
rect -893 -5549 -889 -5546
rect -885 -5546 -873 -5542
rect -859 -5546 -851 -5542
rect -885 -5549 -881 -5546
rect -851 -5549 -847 -5546
rect -843 -5546 -831 -5542
rect -817 -5546 -805 -5542
rect -843 -5549 -839 -5546
rect -809 -5549 -805 -5546
rect -801 -5546 -789 -5542
rect -775 -5542 -771 -5525
rect -751 -5528 -747 -5481
rect -751 -5542 -747 -5532
rect -775 -5546 -763 -5542
rect -801 -5549 -797 -5546
rect -767 -5549 -763 -5546
rect -759 -5546 -747 -5542
rect -759 -5549 -755 -5546
rect -926 -5557 -922 -5553
rect -909 -5557 -905 -5553
rect -868 -5557 -864 -5553
rect -826 -5557 -822 -5553
rect -784 -5557 -780 -5553
rect -743 -5557 -739 -5553
rect -926 -5590 -922 -5586
rect -909 -5590 -905 -5586
rect -889 -5590 -885 -5586
rect -868 -5590 -864 -5586
rect -847 -5590 -843 -5586
rect -826 -5590 -822 -5586
rect -805 -5590 -801 -5586
rect -784 -5590 -780 -5586
rect -763 -5590 -759 -5586
rect -743 -5590 -739 -5586
rect -935 -5645 -931 -5598
rect -935 -5666 -931 -5649
rect -917 -5659 -913 -5598
rect -901 -5659 -897 -5598
rect -877 -5638 -873 -5598
rect -877 -5659 -873 -5642
rect -859 -5659 -855 -5598
rect -835 -5645 -831 -5598
rect -835 -5659 -831 -5649
rect -817 -5638 -813 -5598
rect -817 -5659 -813 -5642
rect -793 -5652 -789 -5598
rect -775 -5630 -771 -5598
rect -775 -5638 -771 -5634
rect -793 -5659 -789 -5656
rect -917 -5663 -908 -5659
rect -901 -5663 -893 -5659
rect -917 -5666 -913 -5663
rect -893 -5666 -889 -5663
rect -885 -5663 -873 -5659
rect -859 -5663 -851 -5659
rect -885 -5666 -881 -5663
rect -851 -5666 -847 -5663
rect -843 -5663 -831 -5659
rect -817 -5663 -805 -5659
rect -843 -5666 -839 -5663
rect -809 -5666 -805 -5663
rect -801 -5663 -789 -5659
rect -775 -5659 -771 -5642
rect -751 -5645 -747 -5598
rect -751 -5659 -747 -5649
rect -775 -5663 -763 -5659
rect -801 -5666 -797 -5663
rect -767 -5666 -763 -5663
rect -759 -5663 -747 -5659
rect -759 -5666 -755 -5663
rect -926 -5674 -922 -5670
rect -909 -5674 -905 -5670
rect -868 -5674 -864 -5670
rect -826 -5674 -822 -5670
rect -784 -5674 -780 -5670
rect -743 -5674 -739 -5670
rect -935 -5707 -931 -5703
rect -918 -5707 -914 -5703
rect -927 -5718 -923 -5715
rect -927 -5722 -912 -5718
rect -916 -5761 -912 -5722
rect -916 -5776 -912 -5765
rect -935 -5780 -912 -5776
rect -909 -5752 -905 -5715
rect -737 -5731 -733 -5517
rect -935 -5783 -931 -5780
rect -909 -5783 -905 -5756
rect -918 -5791 -914 -5787
rect -926 -5826 -922 -5822
rect -900 -5826 -896 -5822
rect -883 -5826 -879 -5822
rect -843 -5826 -839 -5822
rect -822 -5826 -818 -5822
rect -805 -5826 -801 -5822
rect -765 -5826 -761 -5822
rect -741 -5826 -737 -5822
rect -704 -5826 -700 -5822
rect -935 -5851 -931 -5834
rect -1255 -5910 -1251 -5906
rect -1211 -5910 -1207 -5906
rect -1177 -5910 -1173 -5906
rect -1162 -5920 -1158 -5892
rect -935 -5902 -931 -5855
rect -917 -5844 -913 -5834
rect -917 -5902 -913 -5848
rect -909 -5873 -905 -5834
rect -891 -5866 -887 -5834
rect -909 -5902 -905 -5877
rect -891 -5902 -887 -5870
rect -865 -5858 -861 -5834
rect -865 -5895 -861 -5862
rect -831 -5895 -827 -5834
rect -813 -5851 -809 -5834
rect -883 -5902 -879 -5899
rect -875 -5899 -861 -5895
rect -875 -5902 -871 -5899
rect -847 -5902 -843 -5899
rect -839 -5899 -820 -5895
rect -839 -5902 -835 -5899
rect -813 -5902 -809 -5855
rect -787 -5866 -783 -5834
rect -787 -5895 -783 -5870
rect -753 -5888 -749 -5834
rect -753 -5892 -736 -5888
rect -805 -5902 -801 -5899
rect -796 -5899 -783 -5895
rect -796 -5902 -792 -5899
rect -769 -5902 -765 -5899
rect -745 -5902 -741 -5892
rect -729 -5895 -725 -5834
rect -721 -5888 -717 -5834
rect -695 -5858 -691 -5834
rect -721 -5892 -702 -5888
rect -737 -5899 -720 -5895
rect -737 -5902 -733 -5899
rect -713 -5902 -709 -5892
rect -695 -5902 -691 -5862
rect -926 -5910 -922 -5906
rect -900 -5910 -896 -5906
rect -857 -5910 -853 -5906
rect -822 -5910 -818 -5906
rect -778 -5910 -774 -5906
rect -761 -5910 -757 -5906
rect -725 -5910 -721 -5906
rect -704 -5910 -700 -5906
rect -689 -5917 -685 -5870
rect -595 -5873 -591 -5756
rect -589 -5858 -585 -5449
rect -583 -5521 -579 -5022
rect -558 -5048 -554 -5009
rect -558 -5063 -554 -5052
rect -577 -5067 -554 -5063
rect -551 -5039 -547 -5002
rect -379 -5018 -375 -4803
rect -577 -5070 -573 -5067
rect -551 -5070 -547 -5043
rect -560 -5078 -556 -5074
rect -568 -5113 -564 -5109
rect -542 -5113 -538 -5109
rect -525 -5113 -521 -5109
rect -485 -5113 -481 -5109
rect -464 -5113 -460 -5109
rect -447 -5113 -443 -5109
rect -407 -5113 -403 -5109
rect -383 -5113 -379 -5109
rect -346 -5113 -342 -5109
rect -577 -5138 -573 -5121
rect -577 -5189 -573 -5142
rect -559 -5131 -555 -5121
rect -559 -5189 -555 -5135
rect -551 -5160 -547 -5121
rect -533 -5153 -529 -5121
rect -551 -5189 -547 -5164
rect -533 -5189 -529 -5157
rect -507 -5145 -503 -5121
rect -507 -5182 -503 -5149
rect -473 -5182 -469 -5121
rect -455 -5138 -451 -5121
rect -525 -5189 -521 -5186
rect -517 -5186 -503 -5182
rect -517 -5189 -513 -5186
rect -489 -5189 -485 -5186
rect -481 -5186 -462 -5182
rect -481 -5189 -477 -5186
rect -455 -5189 -451 -5142
rect -429 -5153 -425 -5121
rect -429 -5182 -425 -5157
rect -395 -5175 -391 -5121
rect -395 -5179 -378 -5175
rect -447 -5189 -443 -5186
rect -438 -5186 -425 -5182
rect -438 -5189 -434 -5186
rect -411 -5189 -407 -5186
rect -387 -5189 -383 -5179
rect -371 -5182 -367 -5121
rect -363 -5175 -359 -5121
rect -337 -5144 -333 -5121
rect -363 -5179 -344 -5175
rect -379 -5186 -362 -5182
rect -379 -5189 -375 -5186
rect -355 -5189 -351 -5179
rect -337 -5189 -333 -5148
rect -568 -5197 -564 -5193
rect -542 -5197 -538 -5193
rect -499 -5197 -495 -5193
rect -464 -5197 -460 -5193
rect -420 -5197 -416 -5193
rect -403 -5197 -399 -5193
rect -367 -5197 -363 -5193
rect -346 -5197 -342 -5193
rect -331 -5211 -327 -5157
rect -237 -5160 -233 -5043
rect -231 -5145 -227 -4733
rect -225 -4807 -221 -4303
rect -200 -4329 -196 -4290
rect -200 -4344 -196 -4333
rect -219 -4348 -196 -4344
rect -193 -4320 -189 -4283
rect -21 -4307 -17 -4208
rect -15 -4299 -11 -4084
rect -219 -4351 -215 -4348
rect -193 -4351 -189 -4324
rect -202 -4359 -198 -4355
rect -210 -4394 -206 -4390
rect -184 -4394 -180 -4390
rect -167 -4394 -163 -4390
rect -127 -4394 -123 -4390
rect -106 -4394 -102 -4390
rect -89 -4394 -85 -4390
rect -49 -4394 -45 -4390
rect -25 -4394 -21 -4390
rect 12 -4394 16 -4390
rect -219 -4419 -215 -4402
rect -219 -4470 -215 -4423
rect -201 -4412 -197 -4402
rect -201 -4470 -197 -4416
rect -193 -4441 -189 -4402
rect -175 -4434 -171 -4402
rect -193 -4470 -189 -4445
rect -175 -4470 -171 -4438
rect -149 -4426 -145 -4402
rect -149 -4463 -145 -4430
rect -115 -4463 -111 -4402
rect -97 -4419 -93 -4402
rect -167 -4470 -163 -4467
rect -159 -4467 -145 -4463
rect -159 -4470 -155 -4467
rect -131 -4470 -127 -4467
rect -123 -4467 -104 -4463
rect -123 -4470 -119 -4467
rect -97 -4470 -93 -4423
rect -71 -4434 -67 -4402
rect -71 -4463 -67 -4438
rect -37 -4456 -33 -4402
rect -37 -4460 -20 -4456
rect -89 -4470 -85 -4467
rect -80 -4467 -67 -4463
rect -80 -4470 -76 -4467
rect -53 -4470 -49 -4467
rect -29 -4470 -25 -4460
rect -13 -4463 -9 -4402
rect -5 -4456 -1 -4402
rect 21 -4426 25 -4402
rect -5 -4460 14 -4456
rect -21 -4467 -4 -4463
rect -21 -4470 -17 -4467
rect 3 -4470 7 -4460
rect 21 -4470 25 -4430
rect -210 -4478 -206 -4474
rect -184 -4478 -180 -4474
rect -141 -4478 -137 -4474
rect -106 -4478 -102 -4474
rect -62 -4478 -58 -4474
rect -45 -4478 -41 -4474
rect -9 -4478 -5 -4474
rect 12 -4478 16 -4474
rect 27 -4485 31 -4438
rect 191 -4441 195 -4324
rect 197 -4426 201 -4010
rect 203 -4088 207 -3458
rect 228 -3484 232 -3445
rect 228 -3499 232 -3488
rect 209 -3503 232 -3499
rect 235 -3475 239 -3438
rect 407 -3454 411 -3243
rect 209 -3506 213 -3503
rect 235 -3506 239 -3479
rect 226 -3514 230 -3510
rect 218 -3554 222 -3550
rect 244 -3554 248 -3550
rect 261 -3554 265 -3550
rect 301 -3554 305 -3550
rect 322 -3554 326 -3550
rect 339 -3554 343 -3550
rect 379 -3554 383 -3550
rect 403 -3554 407 -3550
rect 440 -3554 444 -3550
rect 209 -3579 213 -3562
rect 209 -3630 213 -3583
rect 227 -3572 231 -3562
rect 227 -3630 231 -3576
rect 235 -3601 239 -3562
rect 253 -3594 257 -3562
rect 235 -3630 239 -3605
rect 253 -3630 257 -3598
rect 279 -3586 283 -3562
rect 279 -3623 283 -3590
rect 313 -3623 317 -3562
rect 331 -3579 335 -3562
rect 261 -3630 265 -3627
rect 269 -3627 283 -3623
rect 269 -3630 273 -3627
rect 297 -3630 301 -3627
rect 305 -3627 324 -3623
rect 305 -3630 309 -3627
rect 331 -3630 335 -3583
rect 357 -3594 361 -3562
rect 357 -3623 361 -3598
rect 391 -3616 395 -3562
rect 391 -3620 408 -3616
rect 339 -3630 343 -3627
rect 348 -3627 361 -3623
rect 348 -3630 352 -3627
rect 375 -3630 379 -3627
rect 399 -3630 403 -3620
rect 415 -3623 419 -3562
rect 423 -3616 427 -3562
rect 449 -3586 453 -3562
rect 423 -3620 442 -3616
rect 407 -3627 424 -3623
rect 407 -3630 411 -3627
rect 431 -3630 435 -3620
rect 449 -3630 453 -3590
rect 218 -3638 222 -3634
rect 244 -3638 248 -3634
rect 287 -3638 291 -3634
rect 322 -3638 326 -3634
rect 366 -3638 370 -3634
rect 383 -3638 387 -3634
rect 419 -3638 423 -3634
rect 440 -3638 444 -3634
rect 455 -3652 459 -3598
rect 547 -3601 551 -3479
rect 553 -3586 557 -3173
rect 559 -3247 563 -2752
rect 584 -2778 588 -2739
rect 584 -2793 588 -2782
rect 565 -2797 588 -2793
rect 591 -2769 595 -2732
rect 763 -2748 767 -2543
rect 565 -2800 569 -2797
rect 591 -2800 595 -2773
rect 582 -2808 586 -2804
rect 574 -2843 578 -2839
rect 600 -2843 604 -2839
rect 617 -2843 621 -2839
rect 657 -2843 661 -2839
rect 678 -2843 682 -2839
rect 695 -2843 699 -2839
rect 735 -2843 739 -2839
rect 759 -2843 763 -2839
rect 796 -2843 800 -2839
rect 565 -2868 569 -2851
rect 565 -2919 569 -2872
rect 583 -2861 587 -2851
rect 583 -2919 587 -2865
rect 591 -2890 595 -2851
rect 609 -2883 613 -2851
rect 591 -2919 595 -2894
rect 609 -2919 613 -2887
rect 635 -2875 639 -2851
rect 635 -2912 639 -2879
rect 669 -2912 673 -2851
rect 687 -2868 691 -2851
rect 617 -2919 621 -2916
rect 625 -2916 639 -2912
rect 625 -2919 629 -2916
rect 653 -2919 657 -2916
rect 661 -2916 680 -2912
rect 661 -2919 665 -2916
rect 687 -2919 691 -2872
rect 713 -2883 717 -2851
rect 713 -2912 717 -2887
rect 747 -2905 751 -2851
rect 747 -2909 764 -2905
rect 695 -2919 699 -2916
rect 704 -2916 717 -2912
rect 704 -2919 708 -2916
rect 731 -2919 735 -2916
rect 755 -2919 759 -2909
rect 771 -2912 775 -2851
rect 779 -2905 783 -2851
rect 805 -2875 809 -2851
rect 779 -2909 798 -2905
rect 763 -2916 780 -2912
rect 763 -2919 767 -2916
rect 787 -2919 791 -2909
rect 805 -2919 809 -2879
rect 574 -2927 578 -2923
rect 600 -2927 604 -2923
rect 643 -2927 647 -2923
rect 678 -2927 682 -2923
rect 722 -2927 726 -2923
rect 739 -2927 743 -2923
rect 775 -2927 779 -2923
rect 796 -2927 800 -2923
rect 811 -2934 815 -2887
rect 945 -2890 949 -2773
rect 951 -2875 955 -2464
rect 957 -2547 961 -2002
rect 982 -2028 986 -1989
rect 982 -2043 986 -2032
rect 963 -2047 986 -2043
rect 989 -2019 993 -1982
rect 1161 -1998 1165 -1791
rect 1211 -1788 1215 -1755
rect 1211 -1823 1215 -1792
rect 1203 -1831 1207 -1827
rect 1203 -1862 1207 -1858
rect 1211 -1903 1215 -1870
rect 1211 -1938 1215 -1907
rect 1203 -1946 1207 -1942
rect 963 -2050 967 -2047
rect 989 -2050 993 -2023
rect 980 -2058 984 -2054
rect 972 -2093 976 -2089
rect 998 -2093 1002 -2089
rect 1015 -2093 1019 -2089
rect 1055 -2093 1059 -2089
rect 1076 -2093 1080 -2089
rect 1093 -2093 1097 -2089
rect 1133 -2093 1137 -2089
rect 1157 -2093 1161 -2089
rect 1194 -2093 1198 -2089
rect 963 -2118 967 -2101
rect 963 -2169 967 -2122
rect 981 -2111 985 -2101
rect 981 -2169 985 -2115
rect 989 -2140 993 -2101
rect 1007 -2133 1011 -2101
rect 989 -2169 993 -2144
rect 1007 -2169 1011 -2137
rect 1033 -2125 1037 -2101
rect 1033 -2162 1037 -2129
rect 1067 -2162 1071 -2101
rect 1085 -2118 1089 -2101
rect 1015 -2169 1019 -2166
rect 1023 -2166 1037 -2162
rect 1023 -2169 1027 -2166
rect 1051 -2169 1055 -2166
rect 1059 -2166 1078 -2162
rect 1059 -2169 1063 -2166
rect 1085 -2169 1089 -2122
rect 1111 -2133 1115 -2101
rect 1111 -2162 1115 -2137
rect 1145 -2155 1149 -2101
rect 1145 -2159 1162 -2155
rect 1093 -2169 1097 -2166
rect 1102 -2166 1115 -2162
rect 1102 -2169 1106 -2166
rect 1129 -2169 1133 -2166
rect 1153 -2169 1157 -2159
rect 1169 -2162 1173 -2101
rect 1177 -2155 1181 -2101
rect 1203 -2123 1207 -2101
rect 1177 -2159 1196 -2155
rect 1161 -2166 1178 -2162
rect 1161 -2169 1165 -2166
rect 1185 -2169 1189 -2159
rect 1203 -2169 1207 -2127
rect 1303 -2125 1307 -2023
rect 972 -2177 976 -2173
rect 998 -2177 1002 -2173
rect 1041 -2177 1045 -2173
rect 1076 -2177 1080 -2173
rect 1120 -2177 1124 -2173
rect 1137 -2177 1141 -2173
rect 1173 -2177 1177 -2173
rect 1194 -2177 1198 -2173
rect 1209 -2191 1213 -2137
rect 1309 -2140 1313 -1722
rect 1315 -1795 1319 -1296
rect 1340 -1322 1344 -1283
rect 1340 -1337 1344 -1326
rect 1321 -1341 1344 -1337
rect 1347 -1313 1351 -1276
rect 1321 -1344 1325 -1341
rect 1347 -1344 1351 -1317
rect 1338 -1352 1342 -1348
rect 1330 -1382 1334 -1378
rect 1347 -1382 1351 -1378
rect 1387 -1382 1391 -1378
rect 1408 -1382 1412 -1378
rect 1321 -1423 1325 -1390
rect 1321 -1458 1325 -1427
rect 1339 -1417 1343 -1390
rect 1339 -1421 1348 -1417
rect 1339 -1458 1343 -1421
rect 1365 -1444 1369 -1390
rect 1365 -1451 1369 -1448
rect 1399 -1451 1403 -1390
rect 1347 -1458 1351 -1455
rect 1356 -1455 1369 -1451
rect 1356 -1458 1360 -1455
rect 1383 -1458 1387 -1455
rect 1391 -1455 1410 -1451
rect 1391 -1458 1395 -1455
rect 1417 -1458 1421 -1390
rect 1330 -1466 1334 -1462
rect 1374 -1466 1378 -1462
rect 1408 -1466 1412 -1462
rect 1417 -1480 1421 -1462
rect 1423 -1487 1427 -1448
rect 1330 -1626 1334 -1622
rect 1347 -1626 1351 -1622
rect 1367 -1626 1371 -1622
rect 1388 -1626 1392 -1622
rect 1409 -1626 1413 -1622
rect 1430 -1626 1434 -1622
rect 1451 -1626 1455 -1622
rect 1472 -1626 1476 -1622
rect 1493 -1626 1497 -1622
rect 1513 -1626 1517 -1622
rect 1321 -1681 1325 -1634
rect 1321 -1702 1325 -1685
rect 1339 -1695 1343 -1634
rect 1355 -1695 1359 -1634
rect 1379 -1674 1383 -1634
rect 1379 -1695 1383 -1678
rect 1397 -1695 1401 -1634
rect 1421 -1681 1425 -1634
rect 1421 -1695 1425 -1685
rect 1439 -1674 1443 -1634
rect 1439 -1695 1443 -1678
rect 1463 -1688 1467 -1634
rect 1481 -1666 1485 -1634
rect 1481 -1674 1485 -1670
rect 1463 -1695 1467 -1692
rect 1339 -1699 1348 -1695
rect 1355 -1699 1363 -1695
rect 1339 -1702 1343 -1699
rect 1363 -1702 1367 -1699
rect 1371 -1699 1383 -1695
rect 1397 -1699 1405 -1695
rect 1371 -1702 1375 -1699
rect 1405 -1702 1409 -1699
rect 1413 -1699 1425 -1695
rect 1439 -1699 1451 -1695
rect 1413 -1702 1417 -1699
rect 1447 -1702 1451 -1699
rect 1455 -1699 1467 -1695
rect 1481 -1695 1485 -1678
rect 1505 -1681 1509 -1634
rect 1505 -1695 1509 -1685
rect 1481 -1699 1493 -1695
rect 1455 -1702 1459 -1699
rect 1489 -1702 1493 -1699
rect 1497 -1699 1509 -1695
rect 1497 -1702 1501 -1699
rect 1330 -1710 1334 -1706
rect 1347 -1710 1351 -1706
rect 1388 -1710 1392 -1706
rect 1430 -1710 1434 -1706
rect 1472 -1710 1476 -1706
rect 1513 -1710 1517 -1706
rect 1519 -1718 1523 -1670
rect 1330 -1747 1334 -1743
rect 1347 -1747 1351 -1743
rect 1367 -1747 1371 -1743
rect 1388 -1747 1392 -1743
rect 1409 -1747 1413 -1743
rect 1430 -1747 1434 -1743
rect 1451 -1747 1455 -1743
rect 1472 -1747 1476 -1743
rect 1493 -1747 1497 -1743
rect 1513 -1747 1517 -1743
rect 1321 -1802 1325 -1755
rect 1321 -1823 1325 -1806
rect 1339 -1816 1343 -1755
rect 1355 -1816 1359 -1755
rect 1379 -1795 1383 -1755
rect 1379 -1816 1383 -1799
rect 1397 -1816 1401 -1755
rect 1421 -1802 1425 -1755
rect 1421 -1816 1425 -1806
rect 1439 -1795 1443 -1755
rect 1439 -1816 1443 -1799
rect 1463 -1809 1467 -1755
rect 1481 -1787 1485 -1755
rect 1481 -1795 1485 -1791
rect 1463 -1816 1467 -1813
rect 1339 -1820 1348 -1816
rect 1355 -1820 1363 -1816
rect 1339 -1823 1343 -1820
rect 1363 -1823 1367 -1820
rect 1371 -1820 1383 -1816
rect 1397 -1820 1405 -1816
rect 1371 -1823 1375 -1820
rect 1405 -1823 1409 -1820
rect 1413 -1820 1425 -1816
rect 1439 -1820 1451 -1816
rect 1413 -1823 1417 -1820
rect 1447 -1823 1451 -1820
rect 1455 -1820 1467 -1816
rect 1481 -1816 1485 -1799
rect 1505 -1802 1509 -1755
rect 1505 -1816 1509 -1806
rect 1481 -1820 1493 -1816
rect 1455 -1823 1459 -1820
rect 1489 -1823 1493 -1820
rect 1497 -1820 1509 -1816
rect 1497 -1823 1501 -1820
rect 1330 -1831 1334 -1827
rect 1347 -1831 1351 -1827
rect 1388 -1831 1392 -1827
rect 1430 -1831 1434 -1827
rect 1472 -1831 1476 -1827
rect 1513 -1831 1517 -1827
rect 1321 -1974 1325 -1970
rect 1338 -1974 1342 -1970
rect 1329 -1985 1333 -1982
rect 1329 -1989 1344 -1985
rect 1315 -2002 1322 -1998
rect 972 -2368 976 -2364
rect 989 -2368 993 -2364
rect 1009 -2368 1013 -2364
rect 1030 -2368 1034 -2364
rect 1051 -2368 1055 -2364
rect 1072 -2368 1076 -2364
rect 1093 -2368 1097 -2364
rect 1114 -2368 1118 -2364
rect 1135 -2368 1139 -2364
rect 1155 -2368 1159 -2364
rect 963 -2423 967 -2376
rect 963 -2444 967 -2427
rect 981 -2437 985 -2376
rect 997 -2437 1001 -2376
rect 1021 -2416 1025 -2376
rect 1021 -2437 1025 -2420
rect 1039 -2437 1043 -2376
rect 1063 -2423 1067 -2376
rect 1063 -2437 1067 -2427
rect 1081 -2416 1085 -2376
rect 1081 -2437 1085 -2420
rect 1105 -2430 1109 -2376
rect 1123 -2408 1127 -2376
rect 1123 -2416 1127 -2412
rect 1105 -2437 1109 -2434
rect 981 -2441 990 -2437
rect 997 -2441 1005 -2437
rect 981 -2444 985 -2441
rect 1005 -2444 1009 -2441
rect 1013 -2441 1025 -2437
rect 1039 -2441 1047 -2437
rect 1013 -2444 1017 -2441
rect 1047 -2444 1051 -2441
rect 1055 -2441 1067 -2437
rect 1081 -2441 1093 -2437
rect 1055 -2444 1059 -2441
rect 1089 -2444 1093 -2441
rect 1097 -2441 1109 -2437
rect 1123 -2437 1127 -2420
rect 1147 -2423 1151 -2376
rect 1147 -2437 1151 -2427
rect 1123 -2441 1135 -2437
rect 1097 -2444 1101 -2441
rect 1131 -2444 1135 -2441
rect 1139 -2441 1151 -2437
rect 1139 -2444 1143 -2441
rect 972 -2452 976 -2448
rect 989 -2452 993 -2448
rect 1030 -2452 1034 -2448
rect 1072 -2452 1076 -2448
rect 1114 -2452 1118 -2448
rect 1155 -2452 1159 -2448
rect 1161 -2460 1165 -2412
rect 1309 -2416 1313 -2195
rect 972 -2499 976 -2495
rect 989 -2499 993 -2495
rect 1009 -2499 1013 -2495
rect 1030 -2499 1034 -2495
rect 1051 -2499 1055 -2495
rect 1072 -2499 1076 -2495
rect 1093 -2499 1097 -2495
rect 1114 -2499 1118 -2495
rect 1135 -2499 1139 -2495
rect 1155 -2499 1159 -2495
rect 963 -2554 967 -2507
rect 963 -2575 967 -2558
rect 981 -2568 985 -2507
rect 997 -2568 1001 -2507
rect 1021 -2547 1025 -2507
rect 1021 -2568 1025 -2551
rect 1039 -2568 1043 -2507
rect 1063 -2554 1067 -2507
rect 1063 -2568 1067 -2558
rect 1081 -2547 1085 -2507
rect 1081 -2568 1085 -2551
rect 1105 -2561 1109 -2507
rect 1123 -2539 1127 -2507
rect 1123 -2547 1127 -2543
rect 1105 -2568 1109 -2565
rect 981 -2572 990 -2568
rect 997 -2572 1005 -2568
rect 981 -2575 985 -2572
rect 1005 -2575 1009 -2572
rect 1013 -2572 1025 -2568
rect 1039 -2572 1047 -2568
rect 1013 -2575 1017 -2572
rect 1047 -2575 1051 -2572
rect 1055 -2572 1067 -2568
rect 1081 -2572 1093 -2568
rect 1055 -2575 1059 -2572
rect 1089 -2575 1093 -2572
rect 1097 -2572 1109 -2568
rect 1123 -2568 1127 -2551
rect 1147 -2554 1151 -2507
rect 1147 -2568 1151 -2558
rect 1123 -2572 1135 -2568
rect 1097 -2575 1101 -2572
rect 1131 -2575 1135 -2572
rect 1139 -2572 1151 -2568
rect 1139 -2575 1143 -2572
rect 972 -2583 976 -2579
rect 989 -2583 993 -2579
rect 1030 -2583 1034 -2579
rect 1072 -2583 1076 -2579
rect 1114 -2583 1118 -2579
rect 1155 -2583 1159 -2579
rect 963 -2724 967 -2720
rect 980 -2724 984 -2720
rect 971 -2735 975 -2732
rect 971 -2739 986 -2735
rect 957 -2752 964 -2748
rect 841 -2962 845 -2958
rect 849 -3003 853 -2978
rect 849 -3034 853 -3007
rect 841 -3046 845 -3042
rect 574 -3078 578 -3074
rect 591 -3078 595 -3074
rect 611 -3078 615 -3074
rect 632 -3078 636 -3074
rect 653 -3078 657 -3074
rect 674 -3078 678 -3074
rect 695 -3078 699 -3074
rect 716 -3078 720 -3074
rect 737 -3078 741 -3074
rect 757 -3078 761 -3074
rect 565 -3133 569 -3086
rect 565 -3154 569 -3137
rect 583 -3147 587 -3086
rect 599 -3147 603 -3086
rect 623 -3126 627 -3086
rect 623 -3147 627 -3130
rect 641 -3147 645 -3086
rect 665 -3133 669 -3086
rect 665 -3147 669 -3137
rect 683 -3126 687 -3086
rect 683 -3147 687 -3130
rect 707 -3140 711 -3086
rect 725 -3118 729 -3086
rect 725 -3126 729 -3122
rect 707 -3147 711 -3144
rect 583 -3151 592 -3147
rect 599 -3151 607 -3147
rect 583 -3154 587 -3151
rect 607 -3154 611 -3151
rect 615 -3151 627 -3147
rect 641 -3151 649 -3147
rect 615 -3154 619 -3151
rect 649 -3154 653 -3151
rect 657 -3151 669 -3147
rect 683 -3151 695 -3147
rect 657 -3154 661 -3151
rect 691 -3154 695 -3151
rect 699 -3151 711 -3147
rect 725 -3147 729 -3130
rect 749 -3133 753 -3086
rect 749 -3147 753 -3137
rect 725 -3151 737 -3147
rect 699 -3154 703 -3151
rect 733 -3154 737 -3151
rect 741 -3151 753 -3147
rect 741 -3154 745 -3151
rect 574 -3162 578 -3158
rect 591 -3162 595 -3158
rect 632 -3162 636 -3158
rect 674 -3162 678 -3158
rect 716 -3162 720 -3158
rect 757 -3162 761 -3158
rect 763 -3169 767 -3122
rect 951 -3126 955 -2938
rect 574 -3199 578 -3195
rect 591 -3199 595 -3195
rect 611 -3199 615 -3195
rect 632 -3199 636 -3195
rect 653 -3199 657 -3195
rect 674 -3199 678 -3195
rect 695 -3199 699 -3195
rect 716 -3199 720 -3195
rect 737 -3199 741 -3195
rect 757 -3199 761 -3195
rect 565 -3254 569 -3207
rect 565 -3275 569 -3258
rect 583 -3268 587 -3207
rect 599 -3268 603 -3207
rect 623 -3247 627 -3207
rect 623 -3268 627 -3251
rect 641 -3268 645 -3207
rect 665 -3254 669 -3207
rect 665 -3268 669 -3258
rect 683 -3247 687 -3207
rect 683 -3268 687 -3251
rect 707 -3261 711 -3207
rect 725 -3239 729 -3207
rect 725 -3247 729 -3243
rect 707 -3268 711 -3265
rect 583 -3272 592 -3268
rect 599 -3272 607 -3268
rect 583 -3275 587 -3272
rect 607 -3275 611 -3272
rect 615 -3272 627 -3268
rect 641 -3272 649 -3268
rect 615 -3275 619 -3272
rect 649 -3275 653 -3272
rect 657 -3272 669 -3268
rect 683 -3272 695 -3268
rect 657 -3275 661 -3272
rect 691 -3275 695 -3272
rect 699 -3272 711 -3268
rect 725 -3268 729 -3251
rect 749 -3254 753 -3207
rect 749 -3268 753 -3258
rect 725 -3272 737 -3268
rect 699 -3275 703 -3272
rect 733 -3275 737 -3272
rect 741 -3272 753 -3268
rect 741 -3275 745 -3272
rect 574 -3283 578 -3279
rect 591 -3283 595 -3279
rect 632 -3283 636 -3279
rect 674 -3283 678 -3279
rect 716 -3283 720 -3279
rect 757 -3283 761 -3279
rect 565 -3430 569 -3426
rect 582 -3430 586 -3426
rect 573 -3441 577 -3438
rect 573 -3445 588 -3441
rect 559 -3458 566 -3454
rect 218 -3915 222 -3911
rect 235 -3915 239 -3911
rect 255 -3915 259 -3911
rect 276 -3915 280 -3911
rect 297 -3915 301 -3911
rect 318 -3915 322 -3911
rect 339 -3915 343 -3911
rect 360 -3915 364 -3911
rect 381 -3915 385 -3911
rect 401 -3915 405 -3911
rect 209 -3970 213 -3923
rect 209 -3991 213 -3974
rect 227 -3984 231 -3923
rect 243 -3984 247 -3923
rect 267 -3963 271 -3923
rect 267 -3984 271 -3967
rect 285 -3984 289 -3923
rect 309 -3970 313 -3923
rect 309 -3984 313 -3974
rect 327 -3963 331 -3923
rect 327 -3984 331 -3967
rect 351 -3977 355 -3923
rect 369 -3955 373 -3923
rect 369 -3963 373 -3959
rect 351 -3984 355 -3981
rect 227 -3988 236 -3984
rect 243 -3988 251 -3984
rect 227 -3991 231 -3988
rect 251 -3991 255 -3988
rect 259 -3988 271 -3984
rect 285 -3988 293 -3984
rect 259 -3991 263 -3988
rect 293 -3991 297 -3988
rect 301 -3988 313 -3984
rect 327 -3988 339 -3984
rect 301 -3991 305 -3988
rect 335 -3991 339 -3988
rect 343 -3988 355 -3984
rect 369 -3984 373 -3967
rect 393 -3970 397 -3923
rect 393 -3984 397 -3974
rect 369 -3988 381 -3984
rect 343 -3991 347 -3988
rect 377 -3991 381 -3988
rect 385 -3988 397 -3984
rect 385 -3991 389 -3988
rect 218 -3999 222 -3995
rect 235 -3999 239 -3995
rect 276 -3999 280 -3995
rect 318 -3999 322 -3995
rect 360 -3999 364 -3995
rect 401 -3999 405 -3995
rect 407 -4006 411 -3959
rect 553 -3963 557 -3656
rect 218 -4040 222 -4036
rect 235 -4040 239 -4036
rect 255 -4040 259 -4036
rect 276 -4040 280 -4036
rect 297 -4040 301 -4036
rect 318 -4040 322 -4036
rect 339 -4040 343 -4036
rect 360 -4040 364 -4036
rect 381 -4040 385 -4036
rect 401 -4040 405 -4036
rect 209 -4095 213 -4048
rect 209 -4116 213 -4099
rect 227 -4109 231 -4048
rect 243 -4109 247 -4048
rect 267 -4088 271 -4048
rect 267 -4109 271 -4092
rect 285 -4109 289 -4048
rect 309 -4095 313 -4048
rect 309 -4109 313 -4099
rect 327 -4088 331 -4048
rect 327 -4109 331 -4092
rect 351 -4102 355 -4048
rect 369 -4080 373 -4048
rect 369 -4088 373 -4084
rect 351 -4109 355 -4106
rect 227 -4113 236 -4109
rect 243 -4113 251 -4109
rect 227 -4116 231 -4113
rect 251 -4116 255 -4113
rect 259 -4113 271 -4109
rect 285 -4113 293 -4109
rect 259 -4116 263 -4113
rect 293 -4116 297 -4113
rect 301 -4113 313 -4109
rect 327 -4113 339 -4109
rect 301 -4116 305 -4113
rect 335 -4116 339 -4113
rect 343 -4113 355 -4109
rect 369 -4109 373 -4092
rect 393 -4095 397 -4048
rect 393 -4109 397 -4099
rect 369 -4113 381 -4109
rect 343 -4116 347 -4113
rect 377 -4116 381 -4113
rect 385 -4113 397 -4109
rect 385 -4116 389 -4113
rect 218 -4124 222 -4120
rect 235 -4124 239 -4120
rect 276 -4124 280 -4120
rect 318 -4124 322 -4120
rect 360 -4124 364 -4120
rect 401 -4124 405 -4120
rect 209 -4275 213 -4271
rect 226 -4275 230 -4271
rect 217 -4286 221 -4283
rect 217 -4290 232 -4286
rect 203 -4303 210 -4299
rect -210 -4638 -206 -4634
rect -193 -4638 -189 -4634
rect -173 -4638 -169 -4634
rect -152 -4638 -148 -4634
rect -131 -4638 -127 -4634
rect -110 -4638 -106 -4634
rect -89 -4638 -85 -4634
rect -68 -4638 -64 -4634
rect -47 -4638 -43 -4634
rect -27 -4638 -23 -4634
rect -219 -4693 -215 -4646
rect -219 -4714 -215 -4697
rect -201 -4707 -197 -4646
rect -185 -4707 -181 -4646
rect -161 -4686 -157 -4646
rect -161 -4707 -157 -4690
rect -143 -4707 -139 -4646
rect -119 -4693 -115 -4646
rect -119 -4707 -115 -4697
rect -101 -4686 -97 -4646
rect -101 -4707 -97 -4690
rect -77 -4700 -73 -4646
rect -59 -4678 -55 -4646
rect -59 -4686 -55 -4682
rect -77 -4707 -73 -4704
rect -201 -4711 -192 -4707
rect -185 -4711 -177 -4707
rect -201 -4714 -197 -4711
rect -177 -4714 -173 -4711
rect -169 -4711 -157 -4707
rect -143 -4711 -135 -4707
rect -169 -4714 -165 -4711
rect -135 -4714 -131 -4711
rect -127 -4711 -115 -4707
rect -101 -4711 -89 -4707
rect -127 -4714 -123 -4711
rect -93 -4714 -89 -4711
rect -85 -4711 -73 -4707
rect -59 -4707 -55 -4690
rect -35 -4693 -31 -4646
rect -35 -4707 -31 -4697
rect -59 -4711 -47 -4707
rect -85 -4714 -81 -4711
rect -51 -4714 -47 -4711
rect -43 -4711 -31 -4707
rect -43 -4714 -39 -4711
rect -210 -4722 -206 -4718
rect -193 -4722 -189 -4718
rect -152 -4722 -148 -4718
rect -110 -4722 -106 -4718
rect -68 -4722 -64 -4718
rect -27 -4722 -23 -4718
rect -21 -4729 -17 -4682
rect 197 -4686 201 -4489
rect -210 -4759 -206 -4755
rect -193 -4759 -189 -4755
rect -173 -4759 -169 -4755
rect -152 -4759 -148 -4755
rect -131 -4759 -127 -4755
rect -110 -4759 -106 -4755
rect -89 -4759 -85 -4755
rect -68 -4759 -64 -4755
rect -47 -4759 -43 -4755
rect -27 -4759 -23 -4755
rect 90 -4759 94 -4755
rect -219 -4814 -215 -4767
rect -219 -4835 -215 -4818
rect -201 -4828 -197 -4767
rect -185 -4828 -181 -4767
rect -161 -4807 -157 -4767
rect -161 -4828 -157 -4811
rect -143 -4828 -139 -4767
rect -119 -4814 -115 -4767
rect -119 -4828 -115 -4818
rect -101 -4807 -97 -4767
rect -101 -4828 -97 -4811
rect -77 -4821 -73 -4767
rect -59 -4799 -55 -4767
rect -59 -4807 -55 -4803
rect -77 -4828 -73 -4825
rect -201 -4832 -192 -4828
rect -185 -4832 -177 -4828
rect -201 -4835 -197 -4832
rect -177 -4835 -173 -4832
rect -169 -4832 -157 -4828
rect -143 -4832 -135 -4828
rect -169 -4835 -165 -4832
rect -135 -4835 -131 -4832
rect -127 -4832 -115 -4828
rect -101 -4832 -89 -4828
rect -127 -4835 -123 -4832
rect -93 -4835 -89 -4832
rect -85 -4832 -73 -4828
rect -59 -4828 -55 -4811
rect -35 -4814 -31 -4767
rect -35 -4828 -31 -4818
rect -59 -4832 -47 -4828
rect -85 -4835 -81 -4832
rect -51 -4835 -47 -4832
rect -43 -4832 -31 -4828
rect -43 -4835 -39 -4832
rect -210 -4843 -206 -4839
rect -193 -4843 -189 -4839
rect -152 -4843 -148 -4839
rect -110 -4843 -106 -4839
rect -68 -4843 -64 -4839
rect -27 -4843 -23 -4839
rect -210 -4877 -206 -4873
rect -193 -4877 -189 -4873
rect -173 -4877 -169 -4873
rect -152 -4877 -148 -4873
rect -131 -4877 -127 -4873
rect -110 -4877 -106 -4873
rect -89 -4877 -85 -4873
rect -68 -4877 -64 -4873
rect -47 -4877 -43 -4873
rect -27 -4877 -23 -4873
rect -219 -4932 -215 -4885
rect -219 -4953 -215 -4936
rect -201 -4946 -197 -4885
rect -185 -4946 -181 -4885
rect -161 -4925 -157 -4885
rect -161 -4946 -157 -4929
rect -143 -4946 -139 -4885
rect -119 -4932 -115 -4885
rect -119 -4946 -115 -4936
rect -101 -4925 -97 -4885
rect -101 -4946 -97 -4929
rect -77 -4939 -73 -4885
rect -59 -4917 -55 -4885
rect -59 -4925 -55 -4921
rect -77 -4946 -73 -4943
rect -201 -4950 -192 -4946
rect -185 -4950 -177 -4946
rect -201 -4953 -197 -4950
rect -177 -4953 -173 -4950
rect -169 -4950 -157 -4946
rect -143 -4950 -135 -4946
rect -169 -4953 -165 -4950
rect -135 -4953 -131 -4950
rect -127 -4950 -115 -4946
rect -101 -4950 -89 -4946
rect -127 -4953 -123 -4950
rect -93 -4953 -89 -4950
rect -85 -4950 -73 -4946
rect -59 -4946 -55 -4929
rect -35 -4932 -31 -4885
rect -35 -4946 -31 -4936
rect -59 -4950 -47 -4946
rect -85 -4953 -81 -4950
rect -51 -4953 -47 -4950
rect -43 -4950 -31 -4946
rect -43 -4953 -39 -4950
rect -210 -4961 -206 -4957
rect -193 -4961 -189 -4957
rect -152 -4961 -148 -4957
rect -110 -4961 -106 -4957
rect -68 -4961 -64 -4957
rect -27 -4961 -23 -4957
rect -219 -4994 -215 -4990
rect -202 -4994 -198 -4990
rect -211 -5005 -207 -5002
rect -211 -5009 -196 -5005
rect -225 -5022 -218 -5018
rect -568 -5353 -564 -5349
rect -551 -5353 -547 -5349
rect -531 -5353 -527 -5349
rect -510 -5353 -506 -5349
rect -489 -5353 -485 -5349
rect -468 -5353 -464 -5349
rect -447 -5353 -443 -5349
rect -426 -5353 -422 -5349
rect -405 -5353 -401 -5349
rect -385 -5353 -381 -5349
rect -327 -5353 -323 -5349
rect -577 -5408 -573 -5361
rect -577 -5429 -573 -5412
rect -559 -5422 -555 -5361
rect -543 -5422 -539 -5361
rect -519 -5401 -515 -5361
rect -519 -5422 -515 -5405
rect -501 -5422 -497 -5361
rect -477 -5408 -473 -5361
rect -477 -5422 -473 -5412
rect -459 -5401 -455 -5361
rect -459 -5422 -455 -5405
rect -435 -5415 -431 -5361
rect -417 -5393 -413 -5361
rect -417 -5401 -413 -5397
rect -435 -5422 -431 -5419
rect -559 -5426 -550 -5422
rect -543 -5426 -535 -5422
rect -559 -5429 -555 -5426
rect -535 -5429 -531 -5426
rect -527 -5426 -515 -5422
rect -501 -5426 -493 -5422
rect -527 -5429 -523 -5426
rect -493 -5429 -489 -5426
rect -485 -5426 -473 -5422
rect -459 -5426 -447 -5422
rect -485 -5429 -481 -5426
rect -451 -5429 -447 -5426
rect -443 -5426 -431 -5422
rect -417 -5422 -413 -5405
rect -393 -5408 -389 -5361
rect -393 -5422 -389 -5412
rect -417 -5426 -405 -5422
rect -443 -5429 -439 -5426
rect -409 -5429 -405 -5426
rect -401 -5426 -389 -5422
rect -401 -5429 -397 -5426
rect -568 -5437 -564 -5433
rect -551 -5437 -547 -5433
rect -510 -5437 -506 -5433
rect -468 -5437 -464 -5433
rect -426 -5437 -422 -5433
rect -385 -5437 -381 -5433
rect -379 -5445 -375 -5397
rect -319 -5396 -315 -5361
rect -319 -5429 -315 -5400
rect -231 -5401 -227 -5215
rect -327 -5437 -323 -5433
rect -568 -5473 -564 -5469
rect -551 -5473 -547 -5469
rect -531 -5473 -527 -5469
rect -510 -5473 -506 -5469
rect -489 -5473 -485 -5469
rect -468 -5473 -464 -5469
rect -447 -5473 -443 -5469
rect -426 -5473 -422 -5469
rect -405 -5473 -401 -5469
rect -385 -5473 -381 -5469
rect -327 -5473 -323 -5469
rect -577 -5528 -573 -5481
rect -577 -5549 -573 -5532
rect -559 -5542 -555 -5481
rect -543 -5542 -539 -5481
rect -519 -5521 -515 -5481
rect -519 -5542 -515 -5525
rect -501 -5542 -497 -5481
rect -477 -5528 -473 -5481
rect -477 -5542 -473 -5532
rect -459 -5521 -455 -5481
rect -459 -5542 -455 -5525
rect -435 -5535 -431 -5481
rect -417 -5513 -413 -5481
rect -417 -5521 -413 -5517
rect -435 -5542 -431 -5539
rect -559 -5546 -550 -5542
rect -543 -5546 -535 -5542
rect -559 -5549 -555 -5546
rect -535 -5549 -531 -5546
rect -527 -5546 -515 -5542
rect -501 -5546 -493 -5542
rect -527 -5549 -523 -5546
rect -493 -5549 -489 -5546
rect -485 -5546 -473 -5542
rect -459 -5546 -447 -5542
rect -485 -5549 -481 -5546
rect -451 -5549 -447 -5546
rect -443 -5546 -431 -5542
rect -417 -5542 -413 -5525
rect -393 -5528 -389 -5481
rect -393 -5542 -389 -5532
rect -417 -5546 -405 -5542
rect -443 -5549 -439 -5546
rect -409 -5549 -405 -5546
rect -401 -5546 -389 -5542
rect -401 -5549 -397 -5546
rect -568 -5557 -564 -5553
rect -551 -5557 -547 -5553
rect -510 -5557 -506 -5553
rect -468 -5557 -464 -5553
rect -426 -5557 -422 -5553
rect -385 -5557 -381 -5553
rect -568 -5590 -564 -5586
rect -551 -5590 -547 -5586
rect -531 -5590 -527 -5586
rect -510 -5590 -506 -5586
rect -489 -5590 -485 -5586
rect -468 -5590 -464 -5586
rect -447 -5590 -443 -5586
rect -426 -5590 -422 -5586
rect -405 -5590 -401 -5586
rect -385 -5590 -381 -5586
rect -577 -5645 -573 -5598
rect -577 -5666 -573 -5649
rect -559 -5659 -555 -5598
rect -543 -5659 -539 -5598
rect -519 -5638 -515 -5598
rect -519 -5659 -515 -5642
rect -501 -5659 -497 -5598
rect -477 -5645 -473 -5598
rect -477 -5659 -473 -5649
rect -459 -5638 -455 -5598
rect -459 -5659 -455 -5642
rect -435 -5652 -431 -5598
rect -417 -5630 -413 -5598
rect -417 -5638 -413 -5634
rect -435 -5659 -431 -5656
rect -559 -5663 -550 -5659
rect -543 -5663 -535 -5659
rect -559 -5666 -555 -5663
rect -535 -5666 -531 -5663
rect -527 -5663 -515 -5659
rect -501 -5663 -493 -5659
rect -527 -5666 -523 -5663
rect -493 -5666 -489 -5663
rect -485 -5663 -473 -5659
rect -459 -5663 -447 -5659
rect -485 -5666 -481 -5663
rect -451 -5666 -447 -5663
rect -443 -5663 -431 -5659
rect -417 -5659 -413 -5642
rect -393 -5645 -389 -5598
rect -393 -5659 -389 -5649
rect -417 -5663 -405 -5659
rect -443 -5666 -439 -5663
rect -409 -5666 -405 -5663
rect -401 -5663 -389 -5659
rect -401 -5666 -397 -5663
rect -568 -5674 -564 -5670
rect -551 -5674 -547 -5670
rect -510 -5674 -506 -5670
rect -468 -5674 -464 -5670
rect -426 -5674 -422 -5670
rect -385 -5674 -381 -5670
rect -577 -5707 -573 -5703
rect -560 -5707 -556 -5703
rect -569 -5718 -565 -5715
rect -569 -5722 -554 -5718
rect -558 -5761 -554 -5722
rect -558 -5776 -554 -5765
rect -577 -5780 -554 -5776
rect -551 -5752 -547 -5715
rect -379 -5731 -375 -5517
rect -319 -5511 -315 -5481
rect -319 -5549 -315 -5515
rect -327 -5557 -323 -5553
rect -577 -5783 -573 -5780
rect -551 -5783 -547 -5756
rect -560 -5791 -556 -5787
rect -568 -5826 -564 -5822
rect -542 -5826 -538 -5822
rect -525 -5826 -521 -5822
rect -485 -5826 -481 -5822
rect -464 -5826 -460 -5822
rect -447 -5826 -443 -5822
rect -407 -5826 -403 -5822
rect -383 -5826 -379 -5822
rect -346 -5826 -342 -5822
rect -577 -5851 -573 -5834
rect -577 -5902 -573 -5855
rect -559 -5844 -555 -5834
rect -559 -5902 -555 -5848
rect -551 -5873 -547 -5834
rect -533 -5866 -529 -5834
rect -551 -5902 -547 -5877
rect -533 -5902 -529 -5870
rect -507 -5858 -503 -5834
rect -507 -5895 -503 -5862
rect -473 -5895 -469 -5834
rect -455 -5851 -451 -5834
rect -525 -5902 -521 -5899
rect -517 -5899 -503 -5895
rect -517 -5902 -513 -5899
rect -489 -5902 -485 -5899
rect -481 -5899 -462 -5895
rect -481 -5902 -477 -5899
rect -455 -5902 -451 -5855
rect -429 -5866 -425 -5834
rect -429 -5895 -425 -5870
rect -395 -5888 -391 -5834
rect -395 -5892 -378 -5888
rect -447 -5902 -443 -5899
rect -438 -5899 -425 -5895
rect -438 -5902 -434 -5899
rect -411 -5902 -407 -5899
rect -387 -5902 -383 -5892
rect -371 -5895 -367 -5834
rect -363 -5888 -359 -5834
rect -337 -5857 -333 -5834
rect -363 -5892 -344 -5888
rect -379 -5899 -362 -5895
rect -379 -5902 -375 -5899
rect -355 -5902 -351 -5892
rect -337 -5902 -333 -5861
rect -568 -5910 -564 -5906
rect -542 -5910 -538 -5906
rect -499 -5910 -495 -5906
rect -464 -5910 -460 -5906
rect -420 -5910 -416 -5906
rect -403 -5910 -399 -5906
rect -367 -5910 -363 -5906
rect -346 -5910 -342 -5906
rect -331 -5917 -327 -5870
rect -237 -5873 -233 -5756
rect -231 -5858 -227 -5448
rect -225 -5521 -221 -5022
rect -200 -5048 -196 -5009
rect -200 -5063 -196 -5052
rect -219 -5067 -196 -5063
rect -193 -5039 -189 -5002
rect -21 -5018 -17 -4803
rect 98 -4802 102 -4791
rect 98 -4823 102 -4806
rect 90 -4843 94 -4839
rect -219 -5070 -215 -5067
rect -193 -5070 -189 -5043
rect -202 -5078 -198 -5074
rect -210 -5113 -206 -5109
rect -184 -5113 -180 -5109
rect -167 -5113 -163 -5109
rect -127 -5113 -123 -5109
rect -106 -5113 -102 -5109
rect -89 -5113 -85 -5109
rect -49 -5113 -45 -5109
rect -25 -5113 -21 -5109
rect 12 -5113 16 -5109
rect -219 -5138 -215 -5121
rect -219 -5189 -215 -5142
rect -201 -5131 -197 -5121
rect -201 -5189 -197 -5135
rect -193 -5160 -189 -5121
rect -175 -5153 -171 -5121
rect -193 -5189 -189 -5164
rect -175 -5189 -171 -5157
rect -149 -5145 -145 -5121
rect -149 -5182 -145 -5149
rect -115 -5182 -111 -5121
rect -97 -5138 -93 -5121
rect -167 -5189 -163 -5186
rect -159 -5186 -145 -5182
rect -159 -5189 -155 -5186
rect -131 -5189 -127 -5186
rect -123 -5186 -104 -5182
rect -123 -5189 -119 -5186
rect -97 -5189 -93 -5142
rect -71 -5153 -67 -5121
rect -71 -5182 -67 -5157
rect -37 -5175 -33 -5121
rect -37 -5179 -20 -5175
rect -89 -5189 -85 -5186
rect -80 -5186 -67 -5182
rect -80 -5189 -76 -5186
rect -53 -5189 -49 -5186
rect -29 -5189 -25 -5179
rect -13 -5182 -9 -5121
rect -5 -5175 -1 -5121
rect 21 -5145 25 -5121
rect -5 -5179 14 -5175
rect -21 -5186 -4 -5182
rect -21 -5189 -17 -5186
rect 3 -5189 7 -5179
rect 21 -5189 25 -5149
rect -210 -5197 -206 -5193
rect -184 -5197 -180 -5193
rect -141 -5197 -137 -5193
rect -106 -5197 -102 -5193
rect -62 -5197 -58 -5193
rect -45 -5197 -41 -5193
rect -9 -5197 -5 -5193
rect 12 -5197 16 -5193
rect 27 -5204 31 -5157
rect 191 -5160 195 -5043
rect 197 -5145 201 -4735
rect 203 -4807 207 -4303
rect 228 -4329 232 -4290
rect 228 -4344 232 -4333
rect 209 -4348 232 -4344
rect 235 -4320 239 -4283
rect 407 -4299 411 -4084
rect 456 -4164 460 -4160
rect 464 -4201 468 -4172
rect 464 -4240 468 -4205
rect 456 -4248 460 -4244
rect 456 -4275 460 -4271
rect 464 -4316 468 -4283
rect 209 -4351 213 -4348
rect 235 -4351 239 -4324
rect 464 -4351 468 -4320
rect 226 -4359 230 -4355
rect 456 -4359 460 -4355
rect 218 -4394 222 -4390
rect 244 -4394 248 -4390
rect 261 -4394 265 -4390
rect 301 -4394 305 -4390
rect 322 -4394 326 -4390
rect 339 -4394 343 -4390
rect 379 -4394 383 -4390
rect 403 -4394 407 -4390
rect 440 -4394 444 -4390
rect 209 -4419 213 -4402
rect 209 -4470 213 -4423
rect 227 -4412 231 -4402
rect 227 -4470 231 -4416
rect 235 -4441 239 -4402
rect 253 -4434 257 -4402
rect 235 -4470 239 -4445
rect 253 -4470 257 -4438
rect 279 -4426 283 -4402
rect 279 -4463 283 -4430
rect 313 -4463 317 -4402
rect 331 -4419 335 -4402
rect 261 -4470 265 -4467
rect 269 -4467 283 -4463
rect 269 -4470 273 -4467
rect 297 -4470 301 -4467
rect 305 -4467 324 -4463
rect 305 -4470 309 -4467
rect 331 -4470 335 -4423
rect 357 -4434 361 -4402
rect 357 -4463 361 -4438
rect 391 -4456 395 -4402
rect 391 -4460 408 -4456
rect 339 -4470 343 -4467
rect 348 -4467 361 -4463
rect 348 -4470 352 -4467
rect 375 -4470 379 -4467
rect 399 -4470 403 -4460
rect 415 -4463 419 -4402
rect 423 -4456 427 -4402
rect 449 -4426 453 -4402
rect 423 -4460 442 -4456
rect 407 -4467 424 -4463
rect 407 -4470 411 -4467
rect 431 -4470 435 -4460
rect 449 -4470 453 -4430
rect 218 -4478 222 -4474
rect 244 -4478 248 -4474
rect 287 -4478 291 -4474
rect 322 -4478 326 -4474
rect 366 -4478 370 -4474
rect 383 -4478 387 -4474
rect 419 -4478 423 -4474
rect 440 -4478 444 -4474
rect 455 -4492 459 -4438
rect 547 -4441 551 -4324
rect 553 -4426 557 -4011
rect 559 -4088 563 -3458
rect 584 -3484 588 -3445
rect 584 -3499 588 -3488
rect 565 -3503 588 -3499
rect 591 -3475 595 -3438
rect 763 -3454 767 -3243
rect 565 -3506 569 -3503
rect 591 -3506 595 -3479
rect 582 -3514 586 -3510
rect 574 -3554 578 -3550
rect 600 -3554 604 -3550
rect 617 -3554 621 -3550
rect 657 -3554 661 -3550
rect 678 -3554 682 -3550
rect 695 -3554 699 -3550
rect 735 -3554 739 -3550
rect 759 -3554 763 -3550
rect 796 -3554 800 -3550
rect 565 -3579 569 -3562
rect 565 -3630 569 -3583
rect 583 -3572 587 -3562
rect 583 -3630 587 -3576
rect 591 -3601 595 -3562
rect 609 -3594 613 -3562
rect 591 -3630 595 -3605
rect 609 -3630 613 -3598
rect 635 -3586 639 -3562
rect 635 -3623 639 -3590
rect 669 -3623 673 -3562
rect 687 -3579 691 -3562
rect 617 -3630 621 -3627
rect 625 -3627 639 -3623
rect 625 -3630 629 -3627
rect 653 -3630 657 -3627
rect 661 -3627 680 -3623
rect 661 -3630 665 -3627
rect 687 -3630 691 -3583
rect 713 -3594 717 -3562
rect 713 -3623 717 -3598
rect 747 -3616 751 -3562
rect 747 -3620 764 -3616
rect 695 -3630 699 -3627
rect 704 -3627 717 -3623
rect 704 -3630 708 -3627
rect 731 -3630 735 -3627
rect 755 -3630 759 -3620
rect 771 -3623 775 -3562
rect 779 -3616 783 -3562
rect 805 -3586 809 -3562
rect 779 -3620 798 -3616
rect 763 -3627 780 -3623
rect 763 -3630 767 -3627
rect 787 -3630 791 -3620
rect 805 -3630 809 -3590
rect 574 -3638 578 -3634
rect 600 -3638 604 -3634
rect 643 -3638 647 -3634
rect 678 -3638 682 -3634
rect 722 -3638 726 -3634
rect 739 -3638 743 -3634
rect 775 -3638 779 -3634
rect 796 -3638 800 -3634
rect 811 -3645 815 -3598
rect 945 -3601 949 -3479
rect 951 -3586 955 -3173
rect 957 -3247 961 -2752
rect 982 -2778 986 -2739
rect 982 -2793 986 -2782
rect 963 -2797 986 -2793
rect 989 -2769 993 -2732
rect 1161 -2748 1165 -2543
rect 963 -2800 967 -2797
rect 989 -2800 993 -2773
rect 980 -2808 984 -2804
rect 972 -2843 976 -2839
rect 998 -2843 1002 -2839
rect 1015 -2843 1019 -2839
rect 1055 -2843 1059 -2839
rect 1076 -2843 1080 -2839
rect 1093 -2843 1097 -2839
rect 1133 -2843 1137 -2839
rect 1157 -2843 1161 -2839
rect 1194 -2843 1198 -2839
rect 963 -2868 967 -2851
rect 963 -2919 967 -2872
rect 981 -2861 985 -2851
rect 981 -2919 985 -2865
rect 989 -2890 993 -2851
rect 1007 -2883 1011 -2851
rect 989 -2919 993 -2894
rect 1007 -2919 1011 -2887
rect 1033 -2875 1037 -2851
rect 1033 -2912 1037 -2879
rect 1067 -2912 1071 -2851
rect 1085 -2868 1089 -2851
rect 1015 -2919 1019 -2916
rect 1023 -2916 1037 -2912
rect 1023 -2919 1027 -2916
rect 1051 -2919 1055 -2916
rect 1059 -2916 1078 -2912
rect 1059 -2919 1063 -2916
rect 1085 -2919 1089 -2872
rect 1111 -2883 1115 -2851
rect 1111 -2912 1115 -2887
rect 1145 -2905 1149 -2851
rect 1145 -2909 1162 -2905
rect 1093 -2919 1097 -2916
rect 1102 -2916 1115 -2912
rect 1102 -2919 1106 -2916
rect 1129 -2919 1133 -2916
rect 1153 -2919 1157 -2909
rect 1169 -2912 1173 -2851
rect 1177 -2905 1181 -2851
rect 1203 -2873 1207 -2851
rect 1177 -2909 1196 -2905
rect 1161 -2916 1178 -2912
rect 1161 -2919 1165 -2916
rect 1185 -2919 1189 -2909
rect 1203 -2919 1207 -2877
rect 1303 -2875 1307 -2773
rect 972 -2927 976 -2923
rect 998 -2927 1002 -2923
rect 1041 -2927 1045 -2923
rect 1076 -2927 1080 -2923
rect 1120 -2927 1124 -2923
rect 1137 -2927 1141 -2923
rect 1173 -2927 1177 -2923
rect 1194 -2927 1198 -2923
rect 1209 -2941 1213 -2887
rect 1309 -2890 1313 -2464
rect 1315 -2547 1319 -2002
rect 1340 -2028 1344 -1989
rect 1340 -2043 1344 -2032
rect 1321 -2047 1344 -2043
rect 1347 -2019 1351 -1982
rect 1519 -1998 1523 -1791
rect 1321 -2050 1325 -2047
rect 1347 -2050 1351 -2023
rect 1338 -2058 1342 -2054
rect 1330 -2093 1334 -2089
rect 1356 -2093 1360 -2089
rect 1373 -2093 1377 -2089
rect 1413 -2093 1417 -2089
rect 1434 -2093 1438 -2089
rect 1451 -2093 1455 -2089
rect 1491 -2093 1495 -2089
rect 1515 -2093 1519 -2089
rect 1552 -2093 1556 -2089
rect 1321 -2118 1325 -2101
rect 1321 -2169 1325 -2122
rect 1339 -2111 1343 -2101
rect 1339 -2169 1343 -2115
rect 1347 -2140 1351 -2101
rect 1365 -2133 1369 -2101
rect 1347 -2169 1351 -2144
rect 1365 -2169 1369 -2137
rect 1391 -2125 1395 -2101
rect 1391 -2162 1395 -2129
rect 1425 -2162 1429 -2101
rect 1443 -2118 1447 -2101
rect 1373 -2169 1377 -2166
rect 1381 -2166 1395 -2162
rect 1381 -2169 1385 -2166
rect 1409 -2169 1413 -2166
rect 1417 -2166 1436 -2162
rect 1417 -2169 1421 -2166
rect 1443 -2169 1447 -2122
rect 1469 -2133 1473 -2101
rect 1469 -2162 1473 -2137
rect 1503 -2155 1507 -2101
rect 1503 -2159 1520 -2155
rect 1451 -2169 1455 -2166
rect 1460 -2166 1473 -2162
rect 1460 -2169 1464 -2166
rect 1487 -2169 1491 -2166
rect 1511 -2169 1515 -2159
rect 1527 -2162 1531 -2101
rect 1535 -2155 1539 -2101
rect 1535 -2159 1554 -2155
rect 1519 -2166 1536 -2162
rect 1519 -2169 1523 -2166
rect 1543 -2169 1547 -2159
rect 1561 -2169 1565 -2101
rect 1330 -2177 1334 -2173
rect 1356 -2177 1360 -2173
rect 1399 -2177 1403 -2173
rect 1434 -2177 1438 -2173
rect 1478 -2177 1482 -2173
rect 1495 -2177 1499 -2173
rect 1531 -2177 1535 -2173
rect 1552 -2177 1556 -2173
rect 1561 -2191 1565 -2173
rect 1567 -2184 1571 -2137
rect 1330 -2368 1334 -2364
rect 1347 -2368 1351 -2364
rect 1367 -2368 1371 -2364
rect 1388 -2368 1392 -2364
rect 1409 -2368 1413 -2364
rect 1430 -2368 1434 -2364
rect 1451 -2368 1455 -2364
rect 1472 -2368 1476 -2364
rect 1493 -2368 1497 -2364
rect 1513 -2368 1517 -2364
rect 1321 -2423 1325 -2376
rect 1321 -2444 1325 -2427
rect 1339 -2437 1343 -2376
rect 1355 -2437 1359 -2376
rect 1379 -2416 1383 -2376
rect 1379 -2437 1383 -2420
rect 1397 -2437 1401 -2376
rect 1421 -2423 1425 -2376
rect 1421 -2437 1425 -2427
rect 1439 -2416 1443 -2376
rect 1439 -2437 1443 -2420
rect 1463 -2430 1467 -2376
rect 1481 -2408 1485 -2376
rect 1481 -2416 1485 -2412
rect 1463 -2437 1467 -2434
rect 1339 -2441 1348 -2437
rect 1355 -2441 1363 -2437
rect 1339 -2444 1343 -2441
rect 1363 -2444 1367 -2441
rect 1371 -2441 1383 -2437
rect 1397 -2441 1405 -2437
rect 1371 -2444 1375 -2441
rect 1405 -2444 1409 -2441
rect 1413 -2441 1425 -2437
rect 1439 -2441 1451 -2437
rect 1413 -2444 1417 -2441
rect 1447 -2444 1451 -2441
rect 1455 -2441 1467 -2437
rect 1481 -2437 1485 -2420
rect 1505 -2423 1509 -2376
rect 1505 -2437 1509 -2427
rect 1481 -2441 1493 -2437
rect 1455 -2444 1459 -2441
rect 1489 -2444 1493 -2441
rect 1497 -2441 1509 -2437
rect 1497 -2444 1501 -2441
rect 1330 -2452 1334 -2448
rect 1347 -2452 1351 -2448
rect 1388 -2452 1392 -2448
rect 1430 -2452 1434 -2448
rect 1472 -2452 1476 -2448
rect 1513 -2452 1517 -2448
rect 1519 -2460 1523 -2412
rect 1330 -2499 1334 -2495
rect 1347 -2499 1351 -2495
rect 1367 -2499 1371 -2495
rect 1388 -2499 1392 -2495
rect 1409 -2499 1413 -2495
rect 1430 -2499 1434 -2495
rect 1451 -2499 1455 -2495
rect 1472 -2499 1476 -2495
rect 1493 -2499 1497 -2495
rect 1513 -2499 1517 -2495
rect 1321 -2554 1325 -2507
rect 1321 -2575 1325 -2558
rect 1339 -2568 1343 -2507
rect 1355 -2568 1359 -2507
rect 1379 -2547 1383 -2507
rect 1379 -2568 1383 -2551
rect 1397 -2568 1401 -2507
rect 1421 -2554 1425 -2507
rect 1421 -2568 1425 -2558
rect 1439 -2547 1443 -2507
rect 1439 -2568 1443 -2551
rect 1463 -2561 1467 -2507
rect 1481 -2539 1485 -2507
rect 1481 -2547 1485 -2543
rect 1463 -2568 1467 -2565
rect 1339 -2572 1348 -2568
rect 1355 -2572 1363 -2568
rect 1339 -2575 1343 -2572
rect 1363 -2575 1367 -2572
rect 1371 -2572 1383 -2568
rect 1397 -2572 1405 -2568
rect 1371 -2575 1375 -2572
rect 1405 -2575 1409 -2572
rect 1413 -2572 1425 -2568
rect 1439 -2572 1451 -2568
rect 1413 -2575 1417 -2572
rect 1447 -2575 1451 -2572
rect 1455 -2572 1467 -2568
rect 1481 -2568 1485 -2551
rect 1505 -2554 1509 -2507
rect 1505 -2568 1509 -2558
rect 1481 -2572 1493 -2568
rect 1455 -2575 1459 -2572
rect 1489 -2575 1493 -2572
rect 1497 -2572 1509 -2568
rect 1497 -2575 1501 -2572
rect 1330 -2583 1334 -2579
rect 1347 -2583 1351 -2579
rect 1388 -2583 1392 -2579
rect 1430 -2583 1434 -2579
rect 1472 -2583 1476 -2579
rect 1513 -2583 1517 -2579
rect 1321 -2724 1325 -2720
rect 1338 -2724 1342 -2720
rect 1329 -2735 1333 -2732
rect 1329 -2739 1344 -2735
rect 1315 -2752 1322 -2748
rect 1199 -2962 1203 -2958
rect 1207 -3004 1211 -2970
rect 1207 -3038 1211 -3008
rect 1199 -3046 1203 -3042
rect 972 -3078 976 -3074
rect 989 -3078 993 -3074
rect 1009 -3078 1013 -3074
rect 1030 -3078 1034 -3074
rect 1051 -3078 1055 -3074
rect 1072 -3078 1076 -3074
rect 1093 -3078 1097 -3074
rect 1114 -3078 1118 -3074
rect 1135 -3078 1139 -3074
rect 1155 -3078 1159 -3074
rect 1199 -3078 1203 -3074
rect 963 -3133 967 -3086
rect 963 -3154 967 -3137
rect 981 -3147 985 -3086
rect 997 -3147 1001 -3086
rect 1021 -3126 1025 -3086
rect 1021 -3147 1025 -3130
rect 1039 -3147 1043 -3086
rect 1063 -3133 1067 -3086
rect 1063 -3147 1067 -3137
rect 1081 -3126 1085 -3086
rect 1081 -3147 1085 -3130
rect 1105 -3140 1109 -3086
rect 1123 -3118 1127 -3086
rect 1123 -3126 1127 -3122
rect 1105 -3147 1109 -3144
rect 981 -3151 990 -3147
rect 997 -3151 1005 -3147
rect 981 -3154 985 -3151
rect 1005 -3154 1009 -3151
rect 1013 -3151 1025 -3147
rect 1039 -3151 1047 -3147
rect 1013 -3154 1017 -3151
rect 1047 -3154 1051 -3151
rect 1055 -3151 1067 -3147
rect 1081 -3151 1093 -3147
rect 1055 -3154 1059 -3151
rect 1089 -3154 1093 -3151
rect 1097 -3151 1109 -3147
rect 1123 -3147 1127 -3130
rect 1147 -3133 1151 -3086
rect 1147 -3147 1151 -3137
rect 1123 -3151 1135 -3147
rect 1097 -3154 1101 -3151
rect 1131 -3154 1135 -3151
rect 1139 -3151 1151 -3147
rect 1139 -3154 1143 -3151
rect 972 -3162 976 -3158
rect 989 -3162 993 -3158
rect 1030 -3162 1034 -3158
rect 1072 -3162 1076 -3158
rect 1114 -3162 1118 -3158
rect 1155 -3162 1159 -3158
rect 1161 -3169 1165 -3122
rect 1207 -3119 1211 -3086
rect 1207 -3154 1211 -3123
rect 1309 -3126 1313 -2945
rect 1199 -3162 1203 -3158
rect 972 -3199 976 -3195
rect 989 -3199 993 -3195
rect 1009 -3199 1013 -3195
rect 1030 -3199 1034 -3195
rect 1051 -3199 1055 -3195
rect 1072 -3199 1076 -3195
rect 1093 -3199 1097 -3195
rect 1114 -3199 1118 -3195
rect 1135 -3199 1139 -3195
rect 1155 -3199 1159 -3195
rect 963 -3254 967 -3207
rect 963 -3275 967 -3258
rect 981 -3268 985 -3207
rect 997 -3268 1001 -3207
rect 1021 -3247 1025 -3207
rect 1021 -3268 1025 -3251
rect 1039 -3268 1043 -3207
rect 1063 -3254 1067 -3207
rect 1063 -3268 1067 -3258
rect 1081 -3247 1085 -3207
rect 1081 -3268 1085 -3251
rect 1105 -3261 1109 -3207
rect 1123 -3239 1127 -3207
rect 1123 -3247 1127 -3243
rect 1105 -3268 1109 -3265
rect 981 -3272 990 -3268
rect 997 -3272 1005 -3268
rect 981 -3275 985 -3272
rect 1005 -3275 1009 -3272
rect 1013 -3272 1025 -3268
rect 1039 -3272 1047 -3268
rect 1013 -3275 1017 -3272
rect 1047 -3275 1051 -3272
rect 1055 -3272 1067 -3268
rect 1081 -3272 1093 -3268
rect 1055 -3275 1059 -3272
rect 1089 -3275 1093 -3272
rect 1097 -3272 1109 -3268
rect 1123 -3268 1127 -3251
rect 1147 -3254 1151 -3207
rect 1147 -3268 1151 -3258
rect 1123 -3272 1135 -3268
rect 1097 -3275 1101 -3272
rect 1131 -3275 1135 -3272
rect 1139 -3272 1151 -3268
rect 1139 -3275 1143 -3272
rect 972 -3283 976 -3279
rect 989 -3283 993 -3279
rect 1030 -3283 1034 -3279
rect 1072 -3283 1076 -3279
rect 1114 -3283 1118 -3279
rect 1155 -3283 1159 -3279
rect 963 -3430 967 -3426
rect 980 -3430 984 -3426
rect 971 -3441 975 -3438
rect 971 -3445 986 -3441
rect 957 -3458 964 -3454
rect 574 -3915 578 -3911
rect 591 -3915 595 -3911
rect 611 -3915 615 -3911
rect 632 -3915 636 -3911
rect 653 -3915 657 -3911
rect 674 -3915 678 -3911
rect 695 -3915 699 -3911
rect 716 -3915 720 -3911
rect 737 -3915 741 -3911
rect 757 -3915 761 -3911
rect 565 -3970 569 -3923
rect 565 -3991 569 -3974
rect 583 -3984 587 -3923
rect 599 -3984 603 -3923
rect 623 -3963 627 -3923
rect 623 -3984 627 -3967
rect 641 -3984 645 -3923
rect 665 -3970 669 -3923
rect 665 -3984 669 -3974
rect 683 -3963 687 -3923
rect 683 -3984 687 -3967
rect 707 -3977 711 -3923
rect 725 -3955 729 -3923
rect 725 -3963 729 -3959
rect 707 -3984 711 -3981
rect 583 -3988 592 -3984
rect 599 -3988 607 -3984
rect 583 -3991 587 -3988
rect 607 -3991 611 -3988
rect 615 -3988 627 -3984
rect 641 -3988 649 -3984
rect 615 -3991 619 -3988
rect 649 -3991 653 -3988
rect 657 -3988 669 -3984
rect 683 -3988 695 -3984
rect 657 -3991 661 -3988
rect 691 -3991 695 -3988
rect 699 -3988 711 -3984
rect 725 -3984 729 -3967
rect 749 -3970 753 -3923
rect 749 -3984 753 -3974
rect 725 -3988 737 -3984
rect 699 -3991 703 -3988
rect 733 -3991 737 -3988
rect 741 -3988 753 -3984
rect 741 -3991 745 -3988
rect 574 -3999 578 -3995
rect 591 -3999 595 -3995
rect 632 -3999 636 -3995
rect 674 -3999 678 -3995
rect 716 -3999 720 -3995
rect 757 -3999 761 -3995
rect 763 -4007 767 -3959
rect 951 -3963 955 -3649
rect 574 -4040 578 -4036
rect 591 -4040 595 -4036
rect 611 -4040 615 -4036
rect 632 -4040 636 -4036
rect 653 -4040 657 -4036
rect 674 -4040 678 -4036
rect 695 -4040 699 -4036
rect 716 -4040 720 -4036
rect 737 -4040 741 -4036
rect 757 -4040 761 -4036
rect 565 -4095 569 -4048
rect 565 -4116 569 -4099
rect 583 -4109 587 -4048
rect 599 -4109 603 -4048
rect 623 -4088 627 -4048
rect 623 -4109 627 -4092
rect 641 -4109 645 -4048
rect 665 -4095 669 -4048
rect 665 -4109 669 -4099
rect 683 -4088 687 -4048
rect 683 -4109 687 -4092
rect 707 -4102 711 -4048
rect 725 -4080 729 -4048
rect 725 -4088 729 -4084
rect 707 -4109 711 -4106
rect 583 -4113 592 -4109
rect 599 -4113 607 -4109
rect 583 -4116 587 -4113
rect 607 -4116 611 -4113
rect 615 -4113 627 -4109
rect 641 -4113 649 -4109
rect 615 -4116 619 -4113
rect 649 -4116 653 -4113
rect 657 -4113 669 -4109
rect 683 -4113 695 -4109
rect 657 -4116 661 -4113
rect 691 -4116 695 -4113
rect 699 -4113 711 -4109
rect 725 -4109 729 -4092
rect 749 -4095 753 -4048
rect 749 -4109 753 -4099
rect 725 -4113 737 -4109
rect 699 -4116 703 -4113
rect 733 -4116 737 -4113
rect 741 -4113 753 -4109
rect 741 -4116 745 -4113
rect 574 -4124 578 -4120
rect 591 -4124 595 -4120
rect 632 -4124 636 -4120
rect 674 -4124 678 -4120
rect 716 -4124 720 -4120
rect 757 -4124 761 -4120
rect 565 -4275 569 -4271
rect 582 -4275 586 -4271
rect 573 -4286 577 -4283
rect 573 -4290 588 -4286
rect 559 -4303 566 -4299
rect 218 -4638 222 -4634
rect 235 -4638 239 -4634
rect 255 -4638 259 -4634
rect 276 -4638 280 -4634
rect 297 -4638 301 -4634
rect 318 -4638 322 -4634
rect 339 -4638 343 -4634
rect 360 -4638 364 -4634
rect 381 -4638 385 -4634
rect 401 -4638 405 -4634
rect 209 -4693 213 -4646
rect 209 -4714 213 -4697
rect 227 -4707 231 -4646
rect 243 -4707 247 -4646
rect 267 -4686 271 -4646
rect 267 -4707 271 -4690
rect 285 -4707 289 -4646
rect 309 -4693 313 -4646
rect 309 -4707 313 -4697
rect 327 -4686 331 -4646
rect 327 -4707 331 -4690
rect 351 -4700 355 -4646
rect 369 -4678 373 -4646
rect 369 -4686 373 -4682
rect 351 -4707 355 -4704
rect 227 -4711 236 -4707
rect 243 -4711 251 -4707
rect 227 -4714 231 -4711
rect 251 -4714 255 -4711
rect 259 -4711 271 -4707
rect 285 -4711 293 -4707
rect 259 -4714 263 -4711
rect 293 -4714 297 -4711
rect 301 -4711 313 -4707
rect 327 -4711 339 -4707
rect 301 -4714 305 -4711
rect 335 -4714 339 -4711
rect 343 -4711 355 -4707
rect 369 -4707 373 -4690
rect 393 -4693 397 -4646
rect 393 -4707 397 -4697
rect 369 -4711 381 -4707
rect 343 -4714 347 -4711
rect 377 -4714 381 -4711
rect 385 -4711 397 -4707
rect 385 -4714 389 -4711
rect 218 -4722 222 -4718
rect 235 -4722 239 -4718
rect 276 -4722 280 -4718
rect 318 -4722 322 -4718
rect 360 -4722 364 -4718
rect 401 -4722 405 -4718
rect 407 -4731 411 -4682
rect 553 -4686 557 -4496
rect 218 -4759 222 -4755
rect 235 -4759 239 -4755
rect 255 -4759 259 -4755
rect 276 -4759 280 -4755
rect 297 -4759 301 -4755
rect 318 -4759 322 -4755
rect 339 -4759 343 -4755
rect 360 -4759 364 -4755
rect 381 -4759 385 -4755
rect 401 -4759 405 -4755
rect 209 -4814 213 -4767
rect 209 -4835 213 -4818
rect 227 -4828 231 -4767
rect 243 -4828 247 -4767
rect 267 -4807 271 -4767
rect 267 -4828 271 -4811
rect 285 -4828 289 -4767
rect 309 -4814 313 -4767
rect 309 -4828 313 -4818
rect 327 -4807 331 -4767
rect 327 -4828 331 -4811
rect 351 -4821 355 -4767
rect 369 -4799 373 -4767
rect 369 -4807 373 -4803
rect 351 -4828 355 -4825
rect 227 -4832 236 -4828
rect 243 -4832 251 -4828
rect 227 -4835 231 -4832
rect 251 -4835 255 -4832
rect 259 -4832 271 -4828
rect 285 -4832 293 -4828
rect 259 -4835 263 -4832
rect 293 -4835 297 -4832
rect 301 -4832 313 -4828
rect 327 -4832 339 -4828
rect 301 -4835 305 -4832
rect 335 -4835 339 -4832
rect 343 -4832 355 -4828
rect 369 -4828 373 -4811
rect 393 -4814 397 -4767
rect 393 -4828 397 -4818
rect 369 -4832 381 -4828
rect 343 -4835 347 -4832
rect 377 -4835 381 -4832
rect 385 -4832 397 -4828
rect 385 -4835 389 -4832
rect 218 -4843 222 -4839
rect 235 -4843 239 -4839
rect 276 -4843 280 -4839
rect 318 -4843 322 -4839
rect 360 -4843 364 -4839
rect 401 -4843 405 -4839
rect 218 -4877 222 -4873
rect 235 -4877 239 -4873
rect 255 -4877 259 -4873
rect 276 -4877 280 -4873
rect 297 -4877 301 -4873
rect 318 -4877 322 -4873
rect 339 -4877 343 -4873
rect 360 -4877 364 -4873
rect 381 -4877 385 -4873
rect 401 -4877 405 -4873
rect 209 -4932 213 -4885
rect 209 -4953 213 -4936
rect 227 -4946 231 -4885
rect 243 -4946 247 -4885
rect 267 -4925 271 -4885
rect 267 -4946 271 -4929
rect 285 -4946 289 -4885
rect 309 -4932 313 -4885
rect 309 -4946 313 -4936
rect 327 -4925 331 -4885
rect 327 -4946 331 -4929
rect 351 -4939 355 -4885
rect 369 -4917 373 -4885
rect 369 -4925 373 -4921
rect 351 -4946 355 -4943
rect 227 -4950 236 -4946
rect 243 -4950 251 -4946
rect 227 -4953 231 -4950
rect 251 -4953 255 -4950
rect 259 -4950 271 -4946
rect 285 -4950 293 -4946
rect 259 -4953 263 -4950
rect 293 -4953 297 -4950
rect 301 -4950 313 -4946
rect 327 -4950 339 -4946
rect 301 -4953 305 -4950
rect 335 -4953 339 -4950
rect 343 -4950 355 -4946
rect 369 -4946 373 -4929
rect 393 -4932 397 -4885
rect 393 -4946 397 -4936
rect 369 -4950 381 -4946
rect 343 -4953 347 -4950
rect 377 -4953 381 -4950
rect 385 -4950 397 -4946
rect 385 -4953 389 -4950
rect 218 -4961 222 -4957
rect 235 -4961 239 -4957
rect 276 -4961 280 -4957
rect 318 -4961 322 -4957
rect 360 -4961 364 -4957
rect 401 -4961 405 -4957
rect 209 -4994 213 -4990
rect 226 -4994 230 -4990
rect 217 -5005 221 -5002
rect 217 -5009 232 -5005
rect 203 -5022 210 -5018
rect -210 -5353 -206 -5349
rect -193 -5353 -189 -5349
rect -173 -5353 -169 -5349
rect -152 -5353 -148 -5349
rect -131 -5353 -127 -5349
rect -110 -5353 -106 -5349
rect -89 -5353 -85 -5349
rect -68 -5353 -64 -5349
rect -47 -5353 -43 -5349
rect -27 -5353 -23 -5349
rect -219 -5408 -215 -5361
rect -219 -5429 -215 -5412
rect -201 -5422 -197 -5361
rect -185 -5422 -181 -5361
rect -161 -5401 -157 -5361
rect -161 -5422 -157 -5405
rect -143 -5422 -139 -5361
rect -119 -5408 -115 -5361
rect -119 -5422 -115 -5412
rect -101 -5401 -97 -5361
rect -101 -5422 -97 -5405
rect -77 -5415 -73 -5361
rect -59 -5393 -55 -5361
rect -59 -5401 -55 -5397
rect -77 -5422 -73 -5419
rect -201 -5426 -192 -5422
rect -185 -5426 -177 -5422
rect -201 -5429 -197 -5426
rect -177 -5429 -173 -5426
rect -169 -5426 -157 -5422
rect -143 -5426 -135 -5422
rect -169 -5429 -165 -5426
rect -135 -5429 -131 -5426
rect -127 -5426 -115 -5422
rect -101 -5426 -89 -5422
rect -127 -5429 -123 -5426
rect -93 -5429 -89 -5426
rect -85 -5426 -73 -5422
rect -59 -5422 -55 -5405
rect -35 -5408 -31 -5361
rect -35 -5422 -31 -5412
rect -59 -5426 -47 -5422
rect -85 -5429 -81 -5426
rect -51 -5429 -47 -5426
rect -43 -5426 -31 -5422
rect -43 -5429 -39 -5426
rect -210 -5437 -206 -5433
rect -193 -5437 -189 -5433
rect -152 -5437 -148 -5433
rect -110 -5437 -106 -5433
rect -68 -5437 -64 -5433
rect -27 -5437 -23 -5433
rect -21 -5444 -17 -5397
rect 197 -5401 201 -5208
rect -210 -5473 -206 -5469
rect -193 -5473 -189 -5469
rect -173 -5473 -169 -5469
rect -152 -5473 -148 -5469
rect -131 -5473 -127 -5469
rect -110 -5473 -106 -5469
rect -89 -5473 -85 -5469
rect -68 -5473 -64 -5469
rect -47 -5473 -43 -5469
rect -27 -5473 -23 -5469
rect -219 -5528 -215 -5481
rect -219 -5549 -215 -5532
rect -201 -5542 -197 -5481
rect -185 -5542 -181 -5481
rect -161 -5521 -157 -5481
rect -161 -5542 -157 -5525
rect -143 -5542 -139 -5481
rect -119 -5528 -115 -5481
rect -119 -5542 -115 -5532
rect -101 -5521 -97 -5481
rect -101 -5542 -97 -5525
rect -77 -5535 -73 -5481
rect -59 -5513 -55 -5481
rect -59 -5521 -55 -5517
rect -77 -5542 -73 -5539
rect -201 -5546 -192 -5542
rect -185 -5546 -177 -5542
rect -201 -5549 -197 -5546
rect -177 -5549 -173 -5546
rect -169 -5546 -157 -5542
rect -143 -5546 -135 -5542
rect -169 -5549 -165 -5546
rect -135 -5549 -131 -5546
rect -127 -5546 -115 -5542
rect -101 -5546 -89 -5542
rect -127 -5549 -123 -5546
rect -93 -5549 -89 -5546
rect -85 -5546 -73 -5542
rect -59 -5542 -55 -5525
rect -35 -5528 -31 -5481
rect -35 -5542 -31 -5532
rect -59 -5546 -47 -5542
rect -85 -5549 -81 -5546
rect -51 -5549 -47 -5546
rect -43 -5546 -31 -5542
rect -43 -5549 -39 -5546
rect -210 -5557 -206 -5553
rect -193 -5557 -189 -5553
rect -152 -5557 -148 -5553
rect -110 -5557 -106 -5553
rect -68 -5557 -64 -5553
rect -27 -5557 -23 -5553
rect -210 -5590 -206 -5586
rect -193 -5590 -189 -5586
rect -173 -5590 -169 -5586
rect -152 -5590 -148 -5586
rect -131 -5590 -127 -5586
rect -110 -5590 -106 -5586
rect -89 -5590 -85 -5586
rect -68 -5590 -64 -5586
rect -47 -5590 -43 -5586
rect -27 -5590 -23 -5586
rect -219 -5645 -215 -5598
rect -219 -5666 -215 -5649
rect -201 -5659 -197 -5598
rect -185 -5659 -181 -5598
rect -161 -5638 -157 -5598
rect -161 -5659 -157 -5642
rect -143 -5659 -139 -5598
rect -119 -5645 -115 -5598
rect -119 -5659 -115 -5649
rect -101 -5638 -97 -5598
rect -101 -5659 -97 -5642
rect -77 -5652 -73 -5598
rect -59 -5630 -55 -5598
rect -59 -5638 -55 -5634
rect -77 -5659 -73 -5656
rect -201 -5663 -192 -5659
rect -185 -5663 -177 -5659
rect -201 -5666 -197 -5663
rect -177 -5666 -173 -5663
rect -169 -5663 -157 -5659
rect -143 -5663 -135 -5659
rect -169 -5666 -165 -5663
rect -135 -5666 -131 -5663
rect -127 -5663 -115 -5659
rect -101 -5663 -89 -5659
rect -127 -5666 -123 -5663
rect -93 -5666 -89 -5663
rect -85 -5663 -73 -5659
rect -59 -5659 -55 -5642
rect -35 -5645 -31 -5598
rect -35 -5659 -31 -5649
rect -59 -5663 -47 -5659
rect -85 -5666 -81 -5663
rect -51 -5666 -47 -5663
rect -43 -5663 -31 -5659
rect -43 -5666 -39 -5663
rect -210 -5674 -206 -5670
rect -193 -5674 -189 -5670
rect -152 -5674 -148 -5670
rect -110 -5674 -106 -5670
rect -68 -5674 -64 -5670
rect -27 -5674 -23 -5670
rect -219 -5707 -215 -5703
rect -202 -5707 -198 -5703
rect -211 -5718 -207 -5715
rect -211 -5722 -196 -5718
rect -200 -5761 -196 -5722
rect -200 -5776 -196 -5765
rect -219 -5780 -196 -5776
rect -193 -5752 -189 -5715
rect -21 -5731 -17 -5517
rect -219 -5783 -215 -5780
rect -193 -5783 -189 -5756
rect -202 -5791 -198 -5787
rect -210 -5826 -206 -5822
rect -184 -5826 -180 -5822
rect -167 -5826 -163 -5822
rect -127 -5826 -123 -5822
rect -106 -5826 -102 -5822
rect -89 -5826 -85 -5822
rect -49 -5826 -45 -5822
rect -25 -5826 -21 -5822
rect 12 -5826 16 -5822
rect -219 -5851 -215 -5834
rect -219 -5902 -215 -5855
rect -201 -5844 -197 -5834
rect -201 -5902 -197 -5848
rect -193 -5873 -189 -5834
rect -175 -5866 -171 -5834
rect -193 -5902 -189 -5877
rect -175 -5902 -171 -5870
rect -149 -5858 -145 -5834
rect -149 -5895 -145 -5862
rect -115 -5895 -111 -5834
rect -97 -5851 -93 -5834
rect -167 -5902 -163 -5899
rect -159 -5899 -145 -5895
rect -159 -5902 -155 -5899
rect -131 -5902 -127 -5899
rect -123 -5899 -104 -5895
rect -123 -5902 -119 -5899
rect -97 -5902 -93 -5855
rect -71 -5866 -67 -5834
rect -71 -5895 -67 -5870
rect -37 -5888 -33 -5834
rect -37 -5892 -20 -5888
rect -89 -5902 -85 -5899
rect -80 -5899 -67 -5895
rect -80 -5902 -76 -5899
rect -53 -5902 -49 -5899
rect -29 -5902 -25 -5892
rect -13 -5895 -9 -5834
rect -5 -5888 -1 -5834
rect 21 -5858 25 -5834
rect -5 -5892 14 -5888
rect -21 -5899 -4 -5895
rect -21 -5902 -17 -5899
rect 3 -5902 7 -5892
rect 21 -5902 25 -5862
rect -210 -5910 -206 -5906
rect -184 -5910 -180 -5906
rect -141 -5910 -137 -5906
rect -106 -5910 -102 -5906
rect -62 -5910 -58 -5906
rect -45 -5910 -41 -5906
rect -9 -5910 -5 -5906
rect 12 -5910 16 -5906
rect 27 -5917 31 -5870
rect 191 -5873 195 -5756
rect 197 -5858 201 -5448
rect 203 -5521 207 -5022
rect 228 -5048 232 -5009
rect 228 -5063 232 -5052
rect 209 -5067 232 -5063
rect 235 -5039 239 -5002
rect 407 -5026 411 -4921
rect 413 -5018 417 -4803
rect 209 -5070 213 -5067
rect 235 -5070 239 -5043
rect 226 -5078 230 -5074
rect 218 -5113 222 -5109
rect 244 -5113 248 -5109
rect 261 -5113 265 -5109
rect 301 -5113 305 -5109
rect 322 -5113 326 -5109
rect 339 -5113 343 -5109
rect 379 -5113 383 -5109
rect 403 -5113 407 -5109
rect 440 -5113 444 -5109
rect 209 -5138 213 -5121
rect 209 -5189 213 -5142
rect 227 -5131 231 -5121
rect 227 -5189 231 -5135
rect 235 -5160 239 -5121
rect 253 -5153 257 -5121
rect 235 -5189 239 -5164
rect 253 -5189 257 -5157
rect 279 -5145 283 -5121
rect 279 -5182 283 -5149
rect 313 -5182 317 -5121
rect 331 -5138 335 -5121
rect 261 -5189 265 -5186
rect 269 -5186 283 -5182
rect 269 -5189 273 -5186
rect 297 -5189 301 -5186
rect 305 -5186 324 -5182
rect 305 -5189 309 -5186
rect 331 -5189 335 -5142
rect 357 -5153 361 -5121
rect 357 -5182 361 -5157
rect 391 -5175 395 -5121
rect 391 -5179 408 -5175
rect 339 -5189 343 -5186
rect 348 -5186 361 -5182
rect 348 -5189 352 -5186
rect 375 -5189 379 -5186
rect 399 -5189 403 -5179
rect 415 -5182 419 -5121
rect 423 -5175 427 -5121
rect 449 -5145 453 -5121
rect 423 -5179 442 -5175
rect 407 -5186 424 -5182
rect 407 -5189 411 -5186
rect 431 -5189 435 -5179
rect 449 -5189 453 -5149
rect 218 -5197 222 -5193
rect 244 -5197 248 -5193
rect 287 -5197 291 -5193
rect 322 -5197 326 -5193
rect 366 -5197 370 -5193
rect 383 -5197 387 -5193
rect 419 -5197 423 -5193
rect 440 -5197 444 -5193
rect 455 -5211 459 -5157
rect 547 -5160 551 -5043
rect 553 -5145 557 -4734
rect 559 -4807 563 -4303
rect 584 -4329 588 -4290
rect 584 -4344 588 -4333
rect 565 -4348 588 -4344
rect 591 -4320 595 -4283
rect 763 -4299 767 -4084
rect 860 -4275 864 -4271
rect 868 -4317 872 -4291
rect 565 -4351 569 -4348
rect 591 -4351 595 -4324
rect 868 -4347 872 -4321
rect 582 -4359 586 -4355
rect 860 -4359 864 -4355
rect 574 -4394 578 -4390
rect 600 -4394 604 -4390
rect 617 -4394 621 -4390
rect 657 -4394 661 -4390
rect 678 -4394 682 -4390
rect 695 -4394 699 -4390
rect 735 -4394 739 -4390
rect 759 -4394 763 -4390
rect 796 -4394 800 -4390
rect 565 -4419 569 -4402
rect 565 -4470 569 -4423
rect 583 -4412 587 -4402
rect 583 -4470 587 -4416
rect 591 -4441 595 -4402
rect 609 -4434 613 -4402
rect 591 -4470 595 -4445
rect 609 -4470 613 -4438
rect 635 -4426 639 -4402
rect 635 -4463 639 -4430
rect 669 -4463 673 -4402
rect 687 -4419 691 -4402
rect 617 -4470 621 -4467
rect 625 -4467 639 -4463
rect 625 -4470 629 -4467
rect 653 -4470 657 -4467
rect 661 -4467 680 -4463
rect 661 -4470 665 -4467
rect 687 -4470 691 -4423
rect 713 -4434 717 -4402
rect 713 -4463 717 -4438
rect 747 -4456 751 -4402
rect 747 -4460 764 -4456
rect 695 -4470 699 -4467
rect 704 -4467 717 -4463
rect 704 -4470 708 -4467
rect 731 -4470 735 -4467
rect 755 -4470 759 -4460
rect 771 -4463 775 -4402
rect 779 -4456 783 -4402
rect 805 -4426 809 -4402
rect 779 -4460 798 -4456
rect 763 -4467 780 -4463
rect 763 -4470 767 -4467
rect 787 -4470 791 -4460
rect 805 -4470 809 -4430
rect 574 -4478 578 -4474
rect 600 -4478 604 -4474
rect 643 -4478 647 -4474
rect 678 -4478 682 -4474
rect 722 -4478 726 -4474
rect 739 -4478 743 -4474
rect 775 -4478 779 -4474
rect 796 -4478 800 -4474
rect 811 -4485 815 -4438
rect 945 -4441 949 -4324
rect 951 -4426 955 -4010
rect 957 -4088 961 -3458
rect 982 -3484 986 -3445
rect 982 -3499 986 -3488
rect 963 -3503 986 -3499
rect 989 -3475 993 -3438
rect 1161 -3454 1165 -3243
rect 963 -3506 967 -3503
rect 989 -3506 993 -3479
rect 980 -3514 984 -3510
rect 972 -3554 976 -3550
rect 998 -3554 1002 -3550
rect 1015 -3554 1019 -3550
rect 1055 -3554 1059 -3550
rect 1076 -3554 1080 -3550
rect 1093 -3554 1097 -3550
rect 1133 -3554 1137 -3550
rect 1157 -3554 1161 -3550
rect 1194 -3554 1198 -3550
rect 963 -3579 967 -3562
rect 963 -3630 967 -3583
rect 981 -3572 985 -3562
rect 981 -3630 985 -3576
rect 989 -3601 993 -3562
rect 1007 -3594 1011 -3562
rect 989 -3630 993 -3605
rect 1007 -3630 1011 -3598
rect 1033 -3586 1037 -3562
rect 1033 -3623 1037 -3590
rect 1067 -3623 1071 -3562
rect 1085 -3579 1089 -3562
rect 1015 -3630 1019 -3627
rect 1023 -3627 1037 -3623
rect 1023 -3630 1027 -3627
rect 1051 -3630 1055 -3627
rect 1059 -3627 1078 -3623
rect 1059 -3630 1063 -3627
rect 1085 -3630 1089 -3583
rect 1111 -3594 1115 -3562
rect 1111 -3623 1115 -3598
rect 1145 -3616 1149 -3562
rect 1145 -3620 1162 -3616
rect 1093 -3630 1097 -3627
rect 1102 -3627 1115 -3623
rect 1102 -3630 1106 -3627
rect 1129 -3630 1133 -3627
rect 1153 -3630 1157 -3620
rect 1169 -3623 1173 -3562
rect 1177 -3616 1181 -3562
rect 1203 -3584 1207 -3562
rect 1177 -3620 1196 -3616
rect 1161 -3627 1178 -3623
rect 1161 -3630 1165 -3627
rect 1185 -3630 1189 -3620
rect 1203 -3630 1207 -3588
rect 1303 -3586 1307 -3479
rect 972 -3638 976 -3634
rect 998 -3638 1002 -3634
rect 1041 -3638 1045 -3634
rect 1076 -3638 1080 -3634
rect 1120 -3638 1124 -3634
rect 1137 -3638 1141 -3634
rect 1173 -3638 1177 -3634
rect 1194 -3638 1198 -3634
rect 1209 -3652 1213 -3598
rect 1309 -3601 1313 -3174
rect 1315 -3247 1319 -2752
rect 1340 -2778 1344 -2739
rect 1340 -2793 1344 -2782
rect 1321 -2797 1344 -2793
rect 1347 -2769 1351 -2732
rect 1519 -2748 1523 -2543
rect 1321 -2800 1325 -2797
rect 1347 -2800 1351 -2773
rect 1338 -2808 1342 -2804
rect 1330 -2843 1334 -2839
rect 1356 -2843 1360 -2839
rect 1373 -2843 1377 -2839
rect 1413 -2843 1417 -2839
rect 1434 -2843 1438 -2839
rect 1451 -2843 1455 -2839
rect 1491 -2843 1495 -2839
rect 1515 -2843 1519 -2839
rect 1552 -2843 1556 -2839
rect 1321 -2868 1325 -2851
rect 1321 -2919 1325 -2872
rect 1339 -2861 1343 -2851
rect 1339 -2919 1343 -2865
rect 1347 -2890 1351 -2851
rect 1365 -2883 1369 -2851
rect 1347 -2919 1351 -2894
rect 1365 -2919 1369 -2887
rect 1391 -2875 1395 -2851
rect 1391 -2912 1395 -2879
rect 1425 -2912 1429 -2851
rect 1443 -2868 1447 -2851
rect 1373 -2919 1377 -2916
rect 1381 -2916 1395 -2912
rect 1381 -2919 1385 -2916
rect 1409 -2919 1413 -2916
rect 1417 -2916 1436 -2912
rect 1417 -2919 1421 -2916
rect 1443 -2919 1447 -2872
rect 1469 -2883 1473 -2851
rect 1469 -2912 1473 -2887
rect 1503 -2905 1507 -2851
rect 1503 -2909 1520 -2905
rect 1451 -2919 1455 -2916
rect 1460 -2916 1473 -2912
rect 1460 -2919 1464 -2916
rect 1487 -2919 1491 -2916
rect 1511 -2919 1515 -2909
rect 1527 -2912 1531 -2851
rect 1535 -2905 1539 -2851
rect 1535 -2909 1554 -2905
rect 1519 -2916 1536 -2912
rect 1519 -2919 1523 -2916
rect 1543 -2919 1547 -2909
rect 1561 -2919 1565 -2851
rect 1330 -2927 1334 -2923
rect 1356 -2927 1360 -2923
rect 1399 -2927 1403 -2923
rect 1434 -2927 1438 -2923
rect 1478 -2927 1482 -2923
rect 1495 -2927 1499 -2923
rect 1531 -2927 1535 -2923
rect 1552 -2927 1556 -2923
rect 1561 -2941 1565 -2923
rect 1567 -2934 1571 -2887
rect 1330 -3078 1334 -3074
rect 1347 -3078 1351 -3074
rect 1367 -3078 1371 -3074
rect 1388 -3078 1392 -3074
rect 1409 -3078 1413 -3074
rect 1430 -3078 1434 -3074
rect 1451 -3078 1455 -3074
rect 1472 -3078 1476 -3074
rect 1493 -3078 1497 -3074
rect 1513 -3078 1517 -3074
rect 1321 -3133 1325 -3086
rect 1321 -3154 1325 -3137
rect 1339 -3147 1343 -3086
rect 1355 -3147 1359 -3086
rect 1379 -3126 1383 -3086
rect 1379 -3147 1383 -3130
rect 1397 -3147 1401 -3086
rect 1421 -3133 1425 -3086
rect 1421 -3147 1425 -3137
rect 1439 -3126 1443 -3086
rect 1439 -3147 1443 -3130
rect 1463 -3140 1467 -3086
rect 1481 -3118 1485 -3086
rect 1481 -3126 1485 -3122
rect 1463 -3147 1467 -3144
rect 1339 -3151 1348 -3147
rect 1355 -3151 1363 -3147
rect 1339 -3154 1343 -3151
rect 1363 -3154 1367 -3151
rect 1371 -3151 1383 -3147
rect 1397 -3151 1405 -3147
rect 1371 -3154 1375 -3151
rect 1405 -3154 1409 -3151
rect 1413 -3151 1425 -3147
rect 1439 -3151 1451 -3147
rect 1413 -3154 1417 -3151
rect 1447 -3154 1451 -3151
rect 1455 -3151 1467 -3147
rect 1481 -3147 1485 -3130
rect 1505 -3133 1509 -3086
rect 1505 -3147 1509 -3137
rect 1481 -3151 1493 -3147
rect 1455 -3154 1459 -3151
rect 1489 -3154 1493 -3151
rect 1497 -3151 1509 -3147
rect 1497 -3154 1501 -3151
rect 1330 -3162 1334 -3158
rect 1347 -3162 1351 -3158
rect 1388 -3162 1392 -3158
rect 1430 -3162 1434 -3158
rect 1472 -3162 1476 -3158
rect 1513 -3162 1517 -3158
rect 1519 -3170 1523 -3122
rect 1330 -3199 1334 -3195
rect 1347 -3199 1351 -3195
rect 1367 -3199 1371 -3195
rect 1388 -3199 1392 -3195
rect 1409 -3199 1413 -3195
rect 1430 -3199 1434 -3195
rect 1451 -3199 1455 -3195
rect 1472 -3199 1476 -3195
rect 1493 -3199 1497 -3195
rect 1513 -3199 1517 -3195
rect 1321 -3254 1325 -3207
rect 1321 -3275 1325 -3258
rect 1339 -3268 1343 -3207
rect 1355 -3268 1359 -3207
rect 1379 -3247 1383 -3207
rect 1379 -3268 1383 -3251
rect 1397 -3268 1401 -3207
rect 1421 -3254 1425 -3207
rect 1421 -3268 1425 -3258
rect 1439 -3247 1443 -3207
rect 1439 -3268 1443 -3251
rect 1463 -3261 1467 -3207
rect 1481 -3239 1485 -3207
rect 1481 -3247 1485 -3243
rect 1463 -3268 1467 -3265
rect 1339 -3272 1348 -3268
rect 1355 -3272 1363 -3268
rect 1339 -3275 1343 -3272
rect 1363 -3275 1367 -3272
rect 1371 -3272 1383 -3268
rect 1397 -3272 1405 -3268
rect 1371 -3275 1375 -3272
rect 1405 -3275 1409 -3272
rect 1413 -3272 1425 -3268
rect 1439 -3272 1451 -3268
rect 1413 -3275 1417 -3272
rect 1447 -3275 1451 -3272
rect 1455 -3272 1467 -3268
rect 1481 -3268 1485 -3251
rect 1505 -3254 1509 -3207
rect 1505 -3268 1509 -3258
rect 1481 -3272 1493 -3268
rect 1455 -3275 1459 -3272
rect 1489 -3275 1493 -3272
rect 1497 -3272 1509 -3268
rect 1497 -3275 1501 -3272
rect 1330 -3283 1334 -3279
rect 1347 -3283 1351 -3279
rect 1388 -3283 1392 -3279
rect 1430 -3283 1434 -3279
rect 1472 -3283 1476 -3279
rect 1513 -3283 1517 -3279
rect 1321 -3430 1325 -3426
rect 1338 -3430 1342 -3426
rect 1329 -3441 1333 -3438
rect 1329 -3445 1344 -3441
rect 1315 -3458 1322 -3454
rect 972 -3915 976 -3911
rect 989 -3915 993 -3911
rect 1009 -3915 1013 -3911
rect 1030 -3915 1034 -3911
rect 1051 -3915 1055 -3911
rect 1072 -3915 1076 -3911
rect 1093 -3915 1097 -3911
rect 1114 -3915 1118 -3911
rect 1135 -3915 1139 -3911
rect 1155 -3915 1159 -3911
rect 963 -3970 967 -3923
rect 963 -3991 967 -3974
rect 981 -3984 985 -3923
rect 997 -3984 1001 -3923
rect 1021 -3963 1025 -3923
rect 1021 -3984 1025 -3967
rect 1039 -3984 1043 -3923
rect 1063 -3970 1067 -3923
rect 1063 -3984 1067 -3974
rect 1081 -3963 1085 -3923
rect 1081 -3984 1085 -3967
rect 1105 -3977 1109 -3923
rect 1123 -3955 1127 -3923
rect 1123 -3963 1127 -3959
rect 1105 -3984 1109 -3981
rect 981 -3988 990 -3984
rect 997 -3988 1005 -3984
rect 981 -3991 985 -3988
rect 1005 -3991 1009 -3988
rect 1013 -3988 1025 -3984
rect 1039 -3988 1047 -3984
rect 1013 -3991 1017 -3988
rect 1047 -3991 1051 -3988
rect 1055 -3988 1067 -3984
rect 1081 -3988 1093 -3984
rect 1055 -3991 1059 -3988
rect 1089 -3991 1093 -3988
rect 1097 -3988 1109 -3984
rect 1123 -3984 1127 -3967
rect 1147 -3970 1151 -3923
rect 1147 -3984 1151 -3974
rect 1123 -3988 1135 -3984
rect 1097 -3991 1101 -3988
rect 1131 -3991 1135 -3988
rect 1139 -3988 1151 -3984
rect 1139 -3991 1143 -3988
rect 972 -3999 976 -3995
rect 989 -3999 993 -3995
rect 1030 -3999 1034 -3995
rect 1072 -3999 1076 -3995
rect 1114 -3999 1118 -3995
rect 1155 -3999 1159 -3995
rect 1161 -4006 1165 -3959
rect 1309 -3963 1313 -3656
rect 972 -4040 976 -4036
rect 989 -4040 993 -4036
rect 1009 -4040 1013 -4036
rect 1030 -4040 1034 -4036
rect 1051 -4040 1055 -4036
rect 1072 -4040 1076 -4036
rect 1093 -4040 1097 -4036
rect 1114 -4040 1118 -4036
rect 1135 -4040 1139 -4036
rect 1155 -4040 1159 -4036
rect 963 -4095 967 -4048
rect 963 -4116 967 -4099
rect 981 -4109 985 -4048
rect 997 -4109 1001 -4048
rect 1021 -4088 1025 -4048
rect 1021 -4109 1025 -4092
rect 1039 -4109 1043 -4048
rect 1063 -4095 1067 -4048
rect 1063 -4109 1067 -4099
rect 1081 -4088 1085 -4048
rect 1081 -4109 1085 -4092
rect 1105 -4102 1109 -4048
rect 1123 -4080 1127 -4048
rect 1123 -4088 1127 -4084
rect 1105 -4109 1109 -4106
rect 981 -4113 990 -4109
rect 997 -4113 1005 -4109
rect 981 -4116 985 -4113
rect 1005 -4116 1009 -4113
rect 1013 -4113 1025 -4109
rect 1039 -4113 1047 -4109
rect 1013 -4116 1017 -4113
rect 1047 -4116 1051 -4113
rect 1055 -4113 1067 -4109
rect 1081 -4113 1093 -4109
rect 1055 -4116 1059 -4113
rect 1089 -4116 1093 -4113
rect 1097 -4113 1109 -4109
rect 1123 -4109 1127 -4092
rect 1147 -4095 1151 -4048
rect 1147 -4109 1151 -4099
rect 1123 -4113 1135 -4109
rect 1097 -4116 1101 -4113
rect 1131 -4116 1135 -4113
rect 1139 -4113 1151 -4109
rect 1139 -4116 1143 -4113
rect 972 -4124 976 -4120
rect 989 -4124 993 -4120
rect 1030 -4124 1034 -4120
rect 1072 -4124 1076 -4120
rect 1114 -4124 1118 -4120
rect 1155 -4124 1159 -4120
rect 963 -4275 967 -4271
rect 980 -4275 984 -4271
rect 971 -4286 975 -4283
rect 971 -4290 986 -4286
rect 957 -4303 964 -4299
rect 574 -4638 578 -4634
rect 591 -4638 595 -4634
rect 611 -4638 615 -4634
rect 632 -4638 636 -4634
rect 653 -4638 657 -4634
rect 674 -4638 678 -4634
rect 695 -4638 699 -4634
rect 716 -4638 720 -4634
rect 737 -4638 741 -4634
rect 757 -4638 761 -4634
rect 565 -4693 569 -4646
rect 565 -4714 569 -4697
rect 583 -4707 587 -4646
rect 599 -4707 603 -4646
rect 623 -4686 627 -4646
rect 623 -4707 627 -4690
rect 641 -4707 645 -4646
rect 665 -4693 669 -4646
rect 665 -4707 669 -4697
rect 683 -4686 687 -4646
rect 683 -4707 687 -4690
rect 707 -4700 711 -4646
rect 725 -4678 729 -4646
rect 725 -4686 729 -4682
rect 707 -4707 711 -4704
rect 583 -4711 592 -4707
rect 599 -4711 607 -4707
rect 583 -4714 587 -4711
rect 607 -4714 611 -4711
rect 615 -4711 627 -4707
rect 641 -4711 649 -4707
rect 615 -4714 619 -4711
rect 649 -4714 653 -4711
rect 657 -4711 669 -4707
rect 683 -4711 695 -4707
rect 657 -4714 661 -4711
rect 691 -4714 695 -4711
rect 699 -4711 711 -4707
rect 725 -4707 729 -4690
rect 749 -4693 753 -4646
rect 749 -4707 753 -4697
rect 725 -4711 737 -4707
rect 699 -4714 703 -4711
rect 733 -4714 737 -4711
rect 741 -4711 753 -4707
rect 741 -4714 745 -4711
rect 574 -4722 578 -4718
rect 591 -4722 595 -4718
rect 632 -4722 636 -4718
rect 674 -4722 678 -4718
rect 716 -4722 720 -4718
rect 757 -4722 761 -4718
rect 763 -4730 767 -4682
rect 951 -4686 955 -4489
rect 574 -4759 578 -4755
rect 591 -4759 595 -4755
rect 611 -4759 615 -4755
rect 632 -4759 636 -4755
rect 653 -4759 657 -4755
rect 674 -4759 678 -4755
rect 695 -4759 699 -4755
rect 716 -4759 720 -4755
rect 737 -4759 741 -4755
rect 757 -4759 761 -4755
rect 565 -4814 569 -4767
rect 565 -4835 569 -4818
rect 583 -4828 587 -4767
rect 599 -4828 603 -4767
rect 623 -4807 627 -4767
rect 623 -4828 627 -4811
rect 641 -4828 645 -4767
rect 665 -4814 669 -4767
rect 665 -4828 669 -4818
rect 683 -4807 687 -4767
rect 683 -4828 687 -4811
rect 707 -4821 711 -4767
rect 725 -4799 729 -4767
rect 725 -4807 729 -4803
rect 707 -4828 711 -4825
rect 583 -4832 592 -4828
rect 599 -4832 607 -4828
rect 583 -4835 587 -4832
rect 607 -4835 611 -4832
rect 615 -4832 627 -4828
rect 641 -4832 649 -4828
rect 615 -4835 619 -4832
rect 649 -4835 653 -4832
rect 657 -4832 669 -4828
rect 683 -4832 695 -4828
rect 657 -4835 661 -4832
rect 691 -4835 695 -4832
rect 699 -4832 711 -4828
rect 725 -4828 729 -4811
rect 749 -4814 753 -4767
rect 749 -4828 753 -4818
rect 725 -4832 737 -4828
rect 699 -4835 703 -4832
rect 733 -4835 737 -4832
rect 741 -4832 753 -4828
rect 741 -4835 745 -4832
rect 574 -4843 578 -4839
rect 591 -4843 595 -4839
rect 632 -4843 636 -4839
rect 674 -4843 678 -4839
rect 716 -4843 720 -4839
rect 757 -4843 761 -4839
rect 565 -4994 569 -4990
rect 582 -4994 586 -4990
rect 573 -5005 577 -5002
rect 573 -5009 588 -5005
rect 559 -5022 566 -5018
rect 218 -5353 222 -5349
rect 235 -5353 239 -5349
rect 255 -5353 259 -5349
rect 276 -5353 280 -5349
rect 297 -5353 301 -5349
rect 318 -5353 322 -5349
rect 339 -5353 343 -5349
rect 360 -5353 364 -5349
rect 381 -5353 385 -5349
rect 401 -5353 405 -5349
rect 466 -5353 470 -5349
rect 209 -5408 213 -5361
rect 209 -5429 213 -5412
rect 227 -5422 231 -5361
rect 243 -5422 247 -5361
rect 267 -5401 271 -5361
rect 267 -5422 271 -5405
rect 285 -5422 289 -5361
rect 309 -5408 313 -5361
rect 309 -5422 313 -5412
rect 327 -5401 331 -5361
rect 327 -5422 331 -5405
rect 351 -5415 355 -5361
rect 369 -5393 373 -5361
rect 369 -5401 373 -5397
rect 351 -5422 355 -5419
rect 227 -5426 236 -5422
rect 243 -5426 251 -5422
rect 227 -5429 231 -5426
rect 251 -5429 255 -5426
rect 259 -5426 271 -5422
rect 285 -5426 293 -5422
rect 259 -5429 263 -5426
rect 293 -5429 297 -5426
rect 301 -5426 313 -5422
rect 327 -5426 339 -5422
rect 301 -5429 305 -5426
rect 335 -5429 339 -5426
rect 343 -5426 355 -5422
rect 369 -5422 373 -5405
rect 393 -5408 397 -5361
rect 474 -5390 478 -5361
rect 393 -5422 397 -5412
rect 369 -5426 381 -5422
rect 343 -5429 347 -5426
rect 377 -5429 381 -5426
rect 385 -5426 397 -5422
rect 385 -5429 389 -5426
rect 218 -5437 222 -5433
rect 235 -5437 239 -5433
rect 276 -5437 280 -5433
rect 318 -5437 322 -5433
rect 360 -5437 364 -5433
rect 401 -5437 405 -5433
rect 407 -5444 411 -5397
rect 474 -5429 478 -5394
rect 553 -5401 557 -5215
rect 466 -5437 470 -5433
rect 218 -5473 222 -5469
rect 235 -5473 239 -5469
rect 255 -5473 259 -5469
rect 276 -5473 280 -5469
rect 297 -5473 301 -5469
rect 318 -5473 322 -5469
rect 339 -5473 343 -5469
rect 360 -5473 364 -5469
rect 381 -5473 385 -5469
rect 401 -5473 405 -5469
rect 466 -5473 470 -5469
rect 209 -5528 213 -5481
rect 209 -5549 213 -5532
rect 227 -5542 231 -5481
rect 243 -5542 247 -5481
rect 267 -5521 271 -5481
rect 267 -5542 271 -5525
rect 285 -5542 289 -5481
rect 309 -5528 313 -5481
rect 309 -5542 313 -5532
rect 327 -5521 331 -5481
rect 327 -5542 331 -5525
rect 351 -5535 355 -5481
rect 369 -5513 373 -5481
rect 369 -5521 373 -5517
rect 351 -5542 355 -5539
rect 227 -5546 236 -5542
rect 243 -5546 251 -5542
rect 227 -5549 231 -5546
rect 251 -5549 255 -5546
rect 259 -5546 271 -5542
rect 285 -5546 293 -5542
rect 259 -5549 263 -5546
rect 293 -5549 297 -5546
rect 301 -5546 313 -5542
rect 327 -5546 339 -5542
rect 301 -5549 305 -5546
rect 335 -5549 339 -5546
rect 343 -5546 355 -5542
rect 369 -5542 373 -5525
rect 393 -5528 397 -5481
rect 393 -5542 397 -5532
rect 369 -5546 381 -5542
rect 343 -5549 347 -5546
rect 377 -5549 381 -5546
rect 385 -5546 397 -5542
rect 385 -5549 389 -5546
rect 218 -5557 222 -5553
rect 235 -5557 239 -5553
rect 276 -5557 280 -5553
rect 318 -5557 322 -5553
rect 360 -5557 364 -5553
rect 401 -5557 405 -5553
rect 218 -5590 222 -5586
rect 235 -5590 239 -5586
rect 255 -5590 259 -5586
rect 276 -5590 280 -5586
rect 297 -5590 301 -5586
rect 318 -5590 322 -5586
rect 339 -5590 343 -5586
rect 360 -5590 364 -5586
rect 381 -5590 385 -5586
rect 401 -5590 405 -5586
rect 209 -5645 213 -5598
rect 209 -5666 213 -5649
rect 227 -5659 231 -5598
rect 243 -5659 247 -5598
rect 267 -5638 271 -5598
rect 267 -5659 271 -5642
rect 285 -5659 289 -5598
rect 309 -5645 313 -5598
rect 309 -5659 313 -5649
rect 327 -5638 331 -5598
rect 327 -5659 331 -5642
rect 351 -5652 355 -5598
rect 369 -5630 373 -5598
rect 369 -5638 373 -5634
rect 351 -5659 355 -5656
rect 227 -5663 236 -5659
rect 243 -5663 251 -5659
rect 227 -5666 231 -5663
rect 251 -5666 255 -5663
rect 259 -5663 271 -5659
rect 285 -5663 293 -5659
rect 259 -5666 263 -5663
rect 293 -5666 297 -5663
rect 301 -5663 313 -5659
rect 327 -5663 339 -5659
rect 301 -5666 305 -5663
rect 335 -5666 339 -5663
rect 343 -5663 355 -5659
rect 369 -5659 373 -5642
rect 393 -5645 397 -5598
rect 393 -5659 397 -5649
rect 369 -5663 381 -5659
rect 343 -5666 347 -5663
rect 377 -5666 381 -5663
rect 385 -5663 397 -5659
rect 385 -5666 389 -5663
rect 218 -5674 222 -5670
rect 235 -5674 239 -5670
rect 276 -5674 280 -5670
rect 318 -5674 322 -5670
rect 360 -5674 364 -5670
rect 401 -5674 405 -5670
rect 209 -5707 213 -5703
rect 226 -5707 230 -5703
rect 217 -5718 221 -5715
rect 217 -5722 232 -5718
rect 228 -5761 232 -5722
rect 228 -5776 232 -5765
rect 209 -5780 232 -5776
rect 235 -5752 239 -5715
rect 407 -5731 411 -5517
rect 474 -5514 478 -5481
rect 474 -5549 478 -5518
rect 466 -5557 470 -5553
rect 209 -5783 213 -5780
rect 235 -5783 239 -5756
rect 226 -5791 230 -5787
rect 218 -5826 222 -5822
rect 244 -5826 248 -5822
rect 261 -5826 265 -5822
rect 301 -5826 305 -5822
rect 322 -5826 326 -5822
rect 339 -5826 343 -5822
rect 379 -5826 383 -5822
rect 403 -5826 407 -5822
rect 440 -5826 444 -5822
rect 209 -5851 213 -5834
rect 209 -5902 213 -5855
rect 227 -5844 231 -5834
rect 227 -5902 231 -5848
rect 235 -5873 239 -5834
rect 253 -5866 257 -5834
rect 235 -5902 239 -5877
rect 253 -5902 257 -5870
rect 279 -5858 283 -5834
rect 279 -5895 283 -5862
rect 313 -5895 317 -5834
rect 331 -5851 335 -5834
rect 261 -5902 265 -5899
rect 269 -5899 283 -5895
rect 269 -5902 273 -5899
rect 297 -5902 301 -5899
rect 305 -5899 324 -5895
rect 305 -5902 309 -5899
rect 331 -5902 335 -5855
rect 357 -5866 361 -5834
rect 357 -5895 361 -5870
rect 391 -5888 395 -5834
rect 391 -5892 408 -5888
rect 339 -5902 343 -5899
rect 348 -5899 361 -5895
rect 348 -5902 352 -5899
rect 375 -5902 379 -5899
rect 399 -5902 403 -5892
rect 415 -5895 419 -5834
rect 423 -5888 427 -5834
rect 449 -5858 453 -5834
rect 423 -5892 442 -5888
rect 407 -5899 424 -5895
rect 407 -5902 411 -5899
rect 431 -5902 435 -5892
rect 449 -5902 453 -5862
rect 218 -5910 222 -5906
rect 244 -5910 248 -5906
rect 287 -5910 291 -5906
rect 322 -5910 326 -5906
rect 366 -5910 370 -5906
rect 383 -5910 387 -5906
rect 419 -5910 423 -5906
rect 440 -5910 444 -5906
rect 455 -5918 459 -5870
rect 547 -5873 551 -5756
rect 553 -5858 557 -5450
rect 559 -5521 563 -5022
rect 584 -5048 588 -5009
rect 584 -5063 588 -5052
rect 565 -5067 588 -5063
rect 591 -5039 595 -5002
rect 763 -5018 767 -4803
rect 565 -5070 569 -5067
rect 591 -5070 595 -5043
rect 582 -5078 586 -5074
rect 574 -5113 578 -5109
rect 600 -5113 604 -5109
rect 617 -5113 621 -5109
rect 657 -5113 661 -5109
rect 678 -5113 682 -5109
rect 695 -5113 699 -5109
rect 735 -5113 739 -5109
rect 759 -5113 763 -5109
rect 796 -5113 800 -5109
rect 565 -5138 569 -5121
rect 565 -5189 569 -5142
rect 583 -5131 587 -5121
rect 583 -5189 587 -5135
rect 591 -5160 595 -5121
rect 609 -5153 613 -5121
rect 591 -5189 595 -5164
rect 609 -5189 613 -5157
rect 635 -5145 639 -5121
rect 635 -5182 639 -5149
rect 669 -5182 673 -5121
rect 687 -5138 691 -5121
rect 617 -5189 621 -5186
rect 625 -5186 639 -5182
rect 625 -5189 629 -5186
rect 653 -5189 657 -5186
rect 661 -5186 680 -5182
rect 661 -5189 665 -5186
rect 687 -5189 691 -5142
rect 713 -5153 717 -5121
rect 713 -5182 717 -5157
rect 747 -5175 751 -5121
rect 747 -5179 764 -5175
rect 695 -5189 699 -5186
rect 704 -5186 717 -5182
rect 704 -5189 708 -5186
rect 731 -5189 735 -5186
rect 755 -5189 759 -5179
rect 771 -5182 775 -5121
rect 779 -5175 783 -5121
rect 805 -5145 809 -5121
rect 779 -5179 798 -5175
rect 763 -5186 780 -5182
rect 763 -5189 767 -5186
rect 787 -5189 791 -5179
rect 805 -5189 809 -5149
rect 574 -5197 578 -5193
rect 600 -5197 604 -5193
rect 643 -5197 647 -5193
rect 678 -5197 682 -5193
rect 722 -5197 726 -5193
rect 739 -5197 743 -5193
rect 775 -5197 779 -5193
rect 796 -5197 800 -5193
rect 811 -5204 815 -5157
rect 945 -5160 949 -5043
rect 951 -5145 955 -4733
rect 957 -4807 961 -4303
rect 982 -4329 986 -4290
rect 982 -4344 986 -4333
rect 963 -4348 986 -4344
rect 989 -4320 993 -4283
rect 1161 -4299 1165 -4084
rect 1201 -4164 1205 -4160
rect 1209 -4201 1213 -4172
rect 1209 -4240 1213 -4205
rect 1201 -4248 1205 -4244
rect 1201 -4275 1205 -4271
rect 1209 -4316 1213 -4283
rect 963 -4351 967 -4348
rect 989 -4351 993 -4324
rect 1209 -4351 1213 -4320
rect 980 -4359 984 -4355
rect 1201 -4359 1205 -4355
rect 972 -4394 976 -4390
rect 998 -4394 1002 -4390
rect 1015 -4394 1019 -4390
rect 1055 -4394 1059 -4390
rect 1076 -4394 1080 -4390
rect 1093 -4394 1097 -4390
rect 1133 -4394 1137 -4390
rect 1157 -4394 1161 -4390
rect 1194 -4394 1198 -4390
rect 963 -4419 967 -4402
rect 963 -4470 967 -4423
rect 981 -4412 985 -4402
rect 981 -4470 985 -4416
rect 989 -4441 993 -4402
rect 1007 -4434 1011 -4402
rect 989 -4470 993 -4445
rect 1007 -4470 1011 -4438
rect 1033 -4426 1037 -4402
rect 1033 -4463 1037 -4430
rect 1067 -4463 1071 -4402
rect 1085 -4419 1089 -4402
rect 1015 -4470 1019 -4467
rect 1023 -4467 1037 -4463
rect 1023 -4470 1027 -4467
rect 1051 -4470 1055 -4467
rect 1059 -4467 1078 -4463
rect 1059 -4470 1063 -4467
rect 1085 -4470 1089 -4423
rect 1111 -4434 1115 -4402
rect 1111 -4463 1115 -4438
rect 1145 -4456 1149 -4402
rect 1145 -4460 1162 -4456
rect 1093 -4470 1097 -4467
rect 1102 -4467 1115 -4463
rect 1102 -4470 1106 -4467
rect 1129 -4470 1133 -4467
rect 1153 -4470 1157 -4460
rect 1169 -4463 1173 -4402
rect 1177 -4456 1181 -4402
rect 1203 -4424 1207 -4402
rect 1177 -4460 1196 -4456
rect 1161 -4467 1178 -4463
rect 1161 -4470 1165 -4467
rect 1185 -4470 1189 -4460
rect 1203 -4470 1207 -4428
rect 1303 -4426 1307 -4324
rect 972 -4478 976 -4474
rect 998 -4478 1002 -4474
rect 1041 -4478 1045 -4474
rect 1076 -4478 1080 -4474
rect 1120 -4478 1124 -4474
rect 1137 -4478 1141 -4474
rect 1173 -4478 1177 -4474
rect 1194 -4478 1198 -4474
rect 1209 -4492 1213 -4438
rect 1309 -4441 1313 -4010
rect 1315 -4088 1319 -3458
rect 1340 -3484 1344 -3445
rect 1340 -3499 1344 -3488
rect 1321 -3503 1344 -3499
rect 1347 -3475 1351 -3438
rect 1519 -3454 1523 -3243
rect 1321 -3506 1325 -3503
rect 1347 -3506 1351 -3479
rect 1338 -3514 1342 -3510
rect 1330 -3554 1334 -3550
rect 1356 -3554 1360 -3550
rect 1373 -3554 1377 -3550
rect 1413 -3554 1417 -3550
rect 1434 -3554 1438 -3550
rect 1451 -3554 1455 -3550
rect 1491 -3554 1495 -3550
rect 1515 -3554 1519 -3550
rect 1552 -3554 1556 -3550
rect 1321 -3579 1325 -3562
rect 1321 -3630 1325 -3583
rect 1339 -3572 1343 -3562
rect 1339 -3630 1343 -3576
rect 1347 -3601 1351 -3562
rect 1365 -3594 1369 -3562
rect 1347 -3630 1351 -3605
rect 1365 -3630 1369 -3598
rect 1391 -3586 1395 -3562
rect 1391 -3623 1395 -3590
rect 1425 -3623 1429 -3562
rect 1443 -3579 1447 -3562
rect 1373 -3630 1377 -3627
rect 1381 -3627 1395 -3623
rect 1381 -3630 1385 -3627
rect 1409 -3630 1413 -3627
rect 1417 -3627 1436 -3623
rect 1417 -3630 1421 -3627
rect 1443 -3630 1447 -3583
rect 1469 -3594 1473 -3562
rect 1469 -3623 1473 -3598
rect 1503 -3616 1507 -3562
rect 1503 -3620 1520 -3616
rect 1451 -3630 1455 -3627
rect 1460 -3627 1473 -3623
rect 1460 -3630 1464 -3627
rect 1487 -3630 1491 -3627
rect 1511 -3630 1515 -3620
rect 1527 -3623 1531 -3562
rect 1535 -3616 1539 -3562
rect 1535 -3620 1554 -3616
rect 1519 -3627 1536 -3623
rect 1519 -3630 1523 -3627
rect 1543 -3630 1547 -3620
rect 1561 -3630 1565 -3562
rect 1330 -3638 1334 -3634
rect 1356 -3638 1360 -3634
rect 1399 -3638 1403 -3634
rect 1434 -3638 1438 -3634
rect 1478 -3638 1482 -3634
rect 1495 -3638 1499 -3634
rect 1531 -3638 1535 -3634
rect 1552 -3638 1556 -3634
rect 1561 -3652 1565 -3634
rect 1567 -3645 1571 -3598
rect 1330 -3915 1334 -3911
rect 1347 -3915 1351 -3911
rect 1367 -3915 1371 -3911
rect 1388 -3915 1392 -3911
rect 1409 -3915 1413 -3911
rect 1430 -3915 1434 -3911
rect 1451 -3915 1455 -3911
rect 1472 -3915 1476 -3911
rect 1493 -3915 1497 -3911
rect 1513 -3915 1517 -3911
rect 1321 -3970 1325 -3923
rect 1321 -3991 1325 -3974
rect 1339 -3984 1343 -3923
rect 1355 -3984 1359 -3923
rect 1379 -3963 1383 -3923
rect 1379 -3984 1383 -3967
rect 1397 -3984 1401 -3923
rect 1421 -3970 1425 -3923
rect 1421 -3984 1425 -3974
rect 1439 -3963 1443 -3923
rect 1439 -3984 1443 -3967
rect 1463 -3977 1467 -3923
rect 1481 -3955 1485 -3923
rect 1481 -3963 1485 -3959
rect 1463 -3984 1467 -3981
rect 1339 -3988 1348 -3984
rect 1355 -3988 1363 -3984
rect 1339 -3991 1343 -3988
rect 1363 -3991 1367 -3988
rect 1371 -3988 1383 -3984
rect 1397 -3988 1405 -3984
rect 1371 -3991 1375 -3988
rect 1405 -3991 1409 -3988
rect 1413 -3988 1425 -3984
rect 1439 -3988 1451 -3984
rect 1413 -3991 1417 -3988
rect 1447 -3991 1451 -3988
rect 1455 -3988 1467 -3984
rect 1481 -3984 1485 -3967
rect 1505 -3970 1509 -3923
rect 1505 -3984 1509 -3974
rect 1481 -3988 1493 -3984
rect 1455 -3991 1459 -3988
rect 1489 -3991 1493 -3988
rect 1497 -3988 1509 -3984
rect 1497 -3991 1501 -3988
rect 1330 -3999 1334 -3995
rect 1347 -3999 1351 -3995
rect 1388 -3999 1392 -3995
rect 1430 -3999 1434 -3995
rect 1472 -3999 1476 -3995
rect 1513 -3999 1517 -3995
rect 1519 -4006 1523 -3959
rect 1330 -4040 1334 -4036
rect 1347 -4040 1351 -4036
rect 1367 -4040 1371 -4036
rect 1388 -4040 1392 -4036
rect 1409 -4040 1413 -4036
rect 1430 -4040 1434 -4036
rect 1451 -4040 1455 -4036
rect 1472 -4040 1476 -4036
rect 1493 -4040 1497 -4036
rect 1513 -4040 1517 -4036
rect 1321 -4095 1325 -4048
rect 1321 -4116 1325 -4099
rect 1339 -4109 1343 -4048
rect 1355 -4109 1359 -4048
rect 1379 -4088 1383 -4048
rect 1379 -4109 1383 -4092
rect 1397 -4109 1401 -4048
rect 1421 -4095 1425 -4048
rect 1421 -4109 1425 -4099
rect 1439 -4088 1443 -4048
rect 1439 -4109 1443 -4092
rect 1463 -4102 1467 -4048
rect 1481 -4080 1485 -4048
rect 1481 -4088 1485 -4084
rect 1463 -4109 1467 -4106
rect 1339 -4113 1348 -4109
rect 1355 -4113 1363 -4109
rect 1339 -4116 1343 -4113
rect 1363 -4116 1367 -4113
rect 1371 -4113 1383 -4109
rect 1397 -4113 1405 -4109
rect 1371 -4116 1375 -4113
rect 1405 -4116 1409 -4113
rect 1413 -4113 1425 -4109
rect 1439 -4113 1451 -4109
rect 1413 -4116 1417 -4113
rect 1447 -4116 1451 -4113
rect 1455 -4113 1467 -4109
rect 1481 -4109 1485 -4092
rect 1505 -4095 1509 -4048
rect 1505 -4109 1509 -4099
rect 1481 -4113 1493 -4109
rect 1455 -4116 1459 -4113
rect 1489 -4116 1493 -4113
rect 1497 -4113 1509 -4109
rect 1497 -4116 1501 -4113
rect 1330 -4124 1334 -4120
rect 1347 -4124 1351 -4120
rect 1388 -4124 1392 -4120
rect 1430 -4124 1434 -4120
rect 1472 -4124 1476 -4120
rect 1513 -4124 1517 -4120
rect 1321 -4275 1325 -4271
rect 1338 -4275 1342 -4271
rect 1329 -4286 1333 -4283
rect 1329 -4290 1344 -4286
rect 1315 -4303 1322 -4299
rect 972 -4638 976 -4634
rect 989 -4638 993 -4634
rect 1009 -4638 1013 -4634
rect 1030 -4638 1034 -4634
rect 1051 -4638 1055 -4634
rect 1072 -4638 1076 -4634
rect 1093 -4638 1097 -4634
rect 1114 -4638 1118 -4634
rect 1135 -4638 1139 -4634
rect 1155 -4638 1159 -4634
rect 963 -4693 967 -4646
rect 963 -4714 967 -4697
rect 981 -4707 985 -4646
rect 997 -4707 1001 -4646
rect 1021 -4686 1025 -4646
rect 1021 -4707 1025 -4690
rect 1039 -4707 1043 -4646
rect 1063 -4693 1067 -4646
rect 1063 -4707 1067 -4697
rect 1081 -4686 1085 -4646
rect 1081 -4707 1085 -4690
rect 1105 -4700 1109 -4646
rect 1123 -4678 1127 -4646
rect 1123 -4686 1127 -4682
rect 1105 -4707 1109 -4704
rect 981 -4711 990 -4707
rect 997 -4711 1005 -4707
rect 981 -4714 985 -4711
rect 1005 -4714 1009 -4711
rect 1013 -4711 1025 -4707
rect 1039 -4711 1047 -4707
rect 1013 -4714 1017 -4711
rect 1047 -4714 1051 -4711
rect 1055 -4711 1067 -4707
rect 1081 -4711 1093 -4707
rect 1055 -4714 1059 -4711
rect 1089 -4714 1093 -4711
rect 1097 -4711 1109 -4707
rect 1123 -4707 1127 -4690
rect 1147 -4693 1151 -4646
rect 1147 -4707 1151 -4697
rect 1123 -4711 1135 -4707
rect 1097 -4714 1101 -4711
rect 1131 -4714 1135 -4711
rect 1139 -4711 1151 -4707
rect 1139 -4714 1143 -4711
rect 972 -4722 976 -4718
rect 989 -4722 993 -4718
rect 1030 -4722 1034 -4718
rect 1072 -4722 1076 -4718
rect 1114 -4722 1118 -4718
rect 1155 -4722 1159 -4718
rect 1161 -4729 1165 -4682
rect 1309 -4686 1313 -4496
rect 972 -4759 976 -4755
rect 989 -4759 993 -4755
rect 1009 -4759 1013 -4755
rect 1030 -4759 1034 -4755
rect 1051 -4759 1055 -4755
rect 1072 -4759 1076 -4755
rect 1093 -4759 1097 -4755
rect 1114 -4759 1118 -4755
rect 1135 -4759 1139 -4755
rect 1155 -4759 1159 -4755
rect 963 -4814 967 -4767
rect 963 -4835 967 -4818
rect 981 -4828 985 -4767
rect 997 -4828 1001 -4767
rect 1021 -4807 1025 -4767
rect 1021 -4828 1025 -4811
rect 1039 -4828 1043 -4767
rect 1063 -4814 1067 -4767
rect 1063 -4828 1067 -4818
rect 1081 -4807 1085 -4767
rect 1081 -4828 1085 -4811
rect 1105 -4821 1109 -4767
rect 1123 -4799 1127 -4767
rect 1123 -4807 1127 -4803
rect 1105 -4828 1109 -4825
rect 981 -4832 990 -4828
rect 997 -4832 1005 -4828
rect 981 -4835 985 -4832
rect 1005 -4835 1009 -4832
rect 1013 -4832 1025 -4828
rect 1039 -4832 1047 -4828
rect 1013 -4835 1017 -4832
rect 1047 -4835 1051 -4832
rect 1055 -4832 1067 -4828
rect 1081 -4832 1093 -4828
rect 1055 -4835 1059 -4832
rect 1089 -4835 1093 -4832
rect 1097 -4832 1109 -4828
rect 1123 -4828 1127 -4811
rect 1147 -4814 1151 -4767
rect 1147 -4828 1151 -4818
rect 1123 -4832 1135 -4828
rect 1097 -4835 1101 -4832
rect 1131 -4835 1135 -4832
rect 1139 -4832 1151 -4828
rect 1139 -4835 1143 -4832
rect 972 -4843 976 -4839
rect 989 -4843 993 -4839
rect 1030 -4843 1034 -4839
rect 1072 -4843 1076 -4839
rect 1114 -4843 1118 -4839
rect 1155 -4843 1159 -4839
rect 963 -4994 967 -4990
rect 980 -4994 984 -4990
rect 971 -5005 975 -5002
rect 971 -5009 986 -5005
rect 957 -5022 964 -5018
rect 574 -5353 578 -5349
rect 591 -5353 595 -5349
rect 611 -5353 615 -5349
rect 632 -5353 636 -5349
rect 653 -5353 657 -5349
rect 674 -5353 678 -5349
rect 695 -5353 699 -5349
rect 716 -5353 720 -5349
rect 737 -5353 741 -5349
rect 757 -5353 761 -5349
rect 867 -5353 871 -5349
rect 565 -5408 569 -5361
rect 565 -5429 569 -5412
rect 583 -5422 587 -5361
rect 599 -5422 603 -5361
rect 623 -5401 627 -5361
rect 623 -5422 627 -5405
rect 641 -5422 645 -5361
rect 665 -5408 669 -5361
rect 665 -5422 669 -5412
rect 683 -5401 687 -5361
rect 683 -5422 687 -5405
rect 707 -5415 711 -5361
rect 725 -5393 729 -5361
rect 725 -5401 729 -5397
rect 707 -5422 711 -5419
rect 583 -5426 592 -5422
rect 599 -5426 607 -5422
rect 583 -5429 587 -5426
rect 607 -5429 611 -5426
rect 615 -5426 627 -5422
rect 641 -5426 649 -5422
rect 615 -5429 619 -5426
rect 649 -5429 653 -5426
rect 657 -5426 669 -5422
rect 683 -5426 695 -5422
rect 657 -5429 661 -5426
rect 691 -5429 695 -5426
rect 699 -5426 711 -5422
rect 725 -5422 729 -5405
rect 749 -5408 753 -5361
rect 749 -5422 753 -5412
rect 725 -5426 737 -5422
rect 699 -5429 703 -5426
rect 733 -5429 737 -5426
rect 741 -5426 753 -5422
rect 741 -5429 745 -5426
rect 574 -5437 578 -5433
rect 591 -5437 595 -5433
rect 632 -5437 636 -5433
rect 674 -5437 678 -5433
rect 716 -5437 720 -5433
rect 757 -5437 761 -5433
rect 763 -5446 767 -5397
rect 875 -5395 879 -5369
rect 875 -5425 879 -5399
rect 951 -5401 955 -5208
rect 867 -5437 871 -5433
rect 574 -5473 578 -5469
rect 591 -5473 595 -5469
rect 611 -5473 615 -5469
rect 632 -5473 636 -5469
rect 653 -5473 657 -5469
rect 674 -5473 678 -5469
rect 695 -5473 699 -5469
rect 716 -5473 720 -5469
rect 737 -5473 741 -5469
rect 757 -5473 761 -5469
rect 565 -5528 569 -5481
rect 565 -5549 569 -5532
rect 583 -5542 587 -5481
rect 599 -5542 603 -5481
rect 623 -5521 627 -5481
rect 623 -5542 627 -5525
rect 641 -5542 645 -5481
rect 665 -5528 669 -5481
rect 665 -5542 669 -5532
rect 683 -5521 687 -5481
rect 683 -5542 687 -5525
rect 707 -5535 711 -5481
rect 725 -5513 729 -5481
rect 725 -5521 729 -5517
rect 707 -5542 711 -5539
rect 583 -5546 592 -5542
rect 599 -5546 607 -5542
rect 583 -5549 587 -5546
rect 607 -5549 611 -5546
rect 615 -5546 627 -5542
rect 641 -5546 649 -5542
rect 615 -5549 619 -5546
rect 649 -5549 653 -5546
rect 657 -5546 669 -5542
rect 683 -5546 695 -5542
rect 657 -5549 661 -5546
rect 691 -5549 695 -5546
rect 699 -5546 711 -5542
rect 725 -5542 729 -5525
rect 749 -5528 753 -5481
rect 749 -5542 753 -5532
rect 725 -5546 737 -5542
rect 699 -5549 703 -5546
rect 733 -5549 737 -5546
rect 741 -5546 753 -5542
rect 741 -5549 745 -5546
rect 574 -5557 578 -5553
rect 591 -5557 595 -5553
rect 632 -5557 636 -5553
rect 674 -5557 678 -5553
rect 716 -5557 720 -5553
rect 757 -5557 761 -5553
rect 574 -5590 578 -5586
rect 591 -5590 595 -5586
rect 611 -5590 615 -5586
rect 632 -5590 636 -5586
rect 653 -5590 657 -5586
rect 674 -5590 678 -5586
rect 695 -5590 699 -5586
rect 716 -5590 720 -5586
rect 737 -5590 741 -5586
rect 757 -5590 761 -5586
rect 565 -5645 569 -5598
rect 565 -5666 569 -5649
rect 583 -5659 587 -5598
rect 599 -5659 603 -5598
rect 623 -5638 627 -5598
rect 623 -5659 627 -5642
rect 641 -5659 645 -5598
rect 665 -5645 669 -5598
rect 665 -5659 669 -5649
rect 683 -5638 687 -5598
rect 683 -5659 687 -5642
rect 707 -5652 711 -5598
rect 725 -5630 729 -5598
rect 725 -5638 729 -5634
rect 707 -5659 711 -5656
rect 583 -5663 592 -5659
rect 599 -5663 607 -5659
rect 583 -5666 587 -5663
rect 607 -5666 611 -5663
rect 615 -5663 627 -5659
rect 641 -5663 649 -5659
rect 615 -5666 619 -5663
rect 649 -5666 653 -5663
rect 657 -5663 669 -5659
rect 683 -5663 695 -5659
rect 657 -5666 661 -5663
rect 691 -5666 695 -5663
rect 699 -5663 711 -5659
rect 725 -5659 729 -5642
rect 749 -5645 753 -5598
rect 749 -5659 753 -5649
rect 725 -5663 737 -5659
rect 699 -5666 703 -5663
rect 733 -5666 737 -5663
rect 741 -5663 753 -5659
rect 741 -5666 745 -5663
rect 574 -5674 578 -5670
rect 591 -5674 595 -5670
rect 632 -5674 636 -5670
rect 674 -5674 678 -5670
rect 716 -5674 720 -5670
rect 757 -5674 761 -5670
rect 565 -5707 569 -5703
rect 582 -5707 586 -5703
rect 573 -5718 577 -5715
rect 573 -5722 588 -5718
rect 584 -5761 588 -5722
rect 584 -5776 588 -5765
rect 565 -5780 588 -5776
rect 591 -5752 595 -5715
rect 763 -5739 767 -5634
rect 769 -5731 773 -5517
rect 565 -5783 569 -5780
rect 591 -5783 595 -5756
rect 582 -5791 586 -5787
rect 574 -5826 578 -5822
rect 600 -5826 604 -5822
rect 617 -5826 621 -5822
rect 657 -5826 661 -5822
rect 678 -5826 682 -5822
rect 695 -5826 699 -5822
rect 735 -5826 739 -5822
rect 759 -5826 763 -5822
rect 796 -5826 800 -5822
rect 565 -5851 569 -5834
rect 565 -5902 569 -5855
rect 583 -5844 587 -5834
rect 583 -5902 587 -5848
rect 591 -5873 595 -5834
rect 609 -5866 613 -5834
rect 591 -5902 595 -5877
rect 609 -5902 613 -5870
rect 635 -5858 639 -5834
rect 635 -5895 639 -5862
rect 669 -5895 673 -5834
rect 687 -5851 691 -5834
rect 617 -5902 621 -5899
rect 625 -5899 639 -5895
rect 625 -5902 629 -5899
rect 653 -5902 657 -5899
rect 661 -5899 680 -5895
rect 661 -5902 665 -5899
rect 687 -5902 691 -5855
rect 713 -5866 717 -5834
rect 713 -5895 717 -5870
rect 747 -5888 751 -5834
rect 747 -5892 764 -5888
rect 695 -5902 699 -5899
rect 704 -5899 717 -5895
rect 704 -5902 708 -5899
rect 731 -5902 735 -5899
rect 755 -5902 759 -5892
rect 771 -5895 775 -5834
rect 779 -5888 783 -5834
rect 805 -5858 809 -5834
rect 779 -5892 798 -5888
rect 763 -5899 780 -5895
rect 763 -5902 767 -5899
rect 787 -5902 791 -5892
rect 805 -5902 809 -5862
rect 574 -5910 578 -5906
rect 600 -5910 604 -5906
rect 643 -5910 647 -5906
rect 678 -5910 682 -5906
rect 722 -5910 726 -5906
rect 739 -5910 743 -5906
rect 775 -5910 779 -5906
rect 796 -5910 800 -5906
rect 811 -5917 815 -5870
rect 945 -5873 949 -5756
rect 951 -5858 955 -5449
rect 957 -5521 961 -5022
rect 982 -5048 986 -5009
rect 982 -5063 986 -5052
rect 963 -5067 986 -5063
rect 989 -5039 993 -5002
rect 1161 -5018 1165 -4803
rect 963 -5070 967 -5067
rect 989 -5070 993 -5043
rect 980 -5078 984 -5074
rect 972 -5113 976 -5109
rect 998 -5113 1002 -5109
rect 1015 -5113 1019 -5109
rect 1055 -5113 1059 -5109
rect 1076 -5113 1080 -5109
rect 1093 -5113 1097 -5109
rect 1133 -5113 1137 -5109
rect 1157 -5113 1161 -5109
rect 1194 -5113 1198 -5109
rect 963 -5138 967 -5121
rect 963 -5189 967 -5142
rect 981 -5131 985 -5121
rect 981 -5189 985 -5135
rect 989 -5160 993 -5121
rect 1007 -5153 1011 -5121
rect 989 -5189 993 -5164
rect 1007 -5189 1011 -5157
rect 1033 -5145 1037 -5121
rect 1033 -5182 1037 -5149
rect 1067 -5182 1071 -5121
rect 1085 -5138 1089 -5121
rect 1015 -5189 1019 -5186
rect 1023 -5186 1037 -5182
rect 1023 -5189 1027 -5186
rect 1051 -5189 1055 -5186
rect 1059 -5186 1078 -5182
rect 1059 -5189 1063 -5186
rect 1085 -5189 1089 -5142
rect 1111 -5153 1115 -5121
rect 1111 -5182 1115 -5157
rect 1145 -5175 1149 -5121
rect 1145 -5179 1162 -5175
rect 1093 -5189 1097 -5186
rect 1102 -5186 1115 -5182
rect 1102 -5189 1106 -5186
rect 1129 -5189 1133 -5186
rect 1153 -5189 1157 -5179
rect 1169 -5182 1173 -5121
rect 1177 -5175 1181 -5121
rect 1203 -5143 1207 -5121
rect 1177 -5179 1196 -5175
rect 1161 -5186 1178 -5182
rect 1161 -5189 1165 -5186
rect 1185 -5189 1189 -5179
rect 1203 -5189 1207 -5147
rect 1303 -5145 1307 -5043
rect 972 -5197 976 -5193
rect 998 -5197 1002 -5193
rect 1041 -5197 1045 -5193
rect 1076 -5197 1080 -5193
rect 1120 -5197 1124 -5193
rect 1137 -5197 1141 -5193
rect 1173 -5197 1177 -5193
rect 1194 -5197 1198 -5193
rect 1209 -5211 1213 -5157
rect 1309 -5160 1313 -4733
rect 1315 -4807 1319 -4303
rect 1340 -4329 1344 -4290
rect 1340 -4344 1344 -4333
rect 1321 -4348 1344 -4344
rect 1347 -4320 1351 -4283
rect 1519 -4299 1523 -4084
rect 1321 -4351 1325 -4348
rect 1347 -4351 1351 -4324
rect 1338 -4359 1342 -4355
rect 1330 -4394 1334 -4390
rect 1356 -4394 1360 -4390
rect 1373 -4394 1377 -4390
rect 1413 -4394 1417 -4390
rect 1434 -4394 1438 -4390
rect 1451 -4394 1455 -4390
rect 1491 -4394 1495 -4390
rect 1515 -4394 1519 -4390
rect 1552 -4394 1556 -4390
rect 1321 -4419 1325 -4402
rect 1321 -4470 1325 -4423
rect 1339 -4412 1343 -4402
rect 1339 -4470 1343 -4416
rect 1347 -4441 1351 -4402
rect 1365 -4434 1369 -4402
rect 1347 -4470 1351 -4445
rect 1365 -4470 1369 -4438
rect 1391 -4426 1395 -4402
rect 1391 -4463 1395 -4430
rect 1425 -4463 1429 -4402
rect 1443 -4419 1447 -4402
rect 1373 -4470 1377 -4467
rect 1381 -4467 1395 -4463
rect 1381 -4470 1385 -4467
rect 1409 -4470 1413 -4467
rect 1417 -4467 1436 -4463
rect 1417 -4470 1421 -4467
rect 1443 -4470 1447 -4423
rect 1469 -4434 1473 -4402
rect 1469 -4463 1473 -4438
rect 1503 -4456 1507 -4402
rect 1503 -4460 1520 -4456
rect 1451 -4470 1455 -4467
rect 1460 -4467 1473 -4463
rect 1460 -4470 1464 -4467
rect 1487 -4470 1491 -4467
rect 1511 -4470 1515 -4460
rect 1527 -4463 1531 -4402
rect 1535 -4456 1539 -4402
rect 1535 -4460 1554 -4456
rect 1519 -4467 1536 -4463
rect 1519 -4470 1523 -4467
rect 1543 -4470 1547 -4460
rect 1561 -4470 1565 -4402
rect 1330 -4478 1334 -4474
rect 1356 -4478 1360 -4474
rect 1399 -4478 1403 -4474
rect 1434 -4478 1438 -4474
rect 1478 -4478 1482 -4474
rect 1495 -4478 1499 -4474
rect 1531 -4478 1535 -4474
rect 1552 -4478 1556 -4474
rect 1561 -4492 1565 -4474
rect 1567 -4485 1571 -4438
rect 1330 -4638 1334 -4634
rect 1347 -4638 1351 -4634
rect 1367 -4638 1371 -4634
rect 1388 -4638 1392 -4634
rect 1409 -4638 1413 -4634
rect 1430 -4638 1434 -4634
rect 1451 -4638 1455 -4634
rect 1472 -4638 1476 -4634
rect 1493 -4638 1497 -4634
rect 1513 -4638 1517 -4634
rect 1321 -4693 1325 -4646
rect 1321 -4714 1325 -4697
rect 1339 -4707 1343 -4646
rect 1355 -4707 1359 -4646
rect 1379 -4686 1383 -4646
rect 1379 -4707 1383 -4690
rect 1397 -4707 1401 -4646
rect 1421 -4693 1425 -4646
rect 1421 -4707 1425 -4697
rect 1439 -4686 1443 -4646
rect 1439 -4707 1443 -4690
rect 1463 -4700 1467 -4646
rect 1481 -4678 1485 -4646
rect 1481 -4686 1485 -4682
rect 1463 -4707 1467 -4704
rect 1339 -4711 1348 -4707
rect 1355 -4711 1363 -4707
rect 1339 -4714 1343 -4711
rect 1363 -4714 1367 -4711
rect 1371 -4711 1383 -4707
rect 1397 -4711 1405 -4707
rect 1371 -4714 1375 -4711
rect 1405 -4714 1409 -4711
rect 1413 -4711 1425 -4707
rect 1439 -4711 1451 -4707
rect 1413 -4714 1417 -4711
rect 1447 -4714 1451 -4711
rect 1455 -4711 1467 -4707
rect 1481 -4707 1485 -4690
rect 1505 -4693 1509 -4646
rect 1505 -4707 1509 -4697
rect 1481 -4711 1493 -4707
rect 1455 -4714 1459 -4711
rect 1489 -4714 1493 -4711
rect 1497 -4711 1509 -4707
rect 1497 -4714 1501 -4711
rect 1330 -4722 1334 -4718
rect 1347 -4722 1351 -4718
rect 1388 -4722 1392 -4718
rect 1430 -4722 1434 -4718
rect 1472 -4722 1476 -4718
rect 1513 -4722 1517 -4718
rect 1519 -4729 1523 -4682
rect 1330 -4759 1334 -4755
rect 1347 -4759 1351 -4755
rect 1367 -4759 1371 -4755
rect 1388 -4759 1392 -4755
rect 1409 -4759 1413 -4755
rect 1430 -4759 1434 -4755
rect 1451 -4759 1455 -4755
rect 1472 -4759 1476 -4755
rect 1493 -4759 1497 -4755
rect 1513 -4759 1517 -4755
rect 1321 -4814 1325 -4767
rect 1321 -4835 1325 -4818
rect 1339 -4828 1343 -4767
rect 1355 -4828 1359 -4767
rect 1379 -4807 1383 -4767
rect 1379 -4828 1383 -4811
rect 1397 -4828 1401 -4767
rect 1421 -4814 1425 -4767
rect 1421 -4828 1425 -4818
rect 1439 -4807 1443 -4767
rect 1439 -4828 1443 -4811
rect 1463 -4821 1467 -4767
rect 1481 -4799 1485 -4767
rect 1481 -4807 1485 -4803
rect 1463 -4828 1467 -4825
rect 1339 -4832 1348 -4828
rect 1355 -4832 1363 -4828
rect 1339 -4835 1343 -4832
rect 1363 -4835 1367 -4832
rect 1371 -4832 1383 -4828
rect 1397 -4832 1405 -4828
rect 1371 -4835 1375 -4832
rect 1405 -4835 1409 -4832
rect 1413 -4832 1425 -4828
rect 1439 -4832 1451 -4828
rect 1413 -4835 1417 -4832
rect 1447 -4835 1451 -4832
rect 1455 -4832 1467 -4828
rect 1481 -4828 1485 -4811
rect 1505 -4814 1509 -4767
rect 1505 -4828 1509 -4818
rect 1481 -4832 1493 -4828
rect 1455 -4835 1459 -4832
rect 1489 -4835 1493 -4832
rect 1497 -4832 1509 -4828
rect 1497 -4835 1501 -4832
rect 1330 -4843 1334 -4839
rect 1347 -4843 1351 -4839
rect 1388 -4843 1392 -4839
rect 1430 -4843 1434 -4839
rect 1472 -4843 1476 -4839
rect 1513 -4843 1517 -4839
rect 1321 -4994 1325 -4990
rect 1338 -4994 1342 -4990
rect 1329 -5005 1333 -5002
rect 1329 -5009 1344 -5005
rect 1315 -5022 1322 -5018
rect 972 -5353 976 -5349
rect 989 -5353 993 -5349
rect 1009 -5353 1013 -5349
rect 1030 -5353 1034 -5349
rect 1051 -5353 1055 -5349
rect 1072 -5353 1076 -5349
rect 1093 -5353 1097 -5349
rect 1114 -5353 1118 -5349
rect 1135 -5353 1139 -5349
rect 1155 -5353 1159 -5349
rect 1210 -5353 1214 -5349
rect 963 -5408 967 -5361
rect 963 -5429 967 -5412
rect 981 -5422 985 -5361
rect 997 -5422 1001 -5361
rect 1021 -5401 1025 -5361
rect 1021 -5422 1025 -5405
rect 1039 -5422 1043 -5361
rect 1063 -5408 1067 -5361
rect 1063 -5422 1067 -5412
rect 1081 -5401 1085 -5361
rect 1081 -5422 1085 -5405
rect 1105 -5415 1109 -5361
rect 1123 -5393 1127 -5361
rect 1123 -5401 1127 -5397
rect 1105 -5422 1109 -5419
rect 981 -5426 990 -5422
rect 997 -5426 1005 -5422
rect 981 -5429 985 -5426
rect 1005 -5429 1009 -5426
rect 1013 -5426 1025 -5422
rect 1039 -5426 1047 -5422
rect 1013 -5429 1017 -5426
rect 1047 -5429 1051 -5426
rect 1055 -5426 1067 -5422
rect 1081 -5426 1093 -5422
rect 1055 -5429 1059 -5426
rect 1089 -5429 1093 -5426
rect 1097 -5426 1109 -5422
rect 1123 -5422 1127 -5405
rect 1147 -5408 1151 -5361
rect 1147 -5422 1151 -5412
rect 1123 -5426 1135 -5422
rect 1097 -5429 1101 -5426
rect 1131 -5429 1135 -5426
rect 1139 -5426 1151 -5422
rect 1139 -5429 1143 -5426
rect 972 -5437 976 -5433
rect 989 -5437 993 -5433
rect 1030 -5437 1034 -5433
rect 1072 -5437 1076 -5433
rect 1114 -5437 1118 -5433
rect 1155 -5437 1159 -5433
rect 1161 -5445 1165 -5397
rect 1218 -5399 1222 -5361
rect 1218 -5429 1222 -5403
rect 1309 -5401 1313 -5215
rect 1210 -5437 1214 -5433
rect 972 -5473 976 -5469
rect 989 -5473 993 -5469
rect 1009 -5473 1013 -5469
rect 1030 -5473 1034 -5469
rect 1051 -5473 1055 -5469
rect 1072 -5473 1076 -5469
rect 1093 -5473 1097 -5469
rect 1114 -5473 1118 -5469
rect 1135 -5473 1139 -5469
rect 1155 -5473 1159 -5469
rect 1210 -5473 1214 -5469
rect 963 -5528 967 -5481
rect 963 -5549 967 -5532
rect 981 -5542 985 -5481
rect 997 -5542 1001 -5481
rect 1021 -5521 1025 -5481
rect 1021 -5542 1025 -5525
rect 1039 -5542 1043 -5481
rect 1063 -5528 1067 -5481
rect 1063 -5542 1067 -5532
rect 1081 -5521 1085 -5481
rect 1081 -5542 1085 -5525
rect 1105 -5535 1109 -5481
rect 1123 -5513 1127 -5481
rect 1123 -5521 1127 -5517
rect 1105 -5542 1109 -5539
rect 981 -5546 990 -5542
rect 997 -5546 1005 -5542
rect 981 -5549 985 -5546
rect 1005 -5549 1009 -5546
rect 1013 -5546 1025 -5542
rect 1039 -5546 1047 -5542
rect 1013 -5549 1017 -5546
rect 1047 -5549 1051 -5546
rect 1055 -5546 1067 -5542
rect 1081 -5546 1093 -5542
rect 1055 -5549 1059 -5546
rect 1089 -5549 1093 -5546
rect 1097 -5546 1109 -5542
rect 1123 -5542 1127 -5525
rect 1147 -5528 1151 -5481
rect 1147 -5542 1151 -5532
rect 1123 -5546 1135 -5542
rect 1097 -5549 1101 -5546
rect 1131 -5549 1135 -5546
rect 1139 -5546 1151 -5542
rect 1139 -5549 1143 -5546
rect 972 -5557 976 -5553
rect 989 -5557 993 -5553
rect 1030 -5557 1034 -5553
rect 1072 -5557 1076 -5553
rect 1114 -5557 1118 -5553
rect 1155 -5557 1159 -5553
rect 963 -5707 967 -5703
rect 980 -5707 984 -5703
rect 971 -5718 975 -5715
rect 971 -5722 986 -5718
rect 982 -5761 986 -5722
rect 982 -5776 986 -5765
rect 963 -5780 986 -5776
rect 989 -5752 993 -5715
rect 1161 -5731 1165 -5517
rect 1218 -5514 1222 -5481
rect 1218 -5549 1222 -5518
rect 1210 -5557 1214 -5553
rect 963 -5783 967 -5780
rect 989 -5783 993 -5756
rect 980 -5791 984 -5787
rect 972 -5826 976 -5822
rect 998 -5826 1002 -5822
rect 1015 -5826 1019 -5822
rect 1055 -5826 1059 -5822
rect 1076 -5826 1080 -5822
rect 1093 -5826 1097 -5822
rect 1133 -5826 1137 -5822
rect 1157 -5826 1161 -5822
rect 1194 -5826 1198 -5822
rect 963 -5851 967 -5834
rect 963 -5902 967 -5855
rect 981 -5844 985 -5834
rect 981 -5902 985 -5848
rect 989 -5873 993 -5834
rect 1007 -5866 1011 -5834
rect 989 -5902 993 -5877
rect 1007 -5902 1011 -5870
rect 1033 -5858 1037 -5834
rect 1033 -5895 1037 -5862
rect 1067 -5895 1071 -5834
rect 1085 -5851 1089 -5834
rect 1015 -5902 1019 -5899
rect 1023 -5899 1037 -5895
rect 1023 -5902 1027 -5899
rect 1051 -5902 1055 -5899
rect 1059 -5899 1078 -5895
rect 1059 -5902 1063 -5899
rect 1085 -5902 1089 -5855
rect 1111 -5866 1115 -5834
rect 1111 -5895 1115 -5870
rect 1145 -5888 1149 -5834
rect 1145 -5892 1162 -5888
rect 1093 -5902 1097 -5899
rect 1102 -5899 1115 -5895
rect 1102 -5902 1106 -5899
rect 1129 -5902 1133 -5899
rect 1153 -5902 1157 -5892
rect 1169 -5895 1173 -5834
rect 1177 -5888 1181 -5834
rect 1203 -5856 1207 -5834
rect 1177 -5892 1196 -5888
rect 1161 -5899 1178 -5895
rect 1161 -5902 1165 -5899
rect 1185 -5902 1189 -5892
rect 1203 -5902 1207 -5860
rect 1303 -5858 1307 -5756
rect 972 -5910 976 -5906
rect 998 -5910 1002 -5906
rect 1041 -5910 1045 -5906
rect 1076 -5910 1080 -5906
rect 1120 -5910 1124 -5906
rect 1137 -5910 1141 -5906
rect 1173 -5910 1177 -5906
rect 1194 -5910 1198 -5906
rect 1209 -5917 1213 -5870
rect 1309 -5873 1313 -5448
rect 1315 -5521 1319 -5022
rect 1340 -5048 1344 -5009
rect 1340 -5063 1344 -5052
rect 1321 -5067 1344 -5063
rect 1347 -5039 1351 -5002
rect 1519 -5018 1523 -4803
rect 1321 -5070 1325 -5067
rect 1347 -5070 1351 -5043
rect 1338 -5078 1342 -5074
rect 1330 -5113 1334 -5109
rect 1356 -5113 1360 -5109
rect 1373 -5113 1377 -5109
rect 1413 -5113 1417 -5109
rect 1434 -5113 1438 -5109
rect 1451 -5113 1455 -5109
rect 1491 -5113 1495 -5109
rect 1515 -5113 1519 -5109
rect 1552 -5113 1556 -5109
rect 1321 -5138 1325 -5121
rect 1321 -5189 1325 -5142
rect 1339 -5131 1343 -5121
rect 1339 -5189 1343 -5135
rect 1347 -5160 1351 -5121
rect 1365 -5153 1369 -5121
rect 1347 -5189 1351 -5164
rect 1365 -5189 1369 -5157
rect 1391 -5145 1395 -5121
rect 1391 -5182 1395 -5149
rect 1425 -5182 1429 -5121
rect 1443 -5138 1447 -5121
rect 1373 -5189 1377 -5186
rect 1381 -5186 1395 -5182
rect 1381 -5189 1385 -5186
rect 1409 -5189 1413 -5186
rect 1417 -5186 1436 -5182
rect 1417 -5189 1421 -5186
rect 1443 -5189 1447 -5142
rect 1469 -5153 1473 -5121
rect 1469 -5182 1473 -5157
rect 1503 -5175 1507 -5121
rect 1503 -5179 1520 -5175
rect 1451 -5189 1455 -5186
rect 1460 -5186 1473 -5182
rect 1460 -5189 1464 -5186
rect 1487 -5189 1491 -5186
rect 1511 -5189 1515 -5179
rect 1527 -5182 1531 -5121
rect 1535 -5175 1539 -5121
rect 1535 -5179 1554 -5175
rect 1519 -5186 1536 -5182
rect 1519 -5189 1523 -5186
rect 1543 -5189 1547 -5179
rect 1561 -5189 1565 -5121
rect 1330 -5197 1334 -5193
rect 1356 -5197 1360 -5193
rect 1399 -5197 1403 -5193
rect 1434 -5197 1438 -5193
rect 1478 -5197 1482 -5193
rect 1495 -5197 1499 -5193
rect 1531 -5197 1535 -5193
rect 1552 -5197 1556 -5193
rect 1561 -5211 1565 -5193
rect 1567 -5204 1571 -5157
rect 1330 -5353 1334 -5349
rect 1347 -5353 1351 -5349
rect 1367 -5353 1371 -5349
rect 1388 -5353 1392 -5349
rect 1409 -5353 1413 -5349
rect 1430 -5353 1434 -5349
rect 1451 -5353 1455 -5349
rect 1472 -5353 1476 -5349
rect 1493 -5353 1497 -5349
rect 1513 -5353 1517 -5349
rect 1321 -5408 1325 -5361
rect 1321 -5429 1325 -5412
rect 1339 -5422 1343 -5361
rect 1355 -5422 1359 -5361
rect 1379 -5401 1383 -5361
rect 1379 -5422 1383 -5405
rect 1397 -5422 1401 -5361
rect 1421 -5408 1425 -5361
rect 1421 -5422 1425 -5412
rect 1439 -5401 1443 -5361
rect 1439 -5422 1443 -5405
rect 1463 -5415 1467 -5361
rect 1481 -5393 1485 -5361
rect 1481 -5401 1485 -5397
rect 1463 -5422 1467 -5419
rect 1339 -5426 1348 -5422
rect 1355 -5426 1363 -5422
rect 1339 -5429 1343 -5426
rect 1363 -5429 1367 -5426
rect 1371 -5426 1383 -5422
rect 1397 -5426 1405 -5422
rect 1371 -5429 1375 -5426
rect 1405 -5429 1409 -5426
rect 1413 -5426 1425 -5422
rect 1439 -5426 1451 -5422
rect 1413 -5429 1417 -5426
rect 1447 -5429 1451 -5426
rect 1455 -5426 1467 -5422
rect 1481 -5422 1485 -5405
rect 1505 -5408 1509 -5361
rect 1505 -5422 1509 -5412
rect 1481 -5426 1493 -5422
rect 1455 -5429 1459 -5426
rect 1489 -5429 1493 -5426
rect 1497 -5426 1509 -5422
rect 1497 -5429 1501 -5426
rect 1330 -5437 1334 -5433
rect 1347 -5437 1351 -5433
rect 1388 -5437 1392 -5433
rect 1430 -5437 1434 -5433
rect 1472 -5437 1476 -5433
rect 1513 -5437 1517 -5433
rect 1519 -5444 1523 -5397
rect 1330 -5473 1334 -5469
rect 1347 -5473 1351 -5469
rect 1367 -5473 1371 -5469
rect 1388 -5473 1392 -5469
rect 1409 -5473 1413 -5469
rect 1430 -5473 1434 -5469
rect 1451 -5473 1455 -5469
rect 1472 -5473 1476 -5469
rect 1493 -5473 1497 -5469
rect 1513 -5473 1517 -5469
rect 1321 -5528 1325 -5481
rect 1321 -5549 1325 -5532
rect 1339 -5542 1343 -5481
rect 1355 -5542 1359 -5481
rect 1379 -5521 1383 -5481
rect 1379 -5542 1383 -5525
rect 1397 -5542 1401 -5481
rect 1421 -5528 1425 -5481
rect 1421 -5542 1425 -5532
rect 1439 -5521 1443 -5481
rect 1439 -5542 1443 -5525
rect 1463 -5535 1467 -5481
rect 1481 -5513 1485 -5481
rect 1481 -5521 1485 -5517
rect 1463 -5542 1467 -5539
rect 1339 -5546 1348 -5542
rect 1355 -5546 1363 -5542
rect 1339 -5549 1343 -5546
rect 1363 -5549 1367 -5546
rect 1371 -5546 1383 -5542
rect 1397 -5546 1405 -5542
rect 1371 -5549 1375 -5546
rect 1405 -5549 1409 -5546
rect 1413 -5546 1425 -5542
rect 1439 -5546 1451 -5542
rect 1413 -5549 1417 -5546
rect 1447 -5549 1451 -5546
rect 1455 -5546 1467 -5542
rect 1481 -5542 1485 -5525
rect 1505 -5528 1509 -5481
rect 1505 -5542 1509 -5532
rect 1481 -5546 1493 -5542
rect 1455 -5549 1459 -5546
rect 1489 -5549 1493 -5546
rect 1497 -5546 1509 -5542
rect 1497 -5549 1501 -5546
rect 1330 -5557 1334 -5553
rect 1347 -5557 1351 -5553
rect 1388 -5557 1392 -5553
rect 1430 -5557 1434 -5553
rect 1472 -5557 1476 -5553
rect 1513 -5557 1517 -5553
rect 1321 -5707 1325 -5703
rect 1338 -5707 1342 -5703
rect 1329 -5718 1333 -5715
rect 1329 -5722 1344 -5718
rect 1340 -5761 1344 -5722
rect 1340 -5776 1344 -5765
rect 1321 -5780 1344 -5776
rect 1347 -5752 1351 -5715
rect 1519 -5731 1523 -5517
rect 1321 -5783 1325 -5780
rect 1347 -5783 1351 -5756
rect 1338 -5791 1342 -5787
rect 1330 -5826 1334 -5822
rect 1356 -5826 1360 -5822
rect 1373 -5826 1377 -5822
rect 1413 -5826 1417 -5822
rect 1434 -5826 1438 -5822
rect 1451 -5826 1455 -5822
rect 1491 -5826 1495 -5822
rect 1515 -5826 1519 -5822
rect 1552 -5826 1556 -5822
rect 1321 -5851 1325 -5834
rect 1321 -5902 1325 -5855
rect 1339 -5844 1343 -5834
rect 1339 -5902 1343 -5848
rect 1347 -5873 1351 -5834
rect 1365 -5866 1369 -5834
rect 1347 -5902 1351 -5877
rect 1365 -5902 1369 -5870
rect 1391 -5858 1395 -5834
rect 1391 -5895 1395 -5862
rect 1425 -5895 1429 -5834
rect 1443 -5851 1447 -5834
rect 1373 -5902 1377 -5899
rect 1381 -5899 1395 -5895
rect 1381 -5902 1385 -5899
rect 1409 -5902 1413 -5899
rect 1417 -5899 1436 -5895
rect 1417 -5902 1421 -5899
rect 1443 -5902 1447 -5855
rect 1469 -5866 1473 -5834
rect 1469 -5895 1473 -5870
rect 1503 -5888 1507 -5834
rect 1503 -5892 1520 -5888
rect 1451 -5902 1455 -5899
rect 1460 -5899 1473 -5895
rect 1460 -5902 1464 -5899
rect 1487 -5902 1491 -5899
rect 1511 -5902 1515 -5892
rect 1527 -5895 1531 -5834
rect 1535 -5888 1539 -5834
rect 1535 -5892 1554 -5888
rect 1519 -5899 1536 -5895
rect 1519 -5902 1523 -5899
rect 1543 -5902 1547 -5892
rect 1561 -5902 1565 -5834
rect 1330 -5910 1334 -5906
rect 1356 -5910 1360 -5906
rect 1399 -5910 1403 -5906
rect 1434 -5910 1438 -5906
rect 1478 -5910 1482 -5906
rect 1495 -5910 1499 -5906
rect 1531 -5910 1535 -5906
rect 1552 -5910 1556 -5906
rect -1270 -5997 -1266 -5924
rect -1255 -5949 -1251 -5945
rect -1238 -5949 -1234 -5945
rect -1218 -5949 -1214 -5945
rect -1197 -5949 -1193 -5945
rect -1176 -5949 -1172 -5945
rect -1155 -5949 -1151 -5945
rect -1134 -5949 -1130 -5945
rect -1113 -5949 -1109 -5945
rect -1092 -5949 -1088 -5945
rect -1072 -5949 -1068 -5945
rect -1264 -6004 -1260 -5957
rect -1264 -6025 -1260 -6008
rect -1246 -6018 -1242 -5957
rect -1230 -6018 -1226 -5957
rect -1206 -5997 -1202 -5957
rect -1206 -6018 -1202 -6001
rect -1188 -6018 -1184 -5957
rect -1164 -6004 -1160 -5957
rect -1164 -6018 -1160 -6008
rect -1146 -5997 -1142 -5957
rect -1146 -6018 -1142 -6001
rect -1122 -6011 -1118 -5957
rect -1104 -5989 -1100 -5957
rect -1104 -5997 -1100 -5993
rect -1122 -6018 -1118 -6015
rect -1246 -6022 -1237 -6018
rect -1230 -6022 -1222 -6018
rect -1246 -6025 -1242 -6022
rect -1222 -6025 -1218 -6022
rect -1214 -6022 -1202 -6018
rect -1188 -6022 -1180 -6018
rect -1214 -6025 -1210 -6022
rect -1180 -6025 -1176 -6022
rect -1172 -6022 -1160 -6018
rect -1146 -6022 -1134 -6018
rect -1172 -6025 -1168 -6022
rect -1138 -6025 -1134 -6022
rect -1130 -6022 -1118 -6018
rect -1104 -6018 -1100 -6001
rect -1080 -6004 -1076 -5957
rect -941 -5997 -937 -5921
rect -926 -5949 -922 -5945
rect -909 -5949 -905 -5945
rect -889 -5949 -885 -5945
rect -868 -5949 -864 -5945
rect -847 -5949 -843 -5945
rect -826 -5949 -822 -5945
rect -805 -5949 -801 -5945
rect -784 -5949 -780 -5945
rect -763 -5949 -759 -5945
rect -743 -5949 -739 -5945
rect -1080 -6018 -1076 -6008
rect -1104 -6022 -1092 -6018
rect -1130 -6025 -1126 -6022
rect -1096 -6025 -1092 -6022
rect -1088 -6022 -1076 -6018
rect -935 -6004 -931 -5957
rect -1088 -6025 -1084 -6022
rect -935 -6025 -931 -6008
rect -917 -6018 -913 -5957
rect -901 -6018 -897 -5957
rect -877 -5997 -873 -5957
rect -877 -6018 -873 -6001
rect -859 -6018 -855 -5957
rect -835 -6004 -831 -5957
rect -835 -6018 -831 -6008
rect -817 -5997 -813 -5957
rect -817 -6018 -813 -6001
rect -793 -6011 -789 -5957
rect -775 -5989 -771 -5957
rect -775 -5997 -771 -5993
rect -793 -6018 -789 -6015
rect -917 -6022 -908 -6018
rect -901 -6022 -893 -6018
rect -917 -6025 -913 -6022
rect -893 -6025 -889 -6022
rect -885 -6022 -873 -6018
rect -859 -6022 -851 -6018
rect -885 -6025 -881 -6022
rect -851 -6025 -847 -6022
rect -843 -6022 -831 -6018
rect -817 -6022 -805 -6018
rect -843 -6025 -839 -6022
rect -809 -6025 -805 -6022
rect -801 -6022 -789 -6018
rect -775 -6018 -771 -6001
rect -751 -6004 -747 -5957
rect -583 -5997 -579 -5921
rect -568 -5949 -564 -5945
rect -551 -5949 -547 -5945
rect -531 -5949 -527 -5945
rect -510 -5949 -506 -5945
rect -489 -5949 -485 -5945
rect -468 -5949 -464 -5945
rect -447 -5949 -443 -5945
rect -426 -5949 -422 -5945
rect -405 -5949 -401 -5945
rect -385 -5949 -381 -5945
rect -751 -6018 -747 -6008
rect -775 -6022 -763 -6018
rect -801 -6025 -797 -6022
rect -767 -6025 -763 -6022
rect -759 -6022 -747 -6018
rect -577 -6004 -573 -5957
rect -759 -6025 -755 -6022
rect -577 -6025 -573 -6008
rect -559 -6018 -555 -5957
rect -543 -6018 -539 -5957
rect -519 -5997 -515 -5957
rect -519 -6018 -515 -6001
rect -501 -6018 -497 -5957
rect -477 -6004 -473 -5957
rect -477 -6018 -473 -6008
rect -459 -5997 -455 -5957
rect -459 -6018 -455 -6001
rect -435 -6011 -431 -5957
rect -417 -5989 -413 -5957
rect -417 -5997 -413 -5993
rect -435 -6018 -431 -6015
rect -559 -6022 -550 -6018
rect -543 -6022 -535 -6018
rect -559 -6025 -555 -6022
rect -535 -6025 -531 -6022
rect -527 -6022 -515 -6018
rect -501 -6022 -493 -6018
rect -527 -6025 -523 -6022
rect -493 -6025 -489 -6022
rect -485 -6022 -473 -6018
rect -459 -6022 -447 -6018
rect -485 -6025 -481 -6022
rect -451 -6025 -447 -6022
rect -443 -6022 -431 -6018
rect -417 -6018 -413 -6001
rect -393 -6004 -389 -5957
rect -225 -5997 -221 -5921
rect -210 -5949 -206 -5945
rect -193 -5949 -189 -5945
rect -173 -5949 -169 -5945
rect -152 -5949 -148 -5945
rect -131 -5949 -127 -5945
rect -110 -5949 -106 -5945
rect -89 -5949 -85 -5945
rect -68 -5949 -64 -5945
rect -47 -5949 -43 -5945
rect -27 -5949 -23 -5945
rect -393 -6018 -389 -6008
rect -417 -6022 -405 -6018
rect -443 -6025 -439 -6022
rect -409 -6025 -405 -6022
rect -401 -6022 -389 -6018
rect -219 -6004 -215 -5957
rect -401 -6025 -397 -6022
rect -219 -6025 -215 -6008
rect -201 -6018 -197 -5957
rect -185 -6018 -181 -5957
rect -161 -5997 -157 -5957
rect -161 -6018 -157 -6001
rect -143 -6018 -139 -5957
rect -119 -6004 -115 -5957
rect -119 -6018 -115 -6008
rect -101 -5997 -97 -5957
rect -101 -6018 -97 -6001
rect -77 -6011 -73 -5957
rect -59 -5989 -55 -5957
rect -59 -5997 -55 -5993
rect -77 -6018 -73 -6015
rect -201 -6022 -192 -6018
rect -185 -6022 -177 -6018
rect -201 -6025 -197 -6022
rect -177 -6025 -173 -6022
rect -169 -6022 -157 -6018
rect -143 -6022 -135 -6018
rect -169 -6025 -165 -6022
rect -135 -6025 -131 -6022
rect -127 -6022 -115 -6018
rect -101 -6022 -89 -6018
rect -127 -6025 -123 -6022
rect -93 -6025 -89 -6022
rect -85 -6022 -73 -6018
rect -59 -6018 -55 -6001
rect -35 -6004 -31 -5957
rect 203 -5997 207 -5922
rect 218 -5949 222 -5945
rect 235 -5949 239 -5945
rect 255 -5949 259 -5945
rect 276 -5949 280 -5945
rect 297 -5949 301 -5945
rect 318 -5949 322 -5945
rect 339 -5949 343 -5945
rect 360 -5949 364 -5945
rect 381 -5949 385 -5945
rect 401 -5949 405 -5945
rect -35 -6018 -31 -6008
rect -59 -6022 -47 -6018
rect -85 -6025 -81 -6022
rect -51 -6025 -47 -6022
rect -43 -6022 -31 -6018
rect 209 -6004 213 -5957
rect -43 -6025 -39 -6022
rect 209 -6025 213 -6008
rect 227 -6018 231 -5957
rect 243 -6018 247 -5957
rect 267 -5997 271 -5957
rect 267 -6018 271 -6001
rect 285 -6018 289 -5957
rect 309 -6004 313 -5957
rect 309 -6018 313 -6008
rect 327 -5997 331 -5957
rect 327 -6018 331 -6001
rect 351 -6011 355 -5957
rect 369 -5989 373 -5957
rect 369 -5997 373 -5993
rect 351 -6018 355 -6015
rect 227 -6022 236 -6018
rect 243 -6022 251 -6018
rect 227 -6025 231 -6022
rect 251 -6025 255 -6022
rect 259 -6022 271 -6018
rect 285 -6022 293 -6018
rect 259 -6025 263 -6022
rect 293 -6025 297 -6022
rect 301 -6022 313 -6018
rect 327 -6022 339 -6018
rect 301 -6025 305 -6022
rect 335 -6025 339 -6022
rect 343 -6022 355 -6018
rect 369 -6018 373 -6001
rect 393 -6004 397 -5957
rect 559 -5997 563 -5921
rect 574 -5949 578 -5945
rect 591 -5949 595 -5945
rect 611 -5949 615 -5945
rect 632 -5949 636 -5945
rect 653 -5949 657 -5945
rect 674 -5949 678 -5945
rect 695 -5949 699 -5945
rect 716 -5949 720 -5945
rect 737 -5949 741 -5945
rect 757 -5949 761 -5945
rect 393 -6018 397 -6008
rect 369 -6022 381 -6018
rect 343 -6025 347 -6022
rect 377 -6025 381 -6022
rect 385 -6022 397 -6018
rect 565 -6004 569 -5957
rect 385 -6025 389 -6022
rect 565 -6025 569 -6008
rect 583 -6018 587 -5957
rect 599 -6018 603 -5957
rect 623 -5997 627 -5957
rect 623 -6018 627 -6001
rect 641 -6018 645 -5957
rect 665 -6004 669 -5957
rect 665 -6018 669 -6008
rect 683 -5997 687 -5957
rect 683 -6018 687 -6001
rect 707 -6011 711 -5957
rect 725 -5989 729 -5957
rect 725 -5997 729 -5993
rect 707 -6018 711 -6015
rect 583 -6022 592 -6018
rect 599 -6022 607 -6018
rect 583 -6025 587 -6022
rect 607 -6025 611 -6022
rect 615 -6022 627 -6018
rect 641 -6022 649 -6018
rect 615 -6025 619 -6022
rect 649 -6025 653 -6022
rect 657 -6022 669 -6018
rect 683 -6022 695 -6018
rect 657 -6025 661 -6022
rect 691 -6025 695 -6022
rect 699 -6022 711 -6018
rect 725 -6018 729 -6001
rect 749 -6004 753 -5957
rect 957 -5997 961 -5921
rect 972 -5949 976 -5945
rect 989 -5949 993 -5945
rect 1009 -5949 1013 -5945
rect 1030 -5949 1034 -5945
rect 1051 -5949 1055 -5945
rect 1072 -5949 1076 -5945
rect 1093 -5949 1097 -5945
rect 1114 -5949 1118 -5945
rect 1135 -5949 1139 -5945
rect 1155 -5949 1159 -5945
rect 749 -6018 753 -6008
rect 725 -6022 737 -6018
rect 699 -6025 703 -6022
rect 733 -6025 737 -6022
rect 741 -6022 753 -6018
rect 963 -6004 967 -5957
rect 741 -6025 745 -6022
rect 963 -6025 967 -6008
rect 981 -6018 985 -5957
rect 997 -6018 1001 -5957
rect 1021 -5997 1025 -5957
rect 1021 -6018 1025 -6001
rect 1039 -6018 1043 -5957
rect 1063 -6004 1067 -5957
rect 1063 -6018 1067 -6008
rect 1081 -5997 1085 -5957
rect 1081 -6018 1085 -6001
rect 1105 -6011 1109 -5957
rect 1123 -5989 1127 -5957
rect 1123 -5997 1127 -5993
rect 1105 -6018 1109 -6015
rect 981 -6022 990 -6018
rect 997 -6022 1005 -6018
rect 981 -6025 985 -6022
rect 1005 -6025 1009 -6022
rect 1013 -6022 1025 -6018
rect 1039 -6022 1047 -6018
rect 1013 -6025 1017 -6022
rect 1047 -6025 1051 -6022
rect 1055 -6022 1067 -6018
rect 1081 -6022 1093 -6018
rect 1055 -6025 1059 -6022
rect 1089 -6025 1093 -6022
rect 1097 -6022 1109 -6018
rect 1123 -6018 1127 -6001
rect 1147 -6004 1151 -5957
rect 1315 -5997 1319 -5921
rect 1330 -5949 1334 -5945
rect 1347 -5949 1351 -5945
rect 1367 -5949 1371 -5945
rect 1388 -5949 1392 -5945
rect 1409 -5949 1413 -5945
rect 1430 -5949 1434 -5945
rect 1451 -5949 1455 -5945
rect 1472 -5949 1476 -5945
rect 1493 -5949 1497 -5945
rect 1513 -5949 1517 -5945
rect 1147 -6018 1151 -6008
rect 1123 -6022 1135 -6018
rect 1097 -6025 1101 -6022
rect 1131 -6025 1135 -6022
rect 1139 -6022 1151 -6018
rect 1321 -6004 1325 -5957
rect 1139 -6025 1143 -6022
rect 1321 -6025 1325 -6008
rect 1339 -6018 1343 -5957
rect 1355 -6018 1359 -5957
rect 1379 -5997 1383 -5957
rect 1379 -6018 1383 -6001
rect 1397 -6018 1401 -5957
rect 1421 -6004 1425 -5957
rect 1421 -6018 1425 -6008
rect 1439 -5997 1443 -5957
rect 1439 -6018 1443 -6001
rect 1463 -6011 1467 -5957
rect 1481 -5989 1485 -5957
rect 1481 -5997 1485 -5993
rect 1463 -6018 1467 -6015
rect 1339 -6022 1348 -6018
rect 1355 -6022 1363 -6018
rect 1339 -6025 1343 -6022
rect 1363 -6025 1367 -6022
rect 1371 -6022 1383 -6018
rect 1397 -6022 1405 -6018
rect 1371 -6025 1375 -6022
rect 1405 -6025 1409 -6022
rect 1413 -6022 1425 -6018
rect 1439 -6022 1451 -6018
rect 1413 -6025 1417 -6022
rect 1447 -6025 1451 -6022
rect 1455 -6022 1467 -6018
rect 1481 -6018 1485 -6001
rect 1505 -6004 1509 -5957
rect 1505 -6018 1509 -6008
rect 1481 -6022 1493 -6018
rect 1455 -6025 1459 -6022
rect 1489 -6025 1493 -6022
rect 1497 -6022 1509 -6018
rect 1497 -6025 1501 -6022
rect -1255 -6033 -1251 -6029
rect -1238 -6033 -1234 -6029
rect -1197 -6033 -1193 -6029
rect -1155 -6033 -1151 -6029
rect -1113 -6033 -1109 -6029
rect -1072 -6033 -1068 -6029
rect -926 -6033 -922 -6029
rect -909 -6033 -905 -6029
rect -868 -6033 -864 -6029
rect -826 -6033 -822 -6029
rect -784 -6033 -780 -6029
rect -743 -6033 -739 -6029
rect -568 -6033 -564 -6029
rect -551 -6033 -547 -6029
rect -510 -6033 -506 -6029
rect -468 -6033 -464 -6029
rect -426 -6033 -422 -6029
rect -385 -6033 -381 -6029
rect -210 -6033 -206 -6029
rect -193 -6033 -189 -6029
rect -152 -6033 -148 -6029
rect -110 -6033 -106 -6029
rect -68 -6033 -64 -6029
rect -27 -6033 -23 -6029
rect 218 -6033 222 -6029
rect 235 -6033 239 -6029
rect 276 -6033 280 -6029
rect 318 -6033 322 -6029
rect 360 -6033 364 -6029
rect 401 -6033 405 -6029
rect 574 -6033 578 -6029
rect 591 -6033 595 -6029
rect 632 -6033 636 -6029
rect 674 -6033 678 -6029
rect 716 -6033 720 -6029
rect 757 -6033 761 -6029
rect 972 -6033 976 -6029
rect 989 -6033 993 -6029
rect 1030 -6033 1034 -6029
rect 1072 -6033 1076 -6029
rect 1114 -6033 1118 -6029
rect 1155 -6033 1159 -6029
rect 1330 -6033 1334 -6029
rect 1347 -6033 1351 -6029
rect 1388 -6033 1392 -6029
rect 1430 -6033 1434 -6029
rect 1472 -6033 1476 -6029
rect 1513 -6033 1517 -6029
rect 1561 -6040 1565 -5906
rect 1567 -5917 1571 -5870
rect 1315 -6115 1319 -6044
rect 1330 -6067 1334 -6063
rect 1347 -6067 1351 -6063
rect 1367 -6067 1371 -6063
rect 1388 -6067 1392 -6063
rect 1409 -6067 1413 -6063
rect 1430 -6067 1434 -6063
rect 1451 -6067 1455 -6063
rect 1472 -6067 1476 -6063
rect 1493 -6067 1497 -6063
rect 1513 -6067 1517 -6063
rect 1321 -6122 1325 -6075
rect 1321 -6143 1325 -6126
rect 1339 -6136 1343 -6075
rect 1355 -6136 1359 -6075
rect 1379 -6115 1383 -6075
rect 1379 -6136 1383 -6119
rect 1397 -6136 1401 -6075
rect 1421 -6122 1425 -6075
rect 1421 -6136 1425 -6126
rect 1439 -6115 1443 -6075
rect 1439 -6136 1443 -6119
rect 1463 -6129 1467 -6075
rect 1481 -6107 1485 -6075
rect 1481 -6115 1485 -6111
rect 1463 -6136 1467 -6133
rect 1339 -6140 1348 -6136
rect 1355 -6140 1363 -6136
rect 1339 -6143 1343 -6140
rect 1363 -6143 1367 -6140
rect 1371 -6140 1383 -6136
rect 1397 -6140 1405 -6136
rect 1371 -6143 1375 -6140
rect 1405 -6143 1409 -6140
rect 1413 -6140 1425 -6136
rect 1439 -6140 1451 -6136
rect 1413 -6143 1417 -6140
rect 1447 -6143 1451 -6140
rect 1455 -6140 1467 -6136
rect 1481 -6136 1485 -6119
rect 1505 -6122 1509 -6075
rect 1505 -6136 1509 -6126
rect 1481 -6140 1493 -6136
rect 1455 -6143 1459 -6140
rect 1489 -6143 1493 -6140
rect 1497 -6140 1509 -6136
rect 1497 -6143 1501 -6140
rect 1330 -6151 1334 -6147
rect 1347 -6151 1351 -6147
rect 1388 -6151 1392 -6147
rect 1430 -6151 1434 -6147
rect 1472 -6151 1476 -6147
rect 1513 -6151 1517 -6147
<< metal2 >>
rect -1495 -1034 -1337 -1030
rect -1333 -1034 -1320 -1030
rect -1316 -1034 -936 -1030
rect -932 -1034 -919 -1030
rect -915 -1034 -577 -1030
rect -573 -1034 -560 -1030
rect -556 -1034 -219 -1030
rect -215 -1034 -202 -1030
rect -198 -1034 209 -1030
rect 213 -1034 226 -1030
rect 230 -1034 565 -1030
rect 569 -1034 582 -1030
rect 586 -1034 963 -1030
rect 967 -1034 980 -1030
rect 984 -1034 1321 -1030
rect 1325 -1034 1338 -1030
rect 1342 -1034 1617 -1030
rect -1495 -1144 -1433 -1034
rect -1421 -1074 -1325 -1070
rect -1321 -1074 -924 -1070
rect -920 -1074 -565 -1070
rect -561 -1074 -207 -1070
rect -203 -1074 221 -1070
rect 225 -1074 577 -1070
rect 581 -1074 975 -1070
rect 979 -1074 1333 -1070
rect 1337 -1074 1617 -1070
rect -944 -1082 -551 -1078
rect -227 -1082 235 -1078
rect 557 -1082 989 -1078
rect -1262 -1090 -910 -1086
rect -585 -1090 -193 -1086
rect 201 -1090 591 -1086
rect 955 -1090 1347 -1086
rect 1633 -1122 1695 -1030
rect -1421 -1126 -1320 -1122
rect -1316 -1126 -919 -1122
rect -915 -1126 -560 -1122
rect -556 -1126 -202 -1122
rect -198 -1126 226 -1122
rect 230 -1126 582 -1122
rect 586 -1126 980 -1122
rect 984 -1126 1338 -1122
rect 1342 -1126 1695 -1122
rect -1495 -1148 -1251 -1144
rect -1247 -1148 -1234 -1144
rect -1230 -1148 -1214 -1144
rect -1210 -1148 -1193 -1144
rect -1189 -1148 -1172 -1144
rect -1168 -1148 -1151 -1144
rect -1147 -1148 -1130 -1144
rect -1126 -1148 -1109 -1144
rect -1105 -1148 -1088 -1144
rect -1084 -1148 -1068 -1144
rect -1064 -1148 -926 -1144
rect -922 -1148 -909 -1144
rect -905 -1148 -889 -1144
rect -885 -1148 -868 -1144
rect -864 -1148 -847 -1144
rect -843 -1148 -826 -1144
rect -822 -1148 -805 -1144
rect -801 -1148 -784 -1144
rect -780 -1148 -763 -1144
rect -759 -1148 -743 -1144
rect -739 -1148 -568 -1144
rect -564 -1148 -551 -1144
rect -547 -1148 -531 -1144
rect -527 -1148 -510 -1144
rect -506 -1148 -489 -1144
rect -485 -1148 -468 -1144
rect -464 -1148 -447 -1144
rect -443 -1148 -426 -1144
rect -422 -1148 -405 -1144
rect -401 -1148 -385 -1144
rect -381 -1148 -210 -1144
rect -206 -1148 -193 -1144
rect -189 -1148 -173 -1144
rect -169 -1148 -152 -1144
rect -148 -1148 -131 -1144
rect -127 -1148 -110 -1144
rect -106 -1148 -89 -1144
rect -85 -1148 -68 -1144
rect -64 -1148 -47 -1144
rect -43 -1148 -27 -1144
rect -23 -1148 218 -1144
rect 222 -1148 235 -1144
rect 239 -1148 255 -1144
rect 259 -1148 276 -1144
rect 280 -1148 297 -1144
rect 301 -1148 318 -1144
rect 322 -1148 339 -1144
rect 343 -1148 360 -1144
rect 364 -1148 381 -1144
rect 385 -1148 401 -1144
rect 405 -1148 574 -1144
rect 578 -1148 591 -1144
rect 595 -1148 611 -1144
rect 615 -1148 632 -1144
rect 636 -1148 653 -1144
rect 657 -1148 674 -1144
rect 678 -1148 695 -1144
rect 699 -1148 716 -1144
rect 720 -1148 737 -1144
rect 741 -1148 757 -1144
rect 761 -1148 972 -1144
rect 976 -1148 989 -1144
rect 993 -1148 1009 -1144
rect 1013 -1148 1030 -1144
rect 1034 -1148 1051 -1144
rect 1055 -1148 1072 -1144
rect 1076 -1148 1093 -1144
rect 1097 -1148 1114 -1144
rect 1118 -1148 1135 -1144
rect 1139 -1148 1155 -1144
rect 1159 -1148 1617 -1144
rect -1495 -1260 -1433 -1148
rect -1229 -1196 -1195 -1192
rect -1131 -1196 -1111 -1192
rect -1096 -1196 -931 -1192
rect -904 -1196 -870 -1192
rect -806 -1196 -786 -1192
rect -771 -1196 -573 -1192
rect -546 -1196 -512 -1192
rect -448 -1196 -428 -1192
rect -413 -1196 -215 -1192
rect -188 -1196 -154 -1192
rect -90 -1196 -70 -1192
rect -55 -1196 213 -1192
rect 240 -1196 274 -1192
rect 338 -1196 358 -1192
rect 373 -1196 569 -1192
rect 596 -1196 630 -1192
rect 694 -1196 714 -1192
rect 729 -1196 967 -1192
rect 994 -1196 1028 -1192
rect 1092 -1196 1112 -1192
rect 1127 -1196 1163 -1192
rect -935 -1200 -931 -1196
rect -577 -1200 -573 -1196
rect -219 -1200 -215 -1196
rect 209 -1200 213 -1196
rect 565 -1200 569 -1196
rect 963 -1200 967 -1196
rect -1307 -1204 -1253 -1200
rect -1249 -1204 -1219 -1200
rect -1198 -1204 -1167 -1200
rect -1138 -1204 -1107 -1200
rect -1096 -1204 -1069 -1200
rect -935 -1204 -928 -1200
rect -924 -1204 -894 -1200
rect -873 -1204 -842 -1200
rect -813 -1204 -782 -1200
rect -771 -1204 -744 -1200
rect -577 -1204 -570 -1200
rect -566 -1204 -536 -1200
rect -515 -1204 -484 -1200
rect -455 -1204 -424 -1200
rect -413 -1204 -386 -1200
rect -219 -1204 -212 -1200
rect -208 -1204 -178 -1200
rect -157 -1204 -126 -1200
rect -97 -1204 -66 -1200
rect -55 -1204 -28 -1200
rect 209 -1204 216 -1200
rect 220 -1204 250 -1200
rect 271 -1204 302 -1200
rect 331 -1204 362 -1200
rect 373 -1204 400 -1200
rect 565 -1204 572 -1200
rect 576 -1204 606 -1200
rect 627 -1204 658 -1200
rect 687 -1204 718 -1200
rect 729 -1204 756 -1200
rect 963 -1204 970 -1200
rect 974 -1204 1004 -1200
rect 1025 -1204 1056 -1200
rect 1085 -1204 1116 -1200
rect 1127 -1204 1154 -1200
rect -1256 -1211 -1209 -1207
rect -1173 -1211 -1160 -1207
rect -1156 -1211 -1125 -1207
rect -1089 -1211 -1076 -1207
rect -1072 -1211 -1060 -1207
rect -931 -1211 -884 -1207
rect -848 -1211 -835 -1207
rect -831 -1211 -800 -1207
rect -764 -1211 -751 -1207
rect -747 -1211 -735 -1207
rect -573 -1211 -526 -1207
rect -490 -1211 -477 -1207
rect -473 -1211 -442 -1207
rect -406 -1211 -393 -1207
rect -389 -1211 -377 -1207
rect -215 -1211 -168 -1207
rect -132 -1211 -119 -1207
rect -115 -1211 -84 -1207
rect -48 -1211 -35 -1207
rect -31 -1211 -19 -1207
rect 213 -1211 260 -1207
rect 296 -1211 309 -1207
rect 313 -1211 344 -1207
rect 380 -1211 393 -1207
rect 397 -1211 409 -1207
rect 569 -1211 616 -1207
rect 652 -1211 665 -1207
rect 669 -1211 700 -1207
rect 736 -1211 749 -1207
rect 753 -1211 765 -1207
rect 967 -1211 1014 -1207
rect 1050 -1211 1063 -1207
rect 1067 -1211 1098 -1207
rect 1134 -1211 1147 -1207
rect 1151 -1211 1163 -1207
rect -1270 -1218 -1249 -1214
rect -1245 -1218 -1135 -1214
rect -1114 -1218 -1083 -1214
rect -952 -1218 -924 -1214
rect -920 -1218 -810 -1214
rect -789 -1218 -758 -1214
rect -583 -1218 -566 -1214
rect -562 -1218 -452 -1214
rect -431 -1218 -400 -1214
rect -236 -1218 -208 -1214
rect -204 -1218 -94 -1214
rect -73 -1218 -42 -1214
rect 202 -1218 220 -1214
rect 224 -1218 334 -1214
rect 355 -1218 386 -1214
rect 540 -1218 576 -1214
rect 580 -1218 690 -1214
rect 711 -1218 742 -1214
rect 956 -1218 974 -1214
rect 978 -1218 1088 -1214
rect 1109 -1218 1140 -1214
rect -1214 -1225 -1191 -1221
rect -1172 -1225 -1153 -1221
rect -889 -1225 -866 -1221
rect -847 -1225 -828 -1221
rect -531 -1225 -508 -1221
rect -489 -1225 -470 -1221
rect -173 -1225 -150 -1221
rect -131 -1225 -112 -1221
rect 255 -1225 278 -1221
rect 297 -1225 316 -1221
rect 611 -1225 634 -1221
rect 653 -1225 672 -1221
rect 1009 -1225 1032 -1221
rect 1051 -1225 1070 -1221
rect 1633 -1236 1695 -1126
rect -1421 -1240 -1251 -1236
rect -1247 -1240 -1234 -1236
rect -1230 -1240 -1193 -1236
rect -1189 -1240 -1151 -1236
rect -1147 -1240 -1109 -1236
rect -1105 -1240 -1068 -1236
rect -1064 -1240 -926 -1236
rect -922 -1240 -909 -1236
rect -905 -1240 -868 -1236
rect -864 -1240 -826 -1236
rect -822 -1240 -784 -1236
rect -780 -1240 -743 -1236
rect -739 -1240 -568 -1236
rect -564 -1240 -551 -1236
rect -547 -1240 -510 -1236
rect -506 -1240 -468 -1236
rect -464 -1240 -426 -1236
rect -422 -1240 -385 -1236
rect -381 -1240 -210 -1236
rect -206 -1240 -193 -1236
rect -189 -1240 -152 -1236
rect -148 -1240 -110 -1236
rect -106 -1240 -68 -1236
rect -64 -1240 -27 -1236
rect -23 -1240 218 -1236
rect 222 -1240 235 -1236
rect 239 -1240 276 -1236
rect 280 -1240 318 -1236
rect 322 -1240 360 -1236
rect 364 -1240 401 -1236
rect 405 -1240 574 -1236
rect 578 -1240 591 -1236
rect 595 -1240 632 -1236
rect 636 -1240 674 -1236
rect 678 -1240 716 -1236
rect 720 -1240 757 -1236
rect 761 -1240 972 -1236
rect 976 -1240 989 -1236
rect 993 -1240 1030 -1236
rect 1034 -1240 1072 -1236
rect 1076 -1240 1114 -1236
rect 1118 -1240 1155 -1236
rect 1159 -1240 1695 -1236
rect -1495 -1264 -1339 -1260
rect -1335 -1264 -1322 -1260
rect -1318 -1264 -935 -1260
rect -931 -1264 -918 -1260
rect -914 -1264 -577 -1260
rect -573 -1264 -560 -1260
rect -556 -1264 -219 -1260
rect -215 -1264 -202 -1260
rect -198 -1264 209 -1260
rect 213 -1264 226 -1260
rect 230 -1264 565 -1260
rect 569 -1264 582 -1260
rect 586 -1264 963 -1260
rect 967 -1264 980 -1260
rect 984 -1264 1321 -1260
rect 1325 -1264 1338 -1260
rect 1342 -1264 1617 -1260
rect -1495 -1374 -1433 -1264
rect -1421 -1304 -1327 -1300
rect -1323 -1304 -923 -1300
rect -919 -1304 -565 -1300
rect -561 -1304 -207 -1300
rect -203 -1304 221 -1300
rect 225 -1304 577 -1300
rect 581 -1304 975 -1300
rect 979 -1304 1333 -1300
rect 1337 -1304 1617 -1300
rect -950 -1317 -909 -1313
rect -591 -1317 -551 -1313
rect -233 -1317 -193 -1313
rect 195 -1317 235 -1313
rect 551 -1317 591 -1313
rect 949 -1317 989 -1313
rect 1313 -1317 1347 -1313
rect 1633 -1352 1695 -1240
rect -1421 -1356 -1322 -1352
rect -1318 -1356 -918 -1352
rect -914 -1356 -560 -1352
rect -556 -1356 -202 -1352
rect -198 -1356 226 -1352
rect 230 -1356 582 -1352
rect 586 -1356 980 -1352
rect 984 -1356 1338 -1352
rect 1342 -1356 1695 -1352
rect -1495 -1378 -1251 -1374
rect -1247 -1378 -1234 -1374
rect -1230 -1378 -1194 -1374
rect -1190 -1378 -1173 -1374
rect -1169 -1378 -926 -1374
rect -922 -1378 -900 -1374
rect -896 -1378 -883 -1374
rect -879 -1378 -843 -1374
rect -839 -1378 -822 -1374
rect -818 -1378 -805 -1374
rect -801 -1378 -765 -1374
rect -761 -1378 -741 -1374
rect -737 -1378 -704 -1374
rect -700 -1378 -568 -1374
rect -564 -1378 -542 -1374
rect -538 -1378 -525 -1374
rect -521 -1378 -485 -1374
rect -481 -1378 -464 -1374
rect -460 -1378 -447 -1374
rect -443 -1378 -407 -1374
rect -403 -1378 -383 -1374
rect -379 -1378 -346 -1374
rect -342 -1378 -210 -1374
rect -206 -1378 -184 -1374
rect -180 -1378 -167 -1374
rect -163 -1378 -127 -1374
rect -123 -1378 -106 -1374
rect -102 -1378 -89 -1374
rect -85 -1378 -49 -1374
rect -45 -1378 -25 -1374
rect -21 -1378 12 -1374
rect 16 -1378 218 -1374
rect 222 -1378 244 -1374
rect 248 -1378 261 -1374
rect 265 -1378 301 -1374
rect 305 -1378 322 -1374
rect 326 -1378 339 -1374
rect 343 -1378 379 -1374
rect 383 -1378 403 -1374
rect 407 -1378 440 -1374
rect 444 -1378 574 -1374
rect 578 -1378 600 -1374
rect 604 -1378 617 -1374
rect 621 -1378 657 -1374
rect 661 -1378 678 -1374
rect 682 -1378 695 -1374
rect 699 -1378 735 -1374
rect 739 -1378 759 -1374
rect 763 -1378 796 -1374
rect 800 -1378 972 -1374
rect 976 -1378 998 -1374
rect 1002 -1378 1015 -1374
rect 1019 -1378 1055 -1374
rect 1059 -1378 1076 -1374
rect 1080 -1378 1093 -1374
rect 1097 -1378 1133 -1374
rect 1137 -1378 1157 -1374
rect 1161 -1378 1194 -1374
rect 1198 -1378 1330 -1374
rect 1334 -1378 1347 -1374
rect 1351 -1378 1387 -1374
rect 1391 -1378 1408 -1374
rect 1412 -1378 1617 -1374
rect -1495 -1497 -1433 -1378
rect -210 -1382 -206 -1378
rect -184 -1382 -180 -1378
rect -167 -1382 -163 -1378
rect -127 -1382 -123 -1378
rect -106 -1382 -102 -1378
rect -89 -1382 -85 -1378
rect -49 -1382 -45 -1378
rect -25 -1382 -21 -1378
rect 12 -1382 16 -1378
rect 218 -1382 222 -1378
rect 244 -1382 248 -1378
rect 261 -1382 265 -1378
rect 301 -1382 305 -1378
rect 322 -1382 326 -1378
rect 339 -1382 343 -1378
rect 379 -1382 383 -1378
rect 403 -1382 407 -1378
rect 440 -1382 444 -1378
rect 574 -1382 578 -1378
rect 600 -1382 604 -1378
rect 617 -1382 621 -1378
rect 657 -1382 661 -1378
rect 678 -1382 682 -1378
rect 695 -1382 699 -1378
rect 735 -1382 739 -1378
rect 759 -1382 763 -1378
rect 796 -1382 800 -1378
rect 972 -1382 976 -1378
rect 998 -1382 1002 -1378
rect 1015 -1382 1019 -1378
rect 1055 -1382 1059 -1378
rect 1076 -1382 1080 -1378
rect 1093 -1382 1097 -1378
rect 1133 -1382 1137 -1378
rect 1157 -1382 1161 -1378
rect 1194 -1382 1198 -1378
rect -920 -1397 -858 -1393
rect -854 -1397 -824 -1393
rect -776 -1397 -746 -1393
rect -562 -1397 -500 -1393
rect -496 -1397 -466 -1393
rect -418 -1397 -388 -1393
rect -204 -1397 -142 -1393
rect -138 -1397 -108 -1393
rect -60 -1397 -30 -1393
rect 224 -1397 286 -1393
rect 290 -1397 320 -1393
rect 368 -1397 398 -1393
rect 580 -1397 642 -1393
rect 646 -1397 676 -1393
rect 724 -1397 754 -1393
rect 978 -1397 1040 -1393
rect 1044 -1397 1074 -1393
rect 1122 -1397 1152 -1393
rect -913 -1404 -882 -1400
rect -555 -1404 -524 -1400
rect -197 -1404 -166 -1400
rect 231 -1404 262 -1400
rect 587 -1404 618 -1400
rect 985 -1404 1016 -1400
rect -931 -1411 -848 -1407
rect -809 -1411 -706 -1407
rect -573 -1411 -490 -1407
rect -451 -1411 -348 -1407
rect -215 -1411 -132 -1407
rect -93 -1411 10 -1407
rect 213 -1411 296 -1407
rect 335 -1411 438 -1407
rect 569 -1411 652 -1407
rect 691 -1411 794 -1407
rect 967 -1411 1050 -1407
rect 1089 -1411 1192 -1407
rect -944 -1418 -928 -1414
rect -894 -1418 -865 -1414
rect -861 -1418 -780 -1414
rect -691 -1418 -592 -1414
rect -585 -1418 -570 -1414
rect -536 -1418 -507 -1414
rect -503 -1418 -422 -1414
rect -333 -1418 -234 -1414
rect -227 -1418 -212 -1414
rect -178 -1418 -149 -1414
rect -145 -1418 -64 -1414
rect 25 -1418 194 -1414
rect 201 -1418 216 -1414
rect 250 -1418 279 -1414
rect 283 -1418 364 -1414
rect 453 -1418 550 -1414
rect 557 -1418 572 -1414
rect 606 -1418 635 -1414
rect 639 -1418 720 -1414
rect 809 -1418 948 -1414
rect 955 -1418 970 -1414
rect 1004 -1418 1033 -1414
rect 1037 -1418 1118 -1414
rect -596 -1422 -592 -1418
rect -238 -1422 -234 -1418
rect 190 -1422 194 -1418
rect 546 -1422 550 -1418
rect 944 -1422 948 -1418
rect -1256 -1427 -1199 -1423
rect -1160 -1426 -902 -1422
rect -887 -1426 -804 -1422
rect -783 -1426 -689 -1422
rect -596 -1426 -544 -1422
rect -529 -1426 -446 -1422
rect -425 -1426 -331 -1422
rect -238 -1426 -186 -1422
rect -171 -1426 -88 -1422
rect -67 -1426 27 -1422
rect 190 -1426 242 -1422
rect 257 -1426 340 -1422
rect 361 -1426 455 -1422
rect 546 -1426 598 -1422
rect 613 -1426 696 -1422
rect 717 -1426 811 -1422
rect 944 -1426 996 -1422
rect 1011 -1426 1094 -1422
rect 1115 -1426 1209 -1422
rect 1325 -1427 1382 -1423
rect -1262 -1434 -1249 -1430
rect -1245 -1434 -1209 -1430
rect -1205 -1434 -1189 -1430
rect -950 -1433 -924 -1429
rect -905 -1433 -776 -1429
rect -591 -1433 -566 -1429
rect -547 -1433 -418 -1429
rect -233 -1433 -208 -1429
rect -189 -1433 -60 -1429
rect 195 -1433 220 -1429
rect 239 -1433 368 -1429
rect 551 -1433 576 -1429
rect 595 -1433 724 -1429
rect 949 -1433 974 -1429
rect 993 -1433 1122 -1429
rect 1207 -1434 1332 -1430
rect 1336 -1434 1372 -1430
rect 1376 -1434 1392 -1430
rect -1309 -1441 -1253 -1437
rect -1249 -1441 -1223 -1437
rect -1219 -1441 -1175 -1437
rect -898 -1440 -794 -1436
rect -790 -1440 -760 -1436
rect -540 -1440 -436 -1436
rect -432 -1440 -402 -1436
rect -182 -1440 -78 -1436
rect -74 -1440 -44 -1436
rect 246 -1440 350 -1436
rect 354 -1440 384 -1436
rect 602 -1440 706 -1436
rect 710 -1440 740 -1436
rect 1000 -1440 1104 -1436
rect 1108 -1440 1138 -1436
rect 1313 -1441 1328 -1437
rect 1332 -1441 1358 -1437
rect 1362 -1441 1406 -1437
rect -1212 -1448 -1158 -1444
rect -924 -1447 -872 -1443
rect -868 -1447 -838 -1443
rect -566 -1447 -514 -1443
rect -510 -1447 -480 -1443
rect -208 -1447 -156 -1443
rect -152 -1447 -122 -1443
rect 220 -1447 272 -1443
rect 276 -1447 306 -1443
rect 576 -1447 628 -1443
rect 632 -1447 662 -1443
rect 974 -1447 1026 -1443
rect 1030 -1447 1060 -1443
rect 1369 -1448 1423 -1444
rect -1230 -1455 -1198 -1451
rect -879 -1455 -847 -1451
rect -801 -1455 -769 -1451
rect -521 -1455 -489 -1451
rect -443 -1455 -411 -1451
rect -163 -1455 -131 -1451
rect -167 -1458 -163 -1455
rect -131 -1458 -127 -1455
rect -85 -1455 -53 -1451
rect -89 -1458 -85 -1455
rect -53 -1458 -49 -1455
rect 265 -1455 297 -1451
rect 261 -1458 265 -1455
rect 297 -1458 301 -1455
rect 343 -1455 375 -1451
rect 339 -1458 343 -1455
rect 375 -1458 379 -1455
rect 621 -1455 653 -1451
rect 617 -1458 621 -1455
rect 653 -1458 657 -1455
rect 699 -1455 731 -1451
rect 695 -1458 699 -1455
rect 731 -1458 735 -1455
rect 1019 -1455 1051 -1451
rect 1015 -1458 1019 -1455
rect 1051 -1458 1055 -1455
rect 1097 -1455 1129 -1451
rect 1351 -1455 1383 -1451
rect 1093 -1458 1097 -1455
rect 1129 -1458 1133 -1455
rect -210 -1466 -206 -1462
rect -184 -1466 -180 -1462
rect -141 -1466 -137 -1462
rect -106 -1466 -102 -1462
rect -62 -1466 -58 -1462
rect -45 -1466 -41 -1462
rect -9 -1466 -5 -1462
rect 12 -1466 16 -1462
rect 218 -1466 222 -1462
rect 244 -1466 248 -1462
rect 287 -1466 291 -1462
rect 322 -1466 326 -1462
rect 366 -1466 370 -1462
rect 383 -1466 387 -1462
rect 419 -1466 423 -1462
rect 440 -1466 444 -1462
rect 574 -1466 578 -1462
rect 600 -1466 604 -1462
rect 643 -1466 647 -1462
rect 678 -1466 682 -1462
rect 722 -1466 726 -1462
rect 739 -1466 743 -1462
rect 775 -1466 779 -1462
rect 796 -1466 800 -1462
rect 972 -1466 976 -1462
rect 998 -1466 1002 -1462
rect 1041 -1466 1045 -1462
rect 1076 -1466 1080 -1462
rect 1120 -1466 1124 -1462
rect 1137 -1466 1141 -1462
rect 1173 -1466 1177 -1462
rect 1194 -1466 1198 -1462
rect 1633 -1466 1695 -1356
rect -1421 -1470 -1251 -1466
rect -1247 -1470 -1207 -1466
rect -1203 -1470 -1173 -1466
rect -1169 -1470 -926 -1466
rect -922 -1470 -900 -1466
rect -896 -1470 -857 -1466
rect -853 -1470 -822 -1466
rect -818 -1470 -778 -1466
rect -774 -1470 -761 -1466
rect -757 -1470 -725 -1466
rect -721 -1470 -704 -1466
rect -700 -1470 -568 -1466
rect -564 -1470 -542 -1466
rect -538 -1470 -499 -1466
rect -495 -1470 -464 -1466
rect -460 -1470 -420 -1466
rect -416 -1470 -403 -1466
rect -399 -1470 -367 -1466
rect -363 -1470 -346 -1466
rect -342 -1470 -210 -1466
rect -206 -1470 -184 -1466
rect -180 -1470 -141 -1466
rect -137 -1470 -106 -1466
rect -102 -1470 -62 -1466
rect -58 -1470 -45 -1466
rect -41 -1470 -9 -1466
rect -5 -1470 12 -1466
rect 16 -1470 218 -1466
rect 222 -1470 244 -1466
rect 248 -1470 287 -1466
rect 291 -1470 322 -1466
rect 326 -1470 366 -1466
rect 370 -1470 383 -1466
rect 387 -1470 419 -1466
rect 423 -1470 440 -1466
rect 444 -1470 574 -1466
rect 578 -1470 600 -1466
rect 604 -1470 643 -1466
rect 647 -1470 678 -1466
rect 682 -1470 722 -1466
rect 726 -1470 739 -1466
rect 743 -1470 775 -1466
rect 779 -1470 796 -1466
rect 800 -1470 972 -1466
rect 976 -1470 998 -1466
rect 1002 -1470 1041 -1466
rect 1045 -1470 1076 -1466
rect 1080 -1470 1120 -1466
rect 1124 -1470 1137 -1466
rect 1141 -1470 1173 -1466
rect 1177 -1470 1194 -1466
rect 1198 -1470 1330 -1466
rect 1334 -1470 1374 -1466
rect 1378 -1470 1408 -1466
rect 1412 -1470 1695 -1466
rect -1268 -1477 -689 -1473
rect -1262 -1484 -1158 -1480
rect -944 -1484 -331 -1480
rect -227 -1484 455 -1480
rect 557 -1484 1209 -1480
rect 1313 -1484 1417 -1480
rect -585 -1491 27 -1487
rect 201 -1491 811 -1487
rect 955 -1491 1423 -1487
rect -1495 -1501 -1251 -1497
rect -1247 -1501 -1234 -1497
rect -1230 -1501 -1214 -1497
rect -1210 -1501 -1193 -1497
rect -1189 -1501 -1172 -1497
rect -1168 -1501 -1151 -1497
rect -1147 -1501 -1130 -1497
rect -1126 -1501 -1109 -1497
rect -1105 -1501 -1088 -1497
rect -1084 -1501 -1068 -1497
rect -1064 -1501 -926 -1497
rect -922 -1501 -909 -1497
rect -905 -1501 -889 -1497
rect -885 -1501 -868 -1497
rect -864 -1501 -847 -1497
rect -843 -1501 -826 -1497
rect -822 -1501 -805 -1497
rect -801 -1501 -784 -1497
rect -780 -1501 -763 -1497
rect -759 -1501 -743 -1497
rect -739 -1501 -568 -1497
rect -564 -1501 -551 -1497
rect -547 -1501 -531 -1497
rect -527 -1501 -510 -1497
rect -506 -1501 -489 -1497
rect -485 -1501 -468 -1497
rect -464 -1501 -447 -1497
rect -443 -1501 -426 -1497
rect -422 -1501 -405 -1497
rect -401 -1501 -385 -1497
rect -381 -1501 -210 -1497
rect -206 -1501 -193 -1497
rect -189 -1501 -173 -1497
rect -169 -1501 -152 -1497
rect -148 -1501 -131 -1497
rect -127 -1501 -110 -1497
rect -106 -1501 -89 -1497
rect -85 -1501 -68 -1497
rect -64 -1501 -47 -1497
rect -43 -1501 -27 -1497
rect -23 -1501 218 -1497
rect 222 -1501 235 -1497
rect 239 -1501 255 -1497
rect 259 -1501 276 -1497
rect 280 -1501 297 -1497
rect 301 -1501 318 -1497
rect 322 -1501 339 -1497
rect 343 -1501 360 -1497
rect 364 -1501 381 -1497
rect 385 -1501 401 -1497
rect 405 -1501 574 -1497
rect 578 -1501 591 -1497
rect 595 -1501 611 -1497
rect 615 -1501 632 -1497
rect 636 -1501 653 -1497
rect 657 -1501 674 -1497
rect 678 -1501 695 -1497
rect 699 -1501 716 -1497
rect 720 -1501 737 -1497
rect 741 -1501 757 -1497
rect 761 -1501 972 -1497
rect 976 -1501 989 -1497
rect 993 -1501 1009 -1497
rect 1013 -1501 1030 -1497
rect 1034 -1501 1051 -1497
rect 1055 -1501 1072 -1497
rect 1076 -1501 1093 -1497
rect 1097 -1501 1114 -1497
rect 1118 -1501 1135 -1497
rect 1139 -1501 1155 -1497
rect 1159 -1501 1617 -1497
rect -1495 -1618 -1433 -1501
rect -1229 -1549 -1195 -1545
rect -1131 -1549 -1111 -1545
rect -1096 -1549 -931 -1545
rect -904 -1549 -870 -1545
rect -806 -1549 -786 -1545
rect -771 -1549 -573 -1545
rect -546 -1549 -512 -1545
rect -448 -1549 -428 -1545
rect -413 -1549 -215 -1545
rect -188 -1549 -154 -1545
rect -90 -1549 -70 -1545
rect -55 -1549 213 -1545
rect 240 -1549 274 -1545
rect 338 -1549 358 -1545
rect 373 -1549 569 -1545
rect 596 -1549 630 -1545
rect 694 -1549 714 -1545
rect 729 -1549 967 -1545
rect 994 -1549 1028 -1545
rect 1092 -1549 1112 -1545
rect 1127 -1549 1163 -1545
rect -935 -1553 -931 -1549
rect -577 -1553 -573 -1549
rect -219 -1553 -215 -1549
rect 209 -1553 213 -1549
rect 565 -1553 569 -1549
rect 963 -1553 967 -1549
rect -1262 -1557 -1253 -1553
rect -1249 -1557 -1219 -1553
rect -1198 -1557 -1167 -1553
rect -1138 -1557 -1107 -1553
rect -1096 -1557 -1069 -1553
rect -935 -1557 -928 -1553
rect -924 -1557 -894 -1553
rect -873 -1557 -842 -1553
rect -813 -1557 -782 -1553
rect -771 -1557 -744 -1553
rect -577 -1557 -570 -1553
rect -566 -1557 -536 -1553
rect -515 -1557 -484 -1553
rect -455 -1557 -424 -1553
rect -413 -1557 -386 -1553
rect -219 -1557 -212 -1553
rect -208 -1557 -178 -1553
rect -157 -1557 -126 -1553
rect -97 -1557 -66 -1553
rect -55 -1557 -28 -1553
rect 209 -1557 216 -1553
rect 220 -1557 250 -1553
rect 271 -1557 302 -1553
rect 331 -1557 362 -1553
rect 373 -1557 400 -1553
rect 565 -1557 572 -1553
rect 576 -1557 606 -1553
rect 627 -1557 658 -1553
rect 687 -1557 718 -1553
rect 729 -1557 756 -1553
rect 963 -1557 970 -1553
rect 974 -1557 1004 -1553
rect 1025 -1557 1056 -1553
rect 1085 -1557 1116 -1553
rect 1127 -1557 1154 -1553
rect -1256 -1564 -1209 -1560
rect -1173 -1564 -1160 -1560
rect -1156 -1564 -1125 -1560
rect -1089 -1564 -1076 -1560
rect -1072 -1564 -1060 -1560
rect -931 -1564 -884 -1560
rect -848 -1564 -835 -1560
rect -831 -1564 -800 -1560
rect -764 -1564 -751 -1560
rect -747 -1564 -735 -1560
rect -573 -1564 -526 -1560
rect -490 -1564 -477 -1560
rect -473 -1564 -442 -1560
rect -406 -1564 -393 -1560
rect -389 -1564 -377 -1560
rect -215 -1564 -168 -1560
rect -132 -1564 -119 -1560
rect -115 -1564 -84 -1560
rect -48 -1564 -35 -1560
rect -31 -1564 -19 -1560
rect 213 -1564 260 -1560
rect 296 -1564 309 -1560
rect 313 -1564 344 -1560
rect 380 -1564 393 -1560
rect 397 -1564 409 -1560
rect 569 -1564 616 -1560
rect 652 -1564 665 -1560
rect 669 -1564 700 -1560
rect 736 -1564 749 -1560
rect 753 -1564 765 -1560
rect 967 -1564 1014 -1560
rect 1050 -1564 1063 -1560
rect 1067 -1564 1098 -1560
rect 1134 -1564 1147 -1560
rect 1151 -1564 1163 -1560
rect -1261 -1571 -1249 -1567
rect -1245 -1571 -1135 -1567
rect -1114 -1571 -1083 -1567
rect -942 -1571 -924 -1567
rect -920 -1571 -810 -1567
rect -789 -1571 -758 -1567
rect -584 -1571 -566 -1567
rect -562 -1571 -452 -1567
rect -431 -1571 -400 -1567
rect -226 -1571 -208 -1567
rect -204 -1571 -94 -1567
rect -73 -1571 -42 -1567
rect 198 -1571 199 -1567
rect 203 -1571 220 -1567
rect 224 -1571 334 -1567
rect 355 -1571 386 -1567
rect 557 -1571 576 -1567
rect 580 -1571 690 -1567
rect 711 -1571 742 -1567
rect 955 -1571 974 -1567
rect 978 -1571 1088 -1567
rect 1109 -1571 1140 -1567
rect -1214 -1578 -1191 -1574
rect -1172 -1578 -1153 -1574
rect -889 -1578 -866 -1574
rect -847 -1578 -828 -1574
rect -531 -1578 -508 -1574
rect -489 -1578 -470 -1574
rect -173 -1578 -150 -1574
rect -131 -1578 -112 -1574
rect 255 -1578 278 -1574
rect 297 -1578 316 -1574
rect 611 -1578 634 -1574
rect 653 -1578 672 -1574
rect 1009 -1578 1032 -1574
rect 1051 -1578 1070 -1574
rect 1633 -1589 1695 -1470
rect -1421 -1593 -1251 -1589
rect -1247 -1593 -1234 -1589
rect -1230 -1593 -1193 -1589
rect -1189 -1593 -1151 -1589
rect -1147 -1593 -1109 -1589
rect -1105 -1593 -1068 -1589
rect -1064 -1593 -926 -1589
rect -922 -1593 -909 -1589
rect -905 -1593 -868 -1589
rect -864 -1593 -826 -1589
rect -822 -1593 -784 -1589
rect -780 -1593 -743 -1589
rect -739 -1593 -568 -1589
rect -564 -1593 -551 -1589
rect -547 -1593 -510 -1589
rect -506 -1593 -468 -1589
rect -464 -1593 -426 -1589
rect -422 -1593 -385 -1589
rect -381 -1593 -210 -1589
rect -206 -1593 -193 -1589
rect -189 -1593 -152 -1589
rect -148 -1593 -110 -1589
rect -106 -1593 -68 -1589
rect -64 -1593 -27 -1589
rect -23 -1593 218 -1589
rect 222 -1593 235 -1589
rect 239 -1593 276 -1589
rect 280 -1593 318 -1589
rect 322 -1593 360 -1589
rect 364 -1593 401 -1589
rect 405 -1593 574 -1589
rect 578 -1593 591 -1589
rect 595 -1593 632 -1589
rect 636 -1593 674 -1589
rect 678 -1593 716 -1589
rect 720 -1593 757 -1589
rect 761 -1593 972 -1589
rect 976 -1593 989 -1589
rect 993 -1593 1030 -1589
rect 1034 -1593 1072 -1589
rect 1076 -1593 1114 -1589
rect 1118 -1593 1155 -1589
rect 1159 -1593 1695 -1589
rect -1495 -1622 -1251 -1618
rect -1247 -1622 -1234 -1618
rect -1230 -1622 -1214 -1618
rect -1210 -1622 -1193 -1618
rect -1189 -1622 -1172 -1618
rect -1168 -1622 -1151 -1618
rect -1147 -1622 -1130 -1618
rect -1126 -1622 -1109 -1618
rect -1105 -1622 -1088 -1618
rect -1084 -1622 -1068 -1618
rect -1064 -1622 -926 -1618
rect -922 -1622 -909 -1618
rect -905 -1622 -889 -1618
rect -885 -1622 -868 -1618
rect -864 -1622 -847 -1618
rect -843 -1622 -826 -1618
rect -822 -1622 -805 -1618
rect -801 -1622 -784 -1618
rect -780 -1622 -763 -1618
rect -759 -1622 -743 -1618
rect -739 -1622 -568 -1618
rect -564 -1622 -551 -1618
rect -547 -1622 -531 -1618
rect -527 -1622 -510 -1618
rect -506 -1622 -489 -1618
rect -485 -1622 -468 -1618
rect -464 -1622 -447 -1618
rect -443 -1622 -426 -1618
rect -422 -1622 -405 -1618
rect -401 -1622 -385 -1618
rect -381 -1622 -210 -1618
rect -206 -1622 -193 -1618
rect -189 -1622 -173 -1618
rect -169 -1622 -152 -1618
rect -148 -1622 -131 -1618
rect -127 -1622 -110 -1618
rect -106 -1622 -89 -1618
rect -85 -1622 -68 -1618
rect -64 -1622 -47 -1618
rect -43 -1622 -27 -1618
rect -23 -1622 218 -1618
rect 222 -1622 235 -1618
rect 239 -1622 255 -1618
rect 259 -1622 276 -1618
rect 280 -1622 297 -1618
rect 301 -1622 318 -1618
rect 322 -1622 339 -1618
rect 343 -1622 360 -1618
rect 364 -1622 381 -1618
rect 385 -1622 401 -1618
rect 405 -1622 574 -1618
rect 578 -1622 591 -1618
rect 595 -1622 611 -1618
rect 615 -1622 632 -1618
rect 636 -1622 653 -1618
rect 657 -1622 674 -1618
rect 678 -1622 695 -1618
rect 699 -1622 716 -1618
rect 720 -1622 737 -1618
rect 741 -1622 757 -1618
rect 761 -1622 972 -1618
rect 976 -1622 989 -1618
rect 993 -1622 1009 -1618
rect 1013 -1622 1030 -1618
rect 1034 -1622 1051 -1618
rect 1055 -1622 1072 -1618
rect 1076 -1622 1093 -1618
rect 1097 -1622 1114 -1618
rect 1118 -1622 1135 -1618
rect 1139 -1622 1155 -1618
rect 1159 -1622 1330 -1618
rect 1334 -1622 1347 -1618
rect 1351 -1622 1367 -1618
rect 1371 -1622 1388 -1618
rect 1392 -1622 1409 -1618
rect 1413 -1622 1430 -1618
rect 1434 -1622 1451 -1618
rect 1455 -1622 1472 -1618
rect 1476 -1622 1493 -1618
rect 1497 -1622 1513 -1618
rect 1517 -1622 1617 -1618
rect -1495 -1739 -1433 -1622
rect -1229 -1670 -1195 -1666
rect -1131 -1670 -1111 -1666
rect -1096 -1670 -1062 -1666
rect -904 -1670 -870 -1666
rect -806 -1670 -786 -1666
rect -771 -1670 -737 -1666
rect -546 -1670 -512 -1666
rect -448 -1670 -428 -1666
rect -413 -1670 -379 -1666
rect -188 -1670 -154 -1666
rect -90 -1670 -70 -1666
rect -55 -1670 -21 -1666
rect 240 -1670 274 -1666
rect 338 -1670 358 -1666
rect 373 -1670 407 -1666
rect 596 -1670 630 -1666
rect 694 -1670 714 -1666
rect 729 -1670 763 -1666
rect 994 -1670 1028 -1666
rect 1092 -1670 1112 -1666
rect 1127 -1670 1161 -1666
rect 1352 -1670 1386 -1666
rect 1450 -1670 1470 -1666
rect 1485 -1670 1519 -1666
rect -1268 -1678 -1253 -1674
rect -1249 -1678 -1219 -1674
rect -1198 -1678 -1167 -1674
rect -1138 -1678 -1107 -1674
rect -1096 -1678 -1069 -1674
rect -944 -1678 -928 -1674
rect -924 -1678 -894 -1674
rect -873 -1678 -842 -1674
rect -813 -1678 -782 -1674
rect -771 -1678 -744 -1674
rect -585 -1678 -570 -1674
rect -566 -1678 -536 -1674
rect -515 -1678 -484 -1674
rect -455 -1678 -424 -1674
rect -413 -1678 -386 -1674
rect -227 -1678 -212 -1674
rect -208 -1678 -178 -1674
rect -157 -1678 -126 -1674
rect -97 -1678 -66 -1674
rect -55 -1678 -28 -1674
rect 201 -1678 216 -1674
rect 220 -1678 250 -1674
rect 271 -1678 302 -1674
rect 331 -1678 362 -1674
rect 373 -1678 400 -1674
rect 557 -1678 572 -1674
rect 576 -1678 606 -1674
rect 627 -1678 658 -1674
rect 687 -1678 718 -1674
rect 729 -1678 756 -1674
rect 955 -1678 970 -1674
rect 974 -1678 1004 -1674
rect 1025 -1678 1056 -1674
rect 1085 -1678 1116 -1674
rect 1127 -1678 1154 -1674
rect 1313 -1678 1328 -1674
rect 1332 -1678 1362 -1674
rect 1383 -1678 1414 -1674
rect 1443 -1678 1474 -1674
rect 1485 -1678 1512 -1674
rect -1256 -1685 -1209 -1681
rect -1173 -1685 -1160 -1681
rect -1156 -1685 -1125 -1681
rect -1089 -1685 -1076 -1681
rect -1072 -1685 -1060 -1681
rect -931 -1685 -884 -1681
rect -848 -1685 -835 -1681
rect -831 -1685 -800 -1681
rect -764 -1685 -751 -1681
rect -747 -1685 -735 -1681
rect -573 -1685 -526 -1681
rect -490 -1685 -477 -1681
rect -473 -1685 -442 -1681
rect -406 -1685 -393 -1681
rect -389 -1685 -377 -1681
rect -215 -1685 -168 -1681
rect -132 -1685 -119 -1681
rect -115 -1685 -84 -1681
rect -48 -1685 -35 -1681
rect -31 -1685 -19 -1681
rect 213 -1685 260 -1681
rect 296 -1685 309 -1681
rect 313 -1685 344 -1681
rect 380 -1685 393 -1681
rect 397 -1685 409 -1681
rect 569 -1685 616 -1681
rect 652 -1685 665 -1681
rect 669 -1685 700 -1681
rect 736 -1685 749 -1681
rect 753 -1685 765 -1681
rect 967 -1685 1014 -1681
rect 1050 -1685 1063 -1681
rect 1067 -1685 1098 -1681
rect 1134 -1685 1147 -1681
rect 1151 -1685 1163 -1681
rect 1325 -1685 1372 -1681
rect 1408 -1685 1421 -1681
rect 1425 -1685 1456 -1681
rect 1492 -1685 1505 -1681
rect 1509 -1685 1521 -1681
rect -1266 -1692 -1249 -1688
rect -1245 -1692 -1135 -1688
rect -1114 -1692 -1083 -1688
rect -937 -1692 -924 -1688
rect -920 -1692 -810 -1688
rect -789 -1692 -758 -1688
rect -584 -1692 -566 -1688
rect -562 -1692 -452 -1688
rect -431 -1692 -400 -1688
rect -226 -1692 -208 -1688
rect -204 -1692 -94 -1688
rect -73 -1692 -42 -1688
rect 203 -1692 220 -1688
rect 224 -1692 334 -1688
rect 355 -1692 386 -1688
rect 564 -1692 576 -1688
rect 580 -1692 690 -1688
rect 711 -1692 742 -1688
rect 955 -1692 974 -1688
rect 978 -1692 1088 -1688
rect 1109 -1692 1140 -1688
rect 1315 -1692 1332 -1688
rect 1336 -1692 1446 -1688
rect 1467 -1692 1498 -1688
rect -1214 -1699 -1191 -1695
rect -1172 -1699 -1153 -1695
rect -889 -1699 -866 -1695
rect -847 -1699 -828 -1695
rect -531 -1699 -508 -1695
rect -489 -1699 -470 -1695
rect -173 -1699 -150 -1695
rect -131 -1699 -112 -1695
rect 255 -1699 278 -1695
rect 297 -1699 316 -1695
rect 611 -1699 634 -1695
rect 653 -1699 672 -1695
rect 1009 -1699 1032 -1695
rect 1051 -1699 1070 -1695
rect 1367 -1699 1390 -1695
rect 1409 -1699 1428 -1695
rect 1633 -1710 1695 -1593
rect -1421 -1714 -1251 -1710
rect -1247 -1714 -1234 -1710
rect -1230 -1714 -1193 -1710
rect -1189 -1714 -1151 -1710
rect -1147 -1714 -1109 -1710
rect -1105 -1714 -1068 -1710
rect -1064 -1714 -926 -1710
rect -922 -1714 -909 -1710
rect -905 -1714 -868 -1710
rect -864 -1714 -826 -1710
rect -822 -1714 -784 -1710
rect -780 -1714 -743 -1710
rect -739 -1714 -568 -1710
rect -564 -1714 -551 -1710
rect -547 -1714 -510 -1710
rect -506 -1714 -468 -1710
rect -464 -1714 -426 -1710
rect -422 -1714 -385 -1710
rect -381 -1714 -210 -1710
rect -206 -1714 -193 -1710
rect -189 -1714 -152 -1710
rect -148 -1714 -110 -1710
rect -106 -1714 -68 -1710
rect -64 -1714 -27 -1710
rect -23 -1714 218 -1710
rect 222 -1714 235 -1710
rect 239 -1714 276 -1710
rect 280 -1714 318 -1710
rect 322 -1714 360 -1710
rect 364 -1714 401 -1710
rect 405 -1714 574 -1710
rect 578 -1714 591 -1710
rect 595 -1714 632 -1710
rect 636 -1714 674 -1710
rect 678 -1714 716 -1710
rect 720 -1714 757 -1710
rect 761 -1714 972 -1710
rect 976 -1714 989 -1710
rect 993 -1714 1030 -1710
rect 1034 -1714 1072 -1710
rect 1076 -1714 1114 -1710
rect 1118 -1714 1155 -1710
rect 1159 -1714 1330 -1710
rect 1334 -1714 1347 -1710
rect 1351 -1714 1388 -1710
rect 1392 -1714 1430 -1710
rect 1434 -1714 1472 -1710
rect 1476 -1714 1513 -1710
rect 1517 -1714 1695 -1710
rect -1262 -1721 -1062 -1717
rect -949 -1722 -737 -1718
rect -585 -1722 -379 -1718
rect -227 -1721 -21 -1717
rect 201 -1722 407 -1718
rect 557 -1721 763 -1717
rect 955 -1721 1161 -1717
rect 1313 -1722 1519 -1718
rect -1495 -1743 -1251 -1739
rect -1247 -1743 -1234 -1739
rect -1230 -1743 -1214 -1739
rect -1210 -1743 -1193 -1739
rect -1189 -1743 -1172 -1739
rect -1168 -1743 -1151 -1739
rect -1147 -1743 -1130 -1739
rect -1126 -1743 -1109 -1739
rect -1105 -1743 -1088 -1739
rect -1084 -1743 -1068 -1739
rect -1064 -1743 -1029 -1739
rect -1025 -1743 -926 -1739
rect -922 -1743 -909 -1739
rect -905 -1743 -889 -1739
rect -885 -1743 -868 -1739
rect -864 -1743 -847 -1739
rect -843 -1743 -826 -1739
rect -822 -1743 -805 -1739
rect -801 -1743 -784 -1739
rect -780 -1743 -763 -1739
rect -759 -1743 -743 -1739
rect -739 -1743 -568 -1739
rect -564 -1743 -551 -1739
rect -547 -1743 -531 -1739
rect -527 -1743 -510 -1739
rect -506 -1743 -489 -1739
rect -485 -1743 -468 -1739
rect -464 -1743 -447 -1739
rect -443 -1743 -426 -1739
rect -422 -1743 -405 -1739
rect -401 -1743 -385 -1739
rect -381 -1743 -332 -1739
rect -328 -1743 -210 -1739
rect -206 -1743 -193 -1739
rect -189 -1743 -173 -1739
rect -169 -1743 -152 -1739
rect -148 -1743 -131 -1739
rect -127 -1743 -110 -1739
rect -106 -1743 -89 -1739
rect -85 -1743 -68 -1739
rect -64 -1743 -47 -1739
rect -43 -1743 -27 -1739
rect -23 -1743 218 -1739
rect 222 -1743 235 -1739
rect 239 -1743 255 -1739
rect 259 -1743 276 -1739
rect 280 -1743 297 -1739
rect 301 -1743 318 -1739
rect 322 -1743 339 -1739
rect 343 -1743 360 -1739
rect 364 -1743 381 -1739
rect 385 -1743 401 -1739
rect 405 -1743 464 -1739
rect 468 -1743 574 -1739
rect 578 -1743 591 -1739
rect 595 -1743 611 -1739
rect 615 -1743 632 -1739
rect 636 -1743 653 -1739
rect 657 -1743 674 -1739
rect 678 -1743 695 -1739
rect 699 -1743 716 -1739
rect 720 -1743 737 -1739
rect 741 -1743 757 -1739
rect 761 -1743 972 -1739
rect 976 -1743 989 -1739
rect 993 -1743 1009 -1739
rect 1013 -1743 1030 -1739
rect 1034 -1743 1051 -1739
rect 1055 -1743 1072 -1739
rect 1076 -1743 1093 -1739
rect 1097 -1743 1114 -1739
rect 1118 -1743 1135 -1739
rect 1139 -1743 1155 -1739
rect 1159 -1743 1203 -1739
rect 1207 -1743 1330 -1739
rect 1334 -1743 1347 -1739
rect 1351 -1743 1367 -1739
rect 1371 -1743 1388 -1739
rect 1392 -1743 1409 -1739
rect 1413 -1743 1430 -1739
rect 1434 -1743 1451 -1739
rect 1455 -1743 1472 -1739
rect 1476 -1743 1493 -1739
rect 1497 -1743 1513 -1739
rect 1517 -1743 1617 -1739
rect -1495 -1854 -1433 -1743
rect -1229 -1791 -1195 -1787
rect -1131 -1791 -1111 -1787
rect -1096 -1791 -1056 -1787
rect -1017 -1792 -1013 -1788
rect -904 -1791 -870 -1787
rect -806 -1791 -786 -1787
rect -771 -1791 -737 -1787
rect -546 -1791 -512 -1787
rect -448 -1791 -428 -1787
rect -413 -1791 -379 -1787
rect -320 -1792 -316 -1788
rect -188 -1791 -154 -1787
rect -90 -1791 -70 -1787
rect -55 -1791 -21 -1787
rect 240 -1791 274 -1787
rect 338 -1791 358 -1787
rect 373 -1791 407 -1787
rect 476 -1792 480 -1788
rect 596 -1791 630 -1787
rect 694 -1791 714 -1787
rect 729 -1791 763 -1787
rect 994 -1791 1028 -1787
rect 1092 -1791 1112 -1787
rect 1127 -1791 1161 -1787
rect 1215 -1792 1219 -1788
rect 1352 -1791 1386 -1787
rect 1450 -1791 1470 -1787
rect 1485 -1791 1519 -1787
rect -1345 -1799 -1253 -1795
rect -1249 -1799 -1219 -1795
rect -1198 -1799 -1167 -1795
rect -1138 -1799 -1107 -1795
rect -1096 -1799 -1069 -1795
rect -938 -1799 -928 -1795
rect -924 -1799 -894 -1795
rect -873 -1799 -842 -1795
rect -813 -1799 -782 -1795
rect -771 -1799 -744 -1795
rect -579 -1799 -570 -1795
rect -566 -1799 -536 -1795
rect -515 -1799 -484 -1795
rect -455 -1799 -424 -1795
rect -413 -1799 -386 -1795
rect -221 -1799 -212 -1795
rect -208 -1799 -178 -1795
rect -157 -1799 -126 -1795
rect -97 -1799 -66 -1795
rect -55 -1799 -28 -1795
rect 207 -1799 216 -1795
rect 220 -1799 250 -1795
rect 271 -1799 302 -1795
rect 331 -1799 362 -1795
rect 373 -1799 400 -1795
rect 563 -1799 572 -1795
rect 576 -1799 606 -1795
rect 627 -1799 658 -1795
rect 687 -1799 718 -1795
rect 729 -1799 756 -1795
rect 961 -1799 970 -1795
rect 974 -1799 1004 -1795
rect 1025 -1799 1056 -1795
rect 1085 -1799 1116 -1795
rect 1127 -1799 1154 -1795
rect 1319 -1799 1328 -1795
rect 1332 -1799 1362 -1795
rect 1383 -1799 1414 -1795
rect 1443 -1799 1474 -1795
rect 1485 -1799 1512 -1795
rect -1256 -1806 -1209 -1802
rect -1173 -1806 -1160 -1802
rect -1156 -1806 -1125 -1802
rect -1089 -1806 -1076 -1802
rect -1072 -1806 -1060 -1802
rect -931 -1806 -884 -1802
rect -848 -1806 -835 -1802
rect -831 -1806 -800 -1802
rect -764 -1806 -751 -1802
rect -747 -1806 -735 -1802
rect -573 -1806 -526 -1802
rect -490 -1806 -477 -1802
rect -473 -1806 -442 -1802
rect -406 -1806 -393 -1802
rect -389 -1806 -377 -1802
rect -215 -1806 -168 -1802
rect -132 -1806 -119 -1802
rect -115 -1806 -84 -1802
rect -48 -1806 -35 -1802
rect -31 -1806 -19 -1802
rect 213 -1806 260 -1802
rect 296 -1806 309 -1802
rect 313 -1806 344 -1802
rect 380 -1806 393 -1802
rect 397 -1806 409 -1802
rect 569 -1806 616 -1802
rect 652 -1806 665 -1802
rect 669 -1806 700 -1802
rect 736 -1806 749 -1802
rect 753 -1806 765 -1802
rect 967 -1806 1014 -1802
rect 1050 -1806 1063 -1802
rect 1067 -1806 1098 -1802
rect 1134 -1806 1147 -1802
rect 1151 -1806 1163 -1802
rect 1325 -1806 1372 -1802
rect 1408 -1806 1421 -1802
rect 1425 -1806 1456 -1802
rect 1492 -1806 1505 -1802
rect 1509 -1806 1521 -1802
rect -1266 -1813 -1249 -1809
rect -1245 -1813 -1135 -1809
rect -1114 -1813 -1083 -1809
rect -942 -1813 -924 -1809
rect -920 -1813 -810 -1809
rect -789 -1813 -758 -1809
rect -584 -1813 -566 -1809
rect -562 -1813 -452 -1809
rect -431 -1813 -400 -1809
rect -226 -1813 -208 -1809
rect -204 -1813 -94 -1809
rect -73 -1813 -42 -1809
rect 203 -1813 220 -1809
rect 224 -1813 334 -1809
rect 355 -1813 386 -1809
rect 557 -1813 576 -1809
rect 580 -1813 690 -1809
rect 711 -1813 742 -1809
rect 955 -1813 974 -1809
rect 978 -1813 1088 -1809
rect 1109 -1813 1140 -1809
rect 1308 -1813 1309 -1809
rect 1313 -1813 1332 -1809
rect 1336 -1813 1446 -1809
rect 1467 -1813 1498 -1809
rect -1214 -1820 -1191 -1816
rect -1172 -1820 -1153 -1816
rect -889 -1820 -866 -1816
rect -847 -1820 -828 -1816
rect -531 -1820 -508 -1816
rect -489 -1820 -470 -1816
rect -173 -1820 -150 -1816
rect -131 -1820 -112 -1816
rect 255 -1820 278 -1816
rect 297 -1820 316 -1816
rect 611 -1820 634 -1816
rect 653 -1820 672 -1816
rect 1009 -1820 1032 -1816
rect 1051 -1820 1070 -1816
rect 1367 -1820 1390 -1816
rect 1409 -1820 1428 -1816
rect 1633 -1831 1695 -1714
rect -1421 -1835 -1251 -1831
rect -1247 -1835 -1234 -1831
rect -1230 -1835 -1193 -1831
rect -1189 -1835 -1151 -1831
rect -1147 -1835 -1109 -1831
rect -1105 -1835 -1068 -1831
rect -1064 -1835 -1029 -1831
rect -1025 -1835 -926 -1831
rect -922 -1835 -909 -1831
rect -905 -1835 -868 -1831
rect -864 -1835 -826 -1831
rect -822 -1835 -784 -1831
rect -780 -1835 -743 -1831
rect -739 -1835 -568 -1831
rect -564 -1835 -551 -1831
rect -547 -1835 -510 -1831
rect -506 -1835 -468 -1831
rect -464 -1835 -426 -1831
rect -422 -1835 -385 -1831
rect -381 -1835 -332 -1831
rect -328 -1835 -210 -1831
rect -206 -1835 -193 -1831
rect -189 -1835 -152 -1831
rect -148 -1835 -110 -1831
rect -106 -1835 -68 -1831
rect -64 -1835 -27 -1831
rect -23 -1835 218 -1831
rect 222 -1835 235 -1831
rect 239 -1835 276 -1831
rect 280 -1835 318 -1831
rect 322 -1835 360 -1831
rect 364 -1835 401 -1831
rect 405 -1835 464 -1831
rect 468 -1835 574 -1831
rect 578 -1835 591 -1831
rect 595 -1835 632 -1831
rect 636 -1835 674 -1831
rect 678 -1835 716 -1831
rect 720 -1835 757 -1831
rect 761 -1835 972 -1831
rect 976 -1835 989 -1831
rect 993 -1835 1030 -1831
rect 1034 -1835 1072 -1831
rect 1076 -1835 1114 -1831
rect 1118 -1835 1155 -1831
rect 1159 -1835 1203 -1831
rect 1207 -1835 1330 -1831
rect 1334 -1835 1347 -1831
rect 1351 -1835 1388 -1831
rect 1392 -1835 1430 -1831
rect 1434 -1835 1472 -1831
rect 1476 -1835 1513 -1831
rect 1517 -1835 1695 -1831
rect -1495 -1858 -1251 -1854
rect -1247 -1858 -1234 -1854
rect -1230 -1858 -1214 -1854
rect -1210 -1858 -1193 -1854
rect -1189 -1858 -1172 -1854
rect -1168 -1858 -1151 -1854
rect -1147 -1858 -1130 -1854
rect -1126 -1858 -1109 -1854
rect -1105 -1858 -1088 -1854
rect -1084 -1858 -1068 -1854
rect -1064 -1858 -1029 -1854
rect -1025 -1858 -673 -1854
rect -669 -1858 -332 -1854
rect -328 -1858 464 -1854
rect 468 -1858 841 -1854
rect 845 -1858 1203 -1854
rect 1207 -1858 1617 -1854
rect -1495 -1966 -1433 -1858
rect -1096 -1898 -1062 -1894
rect -1229 -1906 -1195 -1902
rect -1131 -1906 -1111 -1902
rect -1017 -1907 -1013 -1903
rect -661 -1907 -657 -1903
rect -320 -1907 -316 -1903
rect 476 -1907 480 -1903
rect 853 -1907 857 -1903
rect 1215 -1907 1219 -1903
rect -1421 -1914 -1253 -1910
rect -1249 -1914 -1219 -1910
rect -1198 -1914 -1167 -1910
rect -1138 -1914 -1107 -1910
rect -1096 -1914 -1069 -1910
rect -1256 -1921 -1209 -1917
rect -1173 -1921 -1160 -1917
rect -1156 -1921 -1125 -1917
rect -1089 -1921 -1076 -1917
rect -1072 -1921 -1060 -1917
rect -1274 -1928 -1273 -1924
rect -1269 -1928 -1249 -1924
rect -1245 -1928 -1135 -1924
rect -1114 -1928 -1083 -1924
rect -1214 -1935 -1191 -1931
rect -1172 -1935 -1153 -1931
rect 1633 -1946 1695 -1835
rect -1421 -1950 -1251 -1946
rect -1247 -1950 -1234 -1946
rect -1230 -1950 -1193 -1946
rect -1189 -1950 -1151 -1946
rect -1147 -1950 -1109 -1946
rect -1105 -1950 -1068 -1946
rect -1064 -1950 -1029 -1946
rect -1025 -1950 -673 -1946
rect -669 -1950 -332 -1946
rect -328 -1950 464 -1946
rect 468 -1950 841 -1946
rect 845 -1950 1203 -1946
rect 1207 -1950 1695 -1946
rect -1495 -1970 -1339 -1966
rect -1335 -1970 -1322 -1966
rect -1318 -1970 -935 -1966
rect -931 -1970 -918 -1966
rect -914 -1970 -577 -1966
rect -573 -1970 -560 -1966
rect -556 -1970 -219 -1966
rect -215 -1970 -202 -1966
rect -198 -1970 209 -1966
rect 213 -1970 226 -1966
rect 230 -1970 565 -1966
rect 569 -1970 582 -1966
rect 586 -1970 963 -1966
rect 967 -1970 980 -1966
rect 984 -1970 1321 -1966
rect 1325 -1970 1338 -1966
rect 1342 -1970 1617 -1966
rect -1495 -2085 -1433 -1970
rect -1334 -2002 -1056 -1998
rect -930 -2002 -737 -1998
rect -572 -2002 -379 -1998
rect -214 -2002 -21 -1998
rect 214 -2002 407 -1998
rect 570 -2002 763 -1998
rect 968 -2002 1161 -1998
rect 1326 -2002 1519 -1998
rect -1323 -2010 -1062 -2006
rect -1058 -2010 -923 -2006
rect -919 -2010 -565 -2006
rect -561 -2010 -207 -2006
rect -203 -2010 221 -2006
rect 225 -2010 577 -2006
rect 581 -2010 975 -2006
rect 979 -2010 1333 -2006
rect 1337 -2010 1617 -2006
rect -943 -2023 -909 -2019
rect -591 -2023 -551 -2019
rect -233 -2023 -193 -2019
rect 195 -2023 235 -2019
rect 551 -2023 591 -2019
rect 949 -2023 989 -2019
rect 1307 -2023 1347 -2019
rect 1633 -2058 1695 -1950
rect -1421 -2062 -1322 -2058
rect -1318 -2062 -918 -2058
rect -914 -2062 -560 -2058
rect -556 -2062 -202 -2058
rect -198 -2062 226 -2058
rect 230 -2062 582 -2058
rect 586 -2062 980 -2058
rect 984 -2062 1338 -2058
rect 1342 -2062 1695 -2058
rect -1495 -2089 -1251 -2085
rect -1247 -2089 -1234 -2085
rect -1230 -2089 -1194 -2085
rect -1190 -2089 -1173 -2085
rect -1169 -2089 -926 -2085
rect -922 -2089 -900 -2085
rect -896 -2089 -883 -2085
rect -879 -2089 -843 -2085
rect -839 -2089 -822 -2085
rect -818 -2089 -805 -2085
rect -801 -2089 -765 -2085
rect -761 -2089 -741 -2085
rect -737 -2089 -704 -2085
rect -700 -2089 -568 -2085
rect -564 -2089 -542 -2085
rect -538 -2089 -525 -2085
rect -521 -2089 -485 -2085
rect -481 -2089 -464 -2085
rect -460 -2089 -447 -2085
rect -443 -2089 -407 -2085
rect -403 -2089 -383 -2085
rect -379 -2089 -346 -2085
rect -342 -2089 -210 -2085
rect -206 -2089 -184 -2085
rect -180 -2089 -167 -2085
rect -163 -2089 -127 -2085
rect -123 -2089 -106 -2085
rect -102 -2089 -89 -2085
rect -85 -2089 -49 -2085
rect -45 -2089 -25 -2085
rect -21 -2089 12 -2085
rect 16 -2089 218 -2085
rect 222 -2089 244 -2085
rect 248 -2089 261 -2085
rect 265 -2089 301 -2085
rect 305 -2089 322 -2085
rect 326 -2089 339 -2085
rect 343 -2089 379 -2085
rect 383 -2089 403 -2085
rect 407 -2089 440 -2085
rect 444 -2089 574 -2085
rect 578 -2089 600 -2085
rect 604 -2089 617 -2085
rect 621 -2089 657 -2085
rect 661 -2089 678 -2085
rect 682 -2089 695 -2085
rect 699 -2089 735 -2085
rect 739 -2089 759 -2085
rect 763 -2089 796 -2085
rect 800 -2089 972 -2085
rect 976 -2089 998 -2085
rect 1002 -2089 1015 -2085
rect 1019 -2089 1055 -2085
rect 1059 -2089 1076 -2085
rect 1080 -2089 1093 -2085
rect 1097 -2089 1133 -2085
rect 1137 -2089 1157 -2085
rect 1161 -2089 1194 -2085
rect 1198 -2089 1330 -2085
rect 1334 -2089 1356 -2085
rect 1360 -2089 1373 -2085
rect 1377 -2089 1413 -2085
rect 1417 -2089 1434 -2085
rect 1438 -2089 1451 -2085
rect 1455 -2089 1491 -2085
rect 1495 -2089 1515 -2085
rect 1519 -2089 1552 -2085
rect 1556 -2089 1617 -2085
rect -1495 -2229 -1433 -2089
rect -926 -2093 -922 -2089
rect -900 -2093 -896 -2089
rect -883 -2093 -879 -2089
rect -843 -2093 -839 -2089
rect -822 -2093 -818 -2089
rect -805 -2093 -801 -2089
rect -765 -2093 -761 -2089
rect -741 -2093 -737 -2089
rect -704 -2093 -700 -2089
rect -568 -2093 -564 -2089
rect -542 -2093 -538 -2089
rect -525 -2093 -521 -2089
rect -485 -2093 -481 -2089
rect -464 -2093 -460 -2089
rect -447 -2093 -443 -2089
rect -407 -2093 -403 -2089
rect -383 -2093 -379 -2089
rect -346 -2093 -342 -2089
rect -210 -2093 -206 -2089
rect -184 -2093 -180 -2089
rect -167 -2093 -163 -2089
rect -127 -2093 -123 -2089
rect -106 -2093 -102 -2089
rect -89 -2093 -85 -2089
rect -49 -2093 -45 -2089
rect -25 -2093 -21 -2089
rect 12 -2093 16 -2089
rect 218 -2093 222 -2089
rect 244 -2093 248 -2089
rect 261 -2093 265 -2089
rect 301 -2093 305 -2089
rect 322 -2093 326 -2089
rect 339 -2093 343 -2089
rect 379 -2093 383 -2089
rect 403 -2093 407 -2089
rect 440 -2093 444 -2089
rect 574 -2093 578 -2089
rect 600 -2093 604 -2089
rect 617 -2093 621 -2089
rect 657 -2093 661 -2089
rect 678 -2093 682 -2089
rect 695 -2093 699 -2089
rect 735 -2093 739 -2089
rect 759 -2093 763 -2089
rect 796 -2093 800 -2089
rect 972 -2093 976 -2089
rect 998 -2093 1002 -2089
rect 1015 -2093 1019 -2089
rect 1055 -2093 1059 -2089
rect 1076 -2093 1080 -2089
rect 1093 -2093 1097 -2089
rect 1133 -2093 1137 -2089
rect 1157 -2093 1161 -2089
rect 1194 -2093 1198 -2089
rect 1330 -2093 1334 -2089
rect 1356 -2093 1360 -2089
rect 1373 -2093 1377 -2089
rect 1413 -2093 1417 -2089
rect 1434 -2093 1438 -2089
rect 1451 -2093 1455 -2089
rect 1491 -2093 1495 -2089
rect 1515 -2093 1519 -2089
rect 1552 -2093 1556 -2089
rect -920 -2108 -858 -2104
rect -854 -2108 -824 -2104
rect -776 -2108 -746 -2104
rect -562 -2108 -500 -2104
rect -496 -2108 -466 -2104
rect -418 -2108 -388 -2104
rect -204 -2108 -142 -2104
rect -138 -2108 -108 -2104
rect -60 -2108 -30 -2104
rect 224 -2108 286 -2104
rect 290 -2108 320 -2104
rect 368 -2108 398 -2104
rect 580 -2108 642 -2104
rect 646 -2108 676 -2104
rect 724 -2108 754 -2104
rect 978 -2108 1040 -2104
rect 1044 -2108 1074 -2104
rect 1122 -2108 1152 -2104
rect 1336 -2108 1398 -2104
rect 1402 -2108 1432 -2104
rect 1480 -2108 1510 -2104
rect -913 -2115 -882 -2111
rect -555 -2115 -524 -2111
rect -197 -2115 -166 -2111
rect 231 -2115 262 -2111
rect 587 -2115 618 -2111
rect 985 -2115 1016 -2111
rect 1343 -2115 1374 -2111
rect -931 -2122 -848 -2118
rect -809 -2122 -706 -2118
rect -573 -2122 -490 -2118
rect -451 -2122 -348 -2118
rect -215 -2122 -132 -2118
rect -93 -2122 10 -2118
rect 213 -2122 296 -2118
rect 335 -2122 438 -2118
rect 569 -2122 652 -2118
rect 691 -2122 794 -2118
rect 967 -2122 1050 -2118
rect 1089 -2122 1192 -2118
rect 1325 -2122 1408 -2118
rect 1447 -2122 1550 -2118
rect -949 -2129 -928 -2125
rect -894 -2129 -865 -2125
rect -861 -2129 -780 -2125
rect -691 -2129 -592 -2125
rect -585 -2129 -570 -2125
rect -536 -2129 -507 -2125
rect -503 -2129 -422 -2125
rect -333 -2126 -234 -2122
rect -596 -2133 -592 -2129
rect -238 -2133 -234 -2126
rect -227 -2129 -212 -2125
rect -178 -2129 -149 -2125
rect -145 -2129 -64 -2125
rect 25 -2129 194 -2125
rect 201 -2129 216 -2125
rect 250 -2129 279 -2125
rect 283 -2129 364 -2125
rect 453 -2129 550 -2125
rect 557 -2129 572 -2125
rect 606 -2129 635 -2125
rect 639 -2129 720 -2125
rect 809 -2129 948 -2125
rect 955 -2129 970 -2125
rect 1004 -2129 1033 -2125
rect 1037 -2129 1118 -2125
rect 1207 -2127 1300 -2123
rect 190 -2133 194 -2129
rect 546 -2133 550 -2129
rect 944 -2133 948 -2129
rect 1296 -2133 1300 -2127
rect 1307 -2129 1328 -2125
rect 1362 -2129 1391 -2125
rect 1395 -2129 1476 -2125
rect -1256 -2138 -1199 -2134
rect -1160 -2137 -902 -2133
rect -887 -2137 -804 -2133
rect -783 -2137 -689 -2133
rect -596 -2137 -544 -2133
rect -529 -2137 -446 -2133
rect -425 -2137 -331 -2133
rect -238 -2137 -186 -2133
rect -171 -2137 -88 -2133
rect -67 -2137 27 -2133
rect 190 -2137 242 -2133
rect 257 -2137 340 -2133
rect 361 -2137 455 -2133
rect 546 -2137 598 -2133
rect 613 -2137 696 -2133
rect 717 -2137 811 -2133
rect 944 -2137 996 -2133
rect 1011 -2137 1094 -2133
rect 1115 -2137 1209 -2133
rect 1296 -2137 1354 -2133
rect 1369 -2137 1452 -2133
rect 1473 -2137 1567 -2133
rect -1262 -2145 -1249 -2141
rect -1245 -2145 -1209 -2141
rect -1205 -2145 -1189 -2141
rect -943 -2144 -924 -2140
rect -905 -2144 -776 -2140
rect -591 -2144 -566 -2140
rect -547 -2144 -418 -2140
rect -233 -2144 -208 -2140
rect -189 -2144 -60 -2140
rect 195 -2144 220 -2140
rect 239 -2144 368 -2140
rect 551 -2144 576 -2140
rect 595 -2144 724 -2140
rect 949 -2144 974 -2140
rect 993 -2144 1122 -2140
rect 1313 -2144 1332 -2140
rect 1351 -2144 1480 -2140
rect -1309 -2152 -1253 -2148
rect -1249 -2152 -1223 -2148
rect -1219 -2152 -1175 -2148
rect -898 -2151 -794 -2147
rect -790 -2151 -760 -2147
rect -540 -2151 -436 -2147
rect -432 -2151 -402 -2147
rect -182 -2151 -78 -2147
rect -74 -2151 -44 -2147
rect 246 -2151 350 -2147
rect 354 -2151 384 -2147
rect 602 -2151 706 -2147
rect 710 -2151 740 -2147
rect 1000 -2151 1104 -2147
rect 1108 -2151 1138 -2147
rect 1358 -2151 1462 -2147
rect 1466 -2151 1496 -2147
rect -1212 -2159 -1158 -2155
rect -924 -2158 -872 -2154
rect -868 -2158 -838 -2154
rect -566 -2158 -514 -2154
rect -510 -2158 -480 -2154
rect -208 -2158 -156 -2154
rect -152 -2158 -122 -2154
rect 220 -2158 272 -2154
rect 276 -2158 306 -2154
rect 576 -2158 628 -2154
rect 632 -2158 662 -2154
rect 974 -2158 1026 -2154
rect 1030 -2158 1060 -2154
rect 1332 -2158 1384 -2154
rect 1388 -2158 1418 -2154
rect -1230 -2166 -1198 -2162
rect -879 -2166 -847 -2162
rect -883 -2169 -879 -2166
rect -847 -2169 -843 -2166
rect -801 -2166 -769 -2162
rect -805 -2169 -801 -2166
rect -769 -2169 -765 -2166
rect -521 -2166 -489 -2162
rect -525 -2169 -521 -2166
rect -489 -2169 -485 -2166
rect -443 -2166 -411 -2162
rect -447 -2169 -443 -2166
rect -411 -2169 -407 -2166
rect -163 -2166 -131 -2162
rect -167 -2169 -163 -2166
rect -131 -2169 -127 -2166
rect -85 -2166 -53 -2162
rect -89 -2169 -85 -2166
rect -53 -2169 -49 -2166
rect 265 -2166 297 -2162
rect 261 -2169 265 -2166
rect 297 -2169 301 -2166
rect 343 -2166 375 -2162
rect 339 -2169 343 -2166
rect 375 -2169 379 -2166
rect 621 -2166 653 -2162
rect 617 -2169 621 -2166
rect 653 -2169 657 -2166
rect 699 -2166 731 -2162
rect 695 -2169 699 -2166
rect 731 -2169 735 -2166
rect 1019 -2166 1051 -2162
rect 1015 -2169 1019 -2166
rect 1051 -2169 1055 -2166
rect 1097 -2166 1129 -2162
rect 1093 -2169 1097 -2166
rect 1129 -2169 1133 -2166
rect 1377 -2166 1409 -2162
rect 1373 -2169 1377 -2166
rect 1409 -2169 1413 -2166
rect 1455 -2166 1487 -2162
rect 1451 -2169 1455 -2166
rect 1487 -2169 1491 -2166
rect -926 -2177 -922 -2173
rect -900 -2177 -896 -2173
rect -857 -2177 -853 -2173
rect -822 -2177 -818 -2173
rect -778 -2177 -774 -2173
rect -761 -2177 -757 -2173
rect -725 -2177 -721 -2173
rect -704 -2177 -700 -2173
rect -568 -2177 -564 -2173
rect -542 -2177 -538 -2173
rect -499 -2177 -495 -2173
rect -464 -2177 -460 -2173
rect -420 -2177 -416 -2173
rect -403 -2177 -399 -2173
rect -367 -2177 -363 -2173
rect -346 -2177 -342 -2173
rect -210 -2177 -206 -2173
rect -184 -2177 -180 -2173
rect -141 -2177 -137 -2173
rect -106 -2177 -102 -2173
rect -62 -2177 -58 -2173
rect -45 -2177 -41 -2173
rect -9 -2177 -5 -2173
rect 12 -2177 16 -2173
rect 218 -2177 222 -2173
rect 244 -2177 248 -2173
rect 287 -2177 291 -2173
rect 322 -2177 326 -2173
rect 366 -2177 370 -2173
rect 383 -2177 387 -2173
rect 419 -2177 423 -2173
rect 440 -2177 444 -2173
rect 574 -2177 578 -2173
rect 600 -2177 604 -2173
rect 643 -2177 647 -2173
rect 678 -2177 682 -2173
rect 722 -2177 726 -2173
rect 739 -2177 743 -2173
rect 775 -2177 779 -2173
rect 796 -2177 800 -2173
rect 972 -2177 976 -2173
rect 998 -2177 1002 -2173
rect 1041 -2177 1045 -2173
rect 1076 -2177 1080 -2173
rect 1120 -2177 1124 -2173
rect 1137 -2177 1141 -2173
rect 1173 -2177 1177 -2173
rect 1194 -2177 1198 -2173
rect 1330 -2177 1334 -2173
rect 1356 -2177 1360 -2173
rect 1399 -2177 1403 -2173
rect 1434 -2177 1438 -2173
rect 1478 -2177 1482 -2173
rect 1495 -2177 1499 -2173
rect 1531 -2177 1535 -2173
rect 1552 -2177 1556 -2173
rect 1633 -2177 1695 -2062
rect -1421 -2181 -1251 -2177
rect -1247 -2181 -1207 -2177
rect -1203 -2181 -1173 -2177
rect -1169 -2181 -926 -2177
rect -922 -2181 -900 -2177
rect -896 -2181 -857 -2177
rect -853 -2181 -822 -2177
rect -818 -2181 -778 -2177
rect -774 -2181 -761 -2177
rect -757 -2181 -725 -2177
rect -721 -2181 -704 -2177
rect -700 -2181 -568 -2177
rect -564 -2181 -542 -2177
rect -538 -2181 -499 -2177
rect -495 -2181 -464 -2177
rect -460 -2181 -420 -2177
rect -416 -2181 -403 -2177
rect -399 -2181 -367 -2177
rect -363 -2181 -346 -2177
rect -342 -2181 -210 -2177
rect -206 -2181 -184 -2177
rect -180 -2181 -141 -2177
rect -137 -2181 -106 -2177
rect -102 -2181 -62 -2177
rect -58 -2181 -45 -2177
rect -41 -2181 -9 -2177
rect -5 -2181 12 -2177
rect 16 -2181 218 -2177
rect 222 -2181 244 -2177
rect 248 -2181 287 -2177
rect 291 -2181 322 -2177
rect 326 -2181 366 -2177
rect 370 -2181 383 -2177
rect 387 -2181 419 -2177
rect 423 -2181 440 -2177
rect 444 -2181 574 -2177
rect 578 -2181 600 -2177
rect 604 -2181 643 -2177
rect 647 -2181 678 -2177
rect 682 -2181 722 -2177
rect 726 -2181 739 -2177
rect 743 -2181 775 -2177
rect 779 -2181 796 -2177
rect 800 -2181 972 -2177
rect 976 -2181 998 -2177
rect 1002 -2181 1041 -2177
rect 1045 -2181 1076 -2177
rect 1080 -2181 1120 -2177
rect 1124 -2181 1137 -2177
rect 1141 -2181 1173 -2177
rect 1177 -2181 1194 -2177
rect 1198 -2181 1330 -2177
rect 1334 -2181 1356 -2177
rect 1360 -2181 1399 -2177
rect 1403 -2181 1434 -2177
rect 1438 -2181 1478 -2177
rect 1482 -2181 1495 -2177
rect 1499 -2181 1531 -2177
rect 1535 -2181 1552 -2177
rect 1556 -2181 1695 -2177
rect -1272 -2188 -689 -2184
rect -585 -2188 27 -2184
rect 201 -2188 811 -2184
rect 955 -2188 1567 -2184
rect -1266 -2195 -1158 -2191
rect -943 -2195 -331 -2191
rect -227 -2195 455 -2191
rect 557 -2195 1209 -2191
rect 1313 -2195 1561 -2191
rect -1495 -2233 -1255 -2229
rect -1251 -2233 -1238 -2229
rect -1234 -2233 -1218 -2229
rect -1214 -2233 -1197 -2229
rect -1193 -2233 -1176 -2229
rect -1172 -2233 -1155 -2229
rect -1151 -2233 -1134 -2229
rect -1130 -2233 -1113 -2229
rect -1109 -2233 -1092 -2229
rect -1088 -2233 -1072 -2229
rect -1068 -2233 -926 -2229
rect -922 -2233 -909 -2229
rect -905 -2233 -889 -2229
rect -885 -2233 -868 -2229
rect -864 -2233 -847 -2229
rect -843 -2233 -826 -2229
rect -822 -2233 -805 -2229
rect -801 -2233 -784 -2229
rect -780 -2233 -763 -2229
rect -759 -2233 -743 -2229
rect -739 -2233 -568 -2229
rect -564 -2233 -551 -2229
rect -547 -2233 -531 -2229
rect -527 -2233 -510 -2229
rect -506 -2233 -489 -2229
rect -485 -2233 -468 -2229
rect -464 -2233 -447 -2229
rect -443 -2233 -426 -2229
rect -422 -2233 -405 -2229
rect -401 -2233 -385 -2229
rect -381 -2233 -210 -2229
rect -206 -2233 -193 -2229
rect -189 -2233 -173 -2229
rect -169 -2233 -152 -2229
rect -148 -2233 -131 -2229
rect -127 -2233 -110 -2229
rect -106 -2233 -89 -2229
rect -85 -2233 -68 -2229
rect -64 -2233 -47 -2229
rect -43 -2233 -27 -2229
rect -23 -2233 218 -2229
rect 222 -2233 235 -2229
rect 239 -2233 255 -2229
rect 259 -2233 276 -2229
rect 280 -2233 297 -2229
rect 301 -2233 318 -2229
rect 322 -2233 339 -2229
rect 343 -2233 360 -2229
rect 364 -2233 381 -2229
rect 385 -2233 401 -2229
rect 405 -2233 574 -2229
rect 578 -2233 591 -2229
rect 595 -2233 611 -2229
rect 615 -2233 632 -2229
rect 636 -2233 653 -2229
rect 657 -2233 674 -2229
rect 678 -2233 695 -2229
rect 699 -2233 716 -2229
rect 720 -2233 737 -2229
rect 741 -2233 757 -2229
rect 761 -2233 1617 -2229
rect -1495 -2360 -1433 -2233
rect -1233 -2281 -1199 -2277
rect -1135 -2281 -1115 -2277
rect -1100 -2281 -931 -2277
rect -904 -2281 -870 -2277
rect -806 -2281 -786 -2277
rect -771 -2281 -573 -2277
rect -546 -2281 -512 -2277
rect -448 -2281 -428 -2277
rect -413 -2281 -215 -2277
rect -188 -2281 -154 -2277
rect -90 -2281 -70 -2277
rect -55 -2281 213 -2277
rect 240 -2281 274 -2277
rect 338 -2281 358 -2277
rect 373 -2281 569 -2277
rect 596 -2281 630 -2277
rect 694 -2281 714 -2277
rect 729 -2281 765 -2277
rect -935 -2285 -931 -2281
rect -577 -2285 -573 -2281
rect -219 -2285 -215 -2281
rect 209 -2285 213 -2281
rect 565 -2285 569 -2281
rect -1266 -2289 -1257 -2285
rect -1253 -2289 -1223 -2285
rect -1202 -2289 -1171 -2285
rect -1142 -2289 -1111 -2285
rect -1100 -2289 -1073 -2285
rect -935 -2289 -928 -2285
rect -924 -2289 -894 -2285
rect -873 -2289 -842 -2285
rect -813 -2289 -782 -2285
rect -771 -2289 -744 -2285
rect -577 -2289 -570 -2285
rect -566 -2289 -536 -2285
rect -515 -2289 -484 -2285
rect -455 -2289 -424 -2285
rect -413 -2289 -386 -2285
rect -219 -2289 -212 -2285
rect -208 -2289 -178 -2285
rect -157 -2289 -126 -2285
rect -97 -2289 -66 -2285
rect -55 -2289 -28 -2285
rect 209 -2289 216 -2285
rect 220 -2289 250 -2285
rect 271 -2289 302 -2285
rect 331 -2289 362 -2285
rect 373 -2289 400 -2285
rect 565 -2289 572 -2285
rect 576 -2289 606 -2285
rect 627 -2289 658 -2285
rect 687 -2289 718 -2285
rect 729 -2289 756 -2285
rect -1260 -2296 -1213 -2292
rect -1177 -2296 -1164 -2292
rect -1160 -2296 -1129 -2292
rect -1093 -2296 -1080 -2292
rect -1076 -2296 -1064 -2292
rect -931 -2296 -884 -2292
rect -848 -2296 -835 -2292
rect -831 -2296 -800 -2292
rect -764 -2296 -751 -2292
rect -747 -2296 -735 -2292
rect -573 -2296 -526 -2292
rect -490 -2296 -477 -2292
rect -473 -2296 -442 -2292
rect -406 -2296 -393 -2292
rect -389 -2296 -377 -2292
rect -215 -2296 -168 -2292
rect -132 -2296 -119 -2292
rect -115 -2296 -84 -2292
rect -48 -2296 -35 -2292
rect -31 -2296 -19 -2292
rect 213 -2296 260 -2292
rect 296 -2296 309 -2292
rect 313 -2296 344 -2292
rect 380 -2296 393 -2292
rect 397 -2296 409 -2292
rect 569 -2296 616 -2292
rect 652 -2296 665 -2292
rect 669 -2296 700 -2292
rect 736 -2296 749 -2292
rect 753 -2296 765 -2292
rect -1280 -2303 -1253 -2299
rect -1249 -2303 -1139 -2299
rect -1118 -2303 -1087 -2299
rect -950 -2303 -924 -2299
rect -920 -2303 -810 -2299
rect -789 -2303 -758 -2299
rect -591 -2303 -566 -2299
rect -562 -2303 -452 -2299
rect -431 -2303 -400 -2299
rect -235 -2303 -208 -2299
rect -204 -2303 -94 -2299
rect -73 -2303 -42 -2299
rect 196 -2303 220 -2299
rect 224 -2303 334 -2299
rect 355 -2303 386 -2299
rect 547 -2303 576 -2299
rect 580 -2303 690 -2299
rect 711 -2303 742 -2299
rect -1218 -2310 -1195 -2306
rect -1176 -2310 -1157 -2306
rect -889 -2310 -866 -2306
rect -847 -2310 -828 -2306
rect -531 -2310 -508 -2306
rect -489 -2310 -470 -2306
rect -173 -2310 -150 -2306
rect -131 -2310 -112 -2306
rect 255 -2310 278 -2306
rect 297 -2310 316 -2306
rect 611 -2310 634 -2306
rect 653 -2310 672 -2306
rect 1633 -2321 1695 -2181
rect -1421 -2325 -1255 -2321
rect -1251 -2325 -1238 -2321
rect -1234 -2325 -1197 -2321
rect -1193 -2325 -1155 -2321
rect -1151 -2325 -1113 -2321
rect -1109 -2325 -1072 -2321
rect -1068 -2325 -926 -2321
rect -922 -2325 -909 -2321
rect -905 -2325 -868 -2321
rect -864 -2325 -826 -2321
rect -822 -2325 -784 -2321
rect -780 -2325 -743 -2321
rect -739 -2325 -568 -2321
rect -564 -2325 -551 -2321
rect -547 -2325 -510 -2321
rect -506 -2325 -468 -2321
rect -464 -2325 -426 -2321
rect -422 -2325 -385 -2321
rect -381 -2325 -210 -2321
rect -206 -2325 -193 -2321
rect -189 -2325 -152 -2321
rect -148 -2325 -110 -2321
rect -106 -2325 -68 -2321
rect -64 -2325 -27 -2321
rect -23 -2325 218 -2321
rect 222 -2325 235 -2321
rect 239 -2325 276 -2321
rect 280 -2325 318 -2321
rect 322 -2325 360 -2321
rect 364 -2325 401 -2321
rect 405 -2325 574 -2321
rect 578 -2325 591 -2321
rect 595 -2325 632 -2321
rect 636 -2325 674 -2321
rect 678 -2325 716 -2321
rect 720 -2325 757 -2321
rect 761 -2325 1695 -2321
rect -1495 -2364 -1255 -2360
rect -1251 -2364 -1238 -2360
rect -1234 -2364 -1218 -2360
rect -1214 -2364 -1197 -2360
rect -1193 -2364 -1176 -2360
rect -1172 -2364 -1155 -2360
rect -1151 -2364 -1134 -2360
rect -1130 -2364 -1113 -2360
rect -1109 -2364 -1092 -2360
rect -1088 -2364 -1072 -2360
rect -1068 -2364 -926 -2360
rect -922 -2364 -909 -2360
rect -905 -2364 -889 -2360
rect -885 -2364 -868 -2360
rect -864 -2364 -847 -2360
rect -843 -2364 -826 -2360
rect -822 -2364 -805 -2360
rect -801 -2364 -784 -2360
rect -780 -2364 -763 -2360
rect -759 -2364 -743 -2360
rect -739 -2364 -568 -2360
rect -564 -2364 -551 -2360
rect -547 -2364 -531 -2360
rect -527 -2364 -510 -2360
rect -506 -2364 -489 -2360
rect -485 -2364 -468 -2360
rect -464 -2364 -447 -2360
rect -443 -2364 -426 -2360
rect -422 -2364 -405 -2360
rect -401 -2364 -385 -2360
rect -381 -2364 -210 -2360
rect -206 -2364 -193 -2360
rect -189 -2364 -173 -2360
rect -169 -2364 -152 -2360
rect -148 -2364 -131 -2360
rect -127 -2364 -110 -2360
rect -106 -2364 -89 -2360
rect -85 -2364 -68 -2360
rect -64 -2364 -47 -2360
rect -43 -2364 -27 -2360
rect -23 -2364 218 -2360
rect 222 -2364 235 -2360
rect 239 -2364 255 -2360
rect 259 -2364 276 -2360
rect 280 -2364 297 -2360
rect 301 -2364 318 -2360
rect 322 -2364 339 -2360
rect 343 -2364 360 -2360
rect 364 -2364 381 -2360
rect 385 -2364 401 -2360
rect 405 -2364 574 -2360
rect 578 -2364 591 -2360
rect 595 -2364 611 -2360
rect 615 -2364 632 -2360
rect 636 -2364 653 -2360
rect 657 -2364 674 -2360
rect 678 -2364 695 -2360
rect 699 -2364 716 -2360
rect 720 -2364 737 -2360
rect 741 -2364 757 -2360
rect 761 -2364 972 -2360
rect 976 -2364 989 -2360
rect 993 -2364 1009 -2360
rect 1013 -2364 1030 -2360
rect 1034 -2364 1051 -2360
rect 1055 -2364 1072 -2360
rect 1076 -2364 1093 -2360
rect 1097 -2364 1114 -2360
rect 1118 -2364 1135 -2360
rect 1139 -2364 1155 -2360
rect 1159 -2364 1330 -2360
rect 1334 -2364 1347 -2360
rect 1351 -2364 1367 -2360
rect 1371 -2364 1388 -2360
rect 1392 -2364 1409 -2360
rect 1413 -2364 1430 -2360
rect 1434 -2364 1451 -2360
rect 1455 -2364 1472 -2360
rect 1476 -2364 1493 -2360
rect 1497 -2364 1513 -2360
rect 1517 -2364 1617 -2360
rect -1495 -2491 -1433 -2364
rect -1233 -2412 -1199 -2408
rect -1135 -2412 -1115 -2408
rect -1100 -2412 -1066 -2408
rect -904 -2412 -870 -2408
rect -806 -2412 -786 -2408
rect -771 -2412 -737 -2408
rect -546 -2412 -512 -2408
rect -448 -2412 -428 -2408
rect -413 -2412 -379 -2408
rect -188 -2412 -154 -2408
rect -90 -2412 -70 -2408
rect -55 -2412 -21 -2408
rect 240 -2412 274 -2408
rect 338 -2412 358 -2408
rect 373 -2412 407 -2408
rect 596 -2412 630 -2408
rect 694 -2412 714 -2408
rect 729 -2412 763 -2408
rect 994 -2412 1028 -2408
rect 1092 -2412 1112 -2408
rect 1127 -2412 1161 -2408
rect 1352 -2412 1386 -2408
rect 1450 -2412 1470 -2408
rect 1485 -2412 1519 -2408
rect -1272 -2420 -1257 -2416
rect -1253 -2420 -1223 -2416
rect -1202 -2420 -1171 -2416
rect -1142 -2420 -1111 -2416
rect -1100 -2420 -1073 -2416
rect -943 -2420 -928 -2416
rect -924 -2420 -894 -2416
rect -873 -2420 -842 -2416
rect -813 -2420 -782 -2416
rect -771 -2420 -744 -2416
rect -585 -2420 -570 -2416
rect -566 -2420 -536 -2416
rect -515 -2420 -484 -2416
rect -455 -2420 -424 -2416
rect -413 -2420 -386 -2416
rect -227 -2420 -212 -2416
rect -208 -2420 -178 -2416
rect -157 -2420 -126 -2416
rect -97 -2420 -66 -2416
rect -55 -2420 -28 -2416
rect 201 -2420 216 -2416
rect 220 -2420 250 -2416
rect 271 -2420 302 -2416
rect 331 -2420 362 -2416
rect 373 -2420 400 -2416
rect 557 -2420 572 -2416
rect 576 -2420 606 -2416
rect 627 -2420 658 -2416
rect 687 -2420 718 -2416
rect 729 -2420 756 -2416
rect 955 -2420 970 -2416
rect 974 -2420 1004 -2416
rect 1025 -2420 1056 -2416
rect 1085 -2420 1116 -2416
rect 1127 -2420 1154 -2416
rect 1313 -2420 1328 -2416
rect 1332 -2420 1362 -2416
rect 1383 -2420 1414 -2416
rect 1443 -2420 1474 -2416
rect 1485 -2420 1512 -2416
rect -1260 -2427 -1213 -2423
rect -1177 -2427 -1164 -2423
rect -1160 -2427 -1129 -2423
rect -1093 -2427 -1080 -2423
rect -1076 -2427 -1064 -2423
rect -931 -2427 -884 -2423
rect -848 -2427 -835 -2423
rect -831 -2427 -800 -2423
rect -764 -2427 -751 -2423
rect -747 -2427 -735 -2423
rect -573 -2427 -526 -2423
rect -490 -2427 -477 -2423
rect -473 -2427 -442 -2423
rect -406 -2427 -393 -2423
rect -389 -2427 -377 -2423
rect -215 -2427 -168 -2423
rect -132 -2427 -119 -2423
rect -115 -2427 -84 -2423
rect -48 -2427 -35 -2423
rect -31 -2427 -19 -2423
rect 213 -2427 260 -2423
rect 296 -2427 309 -2423
rect 313 -2427 344 -2423
rect 380 -2427 393 -2423
rect 397 -2427 409 -2423
rect 569 -2427 616 -2423
rect 652 -2427 665 -2423
rect 669 -2427 700 -2423
rect 736 -2427 749 -2423
rect 753 -2427 765 -2423
rect 967 -2427 1014 -2423
rect 1050 -2427 1063 -2423
rect 1067 -2427 1098 -2423
rect 1134 -2427 1147 -2423
rect 1151 -2427 1163 -2423
rect 1325 -2427 1372 -2423
rect 1408 -2427 1421 -2423
rect 1425 -2427 1456 -2423
rect 1492 -2427 1505 -2423
rect 1509 -2427 1521 -2423
rect -1285 -2434 -1284 -2430
rect -1280 -2434 -1253 -2430
rect -1249 -2434 -1139 -2430
rect -1118 -2434 -1087 -2430
rect -950 -2434 -924 -2430
rect -920 -2434 -810 -2430
rect -789 -2434 -758 -2430
rect -591 -2434 -566 -2430
rect -562 -2434 -452 -2430
rect -431 -2434 -400 -2430
rect -235 -2434 -208 -2430
rect -204 -2434 -94 -2430
rect -73 -2434 -42 -2430
rect 196 -2434 220 -2430
rect 224 -2434 334 -2430
rect 355 -2434 386 -2430
rect 547 -2434 576 -2430
rect 580 -2434 690 -2430
rect 711 -2434 742 -2430
rect 954 -2434 974 -2430
rect 978 -2434 1088 -2430
rect 1109 -2434 1140 -2430
rect 1306 -2434 1332 -2430
rect 1336 -2434 1446 -2430
rect 1467 -2434 1498 -2430
rect -1218 -2441 -1195 -2437
rect -1176 -2441 -1157 -2437
rect -889 -2441 -866 -2437
rect -847 -2441 -828 -2437
rect -531 -2441 -508 -2437
rect -489 -2441 -470 -2437
rect -173 -2441 -150 -2437
rect -131 -2441 -112 -2437
rect 255 -2441 278 -2437
rect 297 -2441 316 -2437
rect 611 -2441 634 -2437
rect 653 -2441 672 -2437
rect 1009 -2441 1032 -2437
rect 1051 -2441 1070 -2437
rect 1367 -2441 1390 -2437
rect 1409 -2441 1428 -2437
rect 1633 -2452 1695 -2325
rect -1421 -2456 -1255 -2452
rect -1251 -2456 -1238 -2452
rect -1234 -2456 -1197 -2452
rect -1193 -2456 -1155 -2452
rect -1151 -2456 -1113 -2452
rect -1109 -2456 -1072 -2452
rect -1068 -2456 -926 -2452
rect -922 -2456 -909 -2452
rect -905 -2456 -868 -2452
rect -864 -2456 -826 -2452
rect -822 -2456 -784 -2452
rect -780 -2456 -743 -2452
rect -739 -2456 -568 -2452
rect -564 -2456 -551 -2452
rect -547 -2456 -510 -2452
rect -506 -2456 -468 -2452
rect -464 -2456 -426 -2452
rect -422 -2456 -385 -2452
rect -381 -2456 -210 -2452
rect -206 -2456 -193 -2452
rect -189 -2456 -152 -2452
rect -148 -2456 -110 -2452
rect -106 -2456 -68 -2452
rect -64 -2456 -27 -2452
rect -23 -2456 218 -2452
rect 222 -2456 235 -2452
rect 239 -2456 276 -2452
rect 280 -2456 318 -2452
rect 322 -2456 360 -2452
rect 364 -2456 401 -2452
rect 405 -2456 574 -2452
rect 578 -2456 591 -2452
rect 595 -2456 632 -2452
rect 636 -2456 674 -2452
rect 678 -2456 716 -2452
rect 720 -2456 757 -2452
rect 761 -2456 972 -2452
rect 976 -2456 989 -2452
rect 993 -2456 1030 -2452
rect 1034 -2456 1072 -2452
rect 1076 -2456 1114 -2452
rect 1118 -2456 1155 -2452
rect 1159 -2456 1330 -2452
rect 1334 -2456 1347 -2452
rect 1351 -2456 1388 -2452
rect 1392 -2456 1430 -2452
rect 1434 -2456 1472 -2452
rect 1476 -2456 1513 -2452
rect 1517 -2456 1695 -2452
rect -1266 -2464 -1066 -2460
rect -943 -2463 -737 -2459
rect -585 -2464 -379 -2460
rect -227 -2464 -21 -2460
rect 201 -2463 407 -2459
rect 557 -2463 763 -2459
rect 955 -2464 1161 -2460
rect 1313 -2464 1519 -2460
rect -1495 -2495 -1255 -2491
rect -1251 -2495 -1238 -2491
rect -1234 -2495 -1218 -2491
rect -1214 -2495 -1197 -2491
rect -1193 -2495 -1176 -2491
rect -1172 -2495 -1155 -2491
rect -1151 -2495 -1134 -2491
rect -1130 -2495 -1113 -2491
rect -1109 -2495 -1092 -2491
rect -1088 -2495 -1072 -2491
rect -1068 -2495 -926 -2491
rect -922 -2495 -909 -2491
rect -905 -2495 -889 -2491
rect -885 -2495 -868 -2491
rect -864 -2495 -847 -2491
rect -843 -2495 -826 -2491
rect -822 -2495 -805 -2491
rect -801 -2495 -784 -2491
rect -780 -2495 -763 -2491
rect -759 -2495 -743 -2491
rect -739 -2495 -568 -2491
rect -564 -2495 -551 -2491
rect -547 -2495 -531 -2491
rect -527 -2495 -510 -2491
rect -506 -2495 -489 -2491
rect -485 -2495 -468 -2491
rect -464 -2495 -447 -2491
rect -443 -2495 -426 -2491
rect -422 -2495 -405 -2491
rect -401 -2495 -385 -2491
rect -381 -2495 -210 -2491
rect -206 -2495 -193 -2491
rect -189 -2495 -173 -2491
rect -169 -2495 -152 -2491
rect -148 -2495 -131 -2491
rect -127 -2495 -110 -2491
rect -106 -2495 -89 -2491
rect -85 -2495 -68 -2491
rect -64 -2495 -47 -2491
rect -43 -2495 -27 -2491
rect -23 -2495 90 -2491
rect 94 -2495 218 -2491
rect 222 -2495 235 -2491
rect 239 -2495 255 -2491
rect 259 -2495 276 -2491
rect 280 -2495 297 -2491
rect 301 -2495 318 -2491
rect 322 -2495 339 -2491
rect 343 -2495 360 -2491
rect 364 -2495 381 -2491
rect 385 -2495 401 -2491
rect 405 -2495 574 -2491
rect 578 -2495 591 -2491
rect 595 -2495 611 -2491
rect 615 -2495 632 -2491
rect 636 -2495 653 -2491
rect 657 -2495 674 -2491
rect 678 -2495 695 -2491
rect 699 -2495 716 -2491
rect 720 -2495 737 -2491
rect 741 -2495 757 -2491
rect 761 -2495 972 -2491
rect 976 -2495 989 -2491
rect 993 -2495 1009 -2491
rect 1013 -2495 1030 -2491
rect 1034 -2495 1051 -2491
rect 1055 -2495 1072 -2491
rect 1076 -2495 1093 -2491
rect 1097 -2495 1114 -2491
rect 1118 -2495 1135 -2491
rect 1139 -2495 1155 -2491
rect 1159 -2495 1330 -2491
rect 1334 -2495 1347 -2491
rect 1351 -2495 1367 -2491
rect 1371 -2495 1388 -2491
rect 1392 -2495 1409 -2491
rect 1413 -2495 1430 -2491
rect 1434 -2495 1451 -2491
rect 1455 -2495 1472 -2491
rect 1476 -2495 1493 -2491
rect 1497 -2495 1513 -2491
rect 1517 -2495 1617 -2491
rect -1495 -2603 -1433 -2495
rect -1233 -2543 -1199 -2539
rect -1135 -2543 -1115 -2539
rect -1100 -2543 -1066 -2539
rect -904 -2543 -870 -2539
rect -806 -2543 -786 -2539
rect -771 -2543 -731 -2539
rect -546 -2543 -512 -2539
rect -448 -2543 -428 -2539
rect -413 -2543 -379 -2539
rect -188 -2543 -154 -2539
rect -90 -2543 -70 -2539
rect -55 -2543 -21 -2539
rect -1345 -2551 -1257 -2547
rect -1253 -2551 -1223 -2547
rect -1202 -2551 -1171 -2547
rect -1142 -2551 -1111 -2547
rect -1100 -2551 -1073 -2547
rect -937 -2551 -928 -2547
rect -924 -2551 -894 -2547
rect -873 -2551 -842 -2547
rect -813 -2551 -782 -2547
rect -771 -2551 -744 -2547
rect -579 -2551 -570 -2547
rect -566 -2551 -536 -2547
rect -515 -2551 -484 -2547
rect -455 -2551 -424 -2547
rect -413 -2551 -386 -2547
rect -221 -2551 -212 -2547
rect -208 -2551 -178 -2547
rect -157 -2551 -126 -2547
rect -97 -2551 -66 -2547
rect -55 -2551 -28 -2547
rect 102 -2546 106 -2542
rect 240 -2543 274 -2539
rect 338 -2543 358 -2539
rect 373 -2543 407 -2539
rect 596 -2543 630 -2539
rect 694 -2543 714 -2539
rect 729 -2543 763 -2539
rect 994 -2543 1028 -2539
rect 1092 -2543 1112 -2539
rect 1127 -2543 1161 -2539
rect 1352 -2543 1386 -2539
rect 1450 -2543 1470 -2539
rect 1485 -2543 1519 -2539
rect 207 -2551 216 -2547
rect 220 -2551 250 -2547
rect 271 -2551 302 -2547
rect 331 -2551 362 -2547
rect 373 -2551 400 -2547
rect 563 -2551 572 -2547
rect 576 -2551 606 -2547
rect 627 -2551 658 -2547
rect 687 -2551 718 -2547
rect 729 -2551 756 -2547
rect 961 -2551 970 -2547
rect 974 -2551 1004 -2547
rect 1025 -2551 1056 -2547
rect 1085 -2551 1116 -2547
rect 1127 -2551 1154 -2547
rect 1319 -2551 1328 -2547
rect 1332 -2551 1362 -2547
rect 1383 -2551 1414 -2547
rect 1443 -2551 1474 -2547
rect 1485 -2551 1512 -2547
rect -1260 -2558 -1213 -2554
rect -1177 -2558 -1164 -2554
rect -1160 -2558 -1129 -2554
rect -1093 -2558 -1080 -2554
rect -1076 -2558 -1064 -2554
rect -931 -2558 -884 -2554
rect -848 -2558 -835 -2554
rect -831 -2558 -800 -2554
rect -764 -2558 -751 -2554
rect -747 -2558 -735 -2554
rect -573 -2558 -526 -2554
rect -490 -2558 -477 -2554
rect -473 -2558 -442 -2554
rect -406 -2558 -393 -2554
rect -389 -2558 -377 -2554
rect -215 -2558 -168 -2554
rect -132 -2558 -119 -2554
rect -115 -2558 -84 -2554
rect -48 -2558 -35 -2554
rect -31 -2558 -19 -2554
rect 213 -2558 260 -2554
rect 296 -2558 309 -2554
rect 313 -2558 344 -2554
rect 380 -2558 393 -2554
rect 397 -2558 409 -2554
rect 569 -2558 616 -2554
rect 652 -2558 665 -2554
rect 669 -2558 700 -2554
rect 736 -2558 749 -2554
rect 753 -2558 765 -2554
rect 967 -2558 1014 -2554
rect 1050 -2558 1063 -2554
rect 1067 -2558 1098 -2554
rect 1134 -2558 1147 -2554
rect 1151 -2558 1163 -2554
rect 1325 -2558 1372 -2554
rect 1408 -2558 1421 -2554
rect 1425 -2558 1456 -2554
rect 1492 -2558 1505 -2554
rect 1509 -2558 1521 -2554
rect -1271 -2565 -1253 -2561
rect -1249 -2565 -1139 -2561
rect -1118 -2565 -1087 -2561
rect -938 -2565 -924 -2561
rect -920 -2565 -810 -2561
rect -789 -2565 -758 -2561
rect -582 -2565 -566 -2561
rect -562 -2565 -452 -2561
rect -431 -2565 -400 -2561
rect -224 -2565 -208 -2561
rect -204 -2565 -94 -2561
rect -73 -2565 -42 -2561
rect 202 -2565 220 -2561
rect 224 -2565 334 -2561
rect 355 -2565 386 -2561
rect 560 -2565 576 -2561
rect 580 -2565 690 -2561
rect 711 -2565 742 -2561
rect 948 -2565 974 -2561
rect 978 -2565 1088 -2561
rect 1109 -2565 1140 -2561
rect 1312 -2565 1313 -2561
rect 1317 -2565 1332 -2561
rect 1336 -2565 1446 -2561
rect 1467 -2565 1498 -2561
rect -1218 -2572 -1195 -2568
rect -1176 -2572 -1157 -2568
rect -889 -2572 -866 -2568
rect -847 -2572 -828 -2568
rect -531 -2572 -508 -2568
rect -489 -2572 -470 -2568
rect -173 -2572 -150 -2568
rect -131 -2572 -112 -2568
rect 255 -2572 278 -2568
rect 297 -2572 316 -2568
rect 611 -2572 634 -2568
rect 653 -2572 672 -2568
rect 1009 -2572 1032 -2568
rect 1051 -2572 1070 -2568
rect 1367 -2572 1390 -2568
rect 1409 -2572 1428 -2568
rect 1633 -2583 1695 -2456
rect -1421 -2587 -1255 -2583
rect -1251 -2587 -1238 -2583
rect -1234 -2587 -1197 -2583
rect -1193 -2587 -1155 -2583
rect -1151 -2587 -1113 -2583
rect -1109 -2587 -1072 -2583
rect -1068 -2587 -926 -2583
rect -922 -2587 -909 -2583
rect -905 -2587 -868 -2583
rect -864 -2587 -826 -2583
rect -822 -2587 -784 -2583
rect -780 -2587 -743 -2583
rect -739 -2587 -568 -2583
rect -564 -2587 -551 -2583
rect -547 -2587 -510 -2583
rect -506 -2587 -468 -2583
rect -464 -2587 -426 -2583
rect -422 -2587 -385 -2583
rect -381 -2587 -210 -2583
rect -206 -2587 -193 -2583
rect -189 -2587 -152 -2583
rect -148 -2587 -110 -2583
rect -106 -2587 -68 -2583
rect -64 -2587 -27 -2583
rect -23 -2587 90 -2583
rect 94 -2587 218 -2583
rect 222 -2587 235 -2583
rect 239 -2587 276 -2583
rect 280 -2587 318 -2583
rect 322 -2587 360 -2583
rect 364 -2587 401 -2583
rect 405 -2587 574 -2583
rect 578 -2587 591 -2583
rect 595 -2587 632 -2583
rect 636 -2587 674 -2583
rect 678 -2587 716 -2583
rect 720 -2587 757 -2583
rect 761 -2587 972 -2583
rect 976 -2587 989 -2583
rect 993 -2587 1030 -2583
rect 1034 -2587 1072 -2583
rect 1076 -2587 1114 -2583
rect 1118 -2587 1155 -2583
rect 1159 -2587 1330 -2583
rect 1334 -2587 1347 -2583
rect 1351 -2587 1388 -2583
rect 1392 -2587 1430 -2583
rect 1434 -2587 1472 -2583
rect 1476 -2587 1513 -2583
rect 1517 -2587 1695 -2583
rect -1495 -2607 -1255 -2603
rect -1251 -2607 -1238 -2603
rect -1234 -2607 -1218 -2603
rect -1214 -2607 -1197 -2603
rect -1193 -2607 -1176 -2603
rect -1172 -2607 -1155 -2603
rect -1151 -2607 -1134 -2603
rect -1130 -2607 -1113 -2603
rect -1109 -2607 -1092 -2603
rect -1088 -2607 -1072 -2603
rect -1068 -2607 -926 -2603
rect -922 -2607 -909 -2603
rect -905 -2607 -889 -2603
rect -885 -2607 -868 -2603
rect -864 -2607 -847 -2603
rect -843 -2607 -826 -2603
rect -822 -2607 -805 -2603
rect -801 -2607 -784 -2603
rect -780 -2607 -763 -2603
rect -759 -2607 -743 -2603
rect -739 -2607 1617 -2603
rect -1495 -2716 -1433 -2607
rect -1233 -2655 -1199 -2651
rect -1135 -2655 -1115 -2651
rect -1100 -2655 -931 -2651
rect -904 -2655 -870 -2651
rect -806 -2655 -786 -2651
rect -771 -2655 -737 -2651
rect -935 -2659 -931 -2655
rect -1421 -2663 -1257 -2659
rect -1253 -2663 -1223 -2659
rect -1202 -2663 -1171 -2659
rect -1142 -2663 -1111 -2659
rect -1100 -2663 -1073 -2659
rect -935 -2663 -928 -2659
rect -924 -2663 -894 -2659
rect -873 -2663 -842 -2659
rect -813 -2663 -782 -2659
rect -771 -2663 -744 -2659
rect -1260 -2670 -1213 -2666
rect -1177 -2670 -1164 -2666
rect -1160 -2670 -1129 -2666
rect -1093 -2670 -1080 -2666
rect -1076 -2670 -1064 -2666
rect -931 -2670 -884 -2666
rect -848 -2670 -835 -2666
rect -831 -2670 -800 -2666
rect -764 -2670 -751 -2666
rect -747 -2670 -735 -2666
rect -1271 -2677 -1253 -2673
rect -1249 -2677 -1139 -2673
rect -1118 -2677 -1087 -2673
rect -938 -2677 -924 -2673
rect -920 -2677 -810 -2673
rect -789 -2677 -758 -2673
rect -1218 -2684 -1195 -2680
rect -1176 -2684 -1157 -2680
rect -889 -2684 -866 -2680
rect -847 -2684 -828 -2680
rect 1633 -2695 1695 -2587
rect -1421 -2699 -1255 -2695
rect -1251 -2699 -1238 -2695
rect -1234 -2699 -1197 -2695
rect -1193 -2699 -1155 -2695
rect -1151 -2699 -1113 -2695
rect -1109 -2699 -1072 -2695
rect -1068 -2699 -926 -2695
rect -922 -2699 -909 -2695
rect -905 -2699 -868 -2695
rect -864 -2699 -826 -2695
rect -822 -2699 -784 -2695
rect -780 -2699 -743 -2695
rect -739 -2699 1695 -2695
rect -1495 -2720 -1339 -2716
rect -1335 -2720 -1322 -2716
rect -1318 -2720 -935 -2716
rect -931 -2720 -918 -2716
rect -914 -2720 -577 -2716
rect -573 -2720 -560 -2716
rect -556 -2720 -219 -2716
rect -215 -2720 -202 -2716
rect -198 -2720 209 -2716
rect 213 -2720 226 -2716
rect 230 -2720 565 -2716
rect 569 -2720 582 -2716
rect 586 -2720 963 -2716
rect 967 -2720 980 -2716
rect 984 -2720 1321 -2716
rect 1325 -2720 1338 -2716
rect 1342 -2720 1617 -2716
rect -1495 -2835 -1433 -2720
rect -1334 -2752 -1066 -2748
rect -930 -2752 -731 -2748
rect -572 -2752 -379 -2748
rect -214 -2752 -21 -2748
rect 214 -2752 407 -2748
rect 570 -2752 763 -2748
rect 968 -2752 1161 -2748
rect 1326 -2752 1519 -2748
rect -1323 -2760 -923 -2756
rect -919 -2760 -737 -2756
rect -733 -2760 -565 -2756
rect -561 -2760 -207 -2756
rect -203 -2760 221 -2756
rect 225 -2760 577 -2756
rect 581 -2760 975 -2756
rect 979 -2760 1333 -2756
rect 1337 -2760 1617 -2756
rect -949 -2773 -909 -2769
rect -591 -2773 -551 -2769
rect -233 -2773 -193 -2769
rect 195 -2773 235 -2769
rect 551 -2773 591 -2769
rect 949 -2773 989 -2769
rect 1307 -2773 1347 -2769
rect 1633 -2808 1695 -2699
rect -1421 -2812 -1322 -2808
rect -1318 -2812 -918 -2808
rect -914 -2812 -560 -2808
rect -556 -2812 -202 -2808
rect -198 -2812 226 -2808
rect 230 -2812 582 -2808
rect 586 -2812 980 -2808
rect 984 -2812 1338 -2808
rect 1342 -2812 1695 -2808
rect -1495 -2839 -1255 -2835
rect -1251 -2839 -1238 -2835
rect -1234 -2839 -1198 -2835
rect -1194 -2839 -1177 -2835
rect -1173 -2839 -926 -2835
rect -922 -2839 -900 -2835
rect -896 -2839 -883 -2835
rect -879 -2839 -843 -2835
rect -839 -2839 -822 -2835
rect -818 -2839 -805 -2835
rect -801 -2839 -765 -2835
rect -761 -2839 -741 -2835
rect -737 -2839 -704 -2835
rect -700 -2839 -568 -2835
rect -564 -2839 -542 -2835
rect -538 -2839 -525 -2835
rect -521 -2839 -485 -2835
rect -481 -2839 -464 -2835
rect -460 -2839 -447 -2835
rect -443 -2839 -407 -2835
rect -403 -2839 -383 -2835
rect -379 -2839 -346 -2835
rect -342 -2839 -210 -2835
rect -206 -2839 -184 -2835
rect -180 -2839 -167 -2835
rect -163 -2839 -127 -2835
rect -123 -2839 -106 -2835
rect -102 -2839 -89 -2835
rect -85 -2839 -49 -2835
rect -45 -2839 -25 -2835
rect -21 -2839 12 -2835
rect 16 -2839 218 -2835
rect 222 -2839 244 -2835
rect 248 -2839 261 -2835
rect 265 -2839 301 -2835
rect 305 -2839 322 -2835
rect 326 -2839 339 -2835
rect 343 -2839 379 -2835
rect 383 -2839 403 -2835
rect 407 -2839 440 -2835
rect 444 -2839 574 -2835
rect 578 -2839 600 -2835
rect 604 -2839 617 -2835
rect 621 -2839 657 -2835
rect 661 -2839 678 -2835
rect 682 -2839 695 -2835
rect 699 -2839 735 -2835
rect 739 -2839 759 -2835
rect 763 -2839 796 -2835
rect 800 -2839 972 -2835
rect 976 -2839 998 -2835
rect 1002 -2839 1015 -2835
rect 1019 -2839 1055 -2835
rect 1059 -2839 1076 -2835
rect 1080 -2839 1093 -2835
rect 1097 -2839 1133 -2835
rect 1137 -2839 1157 -2835
rect 1161 -2839 1194 -2835
rect 1198 -2839 1330 -2835
rect 1334 -2839 1356 -2835
rect 1360 -2839 1373 -2835
rect 1377 -2839 1413 -2835
rect 1417 -2839 1434 -2835
rect 1438 -2839 1451 -2835
rect 1455 -2839 1491 -2835
rect 1495 -2839 1515 -2835
rect 1519 -2839 1552 -2835
rect 1556 -2839 1617 -2835
rect -1495 -2954 -1433 -2839
rect -926 -2843 -922 -2839
rect -900 -2843 -896 -2839
rect -883 -2843 -879 -2839
rect -843 -2843 -839 -2839
rect -822 -2843 -818 -2839
rect -805 -2843 -801 -2839
rect -765 -2843 -761 -2839
rect -741 -2843 -737 -2839
rect -704 -2843 -700 -2839
rect -568 -2843 -564 -2839
rect -542 -2843 -538 -2839
rect -525 -2843 -521 -2839
rect -485 -2843 -481 -2839
rect -464 -2843 -460 -2839
rect -447 -2843 -443 -2839
rect -407 -2843 -403 -2839
rect -383 -2843 -379 -2839
rect -346 -2843 -342 -2839
rect -210 -2843 -206 -2839
rect -184 -2843 -180 -2839
rect -167 -2843 -163 -2839
rect -127 -2843 -123 -2839
rect -106 -2843 -102 -2839
rect -89 -2843 -85 -2839
rect -49 -2843 -45 -2839
rect -25 -2843 -21 -2839
rect 12 -2843 16 -2839
rect 218 -2843 222 -2839
rect 244 -2843 248 -2839
rect 261 -2843 265 -2839
rect 301 -2843 305 -2839
rect 322 -2843 326 -2839
rect 339 -2843 343 -2839
rect 379 -2843 383 -2839
rect 403 -2843 407 -2839
rect 440 -2843 444 -2839
rect 574 -2843 578 -2839
rect 600 -2843 604 -2839
rect 617 -2843 621 -2839
rect 657 -2843 661 -2839
rect 678 -2843 682 -2839
rect 695 -2843 699 -2839
rect 735 -2843 739 -2839
rect 759 -2843 763 -2839
rect 796 -2843 800 -2839
rect 972 -2843 976 -2839
rect 998 -2843 1002 -2839
rect 1015 -2843 1019 -2839
rect 1055 -2843 1059 -2839
rect 1076 -2843 1080 -2839
rect 1093 -2843 1097 -2839
rect 1133 -2843 1137 -2839
rect 1157 -2843 1161 -2839
rect 1194 -2843 1198 -2839
rect 1330 -2843 1334 -2839
rect 1356 -2843 1360 -2839
rect 1373 -2843 1377 -2839
rect 1413 -2843 1417 -2839
rect 1434 -2843 1438 -2839
rect 1451 -2843 1455 -2839
rect 1491 -2843 1495 -2839
rect 1515 -2843 1519 -2839
rect 1552 -2843 1556 -2839
rect -920 -2858 -858 -2854
rect -854 -2858 -824 -2854
rect -776 -2858 -746 -2854
rect -562 -2858 -500 -2854
rect -496 -2858 -466 -2854
rect -418 -2858 -388 -2854
rect -204 -2858 -142 -2854
rect -138 -2858 -108 -2854
rect -60 -2858 -30 -2854
rect 224 -2858 286 -2854
rect 290 -2858 320 -2854
rect 368 -2858 398 -2854
rect 580 -2858 642 -2854
rect 646 -2858 676 -2854
rect 724 -2858 754 -2854
rect 978 -2858 1040 -2854
rect 1044 -2858 1074 -2854
rect 1122 -2858 1152 -2854
rect 1336 -2858 1398 -2854
rect 1402 -2858 1432 -2854
rect 1480 -2858 1510 -2854
rect -913 -2865 -882 -2861
rect -555 -2865 -524 -2861
rect -197 -2865 -166 -2861
rect 231 -2865 262 -2861
rect 587 -2865 618 -2861
rect 985 -2865 1016 -2861
rect 1343 -2865 1374 -2861
rect -931 -2872 -848 -2868
rect -809 -2872 -706 -2868
rect -573 -2872 -490 -2868
rect -451 -2872 -348 -2868
rect -215 -2872 -132 -2868
rect -93 -2872 10 -2868
rect 213 -2872 296 -2868
rect 335 -2872 438 -2868
rect 569 -2872 652 -2868
rect 691 -2872 794 -2868
rect 967 -2872 1050 -2868
rect 1089 -2872 1192 -2868
rect 1325 -2872 1408 -2868
rect 1447 -2872 1550 -2868
rect -949 -2879 -928 -2875
rect -894 -2879 -865 -2875
rect -861 -2879 -780 -2875
rect -691 -2879 -592 -2875
rect -585 -2879 -570 -2875
rect -536 -2879 -507 -2875
rect -503 -2879 -422 -2875
rect -333 -2878 -234 -2874
rect -596 -2883 -592 -2879
rect -238 -2883 -234 -2878
rect -227 -2879 -212 -2875
rect -178 -2879 -149 -2875
rect -145 -2879 -64 -2875
rect 25 -2879 194 -2875
rect 201 -2879 216 -2875
rect 250 -2879 279 -2875
rect 283 -2879 364 -2875
rect 453 -2879 550 -2875
rect 557 -2879 572 -2875
rect 606 -2879 635 -2875
rect 639 -2879 720 -2875
rect 809 -2879 948 -2875
rect 955 -2879 970 -2875
rect 1004 -2879 1033 -2875
rect 1037 -2879 1118 -2875
rect 1207 -2877 1300 -2873
rect 190 -2883 194 -2879
rect 546 -2883 550 -2879
rect 944 -2883 948 -2879
rect 1296 -2883 1300 -2877
rect 1307 -2879 1328 -2875
rect 1362 -2879 1391 -2875
rect 1395 -2879 1476 -2875
rect -1260 -2888 -1203 -2884
rect -1164 -2887 -902 -2883
rect -887 -2887 -804 -2883
rect -783 -2887 -689 -2883
rect -596 -2887 -544 -2883
rect -529 -2887 -446 -2883
rect -425 -2887 -331 -2883
rect -238 -2887 -186 -2883
rect -171 -2887 -88 -2883
rect -67 -2887 27 -2883
rect 190 -2887 242 -2883
rect 257 -2887 340 -2883
rect 361 -2887 455 -2883
rect 546 -2887 598 -2883
rect 613 -2887 696 -2883
rect 717 -2887 811 -2883
rect 944 -2887 996 -2883
rect 1011 -2887 1094 -2883
rect 1115 -2887 1209 -2883
rect 1296 -2887 1354 -2883
rect 1369 -2887 1452 -2883
rect 1473 -2887 1567 -2883
rect -1266 -2895 -1253 -2891
rect -1249 -2895 -1213 -2891
rect -1209 -2895 -1193 -2891
rect -943 -2894 -924 -2890
rect -905 -2894 -776 -2890
rect -591 -2894 -566 -2890
rect -547 -2894 -418 -2890
rect -233 -2894 -208 -2890
rect -189 -2894 -60 -2890
rect 195 -2894 220 -2890
rect 239 -2894 368 -2890
rect 551 -2894 576 -2890
rect 595 -2894 724 -2890
rect 949 -2894 974 -2890
rect 993 -2894 1122 -2890
rect 1313 -2894 1332 -2890
rect 1351 -2894 1480 -2890
rect -1309 -2902 -1257 -2898
rect -1253 -2902 -1227 -2898
rect -1223 -2902 -1179 -2898
rect -898 -2901 -794 -2897
rect -790 -2901 -760 -2897
rect -540 -2901 -436 -2897
rect -432 -2901 -402 -2897
rect -182 -2901 -78 -2897
rect -74 -2901 -44 -2897
rect 246 -2901 350 -2897
rect 354 -2901 384 -2897
rect 602 -2901 706 -2897
rect 710 -2901 740 -2897
rect 1000 -2901 1104 -2897
rect 1108 -2901 1138 -2897
rect 1358 -2901 1462 -2897
rect 1466 -2901 1496 -2897
rect -1216 -2909 -1162 -2905
rect -924 -2908 -872 -2904
rect -868 -2908 -838 -2904
rect -566 -2908 -514 -2904
rect -510 -2908 -480 -2904
rect -208 -2908 -156 -2904
rect -152 -2908 -122 -2904
rect 220 -2908 272 -2904
rect 276 -2908 306 -2904
rect 576 -2908 628 -2904
rect 632 -2908 662 -2904
rect 974 -2908 1026 -2904
rect 1030 -2908 1060 -2904
rect 1332 -2908 1384 -2904
rect 1388 -2908 1418 -2904
rect -1234 -2916 -1202 -2912
rect -879 -2916 -847 -2912
rect -883 -2919 -879 -2916
rect -847 -2919 -843 -2916
rect -801 -2916 -769 -2912
rect -805 -2919 -801 -2916
rect -769 -2919 -765 -2916
rect -521 -2916 -489 -2912
rect -525 -2919 -521 -2916
rect -489 -2919 -485 -2916
rect -443 -2916 -411 -2912
rect -447 -2919 -443 -2916
rect -411 -2919 -407 -2916
rect -163 -2916 -131 -2912
rect -167 -2919 -163 -2916
rect -131 -2919 -127 -2916
rect -85 -2916 -53 -2912
rect -89 -2919 -85 -2916
rect -53 -2919 -49 -2916
rect 265 -2916 297 -2912
rect 261 -2919 265 -2916
rect 297 -2919 301 -2916
rect 343 -2916 375 -2912
rect 339 -2919 343 -2916
rect 375 -2919 379 -2916
rect 621 -2916 653 -2912
rect 617 -2919 621 -2916
rect 653 -2919 657 -2916
rect 699 -2916 731 -2912
rect 695 -2919 699 -2916
rect 731 -2919 735 -2916
rect 1019 -2916 1051 -2912
rect 1015 -2919 1019 -2916
rect 1051 -2919 1055 -2916
rect 1097 -2916 1129 -2912
rect 1093 -2919 1097 -2916
rect 1129 -2919 1133 -2916
rect 1377 -2916 1409 -2912
rect 1373 -2919 1377 -2916
rect 1409 -2919 1413 -2916
rect 1455 -2916 1487 -2912
rect 1451 -2919 1455 -2916
rect 1487 -2919 1491 -2916
rect -926 -2927 -922 -2923
rect -900 -2927 -896 -2923
rect -857 -2927 -853 -2923
rect -822 -2927 -818 -2923
rect -778 -2927 -774 -2923
rect -761 -2927 -757 -2923
rect -725 -2927 -721 -2923
rect -704 -2927 -700 -2923
rect -568 -2927 -564 -2923
rect -542 -2927 -538 -2923
rect -499 -2927 -495 -2923
rect -464 -2927 -460 -2923
rect -420 -2927 -416 -2923
rect -403 -2927 -399 -2923
rect -367 -2927 -363 -2923
rect -346 -2927 -342 -2923
rect -210 -2927 -206 -2923
rect -184 -2927 -180 -2923
rect -141 -2927 -137 -2923
rect -106 -2927 -102 -2923
rect -62 -2927 -58 -2923
rect -45 -2927 -41 -2923
rect -9 -2927 -5 -2923
rect 12 -2927 16 -2923
rect 218 -2927 222 -2923
rect 244 -2927 248 -2923
rect 287 -2927 291 -2923
rect 322 -2927 326 -2923
rect 366 -2927 370 -2923
rect 383 -2927 387 -2923
rect 419 -2927 423 -2923
rect 440 -2927 444 -2923
rect 574 -2927 578 -2923
rect 600 -2927 604 -2923
rect 643 -2927 647 -2923
rect 678 -2927 682 -2923
rect 722 -2927 726 -2923
rect 739 -2927 743 -2923
rect 775 -2927 779 -2923
rect 796 -2927 800 -2923
rect 972 -2927 976 -2923
rect 998 -2927 1002 -2923
rect 1041 -2927 1045 -2923
rect 1076 -2927 1080 -2923
rect 1120 -2927 1124 -2923
rect 1137 -2927 1141 -2923
rect 1173 -2927 1177 -2923
rect 1194 -2927 1198 -2923
rect 1330 -2927 1334 -2923
rect 1356 -2927 1360 -2923
rect 1399 -2927 1403 -2923
rect 1434 -2927 1438 -2923
rect 1478 -2927 1482 -2923
rect 1495 -2927 1499 -2923
rect 1531 -2927 1535 -2923
rect 1552 -2927 1556 -2923
rect 1633 -2927 1695 -2812
rect -1421 -2931 -1255 -2927
rect -1251 -2931 -1211 -2927
rect -1207 -2931 -1177 -2927
rect -1173 -2931 -926 -2927
rect -922 -2931 -900 -2927
rect -896 -2931 -857 -2927
rect -853 -2931 -822 -2927
rect -818 -2931 -778 -2927
rect -774 -2931 -761 -2927
rect -757 -2931 -725 -2927
rect -721 -2931 -704 -2927
rect -700 -2931 -568 -2927
rect -564 -2931 -542 -2927
rect -538 -2931 -499 -2927
rect -495 -2931 -464 -2927
rect -460 -2931 -420 -2927
rect -416 -2931 -403 -2927
rect -399 -2931 -367 -2927
rect -363 -2931 -346 -2927
rect -342 -2931 -210 -2927
rect -206 -2931 -184 -2927
rect -180 -2931 -141 -2927
rect -137 -2931 -106 -2927
rect -102 -2931 -62 -2927
rect -58 -2931 -45 -2927
rect -41 -2931 -9 -2927
rect -5 -2931 12 -2927
rect 16 -2931 218 -2927
rect 222 -2931 244 -2927
rect 248 -2931 287 -2927
rect 291 -2931 322 -2927
rect 326 -2931 366 -2927
rect 370 -2931 383 -2927
rect 387 -2931 419 -2927
rect 423 -2931 440 -2927
rect 444 -2931 574 -2927
rect 578 -2931 600 -2927
rect 604 -2931 643 -2927
rect 647 -2931 678 -2927
rect 682 -2931 722 -2927
rect 726 -2931 739 -2927
rect 743 -2931 775 -2927
rect 779 -2931 796 -2927
rect 800 -2931 972 -2927
rect 976 -2931 998 -2927
rect 1002 -2931 1041 -2927
rect 1045 -2931 1076 -2927
rect 1080 -2931 1120 -2927
rect 1124 -2931 1137 -2927
rect 1141 -2931 1173 -2927
rect 1177 -2931 1194 -2927
rect 1198 -2931 1330 -2927
rect 1334 -2931 1356 -2927
rect 1360 -2931 1399 -2927
rect 1403 -2931 1434 -2927
rect 1438 -2931 1478 -2927
rect 1482 -2931 1495 -2927
rect 1499 -2931 1531 -2927
rect 1535 -2931 1552 -2927
rect 1556 -2931 1695 -2927
rect -1272 -2938 -689 -2934
rect -585 -2938 27 -2934
rect 201 -2938 811 -2934
rect 955 -2938 1567 -2934
rect -1266 -2946 -1162 -2942
rect -943 -2945 -331 -2941
rect -227 -2945 455 -2941
rect 557 -2945 1209 -2941
rect 1313 -2945 1561 -2941
rect -1495 -2958 -1255 -2954
rect -1251 -2958 -1238 -2954
rect -1234 -2958 -1218 -2954
rect -1214 -2958 -1197 -2954
rect -1193 -2958 -1176 -2954
rect -1172 -2958 -1155 -2954
rect -1151 -2958 -1134 -2954
rect -1130 -2958 -1113 -2954
rect -1109 -2958 -1092 -2954
rect -1088 -2958 -1072 -2954
rect -1068 -2958 -1026 -2954
rect -1022 -2958 -926 -2954
rect -922 -2958 -909 -2954
rect -905 -2958 -889 -2954
rect -885 -2958 -868 -2954
rect -864 -2958 -847 -2954
rect -843 -2958 -826 -2954
rect -822 -2958 -805 -2954
rect -801 -2958 -784 -2954
rect -780 -2958 -763 -2954
rect -759 -2958 -743 -2954
rect -739 -2958 -672 -2954
rect -668 -2958 -568 -2954
rect -564 -2958 -551 -2954
rect -547 -2958 -531 -2954
rect -527 -2958 -510 -2954
rect -506 -2958 -489 -2954
rect -485 -2958 -468 -2954
rect -464 -2958 -447 -2954
rect -443 -2958 -426 -2954
rect -422 -2958 -405 -2954
rect -401 -2958 -385 -2954
rect -381 -2958 -329 -2954
rect -325 -2958 -210 -2954
rect -206 -2958 -193 -2954
rect -189 -2958 -173 -2954
rect -169 -2958 -152 -2954
rect -148 -2958 -131 -2954
rect -127 -2958 -110 -2954
rect -106 -2958 -89 -2954
rect -85 -2958 -68 -2954
rect -64 -2958 -47 -2954
rect -43 -2958 -27 -2954
rect -23 -2958 218 -2954
rect 222 -2958 235 -2954
rect 239 -2958 255 -2954
rect 259 -2958 276 -2954
rect 280 -2958 297 -2954
rect 301 -2958 318 -2954
rect 322 -2958 339 -2954
rect 343 -2958 360 -2954
rect 364 -2958 381 -2954
rect 385 -2958 401 -2954
rect 405 -2958 472 -2954
rect 476 -2958 841 -2954
rect 845 -2958 1199 -2954
rect 1203 -2958 1617 -2954
rect -1495 -3070 -1433 -2958
rect -1100 -2979 -931 -2975
rect -1233 -3006 -1199 -3002
rect -1135 -3006 -1115 -3002
rect -1266 -3014 -1257 -3010
rect -1253 -3014 -1223 -3010
rect -1202 -3014 -1171 -3010
rect -1142 -3014 -1111 -3010
rect -1100 -3014 -1073 -3010
rect -1014 -3008 -1010 -3004
rect -935 -3010 -931 -2979
rect -413 -2980 -215 -2976
rect -771 -2996 -573 -2992
rect -904 -3006 -870 -3002
rect -806 -3006 -786 -3002
rect -660 -3007 -656 -3003
rect -577 -3010 -573 -2996
rect -546 -3006 -512 -3002
rect -448 -3006 -428 -3002
rect -935 -3014 -928 -3010
rect -924 -3014 -894 -3010
rect -873 -3014 -842 -3010
rect -813 -3014 -782 -3010
rect -771 -3014 -744 -3010
rect -577 -3014 -570 -3010
rect -566 -3014 -536 -3010
rect -515 -3014 -484 -3010
rect -455 -3014 -424 -3010
rect -413 -3014 -386 -3010
rect -317 -3009 -313 -3005
rect -219 -3010 -215 -2980
rect -188 -3006 -154 -3002
rect -90 -3006 -70 -3002
rect -55 -3006 213 -3002
rect 240 -3006 274 -3002
rect 338 -3006 358 -3002
rect 373 -3006 409 -3002
rect 209 -3010 213 -3006
rect 484 -3007 488 -3003
rect 853 -3007 857 -3003
rect -219 -3014 -212 -3010
rect -208 -3014 -178 -3010
rect -157 -3014 -126 -3010
rect -97 -3014 -66 -3010
rect -55 -3014 -28 -3010
rect 209 -3014 216 -3010
rect 220 -3014 250 -3010
rect 271 -3014 302 -3010
rect 331 -3014 362 -3010
rect 373 -3014 400 -3010
rect 1211 -3008 1215 -3004
rect -1260 -3021 -1213 -3017
rect -1177 -3021 -1164 -3017
rect -1160 -3021 -1129 -3017
rect -1093 -3021 -1080 -3017
rect -1076 -3021 -1064 -3017
rect -931 -3021 -884 -3017
rect -848 -3021 -835 -3017
rect -831 -3021 -800 -3017
rect -764 -3021 -751 -3017
rect -747 -3021 -735 -3017
rect -573 -3021 -526 -3017
rect -490 -3021 -477 -3017
rect -473 -3021 -442 -3017
rect -406 -3021 -393 -3017
rect -389 -3021 -377 -3017
rect -215 -3021 -168 -3017
rect -132 -3021 -119 -3017
rect -115 -3021 -84 -3017
rect -48 -3021 -35 -3017
rect -31 -3021 -19 -3017
rect 213 -3021 260 -3017
rect 296 -3021 309 -3017
rect 313 -3021 344 -3017
rect 380 -3021 393 -3017
rect 397 -3021 409 -3017
rect -1268 -3028 -1267 -3024
rect -1263 -3028 -1253 -3024
rect -1249 -3028 -1139 -3024
rect -1118 -3028 -1087 -3024
rect -936 -3028 -924 -3024
rect -920 -3028 -810 -3024
rect -789 -3028 -758 -3024
rect -586 -3028 -566 -3024
rect -562 -3028 -452 -3024
rect -431 -3028 -400 -3024
rect -223 -3028 -208 -3024
rect -204 -3028 -94 -3024
rect -73 -3028 -42 -3024
rect 194 -3028 195 -3024
rect 199 -3028 220 -3024
rect 224 -3028 334 -3024
rect 355 -3028 386 -3024
rect -1218 -3035 -1195 -3031
rect -1176 -3035 -1157 -3031
rect -889 -3035 -866 -3031
rect -847 -3035 -828 -3031
rect -531 -3035 -508 -3031
rect -489 -3035 -470 -3031
rect -173 -3035 -150 -3031
rect -131 -3035 -112 -3031
rect 255 -3035 278 -3031
rect 297 -3035 316 -3031
rect 1633 -3046 1695 -2931
rect -1421 -3050 -1255 -3046
rect -1251 -3050 -1238 -3046
rect -1234 -3050 -1197 -3046
rect -1193 -3050 -1155 -3046
rect -1151 -3050 -1113 -3046
rect -1109 -3050 -1072 -3046
rect -1068 -3050 -1026 -3046
rect -1022 -3050 -926 -3046
rect -922 -3050 -909 -3046
rect -905 -3050 -868 -3046
rect -864 -3050 -826 -3046
rect -822 -3050 -784 -3046
rect -780 -3050 -743 -3046
rect -739 -3050 -672 -3046
rect -668 -3050 -568 -3046
rect -564 -3050 -551 -3046
rect -547 -3050 -510 -3046
rect -506 -3050 -468 -3046
rect -464 -3050 -426 -3046
rect -422 -3050 -385 -3046
rect -381 -3050 -329 -3046
rect -325 -3050 -210 -3046
rect -206 -3050 -193 -3046
rect -189 -3050 -152 -3046
rect -148 -3050 -110 -3046
rect -106 -3050 -68 -3046
rect -64 -3050 -27 -3046
rect -23 -3050 218 -3046
rect 222 -3050 235 -3046
rect 239 -3050 276 -3046
rect 280 -3050 318 -3046
rect 322 -3050 360 -3046
rect 364 -3050 401 -3046
rect 405 -3050 472 -3046
rect 476 -3050 841 -3046
rect 845 -3050 1199 -3046
rect 1203 -3050 1695 -3046
rect -1495 -3074 -1255 -3070
rect -1251 -3074 -1238 -3070
rect -1234 -3074 -1218 -3070
rect -1214 -3074 -1197 -3070
rect -1193 -3074 -1176 -3070
rect -1172 -3074 -1155 -3070
rect -1151 -3074 -1134 -3070
rect -1130 -3074 -1113 -3070
rect -1109 -3074 -1092 -3070
rect -1088 -3074 -1072 -3070
rect -1068 -3074 -1026 -3070
rect -1022 -3074 -926 -3070
rect -922 -3074 -909 -3070
rect -905 -3074 -889 -3070
rect -885 -3074 -868 -3070
rect -864 -3074 -847 -3070
rect -843 -3074 -826 -3070
rect -822 -3074 -805 -3070
rect -801 -3074 -784 -3070
rect -780 -3074 -763 -3070
rect -759 -3074 -743 -3070
rect -739 -3074 -568 -3070
rect -564 -3074 -551 -3070
rect -547 -3074 -531 -3070
rect -527 -3074 -510 -3070
rect -506 -3074 -489 -3070
rect -485 -3074 -468 -3070
rect -464 -3074 -447 -3070
rect -443 -3074 -426 -3070
rect -422 -3074 -405 -3070
rect -401 -3074 -385 -3070
rect -381 -3074 -329 -3070
rect -325 -3074 -210 -3070
rect -206 -3074 -193 -3070
rect -189 -3074 -173 -3070
rect -169 -3074 -152 -3070
rect -148 -3074 -131 -3070
rect -127 -3074 -110 -3070
rect -106 -3074 -89 -3070
rect -85 -3074 -68 -3070
rect -64 -3074 -47 -3070
rect -43 -3074 -27 -3070
rect -23 -3074 218 -3070
rect 222 -3074 235 -3070
rect 239 -3074 255 -3070
rect 259 -3074 276 -3070
rect 280 -3074 297 -3070
rect 301 -3074 318 -3070
rect 322 -3074 339 -3070
rect 343 -3074 360 -3070
rect 364 -3074 381 -3070
rect 385 -3074 401 -3070
rect 405 -3074 472 -3070
rect 476 -3074 574 -3070
rect 578 -3074 591 -3070
rect 595 -3074 611 -3070
rect 615 -3074 632 -3070
rect 636 -3074 653 -3070
rect 657 -3074 674 -3070
rect 678 -3074 695 -3070
rect 699 -3074 716 -3070
rect 720 -3074 737 -3070
rect 741 -3074 757 -3070
rect 761 -3074 972 -3070
rect 976 -3074 989 -3070
rect 993 -3074 1009 -3070
rect 1013 -3074 1030 -3070
rect 1034 -3074 1051 -3070
rect 1055 -3074 1072 -3070
rect 1076 -3074 1093 -3070
rect 1097 -3074 1114 -3070
rect 1118 -3074 1135 -3070
rect 1139 -3074 1155 -3070
rect 1159 -3074 1199 -3070
rect 1203 -3074 1330 -3070
rect 1334 -3074 1347 -3070
rect 1351 -3074 1367 -3070
rect 1371 -3074 1388 -3070
rect 1392 -3074 1409 -3070
rect 1413 -3074 1430 -3070
rect 1434 -3074 1451 -3070
rect 1455 -3074 1472 -3070
rect 1476 -3074 1493 -3070
rect 1497 -3074 1513 -3070
rect 1517 -3074 1617 -3070
rect -1495 -3191 -1433 -3074
rect -1233 -3122 -1199 -3118
rect -1135 -3122 -1115 -3118
rect -1100 -3122 -1066 -3118
rect -1014 -3123 -1010 -3119
rect -904 -3122 -870 -3118
rect -806 -3122 -786 -3118
rect -771 -3122 -737 -3118
rect -546 -3122 -512 -3118
rect -448 -3122 -428 -3118
rect -413 -3122 -379 -3118
rect -1272 -3130 -1257 -3126
rect -1253 -3130 -1223 -3126
rect -1202 -3130 -1171 -3126
rect -1142 -3130 -1111 -3126
rect -1100 -3130 -1073 -3126
rect -943 -3130 -928 -3126
rect -924 -3130 -894 -3126
rect -873 -3130 -842 -3126
rect -813 -3130 -782 -3126
rect -771 -3130 -744 -3126
rect -585 -3130 -570 -3126
rect -566 -3130 -536 -3126
rect -515 -3130 -484 -3126
rect -455 -3130 -424 -3126
rect -413 -3130 -386 -3126
rect -317 -3124 -313 -3120
rect -188 -3122 -154 -3118
rect -90 -3122 -70 -3118
rect -55 -3122 -21 -3118
rect 240 -3122 274 -3118
rect 338 -3122 358 -3118
rect 373 -3122 407 -3118
rect 484 -3123 488 -3119
rect 596 -3122 630 -3118
rect 694 -3122 714 -3118
rect 729 -3122 763 -3118
rect 994 -3122 1028 -3118
rect 1092 -3122 1112 -3118
rect 1127 -3122 1161 -3118
rect 1211 -3123 1215 -3119
rect 1352 -3122 1386 -3118
rect 1450 -3122 1470 -3118
rect 1485 -3122 1519 -3118
rect -227 -3130 -212 -3126
rect -208 -3130 -178 -3126
rect -157 -3130 -126 -3126
rect -97 -3130 -66 -3126
rect -55 -3130 -28 -3126
rect 201 -3130 216 -3126
rect 220 -3130 250 -3126
rect 271 -3130 302 -3126
rect 331 -3130 362 -3126
rect 373 -3130 400 -3126
rect 557 -3130 572 -3126
rect 576 -3130 606 -3126
rect 627 -3130 658 -3126
rect 687 -3130 718 -3126
rect 729 -3130 756 -3126
rect 955 -3130 970 -3126
rect 974 -3130 1004 -3126
rect 1025 -3130 1056 -3126
rect 1085 -3130 1116 -3126
rect 1127 -3130 1154 -3126
rect 1313 -3130 1328 -3126
rect 1332 -3130 1362 -3126
rect 1383 -3130 1414 -3126
rect 1443 -3130 1474 -3126
rect 1485 -3130 1512 -3126
rect -1260 -3137 -1213 -3133
rect -1177 -3137 -1164 -3133
rect -1160 -3137 -1129 -3133
rect -1093 -3137 -1080 -3133
rect -1076 -3137 -1064 -3133
rect -931 -3137 -884 -3133
rect -848 -3137 -835 -3133
rect -831 -3137 -800 -3133
rect -764 -3137 -751 -3133
rect -747 -3137 -735 -3133
rect -573 -3137 -526 -3133
rect -490 -3137 -477 -3133
rect -473 -3137 -442 -3133
rect -406 -3137 -393 -3133
rect -389 -3137 -377 -3133
rect -215 -3137 -168 -3133
rect -132 -3137 -119 -3133
rect -115 -3137 -84 -3133
rect -48 -3137 -35 -3133
rect -31 -3137 -19 -3133
rect 213 -3137 260 -3133
rect 296 -3137 309 -3133
rect 313 -3137 344 -3133
rect 380 -3137 393 -3133
rect 397 -3137 409 -3133
rect 569 -3137 616 -3133
rect 652 -3137 665 -3133
rect 669 -3137 700 -3133
rect 736 -3137 749 -3133
rect 753 -3137 765 -3133
rect 967 -3137 1014 -3133
rect 1050 -3137 1063 -3133
rect 1067 -3137 1098 -3133
rect 1134 -3137 1147 -3133
rect 1151 -3137 1163 -3133
rect 1325 -3137 1372 -3133
rect 1408 -3137 1421 -3133
rect 1425 -3137 1456 -3133
rect 1492 -3137 1505 -3133
rect 1509 -3137 1521 -3133
rect -1274 -3144 -1253 -3140
rect -1249 -3144 -1139 -3140
rect -1118 -3144 -1087 -3140
rect -936 -3144 -924 -3140
rect -920 -3144 -810 -3140
rect -789 -3144 -758 -3140
rect -585 -3144 -584 -3140
rect -580 -3144 -566 -3140
rect -562 -3144 -452 -3140
rect -431 -3144 -400 -3140
rect -221 -3144 -208 -3140
rect -204 -3144 -94 -3140
rect -73 -3144 -42 -3140
rect 200 -3144 201 -3140
rect 205 -3144 220 -3140
rect 224 -3144 334 -3140
rect 355 -3144 386 -3140
rect 562 -3144 576 -3140
rect 580 -3144 690 -3140
rect 711 -3144 742 -3140
rect 958 -3144 974 -3140
rect 978 -3144 1088 -3140
rect 1109 -3144 1140 -3140
rect 1318 -3144 1332 -3140
rect 1336 -3144 1446 -3140
rect 1467 -3144 1498 -3140
rect -1218 -3151 -1195 -3147
rect -1176 -3151 -1157 -3147
rect -889 -3151 -866 -3147
rect -847 -3151 -828 -3147
rect -531 -3151 -508 -3147
rect -489 -3151 -470 -3147
rect -173 -3151 -150 -3147
rect -131 -3151 -112 -3147
rect 255 -3151 278 -3147
rect 297 -3151 316 -3147
rect 611 -3151 634 -3147
rect 653 -3151 672 -3147
rect 1009 -3151 1032 -3147
rect 1051 -3151 1070 -3147
rect 1367 -3151 1390 -3147
rect 1409 -3151 1428 -3147
rect 1633 -3162 1695 -3050
rect -1421 -3166 -1255 -3162
rect -1251 -3166 -1238 -3162
rect -1234 -3166 -1197 -3162
rect -1193 -3166 -1155 -3162
rect -1151 -3166 -1113 -3162
rect -1109 -3166 -1072 -3162
rect -1068 -3166 -1026 -3162
rect -1022 -3166 -926 -3162
rect -922 -3166 -909 -3162
rect -905 -3166 -868 -3162
rect -864 -3166 -826 -3162
rect -822 -3166 -784 -3162
rect -780 -3166 -743 -3162
rect -739 -3166 -568 -3162
rect -564 -3166 -551 -3162
rect -547 -3166 -510 -3162
rect -506 -3166 -468 -3162
rect -464 -3166 -426 -3162
rect -422 -3166 -385 -3162
rect -381 -3166 -329 -3162
rect -325 -3166 -210 -3162
rect -206 -3166 -193 -3162
rect -189 -3166 -152 -3162
rect -148 -3166 -110 -3162
rect -106 -3166 -68 -3162
rect -64 -3166 -27 -3162
rect -23 -3166 218 -3162
rect 222 -3166 235 -3162
rect 239 -3166 276 -3162
rect 280 -3166 318 -3162
rect 322 -3166 360 -3162
rect 364 -3166 401 -3162
rect 405 -3166 472 -3162
rect 476 -3166 574 -3162
rect 578 -3166 591 -3162
rect 595 -3166 632 -3162
rect 636 -3166 674 -3162
rect 678 -3166 716 -3162
rect 720 -3166 757 -3162
rect 761 -3166 972 -3162
rect 976 -3166 989 -3162
rect 993 -3166 1030 -3162
rect 1034 -3166 1072 -3162
rect 1076 -3166 1114 -3162
rect 1118 -3166 1155 -3162
rect 1159 -3166 1199 -3162
rect 1203 -3166 1330 -3162
rect 1334 -3166 1347 -3162
rect 1351 -3166 1388 -3162
rect 1392 -3166 1430 -3162
rect 1434 -3166 1472 -3162
rect 1476 -3166 1513 -3162
rect 1517 -3166 1695 -3162
rect -1266 -3174 -1066 -3170
rect -943 -3174 -737 -3170
rect -585 -3173 -379 -3169
rect -227 -3174 -21 -3170
rect 201 -3173 407 -3169
rect 557 -3173 763 -3169
rect 955 -3173 1161 -3169
rect 1313 -3174 1519 -3170
rect -1495 -3195 -1255 -3191
rect -1251 -3195 -1238 -3191
rect -1234 -3195 -1218 -3191
rect -1214 -3195 -1197 -3191
rect -1193 -3195 -1176 -3191
rect -1172 -3195 -1155 -3191
rect -1151 -3195 -1134 -3191
rect -1130 -3195 -1113 -3191
rect -1109 -3195 -1092 -3191
rect -1088 -3195 -1072 -3191
rect -1068 -3195 -926 -3191
rect -922 -3195 -909 -3191
rect -905 -3195 -889 -3191
rect -885 -3195 -868 -3191
rect -864 -3195 -847 -3191
rect -843 -3195 -826 -3191
rect -822 -3195 -805 -3191
rect -801 -3195 -784 -3191
rect -780 -3195 -763 -3191
rect -759 -3195 -743 -3191
rect -739 -3195 -568 -3191
rect -564 -3195 -551 -3191
rect -547 -3195 -531 -3191
rect -527 -3195 -510 -3191
rect -506 -3195 -489 -3191
rect -485 -3195 -468 -3191
rect -464 -3195 -447 -3191
rect -443 -3195 -426 -3191
rect -422 -3195 -405 -3191
rect -401 -3195 -385 -3191
rect -381 -3195 -210 -3191
rect -206 -3195 -193 -3191
rect -189 -3195 -173 -3191
rect -169 -3195 -152 -3191
rect -148 -3195 -131 -3191
rect -127 -3195 -110 -3191
rect -106 -3195 -89 -3191
rect -85 -3195 -68 -3191
rect -64 -3195 -47 -3191
rect -43 -3195 -27 -3191
rect -23 -3195 218 -3191
rect 222 -3195 235 -3191
rect 239 -3195 255 -3191
rect 259 -3195 276 -3191
rect 280 -3195 297 -3191
rect 301 -3195 318 -3191
rect 322 -3195 339 -3191
rect 343 -3195 360 -3191
rect 364 -3195 381 -3191
rect 385 -3195 401 -3191
rect 405 -3195 574 -3191
rect 578 -3195 591 -3191
rect 595 -3195 611 -3191
rect 615 -3195 632 -3191
rect 636 -3195 653 -3191
rect 657 -3195 674 -3191
rect 678 -3195 695 -3191
rect 699 -3195 716 -3191
rect 720 -3195 737 -3191
rect 741 -3195 757 -3191
rect 761 -3195 972 -3191
rect 976 -3195 989 -3191
rect 993 -3195 1009 -3191
rect 1013 -3195 1030 -3191
rect 1034 -3195 1051 -3191
rect 1055 -3195 1072 -3191
rect 1076 -3195 1093 -3191
rect 1097 -3195 1114 -3191
rect 1118 -3195 1135 -3191
rect 1139 -3195 1155 -3191
rect 1159 -3195 1330 -3191
rect 1334 -3195 1347 -3191
rect 1351 -3195 1367 -3191
rect 1371 -3195 1388 -3191
rect 1392 -3195 1409 -3191
rect 1413 -3195 1430 -3191
rect 1434 -3195 1451 -3191
rect 1455 -3195 1472 -3191
rect 1476 -3195 1493 -3191
rect 1497 -3195 1513 -3191
rect 1517 -3195 1617 -3191
rect -1495 -3305 -1433 -3195
rect -1233 -3243 -1199 -3239
rect -1135 -3243 -1115 -3239
rect -1100 -3243 -1066 -3239
rect -904 -3243 -870 -3239
rect -806 -3243 -786 -3239
rect -771 -3243 -737 -3239
rect -546 -3243 -512 -3239
rect -448 -3243 -428 -3239
rect -413 -3243 -373 -3239
rect -188 -3243 -154 -3239
rect -90 -3243 -70 -3239
rect -55 -3243 -21 -3239
rect 240 -3243 274 -3239
rect 338 -3243 358 -3239
rect 373 -3243 407 -3239
rect 596 -3243 630 -3239
rect 694 -3243 714 -3239
rect 729 -3243 763 -3239
rect 994 -3243 1028 -3239
rect 1092 -3243 1112 -3239
rect 1127 -3243 1161 -3239
rect 1352 -3243 1386 -3239
rect 1450 -3243 1470 -3239
rect 1485 -3243 1519 -3239
rect -1345 -3251 -1257 -3247
rect -1253 -3251 -1223 -3247
rect -1202 -3251 -1171 -3247
rect -1142 -3251 -1111 -3247
rect -1100 -3251 -1073 -3247
rect -937 -3251 -928 -3247
rect -924 -3251 -894 -3247
rect -873 -3251 -842 -3247
rect -813 -3251 -782 -3247
rect -771 -3251 -744 -3247
rect -579 -3251 -570 -3247
rect -566 -3251 -536 -3247
rect -515 -3251 -484 -3247
rect -455 -3251 -424 -3247
rect -413 -3251 -386 -3247
rect -221 -3251 -212 -3247
rect -208 -3251 -178 -3247
rect -157 -3251 -126 -3247
rect -97 -3251 -66 -3247
rect -55 -3251 -28 -3247
rect 207 -3251 216 -3247
rect 220 -3251 250 -3247
rect 271 -3251 302 -3247
rect 331 -3251 362 -3247
rect 373 -3251 400 -3247
rect 563 -3251 572 -3247
rect 576 -3251 606 -3247
rect 627 -3251 658 -3247
rect 687 -3251 718 -3247
rect 729 -3251 756 -3247
rect 961 -3251 970 -3247
rect 974 -3251 1004 -3247
rect 1025 -3251 1056 -3247
rect 1085 -3251 1116 -3247
rect 1127 -3251 1154 -3247
rect 1319 -3251 1328 -3247
rect 1332 -3251 1362 -3247
rect 1383 -3251 1414 -3247
rect 1443 -3251 1474 -3247
rect 1485 -3251 1512 -3247
rect -1260 -3258 -1213 -3254
rect -1177 -3258 -1164 -3254
rect -1160 -3258 -1129 -3254
rect -1093 -3258 -1080 -3254
rect -1076 -3258 -1064 -3254
rect -931 -3258 -884 -3254
rect -848 -3258 -835 -3254
rect -831 -3258 -800 -3254
rect -764 -3258 -751 -3254
rect -747 -3258 -735 -3254
rect -573 -3258 -526 -3254
rect -490 -3258 -477 -3254
rect -473 -3258 -442 -3254
rect -406 -3258 -393 -3254
rect -389 -3258 -377 -3254
rect -215 -3258 -168 -3254
rect -132 -3258 -119 -3254
rect -115 -3258 -84 -3254
rect -48 -3258 -35 -3254
rect -31 -3258 -19 -3254
rect 213 -3258 260 -3254
rect 296 -3258 309 -3254
rect 313 -3258 344 -3254
rect 380 -3258 393 -3254
rect 397 -3258 409 -3254
rect 569 -3258 616 -3254
rect 652 -3258 665 -3254
rect 669 -3258 700 -3254
rect 736 -3258 749 -3254
rect 753 -3258 765 -3254
rect 967 -3258 1014 -3254
rect 1050 -3258 1063 -3254
rect 1067 -3258 1098 -3254
rect 1134 -3258 1147 -3254
rect 1151 -3258 1163 -3254
rect 1325 -3258 1372 -3254
rect 1408 -3258 1421 -3254
rect 1425 -3258 1456 -3254
rect 1492 -3258 1505 -3254
rect 1509 -3258 1521 -3254
rect -1274 -3265 -1253 -3261
rect -1249 -3265 -1139 -3261
rect -1118 -3265 -1087 -3261
rect -936 -3265 -924 -3261
rect -920 -3265 -810 -3261
rect -789 -3265 -758 -3261
rect -580 -3265 -566 -3261
rect -562 -3265 -452 -3261
rect -431 -3265 -400 -3261
rect -221 -3265 -208 -3261
rect -204 -3265 -94 -3261
rect -73 -3265 -42 -3261
rect 205 -3265 220 -3261
rect 224 -3265 334 -3261
rect 355 -3265 386 -3261
rect 562 -3265 576 -3261
rect 580 -3265 690 -3261
rect 711 -3265 742 -3261
rect 958 -3265 974 -3261
rect 978 -3265 1088 -3261
rect 1109 -3265 1140 -3261
rect 1318 -3265 1332 -3261
rect 1336 -3265 1446 -3261
rect 1467 -3265 1498 -3261
rect -1218 -3272 -1195 -3268
rect -1176 -3272 -1157 -3268
rect -889 -3272 -866 -3268
rect -847 -3272 -828 -3268
rect -531 -3272 -508 -3268
rect -489 -3272 -470 -3268
rect -173 -3272 -150 -3268
rect -131 -3272 -112 -3268
rect 255 -3272 278 -3268
rect 297 -3272 316 -3268
rect 611 -3272 634 -3268
rect 653 -3272 672 -3268
rect 1009 -3272 1032 -3268
rect 1051 -3272 1070 -3268
rect 1367 -3272 1390 -3268
rect 1409 -3272 1428 -3268
rect 1633 -3283 1695 -3166
rect -1421 -3287 -1255 -3283
rect -1251 -3287 -1238 -3283
rect -1234 -3287 -1197 -3283
rect -1193 -3287 -1155 -3283
rect -1151 -3287 -1113 -3283
rect -1109 -3287 -1072 -3283
rect -1068 -3287 -926 -3283
rect -922 -3287 -909 -3283
rect -905 -3287 -868 -3283
rect -864 -3287 -826 -3283
rect -822 -3287 -784 -3283
rect -780 -3287 -743 -3283
rect -739 -3287 -568 -3283
rect -564 -3287 -551 -3283
rect -547 -3287 -510 -3283
rect -506 -3287 -468 -3283
rect -464 -3287 -426 -3283
rect -422 -3287 -385 -3283
rect -381 -3287 -210 -3283
rect -206 -3287 -193 -3283
rect -189 -3287 -152 -3283
rect -148 -3287 -110 -3283
rect -106 -3287 -68 -3283
rect -64 -3287 -27 -3283
rect -23 -3287 218 -3283
rect 222 -3287 235 -3283
rect 239 -3287 276 -3283
rect 280 -3287 318 -3283
rect 322 -3287 360 -3283
rect 364 -3287 401 -3283
rect 405 -3287 574 -3283
rect 578 -3287 591 -3283
rect 595 -3287 632 -3283
rect 636 -3287 674 -3283
rect 678 -3287 716 -3283
rect 720 -3287 757 -3283
rect 761 -3287 972 -3283
rect 976 -3287 989 -3283
rect 993 -3287 1030 -3283
rect 1034 -3287 1072 -3283
rect 1076 -3287 1114 -3283
rect 1118 -3287 1155 -3283
rect 1159 -3287 1330 -3283
rect 1334 -3287 1347 -3283
rect 1351 -3287 1388 -3283
rect 1392 -3287 1430 -3283
rect 1434 -3287 1472 -3283
rect 1476 -3287 1513 -3283
rect 1517 -3287 1695 -3283
rect -1495 -3309 -1255 -3305
rect -1251 -3309 -1238 -3305
rect -1234 -3309 -1218 -3305
rect -1214 -3309 -1197 -3305
rect -1193 -3309 -1176 -3305
rect -1172 -3309 -1155 -3305
rect -1151 -3309 -1134 -3305
rect -1130 -3309 -1113 -3305
rect -1109 -3309 -1092 -3305
rect -1088 -3309 -1072 -3305
rect -1068 -3309 -926 -3305
rect -922 -3309 -909 -3305
rect -905 -3309 -889 -3305
rect -885 -3309 -868 -3305
rect -864 -3309 -847 -3305
rect -843 -3309 -826 -3305
rect -822 -3309 -805 -3305
rect -801 -3309 -784 -3305
rect -780 -3309 -763 -3305
rect -759 -3309 -743 -3305
rect -739 -3309 -568 -3305
rect -564 -3309 -551 -3305
rect -547 -3309 -531 -3305
rect -527 -3309 -510 -3305
rect -506 -3309 -489 -3305
rect -485 -3309 -468 -3305
rect -464 -3309 -447 -3305
rect -443 -3309 -426 -3305
rect -422 -3309 -405 -3305
rect -401 -3309 -385 -3305
rect -381 -3309 1617 -3305
rect -1495 -3422 -1433 -3309
rect -1233 -3357 -1199 -3353
rect -1135 -3357 -1115 -3353
rect -1100 -3357 -931 -3353
rect -904 -3357 -870 -3353
rect -806 -3357 -786 -3353
rect -771 -3357 -573 -3353
rect -546 -3357 -512 -3353
rect -448 -3357 -428 -3353
rect -413 -3357 -379 -3353
rect -935 -3361 -931 -3357
rect -577 -3361 -573 -3357
rect -1421 -3365 -1257 -3361
rect -1253 -3365 -1223 -3361
rect -1202 -3365 -1171 -3361
rect -1142 -3365 -1111 -3361
rect -1100 -3365 -1073 -3361
rect -935 -3365 -928 -3361
rect -924 -3365 -894 -3361
rect -873 -3365 -842 -3361
rect -813 -3365 -782 -3361
rect -771 -3365 -744 -3361
rect -577 -3365 -570 -3361
rect -566 -3365 -536 -3361
rect -515 -3365 -484 -3361
rect -455 -3365 -424 -3361
rect -413 -3365 -386 -3361
rect -1260 -3372 -1213 -3368
rect -1177 -3372 -1164 -3368
rect -1160 -3372 -1129 -3368
rect -1093 -3372 -1080 -3368
rect -1076 -3372 -1064 -3368
rect -931 -3372 -884 -3368
rect -848 -3372 -835 -3368
rect -831 -3372 -800 -3368
rect -764 -3372 -751 -3368
rect -747 -3372 -735 -3368
rect -573 -3372 -526 -3368
rect -490 -3372 -477 -3368
rect -473 -3372 -442 -3368
rect -406 -3372 -393 -3368
rect -389 -3372 -377 -3368
rect -1279 -3379 -1278 -3375
rect -1274 -3379 -1253 -3375
rect -1249 -3379 -1139 -3375
rect -1118 -3379 -1087 -3375
rect -936 -3379 -924 -3375
rect -920 -3379 -810 -3375
rect -789 -3379 -758 -3375
rect -580 -3379 -566 -3375
rect -562 -3379 -452 -3375
rect -431 -3379 -400 -3375
rect -1218 -3386 -1195 -3382
rect -1176 -3386 -1157 -3382
rect -889 -3386 -866 -3382
rect -847 -3386 -828 -3382
rect -531 -3386 -508 -3382
rect -489 -3386 -470 -3382
rect 1633 -3397 1695 -3287
rect -1421 -3401 -1255 -3397
rect -1251 -3401 -1238 -3397
rect -1234 -3401 -1197 -3397
rect -1193 -3401 -1155 -3397
rect -1151 -3401 -1113 -3397
rect -1109 -3401 -1072 -3397
rect -1068 -3401 -926 -3397
rect -922 -3401 -909 -3397
rect -905 -3401 -868 -3397
rect -864 -3401 -826 -3397
rect -822 -3401 -784 -3397
rect -780 -3401 -743 -3397
rect -739 -3401 -568 -3397
rect -564 -3401 -551 -3397
rect -547 -3401 -510 -3397
rect -506 -3401 -468 -3397
rect -464 -3401 -426 -3397
rect -422 -3401 -385 -3397
rect -381 -3401 1695 -3397
rect -1495 -3426 -1339 -3422
rect -1335 -3426 -1322 -3422
rect -1318 -3426 -935 -3422
rect -931 -3426 -918 -3422
rect -914 -3426 -577 -3422
rect -573 -3426 -560 -3422
rect -556 -3426 -219 -3422
rect -215 -3426 -202 -3422
rect -198 -3426 209 -3422
rect 213 -3426 226 -3422
rect 230 -3426 565 -3422
rect 569 -3426 582 -3422
rect 586 -3426 963 -3422
rect 967 -3426 980 -3422
rect 984 -3426 1321 -3422
rect 1325 -3426 1338 -3422
rect 1342 -3426 1617 -3422
rect -1495 -3546 -1433 -3426
rect -1334 -3458 -1066 -3454
rect -930 -3458 -737 -3454
rect -572 -3458 -373 -3454
rect -214 -3458 -21 -3454
rect 214 -3458 407 -3454
rect 570 -3458 763 -3454
rect 968 -3458 1161 -3454
rect 1326 -3458 1519 -3454
rect -1323 -3466 -923 -3462
rect -919 -3466 -565 -3462
rect -561 -3466 -379 -3462
rect -375 -3466 -207 -3462
rect -203 -3466 221 -3462
rect 225 -3466 577 -3462
rect 581 -3466 975 -3462
rect 979 -3466 1333 -3462
rect 1337 -3466 1617 -3462
rect -949 -3479 -909 -3475
rect -591 -3479 -551 -3475
rect -233 -3479 -193 -3475
rect 195 -3479 235 -3475
rect 551 -3479 591 -3475
rect 949 -3479 989 -3475
rect 1307 -3479 1347 -3475
rect 1633 -3514 1695 -3401
rect -1421 -3518 -1322 -3514
rect -1318 -3518 -918 -3514
rect -914 -3518 -560 -3514
rect -556 -3518 -202 -3514
rect -198 -3518 226 -3514
rect 230 -3518 582 -3514
rect 586 -3518 980 -3514
rect 984 -3518 1338 -3514
rect 1342 -3518 1695 -3514
rect -1495 -3550 -1255 -3546
rect -1251 -3550 -1238 -3546
rect -1234 -3550 -1198 -3546
rect -1194 -3550 -1177 -3546
rect -1173 -3550 -926 -3546
rect -922 -3550 -900 -3546
rect -896 -3550 -883 -3546
rect -879 -3550 -843 -3546
rect -839 -3550 -822 -3546
rect -818 -3550 -805 -3546
rect -801 -3550 -765 -3546
rect -761 -3550 -741 -3546
rect -737 -3550 -704 -3546
rect -700 -3550 -568 -3546
rect -564 -3550 -542 -3546
rect -538 -3550 -525 -3546
rect -521 -3550 -485 -3546
rect -481 -3550 -464 -3546
rect -460 -3550 -447 -3546
rect -443 -3550 -407 -3546
rect -403 -3550 -383 -3546
rect -379 -3550 -346 -3546
rect -342 -3550 -210 -3546
rect -206 -3550 -184 -3546
rect -180 -3550 -167 -3546
rect -163 -3550 -127 -3546
rect -123 -3550 -106 -3546
rect -102 -3550 -89 -3546
rect -85 -3550 -49 -3546
rect -45 -3550 -25 -3546
rect -21 -3550 12 -3546
rect 16 -3550 218 -3546
rect 222 -3550 244 -3546
rect 248 -3550 261 -3546
rect 265 -3550 301 -3546
rect 305 -3550 322 -3546
rect 326 -3550 339 -3546
rect 343 -3550 379 -3546
rect 383 -3550 403 -3546
rect 407 -3550 440 -3546
rect 444 -3550 574 -3546
rect 578 -3550 600 -3546
rect 604 -3550 617 -3546
rect 621 -3550 657 -3546
rect 661 -3550 678 -3546
rect 682 -3550 695 -3546
rect 699 -3550 735 -3546
rect 739 -3550 759 -3546
rect 763 -3550 796 -3546
rect 800 -3550 972 -3546
rect 976 -3550 998 -3546
rect 1002 -3550 1015 -3546
rect 1019 -3550 1055 -3546
rect 1059 -3550 1076 -3546
rect 1080 -3550 1093 -3546
rect 1097 -3550 1133 -3546
rect 1137 -3550 1157 -3546
rect 1161 -3550 1194 -3546
rect 1198 -3550 1330 -3546
rect 1334 -3550 1356 -3546
rect 1360 -3550 1373 -3546
rect 1377 -3550 1413 -3546
rect 1417 -3550 1434 -3546
rect 1438 -3550 1451 -3546
rect 1455 -3550 1491 -3546
rect 1495 -3550 1515 -3546
rect 1519 -3550 1552 -3546
rect 1556 -3550 1617 -3546
rect -1495 -3676 -1433 -3550
rect -926 -3554 -922 -3550
rect -900 -3554 -896 -3550
rect -883 -3554 -879 -3550
rect -843 -3554 -839 -3550
rect -822 -3554 -818 -3550
rect -805 -3554 -801 -3550
rect -765 -3554 -761 -3550
rect -741 -3554 -737 -3550
rect -704 -3554 -700 -3550
rect -568 -3554 -564 -3550
rect -542 -3554 -538 -3550
rect -525 -3554 -521 -3550
rect -485 -3554 -481 -3550
rect -464 -3554 -460 -3550
rect -447 -3554 -443 -3550
rect -407 -3554 -403 -3550
rect -383 -3554 -379 -3550
rect -346 -3554 -342 -3550
rect -210 -3554 -206 -3550
rect -184 -3554 -180 -3550
rect -167 -3554 -163 -3550
rect -127 -3554 -123 -3550
rect -106 -3554 -102 -3550
rect -89 -3554 -85 -3550
rect -49 -3554 -45 -3550
rect -25 -3554 -21 -3550
rect 12 -3554 16 -3550
rect 218 -3554 222 -3550
rect 244 -3554 248 -3550
rect 261 -3554 265 -3550
rect 301 -3554 305 -3550
rect 322 -3554 326 -3550
rect 339 -3554 343 -3550
rect 379 -3554 383 -3550
rect 403 -3554 407 -3550
rect 440 -3554 444 -3550
rect 574 -3554 578 -3550
rect 600 -3554 604 -3550
rect 617 -3554 621 -3550
rect 657 -3554 661 -3550
rect 678 -3554 682 -3550
rect 695 -3554 699 -3550
rect 735 -3554 739 -3550
rect 759 -3554 763 -3550
rect 796 -3554 800 -3550
rect 972 -3554 976 -3550
rect 998 -3554 1002 -3550
rect 1015 -3554 1019 -3550
rect 1055 -3554 1059 -3550
rect 1076 -3554 1080 -3550
rect 1093 -3554 1097 -3550
rect 1133 -3554 1137 -3550
rect 1157 -3554 1161 -3550
rect 1194 -3554 1198 -3550
rect 1330 -3554 1334 -3550
rect 1356 -3554 1360 -3550
rect 1373 -3554 1377 -3550
rect 1413 -3554 1417 -3550
rect 1434 -3554 1438 -3550
rect 1451 -3554 1455 -3550
rect 1491 -3554 1495 -3550
rect 1515 -3554 1519 -3550
rect 1552 -3554 1556 -3550
rect -920 -3569 -858 -3565
rect -854 -3569 -824 -3565
rect -776 -3569 -746 -3565
rect -562 -3569 -500 -3565
rect -496 -3569 -466 -3565
rect -418 -3569 -388 -3565
rect -204 -3569 -142 -3565
rect -138 -3569 -108 -3565
rect -60 -3569 -30 -3565
rect 224 -3569 286 -3565
rect 290 -3569 320 -3565
rect 368 -3569 398 -3565
rect 580 -3569 642 -3565
rect 646 -3569 676 -3565
rect 724 -3569 754 -3565
rect 978 -3569 1040 -3565
rect 1044 -3569 1074 -3565
rect 1122 -3569 1152 -3565
rect 1336 -3569 1398 -3565
rect 1402 -3569 1432 -3565
rect 1480 -3569 1510 -3565
rect -913 -3576 -882 -3572
rect -555 -3576 -524 -3572
rect -197 -3576 -166 -3572
rect 231 -3576 262 -3572
rect 587 -3576 618 -3572
rect 985 -3576 1016 -3572
rect 1343 -3576 1374 -3572
rect -931 -3583 -848 -3579
rect -809 -3583 -706 -3579
rect -573 -3583 -490 -3579
rect -451 -3583 -348 -3579
rect -215 -3583 -132 -3579
rect -93 -3583 10 -3579
rect 213 -3583 296 -3579
rect 335 -3583 438 -3579
rect 569 -3583 652 -3579
rect 691 -3583 794 -3579
rect 967 -3583 1050 -3579
rect 1089 -3583 1192 -3579
rect 1325 -3583 1408 -3579
rect 1447 -3583 1550 -3579
rect -949 -3590 -928 -3586
rect -894 -3590 -865 -3586
rect -861 -3590 -780 -3586
rect -691 -3590 -592 -3586
rect -585 -3590 -570 -3586
rect -536 -3590 -507 -3586
rect -503 -3590 -422 -3586
rect -333 -3589 -234 -3585
rect -596 -3594 -592 -3590
rect -238 -3594 -234 -3589
rect -227 -3590 -212 -3586
rect -178 -3590 -149 -3586
rect -145 -3590 -64 -3586
rect 25 -3590 194 -3586
rect 201 -3590 216 -3586
rect 250 -3590 279 -3586
rect 283 -3590 364 -3586
rect 453 -3590 550 -3586
rect 557 -3590 572 -3586
rect 606 -3590 635 -3586
rect 639 -3590 720 -3586
rect 809 -3590 948 -3586
rect 955 -3590 970 -3586
rect 1004 -3590 1033 -3586
rect 1037 -3590 1118 -3586
rect 1207 -3588 1300 -3584
rect 190 -3594 194 -3590
rect 546 -3594 550 -3590
rect 944 -3594 948 -3590
rect 1296 -3594 1300 -3588
rect 1307 -3590 1328 -3586
rect 1362 -3590 1391 -3586
rect 1395 -3590 1476 -3586
rect -1260 -3599 -1203 -3595
rect -1164 -3598 -902 -3594
rect -887 -3598 -804 -3594
rect -783 -3598 -689 -3594
rect -596 -3598 -544 -3594
rect -529 -3598 -446 -3594
rect -425 -3598 -331 -3594
rect -238 -3598 -186 -3594
rect -171 -3598 -88 -3594
rect -67 -3598 27 -3594
rect 190 -3598 242 -3594
rect 257 -3598 340 -3594
rect 361 -3598 455 -3594
rect 546 -3598 598 -3594
rect 613 -3598 696 -3594
rect 717 -3598 811 -3594
rect 944 -3598 996 -3594
rect 1011 -3598 1094 -3594
rect 1115 -3598 1209 -3594
rect 1296 -3598 1354 -3594
rect 1369 -3598 1452 -3594
rect 1473 -3598 1567 -3594
rect -1266 -3606 -1253 -3602
rect -1249 -3606 -1213 -3602
rect -1209 -3606 -1193 -3602
rect -943 -3605 -924 -3601
rect -905 -3605 -776 -3601
rect -591 -3605 -566 -3601
rect -547 -3605 -418 -3601
rect -233 -3605 -208 -3601
rect -189 -3605 -60 -3601
rect 195 -3605 220 -3601
rect 239 -3605 368 -3601
rect 551 -3605 576 -3601
rect 595 -3605 724 -3601
rect 949 -3605 974 -3601
rect 993 -3605 1122 -3601
rect 1313 -3605 1332 -3601
rect 1351 -3605 1480 -3601
rect -1309 -3613 -1257 -3609
rect -1253 -3613 -1227 -3609
rect -1223 -3613 -1179 -3609
rect -898 -3612 -794 -3608
rect -790 -3612 -760 -3608
rect -540 -3612 -436 -3608
rect -432 -3612 -402 -3608
rect -182 -3612 -78 -3608
rect -74 -3612 -44 -3608
rect 246 -3612 350 -3608
rect 354 -3612 384 -3608
rect 602 -3612 706 -3608
rect 710 -3612 740 -3608
rect 1000 -3612 1104 -3608
rect 1108 -3612 1138 -3608
rect 1358 -3612 1462 -3608
rect 1466 -3612 1496 -3608
rect -1216 -3620 -1162 -3616
rect -924 -3619 -872 -3615
rect -868 -3619 -838 -3615
rect -566 -3619 -514 -3615
rect -510 -3619 -480 -3615
rect -208 -3619 -156 -3615
rect -152 -3619 -122 -3615
rect 220 -3619 272 -3615
rect 276 -3619 306 -3615
rect 576 -3619 628 -3615
rect 632 -3619 662 -3615
rect 974 -3619 1026 -3615
rect 1030 -3619 1060 -3615
rect 1332 -3619 1384 -3615
rect 1388 -3619 1418 -3615
rect -1234 -3627 -1202 -3623
rect -879 -3627 -847 -3623
rect -883 -3630 -879 -3627
rect -847 -3630 -843 -3627
rect -801 -3627 -769 -3623
rect -805 -3630 -801 -3627
rect -769 -3630 -765 -3627
rect -521 -3627 -489 -3623
rect -525 -3630 -521 -3627
rect -489 -3630 -485 -3627
rect -443 -3627 -411 -3623
rect -447 -3630 -443 -3627
rect -411 -3630 -407 -3627
rect -163 -3627 -131 -3623
rect -167 -3630 -163 -3627
rect -131 -3630 -127 -3627
rect -85 -3627 -53 -3623
rect -89 -3630 -85 -3627
rect -53 -3630 -49 -3627
rect 265 -3627 297 -3623
rect 261 -3630 265 -3627
rect 297 -3630 301 -3627
rect 343 -3627 375 -3623
rect 339 -3630 343 -3627
rect 375 -3630 379 -3627
rect 621 -3627 653 -3623
rect 617 -3630 621 -3627
rect 653 -3630 657 -3627
rect 699 -3627 731 -3623
rect 695 -3630 699 -3627
rect 731 -3630 735 -3627
rect 1019 -3627 1051 -3623
rect 1015 -3630 1019 -3627
rect 1051 -3630 1055 -3627
rect 1097 -3627 1129 -3623
rect 1093 -3630 1097 -3627
rect 1129 -3630 1133 -3627
rect 1377 -3627 1409 -3623
rect 1373 -3630 1377 -3627
rect 1409 -3630 1413 -3627
rect 1455 -3627 1487 -3623
rect 1451 -3630 1455 -3627
rect 1487 -3630 1491 -3627
rect -926 -3638 -922 -3634
rect -900 -3638 -896 -3634
rect -857 -3638 -853 -3634
rect -822 -3638 -818 -3634
rect -778 -3638 -774 -3634
rect -761 -3638 -757 -3634
rect -725 -3638 -721 -3634
rect -704 -3638 -700 -3634
rect -568 -3638 -564 -3634
rect -542 -3638 -538 -3634
rect -499 -3638 -495 -3634
rect -464 -3638 -460 -3634
rect -420 -3638 -416 -3634
rect -403 -3638 -399 -3634
rect -367 -3638 -363 -3634
rect -346 -3638 -342 -3634
rect -210 -3638 -206 -3634
rect -184 -3638 -180 -3634
rect -141 -3638 -137 -3634
rect -106 -3638 -102 -3634
rect -62 -3638 -58 -3634
rect -45 -3638 -41 -3634
rect -9 -3638 -5 -3634
rect 12 -3638 16 -3634
rect 218 -3638 222 -3634
rect 244 -3638 248 -3634
rect 287 -3638 291 -3634
rect 322 -3638 326 -3634
rect 366 -3638 370 -3634
rect 383 -3638 387 -3634
rect 419 -3638 423 -3634
rect 440 -3638 444 -3634
rect 574 -3638 578 -3634
rect 600 -3638 604 -3634
rect 643 -3638 647 -3634
rect 678 -3638 682 -3634
rect 722 -3638 726 -3634
rect 739 -3638 743 -3634
rect 775 -3638 779 -3634
rect 796 -3638 800 -3634
rect 972 -3638 976 -3634
rect 998 -3638 1002 -3634
rect 1041 -3638 1045 -3634
rect 1076 -3638 1080 -3634
rect 1120 -3638 1124 -3634
rect 1137 -3638 1141 -3634
rect 1173 -3638 1177 -3634
rect 1194 -3638 1198 -3634
rect 1330 -3638 1334 -3634
rect 1356 -3638 1360 -3634
rect 1399 -3638 1403 -3634
rect 1434 -3638 1438 -3634
rect 1478 -3638 1482 -3634
rect 1495 -3638 1499 -3634
rect 1531 -3638 1535 -3634
rect 1552 -3638 1556 -3634
rect 1633 -3638 1695 -3518
rect -1421 -3642 -1255 -3638
rect -1251 -3642 -1211 -3638
rect -1207 -3642 -1177 -3638
rect -1173 -3642 -926 -3638
rect -922 -3642 -900 -3638
rect -896 -3642 -857 -3638
rect -853 -3642 -822 -3638
rect -818 -3642 -778 -3638
rect -774 -3642 -761 -3638
rect -757 -3642 -725 -3638
rect -721 -3642 -704 -3638
rect -700 -3642 -568 -3638
rect -564 -3642 -542 -3638
rect -538 -3642 -499 -3638
rect -495 -3642 -464 -3638
rect -460 -3642 -420 -3638
rect -416 -3642 -403 -3638
rect -399 -3642 -367 -3638
rect -363 -3642 -346 -3638
rect -342 -3642 -210 -3638
rect -206 -3642 -184 -3638
rect -180 -3642 -141 -3638
rect -137 -3642 -106 -3638
rect -102 -3642 -62 -3638
rect -58 -3642 -45 -3638
rect -41 -3642 -9 -3638
rect -5 -3642 12 -3638
rect 16 -3642 218 -3638
rect 222 -3642 244 -3638
rect 248 -3642 287 -3638
rect 291 -3642 322 -3638
rect 326 -3642 366 -3638
rect 370 -3642 383 -3638
rect 387 -3642 419 -3638
rect 423 -3642 440 -3638
rect 444 -3642 574 -3638
rect 578 -3642 600 -3638
rect 604 -3642 643 -3638
rect 647 -3642 678 -3638
rect 682 -3642 722 -3638
rect 726 -3642 739 -3638
rect 743 -3642 775 -3638
rect 779 -3642 796 -3638
rect 800 -3642 972 -3638
rect 976 -3642 998 -3638
rect 1002 -3642 1041 -3638
rect 1045 -3642 1076 -3638
rect 1080 -3642 1120 -3638
rect 1124 -3642 1137 -3638
rect 1141 -3642 1173 -3638
rect 1177 -3642 1194 -3638
rect 1198 -3642 1330 -3638
rect 1334 -3642 1356 -3638
rect 1360 -3642 1399 -3638
rect 1403 -3642 1434 -3638
rect 1438 -3642 1478 -3638
rect 1482 -3642 1495 -3638
rect 1499 -3642 1531 -3638
rect 1535 -3642 1552 -3638
rect 1556 -3642 1695 -3638
rect -1272 -3649 -689 -3645
rect -585 -3649 27 -3645
rect 201 -3649 811 -3645
rect 955 -3649 1567 -3645
rect -1266 -3656 -1162 -3652
rect -943 -3656 -331 -3652
rect -227 -3656 455 -3652
rect 557 -3656 1209 -3652
rect 1313 -3656 1561 -3652
rect -1495 -3680 -1255 -3676
rect -1251 -3680 -1238 -3676
rect -1234 -3680 -1218 -3676
rect -1214 -3680 -1197 -3676
rect -1193 -3680 -1176 -3676
rect -1172 -3680 -1155 -3676
rect -1151 -3680 -1134 -3676
rect -1130 -3680 -1113 -3676
rect -1109 -3680 -1092 -3676
rect -1088 -3680 -1072 -3676
rect -1068 -3680 -926 -3676
rect -922 -3680 -909 -3676
rect -905 -3680 -889 -3676
rect -885 -3680 -868 -3676
rect -864 -3680 -847 -3676
rect -843 -3680 -826 -3676
rect -822 -3680 -805 -3676
rect -801 -3680 -784 -3676
rect -780 -3680 -763 -3676
rect -759 -3680 -743 -3676
rect -739 -3680 -568 -3676
rect -564 -3680 -551 -3676
rect -547 -3680 -531 -3676
rect -527 -3680 -510 -3676
rect -506 -3680 -489 -3676
rect -485 -3680 -468 -3676
rect -464 -3680 -447 -3676
rect -443 -3680 -426 -3676
rect -422 -3680 -405 -3676
rect -401 -3680 -385 -3676
rect -381 -3680 -210 -3676
rect -206 -3680 -193 -3676
rect -189 -3680 -173 -3676
rect -169 -3680 -152 -3676
rect -148 -3680 -131 -3676
rect -127 -3680 -110 -3676
rect -106 -3680 -89 -3676
rect -85 -3680 -68 -3676
rect -64 -3680 -47 -3676
rect -43 -3680 -27 -3676
rect -23 -3680 1617 -3676
rect -1495 -3791 -1433 -3680
rect -1233 -3728 -1199 -3724
rect -1135 -3728 -1115 -3724
rect -1100 -3728 -931 -3724
rect -904 -3728 -870 -3724
rect -806 -3728 -786 -3724
rect -771 -3728 -573 -3724
rect -546 -3728 -512 -3724
rect -448 -3728 -428 -3724
rect -413 -3728 -215 -3724
rect -188 -3728 -154 -3724
rect -90 -3728 -70 -3724
rect -55 -3728 -19 -3724
rect -935 -3732 -931 -3728
rect -577 -3732 -573 -3728
rect -219 -3732 -215 -3728
rect -1266 -3736 -1257 -3732
rect -1253 -3736 -1223 -3732
rect -1202 -3736 -1171 -3732
rect -1142 -3736 -1111 -3732
rect -1100 -3736 -1073 -3732
rect -935 -3736 -928 -3732
rect -924 -3736 -894 -3732
rect -873 -3736 -842 -3732
rect -813 -3736 -782 -3732
rect -771 -3736 -744 -3732
rect -577 -3736 -570 -3732
rect -566 -3736 -536 -3732
rect -515 -3736 -484 -3732
rect -455 -3736 -424 -3732
rect -413 -3736 -386 -3732
rect -219 -3736 -212 -3732
rect -208 -3736 -178 -3732
rect -157 -3736 -126 -3732
rect -97 -3736 -66 -3732
rect -55 -3736 -28 -3732
rect -1260 -3743 -1213 -3739
rect -1177 -3743 -1164 -3739
rect -1160 -3743 -1129 -3739
rect -1093 -3743 -1080 -3739
rect -1076 -3743 -1064 -3739
rect -931 -3743 -884 -3739
rect -848 -3743 -835 -3739
rect -831 -3743 -800 -3739
rect -764 -3743 -751 -3739
rect -747 -3743 -735 -3739
rect -573 -3743 -526 -3739
rect -490 -3743 -477 -3739
rect -473 -3743 -442 -3739
rect -406 -3743 -393 -3739
rect -389 -3743 -377 -3739
rect -215 -3743 -168 -3739
rect -132 -3743 -119 -3739
rect -115 -3743 -84 -3739
rect -48 -3743 -35 -3739
rect -31 -3743 -19 -3739
rect -1277 -3750 -1253 -3746
rect -1249 -3750 -1139 -3746
rect -1118 -3750 -1087 -3746
rect -941 -3750 -940 -3746
rect -936 -3750 -924 -3746
rect -920 -3750 -810 -3746
rect -789 -3750 -758 -3746
rect -581 -3750 -580 -3746
rect -576 -3750 -566 -3746
rect -562 -3750 -452 -3746
rect -431 -3750 -400 -3746
rect -221 -3750 -208 -3746
rect -204 -3750 -94 -3746
rect -73 -3750 -42 -3746
rect -1218 -3757 -1195 -3753
rect -1176 -3757 -1157 -3753
rect -889 -3757 -866 -3753
rect -847 -3757 -828 -3753
rect -531 -3757 -508 -3753
rect -489 -3757 -470 -3753
rect -173 -3757 -150 -3753
rect -131 -3757 -112 -3753
rect 1633 -3768 1695 -3642
rect -1421 -3772 -1255 -3768
rect -1251 -3772 -1238 -3768
rect -1234 -3772 -1197 -3768
rect -1193 -3772 -1155 -3768
rect -1151 -3772 -1113 -3768
rect -1109 -3772 -1072 -3768
rect -1068 -3772 -926 -3768
rect -922 -3772 -909 -3768
rect -905 -3772 -868 -3768
rect -864 -3772 -826 -3768
rect -822 -3772 -784 -3768
rect -780 -3772 -743 -3768
rect -739 -3772 -568 -3768
rect -564 -3772 -551 -3768
rect -547 -3772 -510 -3768
rect -506 -3772 -468 -3768
rect -464 -3772 -426 -3768
rect -422 -3772 -385 -3768
rect -381 -3772 -210 -3768
rect -206 -3772 -193 -3768
rect -189 -3772 -152 -3768
rect -148 -3772 -110 -3768
rect -106 -3772 -68 -3768
rect -64 -3772 -27 -3768
rect -23 -3772 1695 -3768
rect -1495 -3795 68 -3791
rect 72 -3795 1618 -3791
rect -1607 -3851 -1598 -3837
rect -1495 -3907 -1433 -3795
rect 80 -3846 92 -3842
rect 1633 -3883 1695 -3772
rect -1421 -3887 68 -3883
rect 72 -3887 1695 -3883
rect -1495 -3911 -1255 -3907
rect -1251 -3911 -1238 -3907
rect -1234 -3911 -1218 -3907
rect -1214 -3911 -1197 -3907
rect -1193 -3911 -1176 -3907
rect -1172 -3911 -1155 -3907
rect -1151 -3911 -1134 -3907
rect -1130 -3911 -1113 -3907
rect -1109 -3911 -1092 -3907
rect -1088 -3911 -1072 -3907
rect -1068 -3911 -926 -3907
rect -922 -3911 -909 -3907
rect -905 -3911 -889 -3907
rect -885 -3911 -868 -3907
rect -864 -3911 -847 -3907
rect -843 -3911 -826 -3907
rect -822 -3911 -805 -3907
rect -801 -3911 -784 -3907
rect -780 -3911 -763 -3907
rect -759 -3911 -743 -3907
rect -739 -3911 -568 -3907
rect -564 -3911 -551 -3907
rect -547 -3911 -531 -3907
rect -527 -3911 -510 -3907
rect -506 -3911 -489 -3907
rect -485 -3911 -468 -3907
rect -464 -3911 -447 -3907
rect -443 -3911 -426 -3907
rect -422 -3911 -405 -3907
rect -401 -3911 -385 -3907
rect -381 -3911 -210 -3907
rect -206 -3911 -193 -3907
rect -189 -3911 -173 -3907
rect -169 -3911 -152 -3907
rect -148 -3911 -131 -3907
rect -127 -3911 -110 -3907
rect -106 -3911 -89 -3907
rect -85 -3911 -68 -3907
rect -64 -3911 -47 -3907
rect -43 -3911 -27 -3907
rect -23 -3911 218 -3907
rect 222 -3911 235 -3907
rect 239 -3911 255 -3907
rect 259 -3911 276 -3907
rect 280 -3911 297 -3907
rect 301 -3911 318 -3907
rect 322 -3911 339 -3907
rect 343 -3911 360 -3907
rect 364 -3911 381 -3907
rect 385 -3911 401 -3907
rect 405 -3911 574 -3907
rect 578 -3911 591 -3907
rect 595 -3911 611 -3907
rect 615 -3911 632 -3907
rect 636 -3911 653 -3907
rect 657 -3911 674 -3907
rect 678 -3911 695 -3907
rect 699 -3911 716 -3907
rect 720 -3911 737 -3907
rect 741 -3911 757 -3907
rect 761 -3911 972 -3907
rect 976 -3911 989 -3907
rect 993 -3911 1009 -3907
rect 1013 -3911 1030 -3907
rect 1034 -3911 1051 -3907
rect 1055 -3911 1072 -3907
rect 1076 -3911 1093 -3907
rect 1097 -3911 1114 -3907
rect 1118 -3911 1135 -3907
rect 1139 -3911 1155 -3907
rect 1159 -3911 1330 -3907
rect 1334 -3911 1347 -3907
rect 1351 -3911 1367 -3907
rect 1371 -3911 1388 -3907
rect 1392 -3911 1409 -3907
rect 1413 -3911 1430 -3907
rect 1434 -3911 1451 -3907
rect 1455 -3911 1472 -3907
rect 1476 -3911 1493 -3907
rect 1497 -3911 1513 -3907
rect 1517 -3911 1617 -3907
rect -1495 -4032 -1433 -3911
rect -1233 -3959 -1199 -3955
rect -1135 -3959 -1115 -3955
rect -1100 -3959 -1066 -3955
rect -904 -3959 -870 -3955
rect -806 -3959 -786 -3955
rect -771 -3959 -737 -3955
rect -546 -3959 -512 -3955
rect -448 -3959 -428 -3955
rect -413 -3959 -379 -3955
rect -188 -3959 -154 -3955
rect -90 -3959 -70 -3955
rect -55 -3959 -21 -3955
rect 240 -3959 274 -3955
rect 338 -3959 358 -3955
rect 373 -3959 407 -3955
rect 596 -3959 630 -3955
rect 694 -3959 714 -3955
rect 729 -3959 763 -3955
rect 994 -3959 1028 -3955
rect 1092 -3959 1112 -3955
rect 1127 -3959 1161 -3955
rect 1352 -3959 1386 -3955
rect 1450 -3959 1470 -3955
rect 1485 -3959 1519 -3955
rect -1272 -3967 -1257 -3963
rect -1253 -3967 -1223 -3963
rect -1202 -3967 -1171 -3963
rect -1142 -3967 -1111 -3963
rect -1100 -3967 -1073 -3963
rect -943 -3967 -928 -3963
rect -924 -3967 -894 -3963
rect -873 -3967 -842 -3963
rect -813 -3967 -782 -3963
rect -771 -3967 -744 -3963
rect -585 -3967 -570 -3963
rect -566 -3967 -536 -3963
rect -515 -3967 -484 -3963
rect -455 -3967 -424 -3963
rect -413 -3967 -386 -3963
rect -227 -3967 -212 -3963
rect -208 -3967 -178 -3963
rect -157 -3967 -126 -3963
rect -97 -3967 -66 -3963
rect -55 -3967 -28 -3963
rect 201 -3967 216 -3963
rect 220 -3967 250 -3963
rect 271 -3967 302 -3963
rect 331 -3967 362 -3963
rect 373 -3967 400 -3963
rect 557 -3967 572 -3963
rect 576 -3967 606 -3963
rect 627 -3967 658 -3963
rect 687 -3967 718 -3963
rect 729 -3967 756 -3963
rect 955 -3967 970 -3963
rect 974 -3967 1004 -3963
rect 1025 -3967 1056 -3963
rect 1085 -3967 1116 -3963
rect 1127 -3967 1154 -3963
rect 1313 -3967 1328 -3963
rect 1332 -3967 1362 -3963
rect 1383 -3967 1414 -3963
rect 1443 -3967 1474 -3963
rect 1485 -3967 1512 -3963
rect -1260 -3974 -1213 -3970
rect -1177 -3974 -1164 -3970
rect -1160 -3974 -1129 -3970
rect -1093 -3974 -1080 -3970
rect -1076 -3974 -1064 -3970
rect -931 -3974 -884 -3970
rect -848 -3974 -835 -3970
rect -831 -3974 -800 -3970
rect -764 -3974 -751 -3970
rect -747 -3974 -735 -3970
rect -573 -3974 -526 -3970
rect -490 -3974 -477 -3970
rect -473 -3974 -442 -3970
rect -406 -3974 -393 -3970
rect -389 -3974 -377 -3970
rect -215 -3974 -168 -3970
rect -132 -3974 -119 -3970
rect -115 -3974 -84 -3970
rect -48 -3974 -35 -3970
rect -31 -3974 -19 -3970
rect 213 -3974 260 -3970
rect 296 -3974 309 -3970
rect 313 -3974 344 -3970
rect 380 -3974 393 -3970
rect 397 -3974 409 -3970
rect 569 -3974 616 -3970
rect 652 -3974 665 -3970
rect 669 -3974 700 -3970
rect 736 -3974 749 -3970
rect 753 -3974 765 -3970
rect 967 -3974 1014 -3970
rect 1050 -3974 1063 -3970
rect 1067 -3974 1098 -3970
rect 1134 -3974 1147 -3970
rect 1151 -3974 1163 -3970
rect 1325 -3974 1372 -3970
rect 1408 -3974 1421 -3970
rect 1425 -3974 1456 -3970
rect 1492 -3974 1505 -3970
rect 1509 -3974 1521 -3970
rect -1268 -3981 -1253 -3977
rect -1249 -3981 -1139 -3977
rect -1118 -3981 -1087 -3977
rect -937 -3981 -924 -3977
rect -920 -3981 -810 -3977
rect -789 -3981 -758 -3977
rect -579 -3981 -566 -3977
rect -562 -3981 -452 -3977
rect -431 -3981 -400 -3977
rect -222 -3981 -208 -3977
rect -204 -3981 -94 -3977
rect -73 -3981 -42 -3977
rect 208 -3981 220 -3977
rect 224 -3981 334 -3977
rect 355 -3981 386 -3977
rect 564 -3981 576 -3977
rect 580 -3981 690 -3977
rect 711 -3981 742 -3977
rect 949 -3981 974 -3977
rect 978 -3981 1088 -3977
rect 1109 -3981 1140 -3977
rect 1319 -3981 1332 -3977
rect 1336 -3981 1446 -3977
rect 1467 -3981 1498 -3977
rect -1218 -3988 -1195 -3984
rect -1176 -3988 -1157 -3984
rect -889 -3988 -866 -3984
rect -847 -3988 -828 -3984
rect -531 -3988 -508 -3984
rect -489 -3988 -470 -3984
rect -173 -3988 -150 -3984
rect -131 -3988 -112 -3984
rect 255 -3988 278 -3984
rect 297 -3988 316 -3984
rect 611 -3988 634 -3984
rect 653 -3988 672 -3984
rect 1009 -3988 1032 -3984
rect 1051 -3988 1070 -3984
rect 1367 -3988 1390 -3984
rect 1409 -3988 1428 -3984
rect 1633 -3999 1695 -3887
rect -1421 -4003 -1255 -3999
rect -1251 -4003 -1238 -3999
rect -1234 -4003 -1197 -3999
rect -1193 -4003 -1155 -3999
rect -1151 -4003 -1113 -3999
rect -1109 -4003 -1072 -3999
rect -1068 -4003 -926 -3999
rect -922 -4003 -909 -3999
rect -905 -4003 -868 -3999
rect -864 -4003 -826 -3999
rect -822 -4003 -784 -3999
rect -780 -4003 -743 -3999
rect -739 -4003 -568 -3999
rect -564 -4003 -551 -3999
rect -547 -4003 -510 -3999
rect -506 -4003 -468 -3999
rect -464 -4003 -426 -3999
rect -422 -4003 -385 -3999
rect -381 -4003 -210 -3999
rect -206 -4003 -193 -3999
rect -189 -4003 -152 -3999
rect -148 -4003 -110 -3999
rect -106 -4003 -68 -3999
rect -64 -4003 -27 -3999
rect -23 -4003 218 -3999
rect 222 -4003 235 -3999
rect 239 -4003 276 -3999
rect 280 -4003 318 -3999
rect 322 -4003 360 -3999
rect 364 -4003 401 -3999
rect 405 -4003 574 -3999
rect 578 -4003 591 -3999
rect 595 -4003 632 -3999
rect 636 -4003 674 -3999
rect 678 -4003 716 -3999
rect 720 -4003 757 -3999
rect 761 -4003 972 -3999
rect 976 -4003 989 -3999
rect 993 -4003 1030 -3999
rect 1034 -4003 1072 -3999
rect 1076 -4003 1114 -3999
rect 1118 -4003 1155 -3999
rect 1159 -4003 1330 -3999
rect 1334 -4003 1347 -3999
rect 1351 -4003 1388 -3999
rect 1392 -4003 1430 -3999
rect 1434 -4003 1472 -3999
rect 1476 -4003 1513 -3999
rect 1517 -4003 1695 -3999
rect -1266 -4010 -1066 -4006
rect -943 -4011 -737 -4007
rect -585 -4010 -379 -4006
rect -227 -4010 -21 -4006
rect 201 -4010 407 -4006
rect 557 -4011 763 -4007
rect 955 -4010 1161 -4006
rect 1313 -4010 1519 -4006
rect -1495 -4036 -1255 -4032
rect -1251 -4036 -1238 -4032
rect -1234 -4036 -1218 -4032
rect -1214 -4036 -1197 -4032
rect -1193 -4036 -1176 -4032
rect -1172 -4036 -1155 -4032
rect -1151 -4036 -1134 -4032
rect -1130 -4036 -1113 -4032
rect -1109 -4036 -1092 -4032
rect -1088 -4036 -1072 -4032
rect -1068 -4036 -926 -4032
rect -922 -4036 -909 -4032
rect -905 -4036 -889 -4032
rect -885 -4036 -868 -4032
rect -864 -4036 -847 -4032
rect -843 -4036 -826 -4032
rect -822 -4036 -805 -4032
rect -801 -4036 -784 -4032
rect -780 -4036 -763 -4032
rect -759 -4036 -743 -4032
rect -739 -4036 -568 -4032
rect -564 -4036 -551 -4032
rect -547 -4036 -531 -4032
rect -527 -4036 -510 -4032
rect -506 -4036 -489 -4032
rect -485 -4036 -468 -4032
rect -464 -4036 -447 -4032
rect -443 -4036 -426 -4032
rect -422 -4036 -405 -4032
rect -401 -4036 -385 -4032
rect -381 -4036 -210 -4032
rect -206 -4036 -193 -4032
rect -189 -4036 -173 -4032
rect -169 -4036 -152 -4032
rect -148 -4036 -131 -4032
rect -127 -4036 -110 -4032
rect -106 -4036 -89 -4032
rect -85 -4036 -68 -4032
rect -64 -4036 -47 -4032
rect -43 -4036 -27 -4032
rect -23 -4036 218 -4032
rect 222 -4036 235 -4032
rect 239 -4036 255 -4032
rect 259 -4036 276 -4032
rect 280 -4036 297 -4032
rect 301 -4036 318 -4032
rect 322 -4036 339 -4032
rect 343 -4036 360 -4032
rect 364 -4036 381 -4032
rect 385 -4036 401 -4032
rect 405 -4036 574 -4032
rect 578 -4036 591 -4032
rect 595 -4036 611 -4032
rect 615 -4036 632 -4032
rect 636 -4036 653 -4032
rect 657 -4036 674 -4032
rect 678 -4036 695 -4032
rect 699 -4036 716 -4032
rect 720 -4036 737 -4032
rect 741 -4036 757 -4032
rect 761 -4036 972 -4032
rect 976 -4036 989 -4032
rect 993 -4036 1009 -4032
rect 1013 -4036 1030 -4032
rect 1034 -4036 1051 -4032
rect 1055 -4036 1072 -4032
rect 1076 -4036 1093 -4032
rect 1097 -4036 1114 -4032
rect 1118 -4036 1135 -4032
rect 1139 -4036 1155 -4032
rect 1159 -4036 1330 -4032
rect 1334 -4036 1347 -4032
rect 1351 -4036 1367 -4032
rect 1371 -4036 1388 -4032
rect 1392 -4036 1409 -4032
rect 1413 -4036 1430 -4032
rect 1434 -4036 1451 -4032
rect 1455 -4036 1472 -4032
rect 1476 -4036 1493 -4032
rect 1497 -4036 1513 -4032
rect 1517 -4036 1617 -4032
rect -1495 -4156 -1433 -4036
rect -1233 -4084 -1199 -4080
rect -1135 -4084 -1115 -4080
rect -1100 -4084 -1066 -4080
rect -904 -4084 -870 -4080
rect -806 -4084 -786 -4080
rect -771 -4084 -737 -4080
rect -546 -4084 -512 -4080
rect -448 -4084 -428 -4080
rect -413 -4084 -379 -4080
rect -188 -4084 -154 -4080
rect -90 -4084 -70 -4080
rect -55 -4084 -15 -4080
rect 240 -4084 274 -4080
rect 338 -4084 358 -4080
rect 373 -4084 407 -4080
rect 596 -4084 630 -4080
rect 694 -4084 714 -4080
rect 729 -4084 763 -4080
rect 994 -4084 1028 -4080
rect 1092 -4084 1112 -4080
rect 1127 -4084 1161 -4080
rect 1352 -4084 1386 -4080
rect 1450 -4084 1470 -4080
rect 1485 -4084 1519 -4080
rect -1345 -4092 -1257 -4088
rect -1253 -4092 -1223 -4088
rect -1202 -4092 -1171 -4088
rect -1142 -4092 -1111 -4088
rect -1100 -4092 -1073 -4088
rect -937 -4092 -928 -4088
rect -924 -4092 -894 -4088
rect -873 -4092 -842 -4088
rect -813 -4092 -782 -4088
rect -771 -4092 -744 -4088
rect -579 -4092 -570 -4088
rect -566 -4092 -536 -4088
rect -515 -4092 -484 -4088
rect -455 -4092 -424 -4088
rect -413 -4092 -386 -4088
rect -221 -4092 -212 -4088
rect -208 -4092 -178 -4088
rect -157 -4092 -126 -4088
rect -97 -4092 -66 -4088
rect -55 -4092 -28 -4088
rect 207 -4092 216 -4088
rect 220 -4092 250 -4088
rect 271 -4092 302 -4088
rect 331 -4092 362 -4088
rect 373 -4092 400 -4088
rect 563 -4092 572 -4088
rect 576 -4092 606 -4088
rect 627 -4092 658 -4088
rect 687 -4092 718 -4088
rect 729 -4092 756 -4088
rect 961 -4092 970 -4088
rect 974 -4092 1004 -4088
rect 1025 -4092 1056 -4088
rect 1085 -4092 1116 -4088
rect 1127 -4092 1154 -4088
rect 1319 -4092 1328 -4088
rect 1332 -4092 1362 -4088
rect 1383 -4092 1414 -4088
rect 1443 -4092 1474 -4088
rect 1485 -4092 1512 -4088
rect -1260 -4099 -1213 -4095
rect -1177 -4099 -1164 -4095
rect -1160 -4099 -1129 -4095
rect -1093 -4099 -1080 -4095
rect -1076 -4099 -1064 -4095
rect -931 -4099 -884 -4095
rect -848 -4099 -835 -4095
rect -831 -4099 -800 -4095
rect -764 -4099 -751 -4095
rect -747 -4099 -735 -4095
rect -573 -4099 -526 -4095
rect -490 -4099 -477 -4095
rect -473 -4099 -442 -4095
rect -406 -4099 -393 -4095
rect -389 -4099 -377 -4095
rect -215 -4099 -168 -4095
rect -132 -4099 -119 -4095
rect -115 -4099 -84 -4095
rect -48 -4099 -35 -4095
rect -31 -4099 -19 -4095
rect 213 -4099 260 -4095
rect 296 -4099 309 -4095
rect 313 -4099 344 -4095
rect 380 -4099 393 -4095
rect 397 -4099 409 -4095
rect 569 -4099 616 -4095
rect 652 -4099 665 -4095
rect 669 -4099 700 -4095
rect 736 -4099 749 -4095
rect 753 -4099 765 -4095
rect 967 -4099 1014 -4095
rect 1050 -4099 1063 -4095
rect 1067 -4099 1098 -4095
rect 1134 -4099 1147 -4095
rect 1151 -4099 1163 -4095
rect 1325 -4099 1372 -4095
rect 1408 -4099 1421 -4095
rect 1425 -4099 1456 -4095
rect 1492 -4099 1505 -4095
rect 1509 -4099 1521 -4095
rect -1273 -4106 -1272 -4102
rect -1268 -4106 -1253 -4102
rect -1249 -4106 -1139 -4102
rect -1118 -4106 -1087 -4102
rect -937 -4106 -924 -4102
rect -920 -4106 -810 -4102
rect -789 -4106 -758 -4102
rect -584 -4106 -583 -4102
rect -579 -4106 -566 -4102
rect -562 -4106 -452 -4102
rect -431 -4106 -400 -4102
rect -227 -4106 -226 -4102
rect -222 -4106 -208 -4102
rect -204 -4106 -94 -4102
rect -73 -4106 -42 -4102
rect 208 -4106 220 -4102
rect 224 -4106 334 -4102
rect 355 -4106 386 -4102
rect 564 -4106 576 -4102
rect 580 -4106 690 -4102
rect 711 -4106 742 -4102
rect 944 -4106 945 -4102
rect 949 -4106 974 -4102
rect 978 -4106 1088 -4102
rect 1109 -4106 1140 -4102
rect 1319 -4106 1332 -4102
rect 1336 -4106 1446 -4102
rect 1467 -4106 1498 -4102
rect -1218 -4113 -1195 -4109
rect -1176 -4113 -1157 -4109
rect -889 -4113 -866 -4109
rect -847 -4113 -828 -4109
rect -531 -4113 -508 -4109
rect -489 -4113 -470 -4109
rect -173 -4113 -150 -4109
rect -131 -4113 -112 -4109
rect 255 -4113 278 -4109
rect 297 -4113 316 -4109
rect 611 -4113 634 -4109
rect 653 -4113 672 -4109
rect 1009 -4113 1032 -4109
rect 1051 -4113 1070 -4109
rect 1367 -4113 1390 -4109
rect 1409 -4113 1428 -4109
rect 1633 -4124 1695 -4003
rect -1421 -4128 -1255 -4124
rect -1251 -4128 -1238 -4124
rect -1234 -4128 -1197 -4124
rect -1193 -4128 -1155 -4124
rect -1151 -4128 -1113 -4124
rect -1109 -4128 -1072 -4124
rect -1068 -4128 -926 -4124
rect -922 -4128 -909 -4124
rect -905 -4128 -868 -4124
rect -864 -4128 -826 -4124
rect -822 -4128 -784 -4124
rect -780 -4128 -743 -4124
rect -739 -4128 -568 -4124
rect -564 -4128 -551 -4124
rect -547 -4128 -510 -4124
rect -506 -4128 -468 -4124
rect -464 -4128 -426 -4124
rect -422 -4128 -385 -4124
rect -381 -4128 -210 -4124
rect -206 -4128 -193 -4124
rect -189 -4128 -152 -4124
rect -148 -4128 -110 -4124
rect -106 -4128 -68 -4124
rect -64 -4128 -27 -4124
rect -23 -4128 218 -4124
rect 222 -4128 235 -4124
rect 239 -4128 276 -4124
rect 280 -4128 318 -4124
rect 322 -4128 360 -4124
rect 364 -4128 401 -4124
rect 405 -4128 574 -4124
rect 578 -4128 591 -4124
rect 595 -4128 632 -4124
rect 636 -4128 674 -4124
rect 678 -4128 716 -4124
rect 720 -4128 757 -4124
rect 761 -4128 972 -4124
rect 976 -4128 989 -4124
rect 993 -4128 1030 -4124
rect 1034 -4128 1072 -4124
rect 1076 -4128 1114 -4124
rect 1118 -4128 1155 -4124
rect 1159 -4128 1330 -4124
rect 1334 -4128 1347 -4124
rect 1351 -4128 1388 -4124
rect 1392 -4128 1430 -4124
rect 1434 -4128 1472 -4124
rect 1476 -4128 1513 -4124
rect 1517 -4128 1695 -4124
rect -1495 -4160 -1255 -4156
rect -1251 -4160 -1238 -4156
rect -1234 -4160 -1218 -4156
rect -1214 -4160 -1197 -4156
rect -1193 -4160 -1176 -4156
rect -1172 -4160 -1155 -4156
rect -1151 -4160 -1134 -4156
rect -1130 -4160 -1113 -4156
rect -1109 -4160 -1092 -4156
rect -1088 -4160 -1072 -4156
rect -1068 -4160 -1029 -4156
rect -1025 -4160 -926 -4156
rect -922 -4160 -909 -4156
rect -905 -4160 -889 -4156
rect -885 -4160 -868 -4156
rect -864 -4160 -847 -4156
rect -843 -4160 -826 -4156
rect -822 -4160 -805 -4156
rect -801 -4160 -784 -4156
rect -780 -4160 -763 -4156
rect -759 -4160 -743 -4156
rect -739 -4160 -568 -4156
rect -564 -4160 -551 -4156
rect -547 -4160 -531 -4156
rect -527 -4160 -510 -4156
rect -506 -4160 -489 -4156
rect -485 -4160 -468 -4156
rect -464 -4160 -447 -4156
rect -443 -4160 -426 -4156
rect -422 -4160 -405 -4156
rect -401 -4160 -385 -4156
rect -381 -4160 -332 -4156
rect -328 -4160 -210 -4156
rect -206 -4160 -193 -4156
rect -189 -4160 -173 -4156
rect -169 -4160 -152 -4156
rect -148 -4160 -131 -4156
rect -127 -4160 -110 -4156
rect -106 -4160 -89 -4156
rect -85 -4160 -68 -4156
rect -64 -4160 -47 -4156
rect -43 -4160 -27 -4156
rect -23 -4160 456 -4156
rect 460 -4160 1201 -4156
rect 1205 -4160 1617 -4156
rect -1495 -4267 -1433 -4160
rect -1100 -4183 -931 -4179
rect -1233 -4208 -1199 -4204
rect -1135 -4208 -1115 -4204
rect -1017 -4205 -1013 -4201
rect -935 -4212 -931 -4183
rect -413 -4186 -215 -4182
rect -904 -4208 -870 -4204
rect -806 -4208 -786 -4204
rect -771 -4208 -573 -4204
rect -546 -4208 -512 -4204
rect -448 -4208 -428 -4204
rect -577 -4212 -573 -4208
rect -320 -4207 -316 -4203
rect -219 -4212 -215 -4186
rect -188 -4208 -154 -4204
rect -90 -4208 -70 -4204
rect -55 -4208 -21 -4204
rect 468 -4205 472 -4201
rect 1213 -4205 1217 -4201
rect -1421 -4216 -1257 -4212
rect -1253 -4216 -1223 -4212
rect -1202 -4216 -1171 -4212
rect -1142 -4216 -1111 -4212
rect -1100 -4216 -1073 -4212
rect -935 -4216 -928 -4212
rect -924 -4216 -894 -4212
rect -873 -4216 -842 -4212
rect -813 -4216 -782 -4212
rect -771 -4216 -744 -4212
rect -577 -4216 -570 -4212
rect -566 -4216 -536 -4212
rect -515 -4216 -484 -4212
rect -455 -4216 -424 -4212
rect -413 -4216 -386 -4212
rect -219 -4216 -212 -4212
rect -208 -4216 -178 -4212
rect -157 -4216 -126 -4212
rect -97 -4216 -66 -4212
rect -55 -4216 -28 -4212
rect -1260 -4223 -1213 -4219
rect -1177 -4223 -1164 -4219
rect -1160 -4223 -1129 -4219
rect -1093 -4223 -1080 -4219
rect -1076 -4223 -1064 -4219
rect -931 -4223 -884 -4219
rect -848 -4223 -835 -4219
rect -831 -4223 -800 -4219
rect -764 -4223 -751 -4219
rect -747 -4223 -735 -4219
rect -573 -4223 -526 -4219
rect -490 -4223 -477 -4219
rect -473 -4223 -442 -4219
rect -406 -4223 -393 -4219
rect -389 -4223 -377 -4219
rect -215 -4223 -168 -4219
rect -132 -4223 -119 -4219
rect -115 -4223 -84 -4219
rect -48 -4223 -35 -4219
rect -31 -4223 -19 -4219
rect -1268 -4230 -1253 -4226
rect -1249 -4230 -1139 -4226
rect -1118 -4230 -1087 -4226
rect -937 -4230 -924 -4226
rect -920 -4230 -810 -4226
rect -789 -4230 -758 -4226
rect -584 -4230 -583 -4226
rect -579 -4230 -566 -4226
rect -562 -4230 -452 -4226
rect -431 -4230 -400 -4226
rect -227 -4230 -226 -4226
rect -222 -4230 -208 -4226
rect -204 -4230 -94 -4226
rect -73 -4230 -42 -4226
rect -1218 -4237 -1195 -4233
rect -1176 -4237 -1157 -4233
rect -889 -4237 -866 -4233
rect -847 -4237 -828 -4233
rect -531 -4237 -508 -4233
rect -489 -4237 -470 -4233
rect -173 -4237 -150 -4233
rect -131 -4237 -112 -4233
rect 1633 -4248 1695 -4128
rect -1421 -4252 -1255 -4248
rect -1251 -4252 -1238 -4248
rect -1234 -4252 -1197 -4248
rect -1193 -4252 -1155 -4248
rect -1151 -4252 -1113 -4248
rect -1109 -4252 -1072 -4248
rect -1068 -4252 -1029 -4248
rect -1025 -4252 -926 -4248
rect -922 -4252 -909 -4248
rect -905 -4252 -868 -4248
rect -864 -4252 -826 -4248
rect -822 -4252 -784 -4248
rect -780 -4252 -743 -4248
rect -739 -4252 -568 -4248
rect -564 -4252 -551 -4248
rect -547 -4252 -510 -4248
rect -506 -4252 -468 -4248
rect -464 -4252 -426 -4248
rect -422 -4252 -385 -4248
rect -381 -4252 -332 -4248
rect -328 -4252 -210 -4248
rect -206 -4252 -193 -4248
rect -189 -4252 -152 -4248
rect -148 -4252 -110 -4248
rect -106 -4252 -68 -4248
rect -64 -4252 -27 -4248
rect -23 -4252 456 -4248
rect 460 -4252 1201 -4248
rect 1205 -4252 1695 -4248
rect -1495 -4271 -1339 -4267
rect -1335 -4271 -1322 -4267
rect -1318 -4271 -1029 -4267
rect -1025 -4271 -935 -4267
rect -931 -4271 -918 -4267
rect -914 -4271 -673 -4267
rect -669 -4271 -577 -4267
rect -573 -4271 -560 -4267
rect -556 -4271 -332 -4267
rect -328 -4271 -219 -4267
rect -215 -4271 -202 -4267
rect -198 -4271 209 -4267
rect 213 -4271 226 -4267
rect 230 -4271 456 -4267
rect 460 -4271 565 -4267
rect 569 -4271 582 -4267
rect 586 -4271 860 -4267
rect 864 -4271 963 -4267
rect 967 -4271 980 -4267
rect 984 -4271 1201 -4267
rect 1205 -4271 1321 -4267
rect 1325 -4271 1338 -4267
rect 1342 -4271 1617 -4267
rect -1495 -4386 -1433 -4271
rect -1334 -4303 -1066 -4299
rect -930 -4303 -737 -4299
rect -572 -4303 -379 -4299
rect -214 -4303 -15 -4299
rect 214 -4303 407 -4299
rect 570 -4303 763 -4299
rect 968 -4303 1161 -4299
rect 1326 -4303 1519 -4299
rect -1323 -4311 -923 -4307
rect -919 -4311 -565 -4307
rect -561 -4311 -207 -4307
rect -203 -4311 -21 -4307
rect -17 -4311 221 -4307
rect 225 -4311 577 -4307
rect 581 -4311 975 -4307
rect 979 -4311 1333 -4307
rect 1337 -4311 1617 -4307
rect -1017 -4320 -1013 -4316
rect -949 -4324 -909 -4320
rect -661 -4321 -657 -4317
rect -591 -4324 -551 -4320
rect -320 -4322 -316 -4318
rect -233 -4324 -193 -4320
rect 195 -4324 235 -4320
rect 468 -4320 472 -4316
rect 551 -4324 591 -4320
rect 872 -4321 876 -4317
rect 949 -4324 989 -4320
rect 1213 -4320 1217 -4316
rect 1307 -4324 1347 -4320
rect 1633 -4359 1695 -4252
rect -1421 -4363 -1322 -4359
rect -1318 -4363 -1029 -4359
rect -1025 -4363 -918 -4359
rect -914 -4363 -673 -4359
rect -669 -4363 -560 -4359
rect -556 -4363 -332 -4359
rect -328 -4363 -202 -4359
rect -198 -4363 226 -4359
rect 230 -4363 456 -4359
rect 460 -4363 582 -4359
rect 586 -4363 860 -4359
rect 864 -4363 980 -4359
rect 984 -4363 1201 -4359
rect 1205 -4363 1338 -4359
rect 1342 -4363 1695 -4359
rect -1495 -4390 -1255 -4386
rect -1251 -4390 -1238 -4386
rect -1234 -4390 -1198 -4386
rect -1194 -4390 -1177 -4386
rect -1173 -4390 -926 -4386
rect -922 -4390 -900 -4386
rect -896 -4390 -883 -4386
rect -879 -4390 -843 -4386
rect -839 -4390 -822 -4386
rect -818 -4390 -805 -4386
rect -801 -4390 -765 -4386
rect -761 -4390 -741 -4386
rect -737 -4390 -704 -4386
rect -700 -4390 -568 -4386
rect -564 -4390 -542 -4386
rect -538 -4390 -525 -4386
rect -521 -4390 -485 -4386
rect -481 -4390 -464 -4386
rect -460 -4390 -447 -4386
rect -443 -4390 -407 -4386
rect -403 -4390 -383 -4386
rect -379 -4390 -346 -4386
rect -342 -4390 -210 -4386
rect -206 -4390 -184 -4386
rect -180 -4390 -167 -4386
rect -163 -4390 -127 -4386
rect -123 -4390 -106 -4386
rect -102 -4390 -89 -4386
rect -85 -4390 -49 -4386
rect -45 -4390 -25 -4386
rect -21 -4390 12 -4386
rect 16 -4390 218 -4386
rect 222 -4390 244 -4386
rect 248 -4390 261 -4386
rect 265 -4390 301 -4386
rect 305 -4390 322 -4386
rect 326 -4390 339 -4386
rect 343 -4390 379 -4386
rect 383 -4390 403 -4386
rect 407 -4390 440 -4386
rect 444 -4390 574 -4386
rect 578 -4390 600 -4386
rect 604 -4390 617 -4386
rect 621 -4390 657 -4386
rect 661 -4390 678 -4386
rect 682 -4390 695 -4386
rect 699 -4390 735 -4386
rect 739 -4390 759 -4386
rect 763 -4390 796 -4386
rect 800 -4390 972 -4386
rect 976 -4390 998 -4386
rect 1002 -4390 1015 -4386
rect 1019 -4390 1055 -4386
rect 1059 -4390 1076 -4386
rect 1080 -4390 1093 -4386
rect 1097 -4390 1133 -4386
rect 1137 -4390 1157 -4386
rect 1161 -4390 1194 -4386
rect 1198 -4390 1330 -4386
rect 1334 -4390 1356 -4386
rect 1360 -4390 1373 -4386
rect 1377 -4390 1413 -4386
rect 1417 -4390 1434 -4386
rect 1438 -4390 1451 -4386
rect 1455 -4390 1491 -4386
rect 1495 -4390 1515 -4386
rect 1519 -4390 1552 -4386
rect 1556 -4390 1617 -4386
rect -1495 -4509 -1433 -4390
rect -926 -4394 -922 -4390
rect -900 -4394 -896 -4390
rect -883 -4394 -879 -4390
rect -843 -4394 -839 -4390
rect -822 -4394 -818 -4390
rect -805 -4394 -801 -4390
rect -765 -4394 -761 -4390
rect -741 -4394 -737 -4390
rect -704 -4394 -700 -4390
rect -568 -4394 -564 -4390
rect -542 -4394 -538 -4390
rect -525 -4394 -521 -4390
rect -485 -4394 -481 -4390
rect -464 -4394 -460 -4390
rect -447 -4394 -443 -4390
rect -407 -4394 -403 -4390
rect -383 -4394 -379 -4390
rect -346 -4394 -342 -4390
rect -210 -4394 -206 -4390
rect -184 -4394 -180 -4390
rect -167 -4394 -163 -4390
rect -127 -4394 -123 -4390
rect -106 -4394 -102 -4390
rect -89 -4394 -85 -4390
rect -49 -4394 -45 -4390
rect -25 -4394 -21 -4390
rect 12 -4394 16 -4390
rect 218 -4394 222 -4390
rect 244 -4394 248 -4390
rect 261 -4394 265 -4390
rect 301 -4394 305 -4390
rect 322 -4394 326 -4390
rect 339 -4394 343 -4390
rect 379 -4394 383 -4390
rect 403 -4394 407 -4390
rect 440 -4394 444 -4390
rect 574 -4394 578 -4390
rect 600 -4394 604 -4390
rect 617 -4394 621 -4390
rect 657 -4394 661 -4390
rect 678 -4394 682 -4390
rect 695 -4394 699 -4390
rect 735 -4394 739 -4390
rect 759 -4394 763 -4390
rect 796 -4394 800 -4390
rect 972 -4394 976 -4390
rect 998 -4394 1002 -4390
rect 1015 -4394 1019 -4390
rect 1055 -4394 1059 -4390
rect 1076 -4394 1080 -4390
rect 1093 -4394 1097 -4390
rect 1133 -4394 1137 -4390
rect 1157 -4394 1161 -4390
rect 1194 -4394 1198 -4390
rect 1330 -4394 1334 -4390
rect 1356 -4394 1360 -4390
rect 1373 -4394 1377 -4390
rect 1413 -4394 1417 -4390
rect 1434 -4394 1438 -4390
rect 1451 -4394 1455 -4390
rect 1491 -4394 1495 -4390
rect 1515 -4394 1519 -4390
rect 1552 -4394 1556 -4390
rect -920 -4409 -858 -4405
rect -854 -4409 -824 -4405
rect -776 -4409 -746 -4405
rect -562 -4409 -500 -4405
rect -496 -4409 -466 -4405
rect -418 -4409 -388 -4405
rect -204 -4409 -142 -4405
rect -138 -4409 -108 -4405
rect -60 -4409 -30 -4405
rect 224 -4409 286 -4405
rect 290 -4409 320 -4405
rect 368 -4409 398 -4405
rect 580 -4409 642 -4405
rect 646 -4409 676 -4405
rect 724 -4409 754 -4405
rect 978 -4409 1040 -4405
rect 1044 -4409 1074 -4405
rect 1122 -4409 1152 -4405
rect 1336 -4409 1398 -4405
rect 1402 -4409 1432 -4405
rect 1480 -4409 1510 -4405
rect -913 -4416 -882 -4412
rect -555 -4416 -524 -4412
rect -197 -4416 -166 -4412
rect 231 -4416 262 -4412
rect 587 -4416 618 -4412
rect 985 -4416 1016 -4412
rect 1343 -4416 1374 -4412
rect -931 -4423 -848 -4419
rect -809 -4423 -706 -4419
rect -573 -4423 -490 -4419
rect -451 -4423 -348 -4419
rect -215 -4423 -132 -4419
rect -93 -4423 10 -4419
rect 213 -4423 296 -4419
rect 335 -4423 438 -4419
rect 569 -4423 652 -4419
rect 691 -4423 794 -4419
rect 967 -4423 1050 -4419
rect 1089 -4423 1192 -4419
rect 1325 -4423 1408 -4419
rect 1447 -4423 1550 -4419
rect -949 -4430 -928 -4426
rect -894 -4430 -865 -4426
rect -861 -4430 -780 -4426
rect -691 -4430 -592 -4426
rect -585 -4430 -570 -4426
rect -536 -4430 -507 -4426
rect -503 -4430 -422 -4426
rect -333 -4429 -234 -4425
rect -596 -4434 -592 -4430
rect -238 -4434 -234 -4429
rect -227 -4430 -212 -4426
rect -178 -4430 -149 -4426
rect -145 -4430 -64 -4426
rect 25 -4430 194 -4426
rect 201 -4430 216 -4426
rect 250 -4430 279 -4426
rect 283 -4430 364 -4426
rect 453 -4430 550 -4426
rect 557 -4430 572 -4426
rect 606 -4430 635 -4426
rect 639 -4430 720 -4426
rect 809 -4430 948 -4426
rect 955 -4430 970 -4426
rect 1004 -4430 1033 -4426
rect 1037 -4430 1118 -4426
rect 1207 -4428 1300 -4424
rect 190 -4434 194 -4430
rect 546 -4434 550 -4430
rect 944 -4434 948 -4430
rect 1296 -4434 1300 -4428
rect 1307 -4430 1328 -4426
rect 1362 -4430 1391 -4426
rect 1395 -4430 1476 -4426
rect -1260 -4439 -1203 -4435
rect -1164 -4438 -902 -4434
rect -887 -4438 -804 -4434
rect -783 -4438 -689 -4434
rect -596 -4438 -544 -4434
rect -529 -4438 -446 -4434
rect -425 -4438 -331 -4434
rect -238 -4438 -186 -4434
rect -171 -4438 -88 -4434
rect -67 -4438 27 -4434
rect 190 -4438 242 -4434
rect 257 -4438 340 -4434
rect 361 -4438 455 -4434
rect 546 -4438 598 -4434
rect 613 -4438 696 -4434
rect 717 -4438 811 -4434
rect 944 -4438 996 -4434
rect 1011 -4438 1094 -4434
rect 1115 -4438 1209 -4434
rect 1296 -4438 1354 -4434
rect 1369 -4438 1452 -4434
rect 1473 -4438 1567 -4434
rect -1266 -4446 -1253 -4442
rect -1249 -4446 -1213 -4442
rect -1209 -4446 -1193 -4442
rect -943 -4445 -924 -4441
rect -905 -4445 -776 -4441
rect -591 -4445 -566 -4441
rect -547 -4445 -418 -4441
rect -233 -4445 -208 -4441
rect -189 -4445 -60 -4441
rect 195 -4445 220 -4441
rect 239 -4445 368 -4441
rect 551 -4445 576 -4441
rect 595 -4445 724 -4441
rect 949 -4445 974 -4441
rect 993 -4445 1122 -4441
rect 1313 -4445 1332 -4441
rect 1351 -4445 1480 -4441
rect -1309 -4453 -1257 -4449
rect -1253 -4453 -1227 -4449
rect -1223 -4453 -1179 -4449
rect -898 -4452 -794 -4448
rect -790 -4452 -760 -4448
rect -540 -4452 -436 -4448
rect -432 -4452 -402 -4448
rect -182 -4452 -78 -4448
rect -74 -4452 -44 -4448
rect 246 -4452 350 -4448
rect 354 -4452 384 -4448
rect 602 -4452 706 -4448
rect 710 -4452 740 -4448
rect 1000 -4452 1104 -4448
rect 1108 -4452 1138 -4448
rect 1358 -4452 1462 -4448
rect 1466 -4452 1496 -4448
rect -1216 -4460 -1162 -4456
rect -924 -4459 -872 -4455
rect -868 -4459 -838 -4455
rect -566 -4459 -514 -4455
rect -510 -4459 -480 -4455
rect -208 -4459 -156 -4455
rect -152 -4459 -122 -4455
rect 220 -4459 272 -4455
rect 276 -4459 306 -4455
rect 576 -4459 628 -4455
rect 632 -4459 662 -4455
rect 974 -4459 1026 -4455
rect 1030 -4459 1060 -4455
rect 1332 -4459 1384 -4455
rect 1388 -4459 1418 -4455
rect -1234 -4467 -1202 -4463
rect -879 -4467 -847 -4463
rect -883 -4470 -879 -4467
rect -847 -4470 -843 -4467
rect -801 -4467 -769 -4463
rect -805 -4470 -801 -4467
rect -769 -4470 -765 -4467
rect -521 -4467 -489 -4463
rect -525 -4470 -521 -4467
rect -489 -4470 -485 -4467
rect -443 -4467 -411 -4463
rect -447 -4470 -443 -4467
rect -411 -4470 -407 -4467
rect -163 -4467 -131 -4463
rect -167 -4470 -163 -4467
rect -131 -4470 -127 -4467
rect -85 -4467 -53 -4463
rect -89 -4470 -85 -4467
rect -53 -4470 -49 -4467
rect 265 -4467 297 -4463
rect 261 -4470 265 -4467
rect 297 -4470 301 -4467
rect 343 -4467 375 -4463
rect 339 -4470 343 -4467
rect 375 -4470 379 -4467
rect 621 -4467 653 -4463
rect 617 -4470 621 -4467
rect 653 -4470 657 -4467
rect 699 -4467 731 -4463
rect 695 -4470 699 -4467
rect 731 -4470 735 -4467
rect 1019 -4467 1051 -4463
rect 1015 -4470 1019 -4467
rect 1051 -4470 1055 -4467
rect 1097 -4467 1129 -4463
rect 1093 -4470 1097 -4467
rect 1129 -4470 1133 -4467
rect 1377 -4467 1409 -4463
rect 1373 -4470 1377 -4467
rect 1409 -4470 1413 -4467
rect 1455 -4467 1487 -4463
rect 1451 -4470 1455 -4467
rect 1487 -4470 1491 -4467
rect -926 -4478 -922 -4474
rect -900 -4478 -896 -4474
rect -857 -4478 -853 -4474
rect -822 -4478 -818 -4474
rect -778 -4478 -774 -4474
rect -761 -4478 -757 -4474
rect -725 -4478 -721 -4474
rect -704 -4478 -700 -4474
rect -568 -4478 -564 -4474
rect -542 -4478 -538 -4474
rect -499 -4478 -495 -4474
rect -464 -4478 -460 -4474
rect -420 -4478 -416 -4474
rect -403 -4478 -399 -4474
rect -367 -4478 -363 -4474
rect -346 -4478 -342 -4474
rect -210 -4478 -206 -4474
rect -184 -4478 -180 -4474
rect -141 -4478 -137 -4474
rect -106 -4478 -102 -4474
rect -62 -4478 -58 -4474
rect -45 -4478 -41 -4474
rect -9 -4478 -5 -4474
rect 12 -4478 16 -4474
rect 218 -4478 222 -4474
rect 244 -4478 248 -4474
rect 287 -4478 291 -4474
rect 322 -4478 326 -4474
rect 366 -4478 370 -4474
rect 383 -4478 387 -4474
rect 419 -4478 423 -4474
rect 440 -4478 444 -4474
rect 574 -4478 578 -4474
rect 600 -4478 604 -4474
rect 643 -4478 647 -4474
rect 678 -4478 682 -4474
rect 722 -4478 726 -4474
rect 739 -4478 743 -4474
rect 775 -4478 779 -4474
rect 796 -4478 800 -4474
rect 972 -4478 976 -4474
rect 998 -4478 1002 -4474
rect 1041 -4478 1045 -4474
rect 1076 -4478 1080 -4474
rect 1120 -4478 1124 -4474
rect 1137 -4478 1141 -4474
rect 1173 -4478 1177 -4474
rect 1194 -4478 1198 -4474
rect 1330 -4478 1334 -4474
rect 1356 -4478 1360 -4474
rect 1399 -4478 1403 -4474
rect 1434 -4478 1438 -4474
rect 1478 -4478 1482 -4474
rect 1495 -4478 1499 -4474
rect 1531 -4478 1535 -4474
rect 1552 -4478 1556 -4474
rect 1633 -4478 1695 -4363
rect -1421 -4482 -1255 -4478
rect -1251 -4482 -1211 -4478
rect -1207 -4482 -1177 -4478
rect -1173 -4482 -926 -4478
rect -922 -4482 -900 -4478
rect -896 -4482 -857 -4478
rect -853 -4482 -822 -4478
rect -818 -4482 -778 -4478
rect -774 -4482 -761 -4478
rect -757 -4482 -725 -4478
rect -721 -4482 -704 -4478
rect -700 -4482 -568 -4478
rect -564 -4482 -542 -4478
rect -538 -4482 -499 -4478
rect -495 -4482 -464 -4478
rect -460 -4482 -420 -4478
rect -416 -4482 -403 -4478
rect -399 -4482 -367 -4478
rect -363 -4482 -346 -4478
rect -342 -4482 -210 -4478
rect -206 -4482 -184 -4478
rect -180 -4482 -141 -4478
rect -137 -4482 -106 -4478
rect -102 -4482 -62 -4478
rect -58 -4482 -45 -4478
rect -41 -4482 -9 -4478
rect -5 -4482 12 -4478
rect 16 -4482 218 -4478
rect 222 -4482 244 -4478
rect 248 -4482 287 -4478
rect 291 -4482 322 -4478
rect 326 -4482 366 -4478
rect 370 -4482 383 -4478
rect 387 -4482 419 -4478
rect 423 -4482 440 -4478
rect 444 -4482 574 -4478
rect 578 -4482 600 -4478
rect 604 -4482 643 -4478
rect 647 -4482 678 -4478
rect 682 -4482 722 -4478
rect 726 -4482 739 -4478
rect 743 -4482 775 -4478
rect 779 -4482 796 -4478
rect 800 -4482 972 -4478
rect 976 -4482 998 -4478
rect 1002 -4482 1041 -4478
rect 1045 -4482 1076 -4478
rect 1080 -4482 1120 -4478
rect 1124 -4482 1137 -4478
rect 1141 -4482 1173 -4478
rect 1177 -4482 1194 -4478
rect 1198 -4482 1330 -4478
rect 1334 -4482 1356 -4478
rect 1360 -4482 1399 -4478
rect 1403 -4482 1434 -4478
rect 1438 -4482 1478 -4478
rect 1482 -4482 1495 -4478
rect 1499 -4482 1531 -4478
rect 1535 -4482 1552 -4478
rect 1556 -4482 1695 -4478
rect -1272 -4489 -689 -4485
rect -585 -4489 27 -4485
rect 201 -4489 811 -4485
rect 955 -4489 1567 -4485
rect -1266 -4496 -1162 -4492
rect -943 -4496 -331 -4492
rect -227 -4496 455 -4492
rect 557 -4496 1209 -4492
rect 1313 -4496 1561 -4492
rect -1495 -4513 -1255 -4509
rect -1251 -4513 -1238 -4509
rect -1234 -4513 -1218 -4509
rect -1214 -4513 -1197 -4509
rect -1193 -4513 -1176 -4509
rect -1172 -4513 -1155 -4509
rect -1151 -4513 -1134 -4509
rect -1130 -4513 -1113 -4509
rect -1109 -4513 -1092 -4509
rect -1088 -4513 -1072 -4509
rect -1068 -4513 -926 -4509
rect -922 -4513 -909 -4509
rect -905 -4513 -889 -4509
rect -885 -4513 -868 -4509
rect -864 -4513 -847 -4509
rect -843 -4513 -826 -4509
rect -822 -4513 -805 -4509
rect -801 -4513 -784 -4509
rect -780 -4513 -763 -4509
rect -759 -4513 -743 -4509
rect -739 -4513 -568 -4509
rect -564 -4513 -551 -4509
rect -547 -4513 -531 -4509
rect -527 -4513 -510 -4509
rect -506 -4513 -489 -4509
rect -485 -4513 -468 -4509
rect -464 -4513 -447 -4509
rect -443 -4513 -426 -4509
rect -422 -4513 -405 -4509
rect -401 -4513 -385 -4509
rect -381 -4513 1617 -4509
rect -1495 -4630 -1433 -4513
rect -1233 -4561 -1199 -4557
rect -1135 -4561 -1115 -4557
rect -1100 -4561 -931 -4557
rect -904 -4561 -870 -4557
rect -806 -4561 -786 -4557
rect -771 -4561 -573 -4557
rect -546 -4561 -512 -4557
rect -448 -4561 -428 -4557
rect -413 -4561 -377 -4557
rect -935 -4565 -931 -4561
rect -577 -4565 -573 -4561
rect -1266 -4569 -1257 -4565
rect -1253 -4569 -1223 -4565
rect -1202 -4569 -1171 -4565
rect -1142 -4569 -1111 -4565
rect -1100 -4569 -1073 -4565
rect -935 -4569 -928 -4565
rect -924 -4569 -894 -4565
rect -873 -4569 -842 -4565
rect -813 -4569 -782 -4565
rect -771 -4569 -744 -4565
rect -577 -4569 -570 -4565
rect -566 -4569 -536 -4565
rect -515 -4569 -484 -4565
rect -455 -4569 -424 -4565
rect -413 -4569 -386 -4565
rect -1260 -4576 -1213 -4572
rect -1177 -4576 -1164 -4572
rect -1160 -4576 -1129 -4572
rect -1093 -4576 -1080 -4572
rect -1076 -4576 -1064 -4572
rect -931 -4576 -884 -4572
rect -848 -4576 -835 -4572
rect -831 -4576 -800 -4572
rect -764 -4576 -751 -4572
rect -747 -4576 -735 -4572
rect -573 -4576 -526 -4572
rect -490 -4576 -477 -4572
rect -473 -4576 -442 -4572
rect -406 -4576 -393 -4572
rect -389 -4576 -377 -4572
rect -1267 -4583 -1253 -4579
rect -1249 -4583 -1139 -4579
rect -1118 -4583 -1087 -4579
rect -938 -4583 -924 -4579
rect -920 -4583 -810 -4579
rect -789 -4583 -758 -4579
rect -583 -4583 -566 -4579
rect -562 -4583 -452 -4579
rect -431 -4583 -400 -4579
rect -1218 -4590 -1195 -4586
rect -1176 -4590 -1157 -4586
rect -889 -4590 -866 -4586
rect -847 -4590 -828 -4586
rect -531 -4590 -508 -4586
rect -489 -4590 -470 -4586
rect 1633 -4601 1695 -4482
rect -1421 -4605 -1255 -4601
rect -1251 -4605 -1238 -4601
rect -1234 -4605 -1197 -4601
rect -1193 -4605 -1155 -4601
rect -1151 -4605 -1113 -4601
rect -1109 -4605 -1072 -4601
rect -1068 -4605 -926 -4601
rect -922 -4605 -909 -4601
rect -905 -4605 -868 -4601
rect -864 -4605 -826 -4601
rect -822 -4605 -784 -4601
rect -780 -4605 -743 -4601
rect -739 -4605 -568 -4601
rect -564 -4605 -551 -4601
rect -547 -4605 -510 -4601
rect -506 -4605 -468 -4601
rect -464 -4605 -426 -4601
rect -422 -4605 -385 -4601
rect -381 -4605 1695 -4601
rect -1495 -4634 -1255 -4630
rect -1251 -4634 -1238 -4630
rect -1234 -4634 -1218 -4630
rect -1214 -4634 -1197 -4630
rect -1193 -4634 -1176 -4630
rect -1172 -4634 -1155 -4630
rect -1151 -4634 -1134 -4630
rect -1130 -4634 -1113 -4630
rect -1109 -4634 -1092 -4630
rect -1088 -4634 -1072 -4630
rect -1068 -4634 -926 -4630
rect -922 -4634 -909 -4630
rect -905 -4634 -889 -4630
rect -885 -4634 -868 -4630
rect -864 -4634 -847 -4630
rect -843 -4634 -826 -4630
rect -822 -4634 -805 -4630
rect -801 -4634 -784 -4630
rect -780 -4634 -763 -4630
rect -759 -4634 -743 -4630
rect -739 -4634 -568 -4630
rect -564 -4634 -551 -4630
rect -547 -4634 -531 -4630
rect -527 -4634 -510 -4630
rect -506 -4634 -489 -4630
rect -485 -4634 -468 -4630
rect -464 -4634 -447 -4630
rect -443 -4634 -426 -4630
rect -422 -4634 -405 -4630
rect -401 -4634 -385 -4630
rect -381 -4634 -210 -4630
rect -206 -4634 -193 -4630
rect -189 -4634 -173 -4630
rect -169 -4634 -152 -4630
rect -148 -4634 -131 -4630
rect -127 -4634 -110 -4630
rect -106 -4634 -89 -4630
rect -85 -4634 -68 -4630
rect -64 -4634 -47 -4630
rect -43 -4634 -27 -4630
rect -23 -4634 218 -4630
rect 222 -4634 235 -4630
rect 239 -4634 255 -4630
rect 259 -4634 276 -4630
rect 280 -4634 297 -4630
rect 301 -4634 318 -4630
rect 322 -4634 339 -4630
rect 343 -4634 360 -4630
rect 364 -4634 381 -4630
rect 385 -4634 401 -4630
rect 405 -4634 574 -4630
rect 578 -4634 591 -4630
rect 595 -4634 611 -4630
rect 615 -4634 632 -4630
rect 636 -4634 653 -4630
rect 657 -4634 674 -4630
rect 678 -4634 695 -4630
rect 699 -4634 716 -4630
rect 720 -4634 737 -4630
rect 741 -4634 757 -4630
rect 761 -4634 972 -4630
rect 976 -4634 989 -4630
rect 993 -4634 1009 -4630
rect 1013 -4634 1030 -4630
rect 1034 -4634 1051 -4630
rect 1055 -4634 1072 -4630
rect 1076 -4634 1093 -4630
rect 1097 -4634 1114 -4630
rect 1118 -4634 1135 -4630
rect 1139 -4634 1155 -4630
rect 1159 -4634 1330 -4630
rect 1334 -4634 1347 -4630
rect 1351 -4634 1367 -4630
rect 1371 -4634 1388 -4630
rect 1392 -4634 1409 -4630
rect 1413 -4634 1430 -4630
rect 1434 -4634 1451 -4630
rect 1455 -4634 1472 -4630
rect 1476 -4634 1493 -4630
rect 1497 -4634 1513 -4630
rect 1517 -4634 1617 -4630
rect -1495 -4751 -1433 -4634
rect -1233 -4682 -1199 -4678
rect -1135 -4682 -1115 -4678
rect -1100 -4682 -1066 -4678
rect -904 -4682 -870 -4678
rect -806 -4682 -786 -4678
rect -771 -4682 -737 -4678
rect -546 -4682 -512 -4678
rect -448 -4682 -428 -4678
rect -413 -4682 -379 -4678
rect -188 -4682 -154 -4678
rect -90 -4682 -70 -4678
rect -55 -4682 -21 -4678
rect 240 -4682 274 -4678
rect 338 -4682 358 -4678
rect 373 -4682 407 -4678
rect 596 -4682 630 -4678
rect 694 -4682 714 -4678
rect 729 -4682 763 -4678
rect 994 -4682 1028 -4678
rect 1092 -4682 1112 -4678
rect 1127 -4682 1161 -4678
rect 1352 -4682 1386 -4678
rect 1450 -4682 1470 -4678
rect 1485 -4682 1519 -4678
rect -1272 -4690 -1257 -4686
rect -1253 -4690 -1223 -4686
rect -1202 -4690 -1171 -4686
rect -1142 -4690 -1111 -4686
rect -1100 -4690 -1073 -4686
rect -943 -4690 -928 -4686
rect -924 -4690 -894 -4686
rect -873 -4690 -842 -4686
rect -813 -4690 -782 -4686
rect -771 -4690 -744 -4686
rect -585 -4690 -570 -4686
rect -566 -4690 -536 -4686
rect -515 -4690 -484 -4686
rect -455 -4690 -424 -4686
rect -413 -4690 -386 -4686
rect -227 -4690 -212 -4686
rect -208 -4690 -178 -4686
rect -157 -4690 -126 -4686
rect -97 -4690 -66 -4686
rect -55 -4690 -28 -4686
rect 201 -4690 216 -4686
rect 220 -4690 250 -4686
rect 271 -4690 302 -4686
rect 331 -4690 362 -4686
rect 373 -4690 400 -4686
rect 557 -4690 572 -4686
rect 576 -4690 606 -4686
rect 627 -4690 658 -4686
rect 687 -4690 718 -4686
rect 729 -4690 756 -4686
rect 955 -4690 970 -4686
rect 974 -4690 1004 -4686
rect 1025 -4690 1056 -4686
rect 1085 -4690 1116 -4686
rect 1127 -4690 1154 -4686
rect 1313 -4690 1328 -4686
rect 1332 -4690 1362 -4686
rect 1383 -4690 1414 -4686
rect 1443 -4690 1474 -4686
rect 1485 -4690 1512 -4686
rect -1260 -4697 -1213 -4693
rect -1177 -4697 -1164 -4693
rect -1160 -4697 -1129 -4693
rect -1093 -4697 -1080 -4693
rect -1076 -4697 -1064 -4693
rect -931 -4697 -884 -4693
rect -848 -4697 -835 -4693
rect -831 -4697 -800 -4693
rect -764 -4697 -751 -4693
rect -747 -4697 -735 -4693
rect -573 -4697 -526 -4693
rect -490 -4697 -477 -4693
rect -473 -4697 -442 -4693
rect -406 -4697 -393 -4693
rect -389 -4697 -377 -4693
rect -215 -4697 -168 -4693
rect -132 -4697 -119 -4693
rect -115 -4697 -84 -4693
rect -48 -4697 -35 -4693
rect -31 -4697 -19 -4693
rect 213 -4697 260 -4693
rect 296 -4697 309 -4693
rect 313 -4697 344 -4693
rect 380 -4697 393 -4693
rect 397 -4697 409 -4693
rect 569 -4697 616 -4693
rect 652 -4697 665 -4693
rect 669 -4697 700 -4693
rect 736 -4697 749 -4693
rect 753 -4697 765 -4693
rect 967 -4697 1014 -4693
rect 1050 -4697 1063 -4693
rect 1067 -4697 1098 -4693
rect 1134 -4697 1147 -4693
rect 1151 -4697 1163 -4693
rect 1325 -4697 1372 -4693
rect 1408 -4697 1421 -4693
rect 1425 -4697 1456 -4693
rect 1492 -4697 1505 -4693
rect 1509 -4697 1521 -4693
rect -1268 -4704 -1253 -4700
rect -1249 -4704 -1139 -4700
rect -1118 -4704 -1087 -4700
rect -937 -4704 -924 -4700
rect -920 -4704 -810 -4700
rect -789 -4704 -758 -4700
rect -583 -4704 -566 -4700
rect -562 -4704 -452 -4700
rect -431 -4704 -400 -4700
rect -222 -4704 -208 -4700
rect -204 -4704 -94 -4700
rect -73 -4704 -42 -4700
rect 206 -4704 220 -4700
rect 224 -4704 334 -4700
rect 355 -4704 386 -4700
rect 562 -4704 576 -4700
rect 580 -4704 690 -4700
rect 711 -4704 742 -4700
rect 959 -4704 974 -4700
rect 978 -4704 1088 -4700
rect 1109 -4704 1140 -4700
rect 1319 -4704 1332 -4700
rect 1336 -4704 1446 -4700
rect 1467 -4704 1498 -4700
rect -1218 -4711 -1195 -4707
rect -1176 -4711 -1157 -4707
rect -889 -4711 -866 -4707
rect -847 -4711 -828 -4707
rect -531 -4711 -508 -4707
rect -489 -4711 -470 -4707
rect -173 -4711 -150 -4707
rect -131 -4711 -112 -4707
rect 255 -4711 278 -4707
rect 297 -4711 316 -4707
rect 611 -4711 634 -4707
rect 653 -4711 672 -4707
rect 1009 -4711 1032 -4707
rect 1051 -4711 1070 -4707
rect 1367 -4711 1390 -4707
rect 1409 -4711 1428 -4707
rect 1633 -4722 1695 -4605
rect -1421 -4726 -1255 -4722
rect -1251 -4726 -1238 -4722
rect -1234 -4726 -1197 -4722
rect -1193 -4726 -1155 -4722
rect -1151 -4726 -1113 -4722
rect -1109 -4726 -1072 -4722
rect -1068 -4726 -926 -4722
rect -922 -4726 -909 -4722
rect -905 -4726 -868 -4722
rect -864 -4726 -826 -4722
rect -822 -4726 -784 -4722
rect -780 -4726 -743 -4722
rect -739 -4726 -568 -4722
rect -564 -4726 -551 -4722
rect -547 -4726 -510 -4722
rect -506 -4726 -468 -4722
rect -464 -4726 -426 -4722
rect -422 -4726 -385 -4722
rect -381 -4726 -210 -4722
rect -206 -4726 -193 -4722
rect -189 -4726 -152 -4722
rect -148 -4726 -110 -4722
rect -106 -4726 -68 -4722
rect -64 -4726 -27 -4722
rect -23 -4726 218 -4722
rect 222 -4726 235 -4722
rect 239 -4726 276 -4722
rect 280 -4726 318 -4722
rect 322 -4726 360 -4722
rect 364 -4726 401 -4722
rect 405 -4726 574 -4722
rect 578 -4726 591 -4722
rect 595 -4726 632 -4722
rect 636 -4726 674 -4722
rect 678 -4726 716 -4722
rect 720 -4726 757 -4722
rect 761 -4726 972 -4722
rect 976 -4726 989 -4722
rect 993 -4726 1030 -4722
rect 1034 -4726 1072 -4722
rect 1076 -4726 1114 -4722
rect 1118 -4726 1155 -4722
rect 1159 -4726 1330 -4722
rect 1334 -4726 1347 -4722
rect 1351 -4726 1388 -4722
rect 1392 -4726 1430 -4722
rect 1434 -4726 1472 -4722
rect 1476 -4726 1513 -4722
rect 1517 -4726 1695 -4722
rect -1266 -4734 -1066 -4730
rect -943 -4733 -737 -4729
rect -585 -4733 -379 -4729
rect -227 -4733 -21 -4729
rect 201 -4735 407 -4731
rect 557 -4734 763 -4730
rect 955 -4733 1161 -4729
rect 1313 -4733 1519 -4729
rect -1495 -4755 -1255 -4751
rect -1251 -4755 -1238 -4751
rect -1234 -4755 -1218 -4751
rect -1214 -4755 -1197 -4751
rect -1193 -4755 -1176 -4751
rect -1172 -4755 -1155 -4751
rect -1151 -4755 -1134 -4751
rect -1130 -4755 -1113 -4751
rect -1109 -4755 -1092 -4751
rect -1088 -4755 -1072 -4751
rect -1068 -4755 -926 -4751
rect -922 -4755 -909 -4751
rect -905 -4755 -889 -4751
rect -885 -4755 -868 -4751
rect -864 -4755 -847 -4751
rect -843 -4755 -826 -4751
rect -822 -4755 -805 -4751
rect -801 -4755 -784 -4751
rect -780 -4755 -763 -4751
rect -759 -4755 -743 -4751
rect -739 -4755 -568 -4751
rect -564 -4755 -551 -4751
rect -547 -4755 -531 -4751
rect -527 -4755 -510 -4751
rect -506 -4755 -489 -4751
rect -485 -4755 -468 -4751
rect -464 -4755 -447 -4751
rect -443 -4755 -426 -4751
rect -422 -4755 -405 -4751
rect -401 -4755 -385 -4751
rect -381 -4755 -210 -4751
rect -206 -4755 -193 -4751
rect -189 -4755 -173 -4751
rect -169 -4755 -152 -4751
rect -148 -4755 -131 -4751
rect -127 -4755 -110 -4751
rect -106 -4755 -89 -4751
rect -85 -4755 -68 -4751
rect -64 -4755 -47 -4751
rect -43 -4755 -27 -4751
rect -23 -4755 90 -4751
rect 94 -4755 218 -4751
rect 222 -4755 235 -4751
rect 239 -4755 255 -4751
rect 259 -4755 276 -4751
rect 280 -4755 297 -4751
rect 301 -4755 318 -4751
rect 322 -4755 339 -4751
rect 343 -4755 360 -4751
rect 364 -4755 381 -4751
rect 385 -4755 401 -4751
rect 405 -4755 574 -4751
rect 578 -4755 591 -4751
rect 595 -4755 611 -4751
rect 615 -4755 632 -4751
rect 636 -4755 653 -4751
rect 657 -4755 674 -4751
rect 678 -4755 695 -4751
rect 699 -4755 716 -4751
rect 720 -4755 737 -4751
rect 741 -4755 757 -4751
rect 761 -4755 972 -4751
rect 976 -4755 989 -4751
rect 993 -4755 1009 -4751
rect 1013 -4755 1030 -4751
rect 1034 -4755 1051 -4751
rect 1055 -4755 1072 -4751
rect 1076 -4755 1093 -4751
rect 1097 -4755 1114 -4751
rect 1118 -4755 1135 -4751
rect 1139 -4755 1155 -4751
rect 1159 -4755 1330 -4751
rect 1334 -4755 1347 -4751
rect 1351 -4755 1367 -4751
rect 1371 -4755 1388 -4751
rect 1392 -4755 1409 -4751
rect 1413 -4755 1430 -4751
rect 1434 -4755 1451 -4751
rect 1455 -4755 1472 -4751
rect 1476 -4755 1493 -4751
rect 1497 -4755 1513 -4751
rect 1517 -4755 1617 -4751
rect -1495 -4869 -1433 -4755
rect -1233 -4803 -1199 -4799
rect -1135 -4803 -1115 -4799
rect -1100 -4803 -1066 -4799
rect -904 -4803 -870 -4799
rect -806 -4803 -786 -4799
rect -771 -4803 -737 -4799
rect -546 -4803 -512 -4799
rect -448 -4803 -428 -4799
rect -413 -4803 -379 -4799
rect -188 -4803 -154 -4799
rect -90 -4803 -70 -4799
rect -55 -4803 -21 -4799
rect -1345 -4811 -1257 -4807
rect -1253 -4811 -1223 -4807
rect -1202 -4811 -1171 -4807
rect -1142 -4811 -1111 -4807
rect -1100 -4811 -1073 -4807
rect -937 -4811 -928 -4807
rect -924 -4811 -894 -4807
rect -873 -4811 -842 -4807
rect -813 -4811 -782 -4807
rect -771 -4811 -744 -4807
rect -579 -4811 -570 -4807
rect -566 -4811 -536 -4807
rect -515 -4811 -484 -4807
rect -455 -4811 -424 -4807
rect -413 -4811 -386 -4807
rect -221 -4811 -212 -4807
rect -208 -4811 -178 -4807
rect -157 -4811 -126 -4807
rect -97 -4811 -66 -4807
rect -55 -4811 -28 -4807
rect 102 -4806 106 -4802
rect 240 -4803 274 -4799
rect 338 -4803 358 -4799
rect 373 -4803 413 -4799
rect 596 -4803 630 -4799
rect 694 -4803 714 -4799
rect 729 -4803 763 -4799
rect 994 -4803 1028 -4799
rect 1092 -4803 1112 -4799
rect 1127 -4803 1161 -4799
rect 1352 -4803 1386 -4799
rect 1450 -4803 1470 -4799
rect 1485 -4803 1519 -4799
rect 207 -4811 216 -4807
rect 220 -4811 250 -4807
rect 271 -4811 302 -4807
rect 331 -4811 362 -4807
rect 373 -4811 400 -4807
rect 563 -4811 572 -4807
rect 576 -4811 606 -4807
rect 627 -4811 658 -4807
rect 687 -4811 718 -4807
rect 729 -4811 756 -4807
rect 961 -4811 970 -4807
rect 974 -4811 1004 -4807
rect 1025 -4811 1056 -4807
rect 1085 -4811 1116 -4807
rect 1127 -4811 1154 -4807
rect 1319 -4811 1328 -4807
rect 1332 -4811 1362 -4807
rect 1383 -4811 1414 -4807
rect 1443 -4811 1474 -4807
rect 1485 -4811 1512 -4807
rect -1260 -4818 -1213 -4814
rect -1177 -4818 -1164 -4814
rect -1160 -4818 -1129 -4814
rect -1093 -4818 -1080 -4814
rect -1076 -4818 -1064 -4814
rect -931 -4818 -884 -4814
rect -848 -4818 -835 -4814
rect -831 -4818 -800 -4814
rect -764 -4818 -751 -4814
rect -747 -4818 -735 -4814
rect -573 -4818 -526 -4814
rect -490 -4818 -477 -4814
rect -473 -4818 -442 -4814
rect -406 -4818 -393 -4814
rect -389 -4818 -377 -4814
rect -215 -4818 -168 -4814
rect -132 -4818 -119 -4814
rect -115 -4818 -84 -4814
rect -48 -4818 -35 -4814
rect -31 -4818 -19 -4814
rect 213 -4818 260 -4814
rect 296 -4818 309 -4814
rect 313 -4818 344 -4814
rect 380 -4818 393 -4814
rect 397 -4818 409 -4814
rect 569 -4818 616 -4814
rect 652 -4818 665 -4814
rect 669 -4818 700 -4814
rect 736 -4818 749 -4814
rect 753 -4818 765 -4814
rect 967 -4818 1014 -4814
rect 1050 -4818 1063 -4814
rect 1067 -4818 1098 -4814
rect 1134 -4818 1147 -4814
rect 1151 -4818 1163 -4814
rect 1325 -4818 1372 -4814
rect 1408 -4818 1421 -4814
rect 1425 -4818 1456 -4814
rect 1492 -4818 1505 -4814
rect 1509 -4818 1521 -4814
rect -1268 -4825 -1253 -4821
rect -1249 -4825 -1139 -4821
rect -1118 -4825 -1087 -4821
rect -937 -4825 -924 -4821
rect -920 -4825 -810 -4821
rect -789 -4825 -758 -4821
rect -583 -4825 -566 -4821
rect -562 -4825 -452 -4821
rect -431 -4825 -400 -4821
rect -222 -4825 -208 -4821
rect -204 -4825 -94 -4821
rect -73 -4825 -42 -4821
rect 206 -4825 220 -4821
rect 224 -4825 334 -4821
rect 355 -4825 386 -4821
rect 562 -4825 576 -4821
rect 580 -4825 690 -4821
rect 711 -4825 742 -4821
rect 959 -4825 974 -4821
rect 978 -4825 1088 -4821
rect 1109 -4825 1140 -4821
rect 1319 -4825 1332 -4821
rect 1336 -4825 1446 -4821
rect 1467 -4825 1498 -4821
rect -1218 -4832 -1195 -4828
rect -1176 -4832 -1157 -4828
rect -889 -4832 -866 -4828
rect -847 -4832 -828 -4828
rect -531 -4832 -508 -4828
rect -489 -4832 -470 -4828
rect -173 -4832 -150 -4828
rect -131 -4832 -112 -4828
rect 255 -4832 278 -4828
rect 297 -4832 316 -4828
rect 611 -4832 634 -4828
rect 653 -4832 672 -4828
rect 1009 -4832 1032 -4828
rect 1051 -4832 1070 -4828
rect 1367 -4832 1390 -4828
rect 1409 -4832 1428 -4828
rect 1633 -4843 1695 -4726
rect -1421 -4847 -1255 -4843
rect -1251 -4847 -1238 -4843
rect -1234 -4847 -1197 -4843
rect -1193 -4847 -1155 -4843
rect -1151 -4847 -1113 -4843
rect -1109 -4847 -1072 -4843
rect -1068 -4847 -926 -4843
rect -922 -4847 -909 -4843
rect -905 -4847 -868 -4843
rect -864 -4847 -826 -4843
rect -822 -4847 -784 -4843
rect -780 -4847 -743 -4843
rect -739 -4847 -568 -4843
rect -564 -4847 -551 -4843
rect -547 -4847 -510 -4843
rect -506 -4847 -468 -4843
rect -464 -4847 -426 -4843
rect -422 -4847 -385 -4843
rect -381 -4847 -210 -4843
rect -206 -4847 -193 -4843
rect -189 -4847 -152 -4843
rect -148 -4847 -110 -4843
rect -106 -4847 -68 -4843
rect -64 -4847 -27 -4843
rect -23 -4847 90 -4843
rect 94 -4847 218 -4843
rect 222 -4847 235 -4843
rect 239 -4847 276 -4843
rect 280 -4847 318 -4843
rect 322 -4847 360 -4843
rect 364 -4847 401 -4843
rect 405 -4847 574 -4843
rect 578 -4847 591 -4843
rect 595 -4847 632 -4843
rect 636 -4847 674 -4843
rect 678 -4847 716 -4843
rect 720 -4847 757 -4843
rect 761 -4847 972 -4843
rect 976 -4847 989 -4843
rect 993 -4847 1030 -4843
rect 1034 -4847 1072 -4843
rect 1076 -4847 1114 -4843
rect 1118 -4847 1155 -4843
rect 1159 -4847 1330 -4843
rect 1334 -4847 1347 -4843
rect 1351 -4847 1388 -4843
rect 1392 -4847 1430 -4843
rect 1434 -4847 1472 -4843
rect 1476 -4847 1513 -4843
rect 1517 -4847 1695 -4843
rect -1495 -4873 -1255 -4869
rect -1251 -4873 -1238 -4869
rect -1234 -4873 -1218 -4869
rect -1214 -4873 -1197 -4869
rect -1193 -4873 -1176 -4869
rect -1172 -4873 -1155 -4869
rect -1151 -4873 -1134 -4869
rect -1130 -4873 -1113 -4869
rect -1109 -4873 -1092 -4869
rect -1088 -4873 -1072 -4869
rect -1068 -4873 -926 -4869
rect -922 -4873 -909 -4869
rect -905 -4873 -889 -4869
rect -885 -4873 -868 -4869
rect -864 -4873 -847 -4869
rect -843 -4873 -826 -4869
rect -822 -4873 -805 -4869
rect -801 -4873 -784 -4869
rect -780 -4873 -763 -4869
rect -759 -4873 -743 -4869
rect -739 -4873 -568 -4869
rect -564 -4873 -551 -4869
rect -547 -4873 -531 -4869
rect -527 -4873 -510 -4869
rect -506 -4873 -489 -4869
rect -485 -4873 -468 -4869
rect -464 -4873 -447 -4869
rect -443 -4873 -426 -4869
rect -422 -4873 -405 -4869
rect -401 -4873 -385 -4869
rect -381 -4873 -210 -4869
rect -206 -4873 -193 -4869
rect -189 -4873 -173 -4869
rect -169 -4873 -152 -4869
rect -148 -4873 -131 -4869
rect -127 -4873 -110 -4869
rect -106 -4873 -89 -4869
rect -85 -4873 -68 -4869
rect -64 -4873 -47 -4869
rect -43 -4873 -27 -4869
rect -23 -4873 218 -4869
rect 222 -4873 235 -4869
rect 239 -4873 255 -4869
rect 259 -4873 276 -4869
rect 280 -4873 297 -4869
rect 301 -4873 318 -4869
rect 322 -4873 339 -4869
rect 343 -4873 360 -4869
rect 364 -4873 381 -4869
rect 385 -4873 401 -4869
rect 405 -4873 1617 -4869
rect -1495 -4986 -1433 -4873
rect -1233 -4921 -1199 -4917
rect -1135 -4921 -1115 -4917
rect -1100 -4921 -931 -4917
rect -904 -4921 -870 -4917
rect -806 -4921 -786 -4917
rect -771 -4921 -573 -4917
rect -546 -4921 -512 -4917
rect -448 -4921 -428 -4917
rect -413 -4921 -215 -4917
rect -188 -4921 -154 -4917
rect -90 -4921 -70 -4917
rect -55 -4921 213 -4917
rect 240 -4921 274 -4917
rect 338 -4921 358 -4917
rect 373 -4921 407 -4917
rect -935 -4925 -931 -4921
rect -577 -4925 -573 -4921
rect -219 -4925 -215 -4921
rect 209 -4925 213 -4921
rect -1421 -4929 -1257 -4925
rect -1253 -4929 -1223 -4925
rect -1202 -4929 -1171 -4925
rect -1142 -4929 -1111 -4925
rect -1100 -4929 -1073 -4925
rect -935 -4929 -928 -4925
rect -924 -4929 -894 -4925
rect -873 -4929 -842 -4925
rect -813 -4929 -782 -4925
rect -771 -4929 -744 -4925
rect -577 -4929 -570 -4925
rect -566 -4929 -536 -4925
rect -515 -4929 -484 -4925
rect -455 -4929 -424 -4925
rect -413 -4929 -386 -4925
rect -219 -4929 -212 -4925
rect -208 -4929 -178 -4925
rect -157 -4929 -126 -4925
rect -97 -4929 -66 -4925
rect -55 -4929 -28 -4925
rect 209 -4929 216 -4925
rect 220 -4929 250 -4925
rect 271 -4929 302 -4925
rect 331 -4929 362 -4925
rect 373 -4929 400 -4925
rect -1260 -4936 -1213 -4932
rect -1177 -4936 -1164 -4932
rect -1160 -4936 -1129 -4932
rect -1093 -4936 -1080 -4932
rect -1076 -4936 -1064 -4932
rect -931 -4936 -884 -4932
rect -848 -4936 -835 -4932
rect -831 -4936 -800 -4932
rect -764 -4936 -751 -4932
rect -747 -4936 -735 -4932
rect -573 -4936 -526 -4932
rect -490 -4936 -477 -4932
rect -473 -4936 -442 -4932
rect -406 -4936 -393 -4932
rect -389 -4936 -377 -4932
rect -215 -4936 -168 -4932
rect -132 -4936 -119 -4932
rect -115 -4936 -84 -4932
rect -48 -4936 -35 -4932
rect -31 -4936 -19 -4932
rect 213 -4936 260 -4932
rect 296 -4936 309 -4932
rect 313 -4936 344 -4932
rect 380 -4936 393 -4932
rect 397 -4936 409 -4932
rect -1271 -4943 -1253 -4939
rect -1249 -4943 -1139 -4939
rect -1118 -4943 -1087 -4939
rect -936 -4943 -924 -4939
rect -920 -4943 -810 -4939
rect -789 -4943 -758 -4939
rect -579 -4943 -566 -4939
rect -562 -4943 -452 -4939
rect -431 -4943 -400 -4939
rect -221 -4943 -208 -4939
rect -204 -4943 -94 -4939
rect -73 -4943 -42 -4939
rect 206 -4943 220 -4939
rect 224 -4943 334 -4939
rect 355 -4943 386 -4939
rect -1218 -4950 -1195 -4946
rect -1176 -4950 -1157 -4946
rect -889 -4950 -866 -4946
rect -847 -4950 -828 -4946
rect -531 -4950 -508 -4946
rect -489 -4950 -470 -4946
rect -173 -4950 -150 -4946
rect -131 -4950 -112 -4946
rect 255 -4950 278 -4946
rect 297 -4950 316 -4946
rect 1633 -4961 1695 -4847
rect -1421 -4965 -1255 -4961
rect -1251 -4965 -1238 -4961
rect -1234 -4965 -1197 -4961
rect -1193 -4965 -1155 -4961
rect -1151 -4965 -1113 -4961
rect -1109 -4965 -1072 -4961
rect -1068 -4965 -926 -4961
rect -922 -4965 -909 -4961
rect -905 -4965 -868 -4961
rect -864 -4965 -826 -4961
rect -822 -4965 -784 -4961
rect -780 -4965 -743 -4961
rect -739 -4965 -568 -4961
rect -564 -4965 -551 -4961
rect -547 -4965 -510 -4961
rect -506 -4965 -468 -4961
rect -464 -4965 -426 -4961
rect -422 -4965 -385 -4961
rect -381 -4965 -210 -4961
rect -206 -4965 -193 -4961
rect -189 -4965 -152 -4961
rect -148 -4965 -110 -4961
rect -106 -4965 -68 -4961
rect -64 -4965 -27 -4961
rect -23 -4965 218 -4961
rect 222 -4965 235 -4961
rect 239 -4965 276 -4961
rect 280 -4965 318 -4961
rect 322 -4965 360 -4961
rect 364 -4965 401 -4961
rect 405 -4965 1695 -4961
rect -1495 -4990 -1339 -4986
rect -1335 -4990 -1322 -4986
rect -1318 -4990 -935 -4986
rect -931 -4990 -918 -4986
rect -914 -4990 -577 -4986
rect -573 -4990 -560 -4986
rect -556 -4990 -219 -4986
rect -215 -4990 -202 -4986
rect -198 -4990 209 -4986
rect 213 -4990 226 -4986
rect 230 -4990 565 -4986
rect 569 -4990 582 -4986
rect 586 -4990 963 -4986
rect 967 -4990 980 -4986
rect 984 -4990 1321 -4986
rect 1325 -4990 1338 -4986
rect 1342 -4990 1617 -4986
rect -1495 -5105 -1433 -4990
rect -1334 -5022 -1066 -5018
rect -930 -5022 -737 -5018
rect -572 -5022 -379 -5018
rect -214 -5022 -21 -5018
rect 214 -5022 413 -5018
rect 566 -5022 763 -5018
rect 968 -5022 1161 -5018
rect 1326 -5022 1519 -5018
rect -1323 -5030 -923 -5026
rect -919 -5030 -565 -5026
rect -561 -5030 -207 -5026
rect -203 -5030 221 -5026
rect 225 -5030 407 -5026
rect 411 -5030 577 -5026
rect 581 -5030 975 -5026
rect 979 -5030 1333 -5026
rect 1337 -5030 1617 -5026
rect -949 -5043 -909 -5039
rect -591 -5043 -551 -5039
rect -233 -5043 -193 -5039
rect 195 -5043 235 -5039
rect 551 -5043 591 -5039
rect 949 -5043 989 -5039
rect 1307 -5043 1347 -5039
rect 1633 -5078 1695 -4965
rect -1421 -5082 -1322 -5078
rect -1318 -5082 -918 -5078
rect -914 -5082 -560 -5078
rect -556 -5082 -202 -5078
rect -198 -5082 226 -5078
rect 230 -5082 582 -5078
rect 586 -5082 980 -5078
rect 984 -5082 1338 -5078
rect 1342 -5082 1695 -5078
rect -1495 -5109 -1255 -5105
rect -1251 -5109 -1238 -5105
rect -1234 -5109 -1198 -5105
rect -1194 -5109 -1177 -5105
rect -1173 -5109 -926 -5105
rect -922 -5109 -900 -5105
rect -896 -5109 -883 -5105
rect -879 -5109 -843 -5105
rect -839 -5109 -822 -5105
rect -818 -5109 -805 -5105
rect -801 -5109 -765 -5105
rect -761 -5109 -741 -5105
rect -737 -5109 -704 -5105
rect -700 -5109 -568 -5105
rect -564 -5109 -542 -5105
rect -538 -5109 -525 -5105
rect -521 -5109 -485 -5105
rect -481 -5109 -464 -5105
rect -460 -5109 -447 -5105
rect -443 -5109 -407 -5105
rect -403 -5109 -383 -5105
rect -379 -5109 -346 -5105
rect -342 -5109 -210 -5105
rect -206 -5109 -184 -5105
rect -180 -5109 -167 -5105
rect -163 -5109 -127 -5105
rect -123 -5109 -106 -5105
rect -102 -5109 -89 -5105
rect -85 -5109 -49 -5105
rect -45 -5109 -25 -5105
rect -21 -5109 12 -5105
rect 16 -5109 218 -5105
rect 222 -5109 244 -5105
rect 248 -5109 261 -5105
rect 265 -5109 301 -5105
rect 305 -5109 322 -5105
rect 326 -5109 339 -5105
rect 343 -5109 379 -5105
rect 383 -5109 403 -5105
rect 407 -5109 440 -5105
rect 444 -5109 574 -5105
rect 578 -5109 600 -5105
rect 604 -5109 617 -5105
rect 621 -5109 657 -5105
rect 661 -5109 678 -5105
rect 682 -5109 695 -5105
rect 699 -5109 735 -5105
rect 739 -5109 759 -5105
rect 763 -5109 796 -5105
rect 800 -5109 972 -5105
rect 976 -5109 998 -5105
rect 1002 -5109 1015 -5105
rect 1019 -5109 1055 -5105
rect 1059 -5109 1076 -5105
rect 1080 -5109 1093 -5105
rect 1097 -5109 1133 -5105
rect 1137 -5109 1157 -5105
rect 1161 -5109 1194 -5105
rect 1198 -5109 1330 -5105
rect 1334 -5109 1356 -5105
rect 1360 -5109 1373 -5105
rect 1377 -5109 1413 -5105
rect 1417 -5109 1434 -5105
rect 1438 -5109 1451 -5105
rect 1455 -5109 1491 -5105
rect 1495 -5109 1515 -5105
rect 1519 -5109 1552 -5105
rect 1556 -5109 1617 -5105
rect -1495 -5224 -1433 -5109
rect -926 -5113 -922 -5109
rect -900 -5113 -896 -5109
rect -883 -5113 -879 -5109
rect -843 -5113 -839 -5109
rect -822 -5113 -818 -5109
rect -805 -5113 -801 -5109
rect -765 -5113 -761 -5109
rect -741 -5113 -737 -5109
rect -704 -5113 -700 -5109
rect -568 -5113 -564 -5109
rect -542 -5113 -538 -5109
rect -525 -5113 -521 -5109
rect -485 -5113 -481 -5109
rect -464 -5113 -460 -5109
rect -447 -5113 -443 -5109
rect -407 -5113 -403 -5109
rect -383 -5113 -379 -5109
rect -346 -5113 -342 -5109
rect -210 -5113 -206 -5109
rect -184 -5113 -180 -5109
rect -167 -5113 -163 -5109
rect -127 -5113 -123 -5109
rect -106 -5113 -102 -5109
rect -89 -5113 -85 -5109
rect -49 -5113 -45 -5109
rect -25 -5113 -21 -5109
rect 12 -5113 16 -5109
rect 218 -5113 222 -5109
rect 244 -5113 248 -5109
rect 261 -5113 265 -5109
rect 301 -5113 305 -5109
rect 322 -5113 326 -5109
rect 339 -5113 343 -5109
rect 379 -5113 383 -5109
rect 403 -5113 407 -5109
rect 440 -5113 444 -5109
rect 574 -5113 578 -5109
rect 600 -5113 604 -5109
rect 617 -5113 621 -5109
rect 657 -5113 661 -5109
rect 678 -5113 682 -5109
rect 695 -5113 699 -5109
rect 735 -5113 739 -5109
rect 759 -5113 763 -5109
rect 796 -5113 800 -5109
rect 972 -5113 976 -5109
rect 998 -5113 1002 -5109
rect 1015 -5113 1019 -5109
rect 1055 -5113 1059 -5109
rect 1076 -5113 1080 -5109
rect 1093 -5113 1097 -5109
rect 1133 -5113 1137 -5109
rect 1157 -5113 1161 -5109
rect 1194 -5113 1198 -5109
rect 1330 -5113 1334 -5109
rect 1356 -5113 1360 -5109
rect 1373 -5113 1377 -5109
rect 1413 -5113 1417 -5109
rect 1434 -5113 1438 -5109
rect 1451 -5113 1455 -5109
rect 1491 -5113 1495 -5109
rect 1515 -5113 1519 -5109
rect 1552 -5113 1556 -5109
rect -920 -5128 -858 -5124
rect -854 -5128 -824 -5124
rect -776 -5128 -746 -5124
rect -562 -5128 -500 -5124
rect -496 -5128 -466 -5124
rect -418 -5128 -388 -5124
rect -204 -5128 -142 -5124
rect -138 -5128 -108 -5124
rect -60 -5128 -30 -5124
rect 224 -5128 286 -5124
rect 290 -5128 320 -5124
rect 368 -5128 398 -5124
rect 580 -5128 642 -5124
rect 646 -5128 676 -5124
rect 724 -5128 754 -5124
rect 978 -5128 1040 -5124
rect 1044 -5128 1074 -5124
rect 1122 -5128 1152 -5124
rect 1336 -5128 1398 -5124
rect 1402 -5128 1432 -5124
rect 1480 -5128 1510 -5124
rect -913 -5135 -882 -5131
rect -555 -5135 -524 -5131
rect -197 -5135 -166 -5131
rect 231 -5135 262 -5131
rect 587 -5135 618 -5131
rect 985 -5135 1016 -5131
rect 1343 -5135 1374 -5131
rect -931 -5142 -848 -5138
rect -809 -5142 -706 -5138
rect -573 -5142 -490 -5138
rect -451 -5142 -348 -5138
rect -215 -5142 -132 -5138
rect -93 -5142 10 -5138
rect 213 -5142 296 -5138
rect 335 -5142 438 -5138
rect 569 -5142 652 -5138
rect 691 -5142 794 -5138
rect 967 -5142 1050 -5138
rect 1089 -5142 1192 -5138
rect 1325 -5142 1408 -5138
rect 1447 -5142 1550 -5138
rect -949 -5149 -928 -5145
rect -894 -5149 -865 -5145
rect -861 -5149 -780 -5145
rect -691 -5149 -592 -5145
rect -585 -5149 -570 -5145
rect -536 -5149 -507 -5145
rect -503 -5149 -422 -5145
rect -333 -5148 -234 -5144
rect -596 -5153 -592 -5149
rect -238 -5153 -234 -5148
rect -227 -5149 -212 -5145
rect -178 -5149 -149 -5145
rect -145 -5149 -64 -5145
rect 25 -5149 194 -5145
rect 201 -5149 216 -5145
rect 250 -5149 279 -5145
rect 283 -5149 364 -5145
rect 453 -5149 550 -5145
rect 557 -5149 572 -5145
rect 606 -5149 635 -5145
rect 639 -5149 720 -5145
rect 809 -5149 948 -5145
rect 955 -5149 970 -5145
rect 1004 -5149 1033 -5145
rect 1037 -5149 1118 -5145
rect 1207 -5147 1300 -5143
rect 190 -5153 194 -5149
rect 546 -5153 550 -5149
rect 944 -5153 948 -5149
rect 1296 -5153 1300 -5147
rect 1307 -5149 1328 -5145
rect 1362 -5149 1391 -5145
rect 1395 -5149 1476 -5145
rect -1260 -5158 -1203 -5154
rect -1164 -5157 -902 -5153
rect -887 -5157 -804 -5153
rect -783 -5157 -689 -5153
rect -596 -5157 -544 -5153
rect -529 -5157 -446 -5153
rect -425 -5157 -331 -5153
rect -238 -5157 -186 -5153
rect -171 -5157 -88 -5153
rect -67 -5157 27 -5153
rect 190 -5157 242 -5153
rect 257 -5157 340 -5153
rect 361 -5157 455 -5153
rect 546 -5157 598 -5153
rect 613 -5157 696 -5153
rect 717 -5157 811 -5153
rect 944 -5157 996 -5153
rect 1011 -5157 1094 -5153
rect 1115 -5157 1209 -5153
rect 1296 -5157 1354 -5153
rect 1369 -5157 1452 -5153
rect 1473 -5157 1567 -5153
rect -1266 -5165 -1253 -5161
rect -1249 -5165 -1213 -5161
rect -1209 -5165 -1193 -5161
rect -943 -5164 -924 -5160
rect -905 -5164 -776 -5160
rect -591 -5164 -566 -5160
rect -547 -5164 -418 -5160
rect -233 -5164 -208 -5160
rect -189 -5164 -60 -5160
rect 195 -5164 220 -5160
rect 239 -5164 368 -5160
rect 551 -5164 576 -5160
rect 595 -5164 724 -5160
rect 949 -5164 974 -5160
rect 993 -5164 1122 -5160
rect 1313 -5164 1332 -5160
rect 1351 -5164 1480 -5160
rect -1309 -5172 -1257 -5168
rect -1253 -5172 -1227 -5168
rect -1223 -5172 -1179 -5168
rect -898 -5171 -794 -5167
rect -790 -5171 -760 -5167
rect -540 -5171 -436 -5167
rect -432 -5171 -402 -5167
rect -182 -5171 -78 -5167
rect -74 -5171 -44 -5167
rect 246 -5171 350 -5167
rect 354 -5171 384 -5167
rect 602 -5171 706 -5167
rect 710 -5171 740 -5167
rect 1000 -5171 1104 -5167
rect 1108 -5171 1138 -5167
rect 1358 -5171 1462 -5167
rect 1466 -5171 1496 -5167
rect -1216 -5179 -1162 -5175
rect -924 -5178 -872 -5174
rect -868 -5178 -838 -5174
rect -566 -5178 -514 -5174
rect -510 -5178 -480 -5174
rect -208 -5178 -156 -5174
rect -152 -5178 -122 -5174
rect 220 -5178 272 -5174
rect 276 -5178 306 -5174
rect 576 -5178 628 -5174
rect 632 -5178 662 -5174
rect 974 -5178 1026 -5174
rect 1030 -5178 1060 -5174
rect 1332 -5178 1384 -5174
rect 1388 -5178 1418 -5174
rect -1234 -5186 -1202 -5182
rect -879 -5186 -847 -5182
rect -883 -5189 -879 -5186
rect -847 -5189 -843 -5186
rect -801 -5186 -769 -5182
rect -805 -5189 -801 -5186
rect -769 -5189 -765 -5186
rect -521 -5186 -489 -5182
rect -525 -5189 -521 -5186
rect -489 -5189 -485 -5186
rect -443 -5186 -411 -5182
rect -447 -5189 -443 -5186
rect -411 -5189 -407 -5186
rect -163 -5186 -131 -5182
rect -167 -5189 -163 -5186
rect -131 -5189 -127 -5186
rect -85 -5186 -53 -5182
rect -89 -5189 -85 -5186
rect -53 -5189 -49 -5186
rect 265 -5186 297 -5182
rect 261 -5189 265 -5186
rect 297 -5189 301 -5186
rect 343 -5186 375 -5182
rect 339 -5189 343 -5186
rect 375 -5189 379 -5186
rect 621 -5186 653 -5182
rect 617 -5189 621 -5186
rect 653 -5189 657 -5186
rect 699 -5186 731 -5182
rect 695 -5189 699 -5186
rect 731 -5189 735 -5186
rect 1019 -5186 1051 -5182
rect 1015 -5189 1019 -5186
rect 1051 -5189 1055 -5186
rect 1097 -5186 1129 -5182
rect 1093 -5189 1097 -5186
rect 1129 -5189 1133 -5186
rect 1377 -5186 1409 -5182
rect 1373 -5189 1377 -5186
rect 1409 -5189 1413 -5186
rect 1455 -5186 1487 -5182
rect 1451 -5189 1455 -5186
rect 1487 -5189 1491 -5186
rect -926 -5197 -922 -5193
rect -900 -5197 -896 -5193
rect -857 -5197 -853 -5193
rect -822 -5197 -818 -5193
rect -778 -5197 -774 -5193
rect -761 -5197 -757 -5193
rect -725 -5197 -721 -5193
rect -704 -5197 -700 -5193
rect -568 -5197 -564 -5193
rect -542 -5197 -538 -5193
rect -499 -5197 -495 -5193
rect -464 -5197 -460 -5193
rect -420 -5197 -416 -5193
rect -403 -5197 -399 -5193
rect -367 -5197 -363 -5193
rect -346 -5197 -342 -5193
rect -210 -5197 -206 -5193
rect -184 -5197 -180 -5193
rect -141 -5197 -137 -5193
rect -106 -5197 -102 -5193
rect -62 -5197 -58 -5193
rect -45 -5197 -41 -5193
rect -9 -5197 -5 -5193
rect 12 -5197 16 -5193
rect 218 -5197 222 -5193
rect 244 -5197 248 -5193
rect 287 -5197 291 -5193
rect 322 -5197 326 -5193
rect 366 -5197 370 -5193
rect 383 -5197 387 -5193
rect 419 -5197 423 -5193
rect 440 -5197 444 -5193
rect 574 -5197 578 -5193
rect 600 -5197 604 -5193
rect 643 -5197 647 -5193
rect 678 -5197 682 -5193
rect 722 -5197 726 -5193
rect 739 -5197 743 -5193
rect 775 -5197 779 -5193
rect 796 -5197 800 -5193
rect 972 -5197 976 -5193
rect 998 -5197 1002 -5193
rect 1041 -5197 1045 -5193
rect 1076 -5197 1080 -5193
rect 1120 -5197 1124 -5193
rect 1137 -5197 1141 -5193
rect 1173 -5197 1177 -5193
rect 1194 -5197 1198 -5193
rect 1330 -5197 1334 -5193
rect 1356 -5197 1360 -5193
rect 1399 -5197 1403 -5193
rect 1434 -5197 1438 -5193
rect 1478 -5197 1482 -5193
rect 1495 -5197 1499 -5193
rect 1531 -5197 1535 -5193
rect 1552 -5197 1556 -5193
rect 1633 -5197 1695 -5082
rect -1421 -5201 -1255 -5197
rect -1251 -5201 -1211 -5197
rect -1207 -5201 -1177 -5197
rect -1173 -5201 -926 -5197
rect -922 -5201 -900 -5197
rect -896 -5201 -857 -5197
rect -853 -5201 -822 -5197
rect -818 -5201 -778 -5197
rect -774 -5201 -761 -5197
rect -757 -5201 -725 -5197
rect -721 -5201 -704 -5197
rect -700 -5201 -568 -5197
rect -564 -5201 -542 -5197
rect -538 -5201 -499 -5197
rect -495 -5201 -464 -5197
rect -460 -5201 -420 -5197
rect -416 -5201 -403 -5197
rect -399 -5201 -367 -5197
rect -363 -5201 -346 -5197
rect -342 -5201 -210 -5197
rect -206 -5201 -184 -5197
rect -180 -5201 -141 -5197
rect -137 -5201 -106 -5197
rect -102 -5201 -62 -5197
rect -58 -5201 -45 -5197
rect -41 -5201 -9 -5197
rect -5 -5201 12 -5197
rect 16 -5201 218 -5197
rect 222 -5201 244 -5197
rect 248 -5201 287 -5197
rect 291 -5201 322 -5197
rect 326 -5201 366 -5197
rect 370 -5201 383 -5197
rect 387 -5201 419 -5197
rect 423 -5201 440 -5197
rect 444 -5201 574 -5197
rect 578 -5201 600 -5197
rect 604 -5201 643 -5197
rect 647 -5201 678 -5197
rect 682 -5201 722 -5197
rect 726 -5201 739 -5197
rect 743 -5201 775 -5197
rect 779 -5201 796 -5197
rect 800 -5201 972 -5197
rect 976 -5201 998 -5197
rect 1002 -5201 1041 -5197
rect 1045 -5201 1076 -5197
rect 1080 -5201 1120 -5197
rect 1124 -5201 1137 -5197
rect 1141 -5201 1173 -5197
rect 1177 -5201 1194 -5197
rect 1198 -5201 1330 -5197
rect 1334 -5201 1356 -5197
rect 1360 -5201 1399 -5197
rect 1403 -5201 1434 -5197
rect 1438 -5201 1478 -5197
rect 1482 -5201 1495 -5197
rect 1499 -5201 1531 -5197
rect 1535 -5201 1552 -5197
rect 1556 -5201 1695 -5197
rect -1272 -5208 -689 -5204
rect -585 -5208 27 -5204
rect 201 -5208 811 -5204
rect 955 -5208 1567 -5204
rect -1266 -5216 -1162 -5212
rect -943 -5215 -331 -5211
rect -227 -5215 455 -5211
rect 557 -5215 1209 -5211
rect 1313 -5215 1561 -5211
rect -1495 -5228 -1255 -5224
rect -1251 -5228 -1238 -5224
rect -1234 -5228 -1218 -5224
rect -1214 -5228 -1197 -5224
rect -1193 -5228 -1176 -5224
rect -1172 -5228 -1155 -5224
rect -1151 -5228 -1134 -5224
rect -1130 -5228 -1113 -5224
rect -1109 -5228 -1092 -5224
rect -1088 -5228 -1072 -5224
rect -1068 -5228 -926 -5224
rect -922 -5228 -909 -5224
rect -905 -5228 -889 -5224
rect -885 -5228 -868 -5224
rect -864 -5228 -847 -5224
rect -843 -5228 -826 -5224
rect -822 -5228 -805 -5224
rect -801 -5228 -784 -5224
rect -780 -5228 -763 -5224
rect -759 -5228 -743 -5224
rect -739 -5228 1617 -5224
rect -1495 -5345 -1433 -5228
rect -1233 -5276 -1199 -5272
rect -1135 -5276 -1115 -5272
rect -1100 -5276 -931 -5272
rect -904 -5276 -870 -5272
rect -806 -5276 -786 -5272
rect -771 -5276 -735 -5272
rect -935 -5280 -931 -5276
rect -1266 -5284 -1257 -5280
rect -1253 -5284 -1223 -5280
rect -1202 -5284 -1171 -5280
rect -1142 -5284 -1111 -5280
rect -1100 -5284 -1073 -5280
rect -935 -5284 -928 -5280
rect -924 -5284 -894 -5280
rect -873 -5284 -842 -5280
rect -813 -5284 -782 -5280
rect -771 -5284 -744 -5280
rect -1260 -5291 -1213 -5287
rect -1177 -5291 -1164 -5287
rect -1160 -5291 -1129 -5287
rect -1093 -5291 -1080 -5287
rect -1076 -5291 -1064 -5287
rect -931 -5291 -884 -5287
rect -848 -5291 -835 -5287
rect -831 -5291 -800 -5287
rect -764 -5291 -751 -5287
rect -747 -5291 -735 -5287
rect -1266 -5298 -1253 -5294
rect -1249 -5298 -1139 -5294
rect -1118 -5298 -1087 -5294
rect -938 -5298 -924 -5294
rect -920 -5298 -810 -5294
rect -789 -5298 -758 -5294
rect -1218 -5305 -1195 -5301
rect -1176 -5305 -1157 -5301
rect -889 -5305 -866 -5301
rect -847 -5305 -828 -5301
rect 1633 -5316 1695 -5201
rect -1421 -5320 -1255 -5316
rect -1251 -5320 -1238 -5316
rect -1234 -5320 -1197 -5316
rect -1193 -5320 -1155 -5316
rect -1151 -5320 -1113 -5316
rect -1109 -5320 -1072 -5316
rect -1068 -5320 -926 -5316
rect -922 -5320 -909 -5316
rect -905 -5320 -868 -5316
rect -864 -5320 -826 -5316
rect -822 -5320 -784 -5316
rect -780 -5320 -743 -5316
rect -739 -5320 1695 -5316
rect -1495 -5349 -1255 -5345
rect -1251 -5349 -1238 -5345
rect -1234 -5349 -1218 -5345
rect -1214 -5349 -1197 -5345
rect -1193 -5349 -1176 -5345
rect -1172 -5349 -1155 -5345
rect -1151 -5349 -1134 -5345
rect -1130 -5349 -1113 -5345
rect -1109 -5349 -1092 -5345
rect -1088 -5349 -1072 -5345
rect -1068 -5349 -1026 -5345
rect -1022 -5349 -926 -5345
rect -922 -5349 -909 -5345
rect -905 -5349 -889 -5345
rect -885 -5349 -868 -5345
rect -864 -5349 -847 -5345
rect -843 -5349 -826 -5345
rect -822 -5349 -805 -5345
rect -801 -5349 -784 -5345
rect -780 -5349 -763 -5345
rect -759 -5349 -743 -5345
rect -739 -5349 -673 -5345
rect -669 -5349 -568 -5345
rect -564 -5349 -551 -5345
rect -547 -5349 -531 -5345
rect -527 -5349 -510 -5345
rect -506 -5349 -489 -5345
rect -485 -5349 -468 -5345
rect -464 -5349 -447 -5345
rect -443 -5349 -426 -5345
rect -422 -5349 -405 -5345
rect -401 -5349 -385 -5345
rect -381 -5349 -327 -5345
rect -323 -5349 -210 -5345
rect -206 -5349 -193 -5345
rect -189 -5349 -173 -5345
rect -169 -5349 -152 -5345
rect -148 -5349 -131 -5345
rect -127 -5349 -110 -5345
rect -106 -5349 -89 -5345
rect -85 -5349 -68 -5345
rect -64 -5349 -47 -5345
rect -43 -5349 -27 -5345
rect -23 -5349 218 -5345
rect 222 -5349 235 -5345
rect 239 -5349 255 -5345
rect 259 -5349 276 -5345
rect 280 -5349 297 -5345
rect 301 -5349 318 -5345
rect 322 -5349 339 -5345
rect 343 -5349 360 -5345
rect 364 -5349 381 -5345
rect 385 -5349 401 -5345
rect 405 -5349 466 -5345
rect 470 -5349 574 -5345
rect 578 -5349 591 -5345
rect 595 -5349 611 -5345
rect 615 -5349 632 -5345
rect 636 -5349 653 -5345
rect 657 -5349 674 -5345
rect 678 -5349 695 -5345
rect 699 -5349 716 -5345
rect 720 -5349 737 -5345
rect 741 -5349 757 -5345
rect 761 -5349 867 -5345
rect 871 -5349 972 -5345
rect 976 -5349 989 -5345
rect 993 -5349 1009 -5345
rect 1013 -5349 1030 -5345
rect 1034 -5349 1051 -5345
rect 1055 -5349 1072 -5345
rect 1076 -5349 1093 -5345
rect 1097 -5349 1114 -5345
rect 1118 -5349 1135 -5345
rect 1139 -5349 1155 -5345
rect 1159 -5349 1210 -5345
rect 1214 -5349 1330 -5345
rect 1334 -5349 1347 -5345
rect 1351 -5349 1367 -5345
rect 1371 -5349 1388 -5345
rect 1392 -5349 1409 -5345
rect 1413 -5349 1430 -5345
rect 1434 -5349 1451 -5345
rect 1455 -5349 1472 -5345
rect 1476 -5349 1493 -5345
rect 1497 -5349 1513 -5345
rect 1517 -5349 1617 -5345
rect -1495 -5465 -1433 -5349
rect -1233 -5397 -1199 -5393
rect -1135 -5397 -1115 -5393
rect -1100 -5397 -1066 -5393
rect -1014 -5394 -1010 -5390
rect -904 -5397 -870 -5393
rect -806 -5397 -786 -5393
rect -771 -5397 -737 -5393
rect -1272 -5405 -1257 -5401
rect -1253 -5405 -1223 -5401
rect -1202 -5405 -1171 -5401
rect -1142 -5405 -1111 -5401
rect -1100 -5405 -1073 -5401
rect -943 -5405 -928 -5401
rect -924 -5405 -894 -5401
rect -873 -5405 -842 -5401
rect -813 -5405 -782 -5401
rect -771 -5405 -744 -5401
rect -661 -5399 -657 -5395
rect -546 -5397 -512 -5393
rect -448 -5397 -428 -5393
rect -413 -5397 -379 -5393
rect -585 -5405 -570 -5401
rect -566 -5405 -536 -5401
rect -515 -5405 -484 -5401
rect -455 -5405 -424 -5401
rect -413 -5405 -386 -5401
rect -315 -5400 -311 -5396
rect -188 -5397 -154 -5393
rect -90 -5397 -70 -5393
rect -55 -5397 -21 -5393
rect 240 -5397 274 -5393
rect 338 -5397 358 -5393
rect 373 -5397 407 -5393
rect 478 -5394 482 -5390
rect 596 -5397 630 -5393
rect 694 -5397 714 -5393
rect 729 -5397 763 -5393
rect -227 -5405 -212 -5401
rect -208 -5405 -178 -5401
rect -157 -5405 -126 -5401
rect -97 -5405 -66 -5401
rect -55 -5405 -28 -5401
rect 201 -5405 216 -5401
rect 220 -5405 250 -5401
rect 271 -5405 302 -5401
rect 331 -5405 362 -5401
rect 373 -5405 400 -5401
rect 557 -5405 572 -5401
rect 576 -5405 606 -5401
rect 627 -5405 658 -5401
rect 687 -5405 718 -5401
rect 729 -5405 756 -5401
rect 879 -5399 883 -5395
rect 994 -5397 1028 -5393
rect 1092 -5397 1112 -5393
rect 1127 -5397 1161 -5393
rect 955 -5405 970 -5401
rect 974 -5405 1004 -5401
rect 1025 -5405 1056 -5401
rect 1085 -5405 1116 -5401
rect 1127 -5405 1154 -5401
rect 1352 -5397 1386 -5393
rect 1450 -5397 1470 -5393
rect 1485 -5397 1519 -5393
rect 1222 -5403 1226 -5399
rect 1313 -5405 1328 -5401
rect 1332 -5405 1362 -5401
rect 1383 -5405 1414 -5401
rect 1443 -5405 1474 -5401
rect 1485 -5405 1512 -5401
rect -1260 -5412 -1213 -5408
rect -1177 -5412 -1164 -5408
rect -1160 -5412 -1129 -5408
rect -1093 -5412 -1080 -5408
rect -1076 -5412 -1064 -5408
rect -931 -5412 -884 -5408
rect -848 -5412 -835 -5408
rect -831 -5412 -800 -5408
rect -764 -5412 -751 -5408
rect -747 -5412 -735 -5408
rect -573 -5412 -526 -5408
rect -490 -5412 -477 -5408
rect -473 -5412 -442 -5408
rect -406 -5412 -393 -5408
rect -389 -5412 -377 -5408
rect -215 -5412 -168 -5408
rect -132 -5412 -119 -5408
rect -115 -5412 -84 -5408
rect -48 -5412 -35 -5408
rect -31 -5412 -19 -5408
rect 213 -5412 260 -5408
rect 296 -5412 309 -5408
rect 313 -5412 344 -5408
rect 380 -5412 393 -5408
rect 397 -5412 409 -5408
rect 569 -5412 616 -5408
rect 652 -5412 665 -5408
rect 669 -5412 700 -5408
rect 736 -5412 749 -5408
rect 753 -5412 765 -5408
rect 967 -5412 1014 -5408
rect 1050 -5412 1063 -5408
rect 1067 -5412 1098 -5408
rect 1134 -5412 1147 -5408
rect 1151 -5412 1163 -5408
rect 1325 -5412 1372 -5408
rect 1408 -5412 1421 -5408
rect 1425 -5412 1456 -5408
rect 1492 -5412 1505 -5408
rect 1509 -5412 1521 -5408
rect -1266 -5419 -1253 -5415
rect -1249 -5419 -1139 -5415
rect -1118 -5419 -1087 -5415
rect -938 -5419 -924 -5415
rect -920 -5419 -810 -5415
rect -789 -5419 -758 -5415
rect -581 -5419 -566 -5415
rect -562 -5419 -452 -5415
rect -431 -5419 -400 -5415
rect -222 -5419 -208 -5415
rect -204 -5419 -94 -5415
rect -73 -5419 -42 -5415
rect 209 -5419 220 -5415
rect 224 -5419 334 -5415
rect 355 -5419 386 -5415
rect 561 -5419 576 -5415
rect 580 -5419 690 -5415
rect 711 -5419 742 -5415
rect 956 -5419 974 -5415
rect 978 -5419 1088 -5415
rect 1109 -5419 1140 -5415
rect 1317 -5419 1332 -5415
rect 1336 -5419 1446 -5415
rect 1467 -5419 1498 -5415
rect -1218 -5426 -1195 -5422
rect -1176 -5426 -1157 -5422
rect -889 -5426 -866 -5422
rect -847 -5426 -828 -5422
rect -531 -5426 -508 -5422
rect -489 -5426 -470 -5422
rect -173 -5426 -150 -5422
rect -131 -5426 -112 -5422
rect 255 -5426 278 -5422
rect 297 -5426 316 -5422
rect 611 -5426 634 -5422
rect 653 -5426 672 -5422
rect 1009 -5426 1032 -5422
rect 1051 -5426 1070 -5422
rect 1367 -5426 1390 -5422
rect 1409 -5426 1428 -5422
rect 1633 -5437 1695 -5320
rect -1421 -5441 -1255 -5437
rect -1251 -5441 -1238 -5437
rect -1234 -5441 -1197 -5437
rect -1193 -5441 -1155 -5437
rect -1151 -5441 -1113 -5437
rect -1109 -5441 -1072 -5437
rect -1068 -5441 -1026 -5437
rect -1022 -5441 -926 -5437
rect -922 -5441 -909 -5437
rect -905 -5441 -868 -5437
rect -864 -5441 -826 -5437
rect -822 -5441 -784 -5437
rect -780 -5441 -743 -5437
rect -739 -5441 -673 -5437
rect -669 -5441 -568 -5437
rect -564 -5441 -551 -5437
rect -547 -5441 -510 -5437
rect -506 -5441 -468 -5437
rect -464 -5441 -426 -5437
rect -422 -5441 -385 -5437
rect -381 -5441 -327 -5437
rect -323 -5441 -210 -5437
rect -206 -5441 -193 -5437
rect -189 -5441 -152 -5437
rect -148 -5441 -110 -5437
rect -106 -5441 -68 -5437
rect -64 -5441 -27 -5437
rect -23 -5441 218 -5437
rect 222 -5441 235 -5437
rect 239 -5441 276 -5437
rect 280 -5441 318 -5437
rect 322 -5441 360 -5437
rect 364 -5441 401 -5437
rect 405 -5441 466 -5437
rect 470 -5441 574 -5437
rect 578 -5441 591 -5437
rect 595 -5441 632 -5437
rect 636 -5441 674 -5437
rect 678 -5441 716 -5437
rect 720 -5441 757 -5437
rect 761 -5441 867 -5437
rect 871 -5441 972 -5437
rect 976 -5441 989 -5437
rect 993 -5441 1030 -5437
rect 1034 -5441 1072 -5437
rect 1076 -5441 1114 -5437
rect 1118 -5441 1155 -5437
rect 1159 -5441 1210 -5437
rect 1214 -5441 1330 -5437
rect 1334 -5441 1347 -5437
rect 1351 -5441 1388 -5437
rect 1392 -5441 1430 -5437
rect 1434 -5441 1472 -5437
rect 1476 -5441 1513 -5437
rect 1517 -5441 1695 -5437
rect -1266 -5448 -1066 -5444
rect -943 -5448 -737 -5444
rect -585 -5449 -379 -5445
rect -227 -5448 -21 -5444
rect 201 -5448 407 -5444
rect 557 -5450 763 -5446
rect 955 -5449 1161 -5445
rect 1313 -5448 1519 -5444
rect -1495 -5469 -1255 -5465
rect -1251 -5469 -1238 -5465
rect -1234 -5469 -1218 -5465
rect -1214 -5469 -1197 -5465
rect -1193 -5469 -1176 -5465
rect -1172 -5469 -1155 -5465
rect -1151 -5469 -1134 -5465
rect -1130 -5469 -1113 -5465
rect -1109 -5469 -1092 -5465
rect -1088 -5469 -1072 -5465
rect -1068 -5469 -1026 -5465
rect -1022 -5469 -926 -5465
rect -922 -5469 -909 -5465
rect -905 -5469 -889 -5465
rect -885 -5469 -868 -5465
rect -864 -5469 -847 -5465
rect -843 -5469 -826 -5465
rect -822 -5469 -805 -5465
rect -801 -5469 -784 -5465
rect -780 -5469 -763 -5465
rect -759 -5469 -743 -5465
rect -739 -5469 -568 -5465
rect -564 -5469 -551 -5465
rect -547 -5469 -531 -5465
rect -527 -5469 -510 -5465
rect -506 -5469 -489 -5465
rect -485 -5469 -468 -5465
rect -464 -5469 -447 -5465
rect -443 -5469 -426 -5465
rect -422 -5469 -405 -5465
rect -401 -5469 -385 -5465
rect -381 -5469 -327 -5465
rect -323 -5469 -210 -5465
rect -206 -5469 -193 -5465
rect -189 -5469 -173 -5465
rect -169 -5469 -152 -5465
rect -148 -5469 -131 -5465
rect -127 -5469 -110 -5465
rect -106 -5469 -89 -5465
rect -85 -5469 -68 -5465
rect -64 -5469 -47 -5465
rect -43 -5469 -27 -5465
rect -23 -5469 218 -5465
rect 222 -5469 235 -5465
rect 239 -5469 255 -5465
rect 259 -5469 276 -5465
rect 280 -5469 297 -5465
rect 301 -5469 318 -5465
rect 322 -5469 339 -5465
rect 343 -5469 360 -5465
rect 364 -5469 381 -5465
rect 385 -5469 401 -5465
rect 405 -5469 466 -5465
rect 470 -5469 574 -5465
rect 578 -5469 591 -5465
rect 595 -5469 611 -5465
rect 615 -5469 632 -5465
rect 636 -5469 653 -5465
rect 657 -5469 674 -5465
rect 678 -5469 695 -5465
rect 699 -5469 716 -5465
rect 720 -5469 737 -5465
rect 741 -5469 757 -5465
rect 761 -5469 972 -5465
rect 976 -5469 989 -5465
rect 993 -5469 1009 -5465
rect 1013 -5469 1030 -5465
rect 1034 -5469 1051 -5465
rect 1055 -5469 1072 -5465
rect 1076 -5469 1093 -5465
rect 1097 -5469 1114 -5465
rect 1118 -5469 1135 -5465
rect 1139 -5469 1155 -5465
rect 1159 -5469 1210 -5465
rect 1214 -5469 1330 -5465
rect 1334 -5469 1347 -5465
rect 1351 -5469 1367 -5465
rect 1371 -5469 1388 -5465
rect 1392 -5469 1409 -5465
rect 1413 -5469 1430 -5465
rect 1434 -5469 1451 -5465
rect 1455 -5469 1472 -5465
rect 1476 -5469 1493 -5465
rect 1497 -5469 1513 -5465
rect 1517 -5469 1617 -5465
rect -1495 -5582 -1433 -5469
rect -1233 -5517 -1199 -5513
rect -1135 -5517 -1115 -5513
rect -1100 -5517 -1066 -5513
rect -1345 -5525 -1257 -5521
rect -1253 -5525 -1223 -5521
rect -1202 -5525 -1171 -5521
rect -1142 -5525 -1111 -5521
rect -1100 -5525 -1073 -5521
rect -1014 -5518 -1010 -5514
rect -904 -5517 -870 -5513
rect -806 -5517 -786 -5513
rect -771 -5517 -737 -5513
rect -546 -5517 -512 -5513
rect -448 -5517 -428 -5513
rect -413 -5517 -379 -5513
rect -315 -5515 -311 -5511
rect -188 -5517 -154 -5513
rect -90 -5517 -70 -5513
rect -55 -5517 -21 -5513
rect 240 -5517 274 -5513
rect 338 -5517 358 -5513
rect 373 -5517 407 -5513
rect -937 -5525 -928 -5521
rect -924 -5525 -894 -5521
rect -873 -5525 -842 -5521
rect -813 -5525 -782 -5521
rect -771 -5525 -744 -5521
rect -579 -5525 -570 -5521
rect -566 -5525 -536 -5521
rect -515 -5525 -484 -5521
rect -455 -5525 -424 -5521
rect -413 -5525 -386 -5521
rect -221 -5525 -212 -5521
rect -208 -5525 -178 -5521
rect -157 -5525 -126 -5521
rect -97 -5525 -66 -5521
rect -55 -5525 -28 -5521
rect 207 -5525 216 -5521
rect 220 -5525 250 -5521
rect 271 -5525 302 -5521
rect 331 -5525 362 -5521
rect 373 -5525 400 -5521
rect 478 -5518 482 -5514
rect 596 -5517 630 -5513
rect 694 -5517 714 -5513
rect 729 -5517 769 -5513
rect 994 -5517 1028 -5513
rect 1092 -5517 1112 -5513
rect 1127 -5517 1161 -5513
rect 563 -5525 572 -5521
rect 576 -5525 606 -5521
rect 627 -5525 658 -5521
rect 687 -5525 718 -5521
rect 729 -5525 756 -5521
rect 961 -5525 970 -5521
rect 974 -5525 1004 -5521
rect 1025 -5525 1056 -5521
rect 1085 -5525 1116 -5521
rect 1127 -5525 1154 -5521
rect 1222 -5518 1226 -5514
rect 1352 -5517 1386 -5513
rect 1450 -5517 1470 -5513
rect 1485 -5517 1519 -5513
rect 1319 -5525 1328 -5521
rect 1332 -5525 1362 -5521
rect 1383 -5525 1414 -5521
rect 1443 -5525 1474 -5521
rect 1485 -5525 1512 -5521
rect -1260 -5532 -1213 -5528
rect -1177 -5532 -1164 -5528
rect -1160 -5532 -1129 -5528
rect -1093 -5532 -1080 -5528
rect -1076 -5532 -1064 -5528
rect -931 -5532 -884 -5528
rect -848 -5532 -835 -5528
rect -831 -5532 -800 -5528
rect -764 -5532 -751 -5528
rect -747 -5532 -735 -5528
rect -573 -5532 -526 -5528
rect -490 -5532 -477 -5528
rect -473 -5532 -442 -5528
rect -406 -5532 -393 -5528
rect -389 -5532 -377 -5528
rect -215 -5532 -168 -5528
rect -132 -5532 -119 -5528
rect -115 -5532 -84 -5528
rect -48 -5532 -35 -5528
rect -31 -5532 -19 -5528
rect 213 -5532 260 -5528
rect 296 -5532 309 -5528
rect 313 -5532 344 -5528
rect 380 -5532 393 -5528
rect 397 -5532 409 -5528
rect 569 -5532 616 -5528
rect 652 -5532 665 -5528
rect 669 -5532 700 -5528
rect 736 -5532 749 -5528
rect 753 -5532 765 -5528
rect 967 -5532 1014 -5528
rect 1050 -5532 1063 -5528
rect 1067 -5532 1098 -5528
rect 1134 -5532 1147 -5528
rect 1151 -5532 1163 -5528
rect 1325 -5532 1372 -5528
rect 1408 -5532 1421 -5528
rect 1425 -5532 1456 -5528
rect 1492 -5532 1505 -5528
rect 1509 -5532 1521 -5528
rect -1274 -5539 -1253 -5535
rect -1249 -5539 -1139 -5535
rect -1118 -5539 -1087 -5535
rect -937 -5539 -924 -5535
rect -920 -5539 -810 -5535
rect -789 -5539 -758 -5535
rect -577 -5539 -566 -5535
rect -562 -5539 -452 -5535
rect -431 -5539 -400 -5535
rect -223 -5539 -208 -5535
rect -204 -5539 -94 -5535
rect -73 -5539 -42 -5535
rect 207 -5539 220 -5535
rect 224 -5539 334 -5535
rect 355 -5539 386 -5535
rect 565 -5539 576 -5535
rect 580 -5539 690 -5535
rect 711 -5539 742 -5535
rect 957 -5539 974 -5535
rect 978 -5539 1088 -5535
rect 1109 -5539 1140 -5535
rect 1320 -5539 1332 -5535
rect 1336 -5539 1446 -5535
rect 1467 -5539 1498 -5535
rect -1218 -5546 -1195 -5542
rect -1176 -5546 -1157 -5542
rect -889 -5546 -866 -5542
rect -847 -5546 -828 -5542
rect -531 -5546 -508 -5542
rect -489 -5546 -470 -5542
rect -173 -5546 -150 -5542
rect -131 -5546 -112 -5542
rect 255 -5546 278 -5542
rect 297 -5546 316 -5542
rect 611 -5546 634 -5542
rect 653 -5546 672 -5542
rect 1009 -5546 1032 -5542
rect 1051 -5546 1070 -5542
rect 1367 -5546 1390 -5542
rect 1409 -5546 1428 -5542
rect 1633 -5557 1695 -5441
rect -1421 -5561 -1255 -5557
rect -1251 -5561 -1238 -5557
rect -1234 -5561 -1197 -5557
rect -1193 -5561 -1155 -5557
rect -1151 -5561 -1113 -5557
rect -1109 -5561 -1072 -5557
rect -1068 -5561 -1026 -5557
rect -1022 -5561 -926 -5557
rect -922 -5561 -909 -5557
rect -905 -5561 -868 -5557
rect -864 -5561 -826 -5557
rect -822 -5561 -784 -5557
rect -780 -5561 -743 -5557
rect -739 -5561 -568 -5557
rect -564 -5561 -551 -5557
rect -547 -5561 -510 -5557
rect -506 -5561 -468 -5557
rect -464 -5561 -426 -5557
rect -422 -5561 -385 -5557
rect -381 -5561 -327 -5557
rect -323 -5561 -210 -5557
rect -206 -5561 -193 -5557
rect -189 -5561 -152 -5557
rect -148 -5561 -110 -5557
rect -106 -5561 -68 -5557
rect -64 -5561 -27 -5557
rect -23 -5561 218 -5557
rect 222 -5561 235 -5557
rect 239 -5561 276 -5557
rect 280 -5561 318 -5557
rect 322 -5561 360 -5557
rect 364 -5561 401 -5557
rect 405 -5561 466 -5557
rect 470 -5561 574 -5557
rect 578 -5561 591 -5557
rect 595 -5561 632 -5557
rect 636 -5561 674 -5557
rect 678 -5561 716 -5557
rect 720 -5561 757 -5557
rect 761 -5561 972 -5557
rect 976 -5561 989 -5557
rect 993 -5561 1030 -5557
rect 1034 -5561 1072 -5557
rect 1076 -5561 1114 -5557
rect 1118 -5561 1155 -5557
rect 1159 -5561 1210 -5557
rect 1214 -5561 1330 -5557
rect 1334 -5561 1347 -5557
rect 1351 -5561 1388 -5557
rect 1392 -5561 1430 -5557
rect 1434 -5561 1472 -5557
rect 1476 -5561 1513 -5557
rect 1517 -5561 1695 -5557
rect -1495 -5586 -1255 -5582
rect -1251 -5586 -1238 -5582
rect -1234 -5586 -1218 -5582
rect -1214 -5586 -1197 -5582
rect -1193 -5586 -1176 -5582
rect -1172 -5586 -1155 -5582
rect -1151 -5586 -1134 -5582
rect -1130 -5586 -1113 -5582
rect -1109 -5586 -1092 -5582
rect -1088 -5586 -1072 -5582
rect -1068 -5586 -926 -5582
rect -922 -5586 -909 -5582
rect -905 -5586 -889 -5582
rect -885 -5586 -868 -5582
rect -864 -5586 -847 -5582
rect -843 -5586 -826 -5582
rect -822 -5586 -805 -5582
rect -801 -5586 -784 -5582
rect -780 -5586 -763 -5582
rect -759 -5586 -743 -5582
rect -739 -5586 -568 -5582
rect -564 -5586 -551 -5582
rect -547 -5586 -531 -5582
rect -527 -5586 -510 -5582
rect -506 -5586 -489 -5582
rect -485 -5586 -468 -5582
rect -464 -5586 -447 -5582
rect -443 -5586 -426 -5582
rect -422 -5586 -405 -5582
rect -401 -5586 -385 -5582
rect -381 -5586 -210 -5582
rect -206 -5586 -193 -5582
rect -189 -5586 -173 -5582
rect -169 -5586 -152 -5582
rect -148 -5586 -131 -5582
rect -127 -5586 -110 -5582
rect -106 -5586 -89 -5582
rect -85 -5586 -68 -5582
rect -64 -5586 -47 -5582
rect -43 -5586 -27 -5582
rect -23 -5586 218 -5582
rect 222 -5586 235 -5582
rect 239 -5586 255 -5582
rect 259 -5586 276 -5582
rect 280 -5586 297 -5582
rect 301 -5586 318 -5582
rect 322 -5586 339 -5582
rect 343 -5586 360 -5582
rect 364 -5586 381 -5582
rect 385 -5586 401 -5582
rect 405 -5586 574 -5582
rect 578 -5586 591 -5582
rect 595 -5586 611 -5582
rect 615 -5586 632 -5582
rect 636 -5586 653 -5582
rect 657 -5586 674 -5582
rect 678 -5586 695 -5582
rect 699 -5586 716 -5582
rect 720 -5586 737 -5582
rect 741 -5586 757 -5582
rect 761 -5586 1617 -5582
rect -1495 -5699 -1433 -5586
rect -1233 -5634 -1199 -5630
rect -1135 -5634 -1115 -5630
rect -1100 -5634 -931 -5630
rect -904 -5634 -870 -5630
rect -806 -5634 -786 -5630
rect -771 -5634 -573 -5630
rect -546 -5634 -512 -5630
rect -448 -5634 -428 -5630
rect -413 -5634 -215 -5630
rect -188 -5634 -154 -5630
rect -90 -5634 -70 -5630
rect -55 -5634 213 -5630
rect 240 -5634 274 -5630
rect 338 -5634 358 -5630
rect 373 -5634 569 -5630
rect 596 -5634 630 -5630
rect 694 -5634 714 -5630
rect 729 -5634 763 -5630
rect -935 -5638 -931 -5634
rect -577 -5638 -573 -5634
rect -219 -5638 -215 -5634
rect 209 -5638 213 -5634
rect 565 -5638 569 -5634
rect -1421 -5642 -1257 -5638
rect -1253 -5642 -1223 -5638
rect -1202 -5642 -1171 -5638
rect -1142 -5642 -1111 -5638
rect -1100 -5642 -1073 -5638
rect -935 -5642 -928 -5638
rect -924 -5642 -894 -5638
rect -873 -5642 -842 -5638
rect -813 -5642 -782 -5638
rect -771 -5642 -744 -5638
rect -577 -5642 -570 -5638
rect -566 -5642 -536 -5638
rect -515 -5642 -484 -5638
rect -455 -5642 -424 -5638
rect -413 -5642 -386 -5638
rect -219 -5642 -212 -5638
rect -208 -5642 -178 -5638
rect -157 -5642 -126 -5638
rect -97 -5642 -66 -5638
rect -55 -5642 -28 -5638
rect 209 -5642 216 -5638
rect 220 -5642 250 -5638
rect 271 -5642 302 -5638
rect 331 -5642 362 -5638
rect 373 -5642 400 -5638
rect 565 -5642 572 -5638
rect 576 -5642 606 -5638
rect 627 -5642 658 -5638
rect 687 -5642 718 -5638
rect 729 -5642 756 -5638
rect -1260 -5649 -1213 -5645
rect -1177 -5649 -1164 -5645
rect -1160 -5649 -1129 -5645
rect -1093 -5649 -1080 -5645
rect -1076 -5649 -1064 -5645
rect -931 -5649 -884 -5645
rect -848 -5649 -835 -5645
rect -831 -5649 -800 -5645
rect -764 -5649 -751 -5645
rect -747 -5649 -735 -5645
rect -573 -5649 -526 -5645
rect -490 -5649 -477 -5645
rect -473 -5649 -442 -5645
rect -406 -5649 -393 -5645
rect -389 -5649 -377 -5645
rect -215 -5649 -168 -5645
rect -132 -5649 -119 -5645
rect -115 -5649 -84 -5645
rect -48 -5649 -35 -5645
rect -31 -5649 -19 -5645
rect 213 -5649 260 -5645
rect 296 -5649 309 -5645
rect 313 -5649 344 -5645
rect 380 -5649 393 -5645
rect 397 -5649 409 -5645
rect 569 -5649 616 -5645
rect 652 -5649 665 -5645
rect 669 -5649 700 -5645
rect 736 -5649 749 -5645
rect 753 -5649 765 -5645
rect -1274 -5656 -1253 -5652
rect -1249 -5656 -1139 -5652
rect -1118 -5656 -1087 -5652
rect -937 -5656 -924 -5652
rect -920 -5656 -810 -5652
rect -789 -5656 -758 -5652
rect -577 -5656 -566 -5652
rect -562 -5656 -452 -5652
rect -431 -5656 -400 -5652
rect -223 -5656 -208 -5652
rect -204 -5656 -94 -5652
rect -73 -5656 -42 -5652
rect 207 -5656 220 -5652
rect 224 -5656 334 -5652
rect 355 -5656 386 -5652
rect 565 -5656 576 -5652
rect 580 -5656 690 -5652
rect 711 -5656 742 -5652
rect -1218 -5663 -1195 -5659
rect -1176 -5663 -1157 -5659
rect -889 -5663 -866 -5659
rect -847 -5663 -828 -5659
rect -531 -5663 -508 -5659
rect -489 -5663 -470 -5659
rect -173 -5663 -150 -5659
rect -131 -5663 -112 -5659
rect 255 -5663 278 -5659
rect 297 -5663 316 -5659
rect 611 -5663 634 -5659
rect 653 -5663 672 -5659
rect 1633 -5674 1695 -5561
rect -1421 -5678 -1255 -5674
rect -1251 -5678 -1238 -5674
rect -1234 -5678 -1197 -5674
rect -1193 -5678 -1155 -5674
rect -1151 -5678 -1113 -5674
rect -1109 -5678 -1072 -5674
rect -1068 -5678 -926 -5674
rect -922 -5678 -909 -5674
rect -905 -5678 -868 -5674
rect -864 -5678 -826 -5674
rect -822 -5678 -784 -5674
rect -780 -5678 -743 -5674
rect -739 -5678 -568 -5674
rect -564 -5678 -551 -5674
rect -547 -5678 -510 -5674
rect -506 -5678 -468 -5674
rect -464 -5678 -426 -5674
rect -422 -5678 -385 -5674
rect -381 -5678 -210 -5674
rect -206 -5678 -193 -5674
rect -189 -5678 -152 -5674
rect -148 -5678 -110 -5674
rect -106 -5678 -68 -5674
rect -64 -5678 -27 -5674
rect -23 -5678 218 -5674
rect 222 -5678 235 -5674
rect 239 -5678 276 -5674
rect 280 -5678 318 -5674
rect 322 -5678 360 -5674
rect 364 -5678 401 -5674
rect 405 -5678 574 -5674
rect 578 -5678 591 -5674
rect 595 -5678 632 -5674
rect 636 -5678 674 -5674
rect 678 -5678 716 -5674
rect 720 -5678 757 -5674
rect 761 -5678 1695 -5674
rect -1495 -5703 -1339 -5699
rect -1335 -5703 -1322 -5699
rect -1318 -5703 -935 -5699
rect -931 -5703 -918 -5699
rect -914 -5703 -577 -5699
rect -573 -5703 -560 -5699
rect -556 -5703 -219 -5699
rect -215 -5703 -202 -5699
rect -198 -5703 209 -5699
rect 213 -5703 226 -5699
rect 230 -5703 565 -5699
rect 569 -5703 582 -5699
rect 586 -5703 963 -5699
rect 967 -5703 980 -5699
rect 984 -5703 1321 -5699
rect 1325 -5703 1338 -5699
rect 1342 -5703 1617 -5699
rect -1495 -5818 -1433 -5703
rect -1334 -5735 -1066 -5731
rect -930 -5735 -737 -5731
rect -572 -5735 -379 -5731
rect -214 -5735 -21 -5731
rect 214 -5735 407 -5731
rect 570 -5735 769 -5731
rect 968 -5735 1161 -5731
rect 1326 -5735 1519 -5731
rect -1323 -5743 -923 -5739
rect -919 -5743 -565 -5739
rect -561 -5743 -207 -5739
rect -203 -5743 221 -5739
rect 225 -5743 577 -5739
rect 581 -5743 763 -5739
rect 767 -5743 975 -5739
rect 979 -5743 1333 -5739
rect 1337 -5743 1617 -5739
rect -949 -5756 -909 -5752
rect -591 -5756 -551 -5752
rect -233 -5756 -193 -5752
rect 195 -5756 235 -5752
rect 551 -5756 591 -5752
rect 949 -5756 989 -5752
rect 1307 -5756 1347 -5752
rect 1633 -5791 1695 -5678
rect -1421 -5795 -1322 -5791
rect -1318 -5795 -918 -5791
rect -914 -5795 -560 -5791
rect -556 -5795 -202 -5791
rect -198 -5795 226 -5791
rect 230 -5795 582 -5791
rect 586 -5795 980 -5791
rect 984 -5795 1338 -5791
rect 1342 -5795 1695 -5791
rect -1495 -5822 -1255 -5818
rect -1251 -5822 -1238 -5818
rect -1234 -5822 -1198 -5818
rect -1194 -5822 -1177 -5818
rect -1173 -5822 -926 -5818
rect -922 -5822 -900 -5818
rect -896 -5822 -883 -5818
rect -879 -5822 -843 -5818
rect -839 -5822 -822 -5818
rect -818 -5822 -805 -5818
rect -801 -5822 -765 -5818
rect -761 -5822 -741 -5818
rect -737 -5822 -704 -5818
rect -700 -5822 -568 -5818
rect -564 -5822 -542 -5818
rect -538 -5822 -525 -5818
rect -521 -5822 -485 -5818
rect -481 -5822 -464 -5818
rect -460 -5822 -447 -5818
rect -443 -5822 -407 -5818
rect -403 -5822 -383 -5818
rect -379 -5822 -346 -5818
rect -342 -5822 -210 -5818
rect -206 -5822 -184 -5818
rect -180 -5822 -167 -5818
rect -163 -5822 -127 -5818
rect -123 -5822 -106 -5818
rect -102 -5822 -89 -5818
rect -85 -5822 -49 -5818
rect -45 -5822 -25 -5818
rect -21 -5822 12 -5818
rect 16 -5822 218 -5818
rect 222 -5822 244 -5818
rect 248 -5822 261 -5818
rect 265 -5822 301 -5818
rect 305 -5822 322 -5818
rect 326 -5822 339 -5818
rect 343 -5822 379 -5818
rect 383 -5822 403 -5818
rect 407 -5822 440 -5818
rect 444 -5822 574 -5818
rect 578 -5822 600 -5818
rect 604 -5822 617 -5818
rect 621 -5822 657 -5818
rect 661 -5822 678 -5818
rect 682 -5822 695 -5818
rect 699 -5822 735 -5818
rect 739 -5822 759 -5818
rect 763 -5822 796 -5818
rect 800 -5822 972 -5818
rect 976 -5822 998 -5818
rect 1002 -5822 1015 -5818
rect 1019 -5822 1055 -5818
rect 1059 -5822 1076 -5818
rect 1080 -5822 1093 -5818
rect 1097 -5822 1133 -5818
rect 1137 -5822 1157 -5818
rect 1161 -5822 1194 -5818
rect 1198 -5822 1330 -5818
rect 1334 -5822 1356 -5818
rect 1360 -5822 1373 -5818
rect 1377 -5822 1413 -5818
rect 1417 -5822 1434 -5818
rect 1438 -5822 1451 -5818
rect 1455 -5822 1491 -5818
rect 1495 -5822 1515 -5818
rect 1519 -5822 1552 -5818
rect 1556 -5822 1617 -5818
rect -1495 -5941 -1433 -5822
rect -926 -5826 -922 -5822
rect -900 -5826 -896 -5822
rect -883 -5826 -879 -5822
rect -843 -5826 -839 -5822
rect -822 -5826 -818 -5822
rect -805 -5826 -801 -5822
rect -765 -5826 -761 -5822
rect -741 -5826 -737 -5822
rect -704 -5826 -700 -5822
rect -568 -5826 -564 -5822
rect -542 -5826 -538 -5822
rect -525 -5826 -521 -5822
rect -485 -5826 -481 -5822
rect -464 -5826 -460 -5822
rect -447 -5826 -443 -5822
rect -407 -5826 -403 -5822
rect -383 -5826 -379 -5822
rect -346 -5826 -342 -5822
rect -210 -5826 -206 -5822
rect -184 -5826 -180 -5822
rect -167 -5826 -163 -5822
rect -127 -5826 -123 -5822
rect -106 -5826 -102 -5822
rect -89 -5826 -85 -5822
rect -49 -5826 -45 -5822
rect -25 -5826 -21 -5822
rect 12 -5826 16 -5822
rect 218 -5826 222 -5822
rect 244 -5826 248 -5822
rect 261 -5826 265 -5822
rect 301 -5826 305 -5822
rect 322 -5826 326 -5822
rect 339 -5826 343 -5822
rect 379 -5826 383 -5822
rect 403 -5826 407 -5822
rect 440 -5826 444 -5822
rect 574 -5826 578 -5822
rect 600 -5826 604 -5822
rect 617 -5826 621 -5822
rect 657 -5826 661 -5822
rect 678 -5826 682 -5822
rect 695 -5826 699 -5822
rect 735 -5826 739 -5822
rect 759 -5826 763 -5822
rect 796 -5826 800 -5822
rect 972 -5826 976 -5822
rect 998 -5826 1002 -5822
rect 1015 -5826 1019 -5822
rect 1055 -5826 1059 -5822
rect 1076 -5826 1080 -5822
rect 1093 -5826 1097 -5822
rect 1133 -5826 1137 -5822
rect 1157 -5826 1161 -5822
rect 1194 -5826 1198 -5822
rect 1330 -5826 1334 -5822
rect 1356 -5826 1360 -5822
rect 1373 -5826 1377 -5822
rect 1413 -5826 1417 -5822
rect 1434 -5826 1438 -5822
rect 1451 -5826 1455 -5822
rect 1491 -5826 1495 -5822
rect 1515 -5826 1519 -5822
rect 1552 -5826 1556 -5822
rect -920 -5841 -858 -5837
rect -854 -5841 -824 -5837
rect -776 -5841 -746 -5837
rect -562 -5841 -500 -5837
rect -496 -5841 -466 -5837
rect -418 -5841 -388 -5837
rect -204 -5841 -142 -5837
rect -138 -5841 -108 -5837
rect -60 -5841 -30 -5837
rect 224 -5841 286 -5837
rect 290 -5841 320 -5837
rect 368 -5841 398 -5837
rect 580 -5841 642 -5837
rect 646 -5841 676 -5837
rect 724 -5841 754 -5837
rect 978 -5841 1040 -5837
rect 1044 -5841 1074 -5837
rect 1122 -5841 1152 -5837
rect 1336 -5841 1398 -5837
rect 1402 -5841 1432 -5837
rect 1480 -5841 1510 -5837
rect -913 -5848 -882 -5844
rect -555 -5848 -524 -5844
rect -197 -5848 -166 -5844
rect 231 -5848 262 -5844
rect 587 -5848 618 -5844
rect 985 -5848 1016 -5844
rect 1343 -5848 1374 -5844
rect -931 -5855 -848 -5851
rect -809 -5855 -706 -5851
rect -573 -5855 -490 -5851
rect -451 -5855 -348 -5851
rect -215 -5855 -132 -5851
rect -93 -5855 10 -5851
rect 213 -5855 296 -5851
rect 335 -5855 438 -5851
rect 569 -5855 652 -5851
rect 691 -5855 794 -5851
rect 967 -5855 1050 -5851
rect 1089 -5855 1192 -5851
rect 1325 -5855 1408 -5851
rect 1447 -5855 1550 -5851
rect -949 -5862 -928 -5858
rect -894 -5862 -865 -5858
rect -861 -5862 -780 -5858
rect -691 -5862 -592 -5858
rect -585 -5862 -570 -5858
rect -536 -5862 -507 -5858
rect -503 -5862 -422 -5858
rect -333 -5861 -234 -5857
rect -596 -5866 -592 -5862
rect -238 -5866 -234 -5861
rect -227 -5862 -212 -5858
rect -178 -5862 -149 -5858
rect -145 -5862 -64 -5858
rect 25 -5862 194 -5858
rect 201 -5862 216 -5858
rect 250 -5862 279 -5858
rect 283 -5862 364 -5858
rect 453 -5862 550 -5858
rect 557 -5862 572 -5858
rect 606 -5862 635 -5858
rect 639 -5862 720 -5858
rect 809 -5862 948 -5858
rect 955 -5862 970 -5858
rect 1004 -5862 1033 -5858
rect 1037 -5862 1118 -5858
rect 1207 -5860 1300 -5856
rect 190 -5866 194 -5862
rect 546 -5866 550 -5862
rect 944 -5866 948 -5862
rect 1296 -5866 1300 -5860
rect 1307 -5862 1328 -5858
rect 1362 -5862 1391 -5858
rect 1395 -5862 1476 -5858
rect -1260 -5871 -1203 -5867
rect -1164 -5870 -902 -5866
rect -887 -5870 -804 -5866
rect -783 -5870 -689 -5866
rect -596 -5870 -544 -5866
rect -529 -5870 -446 -5866
rect -425 -5870 -331 -5866
rect -238 -5870 -186 -5866
rect -171 -5870 -88 -5866
rect -67 -5870 27 -5866
rect 190 -5870 242 -5866
rect 257 -5870 340 -5866
rect 361 -5870 455 -5866
rect 546 -5870 598 -5866
rect 613 -5870 696 -5866
rect 717 -5870 811 -5866
rect 944 -5870 996 -5866
rect 1011 -5870 1094 -5866
rect 1115 -5870 1209 -5866
rect 1296 -5870 1354 -5866
rect 1369 -5870 1452 -5866
rect 1473 -5870 1567 -5866
rect -1266 -5878 -1253 -5874
rect -1249 -5878 -1213 -5874
rect -1209 -5878 -1193 -5874
rect -943 -5877 -924 -5873
rect -905 -5877 -776 -5873
rect -591 -5877 -566 -5873
rect -547 -5877 -418 -5873
rect -233 -5877 -208 -5873
rect -189 -5877 -60 -5873
rect 195 -5877 220 -5873
rect 239 -5877 368 -5873
rect 551 -5877 576 -5873
rect 595 -5877 724 -5873
rect 949 -5877 974 -5873
rect 993 -5877 1122 -5873
rect 1313 -5877 1332 -5873
rect 1351 -5877 1480 -5873
rect -1309 -5885 -1257 -5881
rect -1253 -5885 -1227 -5881
rect -1223 -5885 -1179 -5881
rect -898 -5884 -794 -5880
rect -790 -5884 -760 -5880
rect -540 -5884 -436 -5880
rect -432 -5884 -402 -5880
rect -182 -5884 -78 -5880
rect -74 -5884 -44 -5880
rect 246 -5884 350 -5880
rect 354 -5884 384 -5880
rect 602 -5884 706 -5880
rect 710 -5884 740 -5880
rect 1000 -5884 1104 -5880
rect 1108 -5884 1138 -5880
rect 1358 -5884 1462 -5880
rect 1466 -5884 1496 -5880
rect -1216 -5892 -1162 -5888
rect -924 -5891 -872 -5887
rect -868 -5891 -838 -5887
rect -566 -5891 -514 -5887
rect -510 -5891 -480 -5887
rect -208 -5891 -156 -5887
rect -152 -5891 -122 -5887
rect 220 -5891 272 -5887
rect 276 -5891 306 -5887
rect 576 -5891 628 -5887
rect 632 -5891 662 -5887
rect 974 -5891 1026 -5887
rect 1030 -5891 1060 -5887
rect 1332 -5891 1384 -5887
rect 1388 -5891 1418 -5887
rect -1234 -5899 -1202 -5895
rect -879 -5899 -847 -5895
rect -883 -5902 -879 -5899
rect -847 -5902 -843 -5899
rect -801 -5899 -769 -5895
rect -805 -5902 -801 -5899
rect -769 -5902 -765 -5899
rect -521 -5899 -489 -5895
rect -525 -5902 -521 -5899
rect -489 -5902 -485 -5899
rect -443 -5899 -411 -5895
rect -447 -5902 -443 -5899
rect -411 -5902 -407 -5899
rect -163 -5899 -131 -5895
rect -167 -5902 -163 -5899
rect -131 -5902 -127 -5899
rect -85 -5899 -53 -5895
rect -89 -5902 -85 -5899
rect -53 -5902 -49 -5899
rect 265 -5899 297 -5895
rect 261 -5902 265 -5899
rect 297 -5902 301 -5899
rect 343 -5899 375 -5895
rect 339 -5902 343 -5899
rect 375 -5902 379 -5899
rect 621 -5899 653 -5895
rect 617 -5902 621 -5899
rect 653 -5902 657 -5899
rect 699 -5899 731 -5895
rect 695 -5902 699 -5899
rect 731 -5902 735 -5899
rect 1019 -5899 1051 -5895
rect 1015 -5902 1019 -5899
rect 1051 -5902 1055 -5899
rect 1097 -5899 1129 -5895
rect 1093 -5902 1097 -5899
rect 1129 -5902 1133 -5899
rect 1377 -5899 1409 -5895
rect 1373 -5902 1377 -5899
rect 1409 -5902 1413 -5899
rect 1455 -5899 1487 -5895
rect 1451 -5902 1455 -5899
rect 1487 -5902 1491 -5899
rect -926 -5910 -922 -5906
rect -900 -5910 -896 -5906
rect -857 -5910 -853 -5906
rect -822 -5910 -818 -5906
rect -778 -5910 -774 -5906
rect -761 -5910 -757 -5906
rect -725 -5910 -721 -5906
rect -704 -5910 -700 -5906
rect -568 -5910 -564 -5906
rect -542 -5910 -538 -5906
rect -499 -5910 -495 -5906
rect -464 -5910 -460 -5906
rect -420 -5910 -416 -5906
rect -403 -5910 -399 -5906
rect -367 -5910 -363 -5906
rect -346 -5910 -342 -5906
rect -210 -5910 -206 -5906
rect -184 -5910 -180 -5906
rect -141 -5910 -137 -5906
rect -106 -5910 -102 -5906
rect -62 -5910 -58 -5906
rect -45 -5910 -41 -5906
rect -9 -5910 -5 -5906
rect 12 -5910 16 -5906
rect 218 -5910 222 -5906
rect 244 -5910 248 -5906
rect 287 -5910 291 -5906
rect 322 -5910 326 -5906
rect 366 -5910 370 -5906
rect 383 -5910 387 -5906
rect 419 -5910 423 -5906
rect 440 -5910 444 -5906
rect 574 -5910 578 -5906
rect 600 -5910 604 -5906
rect 643 -5910 647 -5906
rect 678 -5910 682 -5906
rect 722 -5910 726 -5906
rect 739 -5910 743 -5906
rect 775 -5910 779 -5906
rect 796 -5910 800 -5906
rect 972 -5910 976 -5906
rect 998 -5910 1002 -5906
rect 1041 -5910 1045 -5906
rect 1076 -5910 1080 -5906
rect 1120 -5910 1124 -5906
rect 1137 -5910 1141 -5906
rect 1173 -5910 1177 -5906
rect 1194 -5910 1198 -5906
rect 1330 -5910 1334 -5906
rect 1356 -5910 1360 -5906
rect 1399 -5910 1403 -5906
rect 1434 -5910 1438 -5906
rect 1478 -5910 1482 -5906
rect 1495 -5910 1499 -5906
rect 1531 -5910 1535 -5906
rect 1552 -5910 1556 -5906
rect 1633 -5910 1695 -5795
rect -1421 -5914 -1255 -5910
rect -1251 -5914 -1211 -5910
rect -1207 -5914 -1177 -5910
rect -1173 -5914 -926 -5910
rect -922 -5914 -900 -5910
rect -896 -5914 -857 -5910
rect -853 -5914 -822 -5910
rect -818 -5914 -778 -5910
rect -774 -5914 -761 -5910
rect -757 -5914 -725 -5910
rect -721 -5914 -704 -5910
rect -700 -5914 -568 -5910
rect -564 -5914 -542 -5910
rect -538 -5914 -499 -5910
rect -495 -5914 -464 -5910
rect -460 -5914 -420 -5910
rect -416 -5914 -403 -5910
rect -399 -5914 -367 -5910
rect -363 -5914 -346 -5910
rect -342 -5914 -210 -5910
rect -206 -5914 -184 -5910
rect -180 -5914 -141 -5910
rect -137 -5914 -106 -5910
rect -102 -5914 -62 -5910
rect -58 -5914 -45 -5910
rect -41 -5914 -9 -5910
rect -5 -5914 12 -5910
rect 16 -5914 218 -5910
rect 222 -5914 244 -5910
rect 248 -5914 287 -5910
rect 291 -5914 322 -5910
rect 326 -5914 366 -5910
rect 370 -5914 383 -5910
rect 387 -5914 419 -5910
rect 423 -5914 440 -5910
rect 444 -5914 574 -5910
rect 578 -5914 600 -5910
rect 604 -5914 643 -5910
rect 647 -5914 678 -5910
rect 682 -5914 722 -5910
rect 726 -5914 739 -5910
rect 743 -5914 775 -5910
rect 779 -5914 796 -5910
rect 800 -5914 972 -5910
rect 976 -5914 998 -5910
rect 1002 -5914 1041 -5910
rect 1045 -5914 1076 -5910
rect 1080 -5914 1120 -5910
rect 1124 -5914 1137 -5910
rect 1141 -5914 1173 -5910
rect 1177 -5914 1194 -5910
rect 1198 -5914 1330 -5910
rect 1334 -5914 1356 -5910
rect 1360 -5914 1399 -5910
rect 1403 -5914 1434 -5910
rect 1438 -5914 1478 -5910
rect 1482 -5914 1495 -5910
rect 1499 -5914 1531 -5910
rect 1535 -5914 1552 -5910
rect 1556 -5914 1695 -5910
rect -1266 -5924 -1162 -5920
rect -937 -5921 -689 -5917
rect -579 -5921 -331 -5917
rect -221 -5921 27 -5917
rect 207 -5922 455 -5918
rect 563 -5921 811 -5917
rect 961 -5921 1209 -5917
rect 1319 -5921 1567 -5917
rect -1495 -5945 -1255 -5941
rect -1251 -5945 -1238 -5941
rect -1234 -5945 -1218 -5941
rect -1214 -5945 -1197 -5941
rect -1193 -5945 -1176 -5941
rect -1172 -5945 -1155 -5941
rect -1151 -5945 -1134 -5941
rect -1130 -5945 -1113 -5941
rect -1109 -5945 -1092 -5941
rect -1088 -5945 -1072 -5941
rect -1068 -5945 -926 -5941
rect -922 -5945 -909 -5941
rect -905 -5945 -889 -5941
rect -885 -5945 -868 -5941
rect -864 -5945 -847 -5941
rect -843 -5945 -826 -5941
rect -822 -5945 -805 -5941
rect -801 -5945 -784 -5941
rect -780 -5945 -763 -5941
rect -759 -5945 -743 -5941
rect -739 -5945 -568 -5941
rect -564 -5945 -551 -5941
rect -547 -5945 -531 -5941
rect -527 -5945 -510 -5941
rect -506 -5945 -489 -5941
rect -485 -5945 -468 -5941
rect -464 -5945 -447 -5941
rect -443 -5945 -426 -5941
rect -422 -5945 -405 -5941
rect -401 -5945 -385 -5941
rect -381 -5945 -210 -5941
rect -206 -5945 -193 -5941
rect -189 -5945 -173 -5941
rect -169 -5945 -152 -5941
rect -148 -5945 -131 -5941
rect -127 -5945 -110 -5941
rect -106 -5945 -89 -5941
rect -85 -5945 -68 -5941
rect -64 -5945 -47 -5941
rect -43 -5945 -27 -5941
rect -23 -5945 218 -5941
rect 222 -5945 235 -5941
rect 239 -5945 255 -5941
rect 259 -5945 276 -5941
rect 280 -5945 297 -5941
rect 301 -5945 318 -5941
rect 322 -5945 339 -5941
rect 343 -5945 360 -5941
rect 364 -5945 381 -5941
rect 385 -5945 401 -5941
rect 405 -5945 574 -5941
rect 578 -5945 591 -5941
rect 595 -5945 611 -5941
rect 615 -5945 632 -5941
rect 636 -5945 653 -5941
rect 657 -5945 674 -5941
rect 678 -5945 695 -5941
rect 699 -5945 716 -5941
rect 720 -5945 737 -5941
rect 741 -5945 757 -5941
rect 761 -5945 972 -5941
rect 976 -5945 989 -5941
rect 993 -5945 1009 -5941
rect 1013 -5945 1030 -5941
rect 1034 -5945 1051 -5941
rect 1055 -5945 1072 -5941
rect 1076 -5945 1093 -5941
rect 1097 -5945 1114 -5941
rect 1118 -5945 1135 -5941
rect 1139 -5945 1155 -5941
rect 1159 -5945 1330 -5941
rect 1334 -5945 1347 -5941
rect 1351 -5945 1367 -5941
rect 1371 -5945 1388 -5941
rect 1392 -5945 1409 -5941
rect 1413 -5945 1430 -5941
rect 1434 -5945 1451 -5941
rect 1455 -5945 1472 -5941
rect 1476 -5945 1493 -5941
rect 1497 -5945 1513 -5941
rect 1517 -5945 1617 -5941
rect -1495 -6059 -1433 -5945
rect -1233 -5993 -1199 -5989
rect -1135 -5993 -1115 -5989
rect -1100 -5993 -1064 -5989
rect -904 -5993 -870 -5989
rect -806 -5993 -786 -5989
rect -771 -5993 -735 -5989
rect -546 -5993 -512 -5989
rect -448 -5993 -428 -5989
rect -413 -5993 -377 -5989
rect -188 -5993 -154 -5989
rect -90 -5993 -70 -5989
rect -55 -5993 -19 -5989
rect 240 -5993 274 -5989
rect 338 -5993 358 -5989
rect 373 -5993 409 -5989
rect 596 -5993 630 -5989
rect 694 -5993 714 -5989
rect 729 -5993 765 -5989
rect 994 -5993 1028 -5989
rect 1092 -5993 1112 -5989
rect 1127 -5993 1163 -5989
rect 1352 -5993 1386 -5989
rect 1450 -5993 1470 -5989
rect 1485 -5993 1521 -5989
rect -1266 -6001 -1257 -5997
rect -1253 -6001 -1223 -5997
rect -1202 -6001 -1171 -5997
rect -1142 -6001 -1111 -5997
rect -1100 -6001 -1073 -5997
rect -937 -6001 -928 -5997
rect -924 -6001 -894 -5997
rect -873 -6001 -842 -5997
rect -813 -6001 -782 -5997
rect -771 -6001 -744 -5997
rect -579 -6001 -570 -5997
rect -566 -6001 -536 -5997
rect -515 -6001 -484 -5997
rect -455 -6001 -424 -5997
rect -413 -6001 -386 -5997
rect -221 -6001 -212 -5997
rect -208 -6001 -178 -5997
rect -157 -6001 -126 -5997
rect -97 -6001 -66 -5997
rect -55 -6001 -28 -5997
rect 207 -6001 216 -5997
rect 220 -6001 250 -5997
rect 271 -6001 302 -5997
rect 331 -6001 362 -5997
rect 373 -6001 400 -5997
rect 563 -6001 572 -5997
rect 576 -6001 606 -5997
rect 627 -6001 658 -5997
rect 687 -6001 718 -5997
rect 729 -6001 756 -5997
rect 961 -6001 970 -5997
rect 974 -6001 1004 -5997
rect 1025 -6001 1056 -5997
rect 1085 -6001 1116 -5997
rect 1127 -6001 1154 -5997
rect 1319 -6001 1328 -5997
rect 1332 -6001 1362 -5997
rect 1383 -6001 1414 -5997
rect 1443 -6001 1474 -5997
rect 1485 -6001 1512 -5997
rect -1260 -6008 -1213 -6004
rect -1177 -6008 -1164 -6004
rect -1160 -6008 -1129 -6004
rect -1093 -6008 -1080 -6004
rect -1076 -6008 -1064 -6004
rect -931 -6008 -884 -6004
rect -848 -6008 -835 -6004
rect -831 -6008 -800 -6004
rect -764 -6008 -751 -6004
rect -747 -6008 -735 -6004
rect -573 -6008 -526 -6004
rect -490 -6008 -477 -6004
rect -473 -6008 -442 -6004
rect -406 -6008 -393 -6004
rect -389 -6008 -377 -6004
rect -215 -6008 -168 -6004
rect -132 -6008 -119 -6004
rect -115 -6008 -84 -6004
rect -48 -6008 -35 -6004
rect -31 -6008 -19 -6004
rect 213 -6008 260 -6004
rect 296 -6008 309 -6004
rect 313 -6008 344 -6004
rect 380 -6008 393 -6004
rect 397 -6008 409 -6004
rect 569 -6008 616 -6004
rect 652 -6008 665 -6004
rect 669 -6008 700 -6004
rect 736 -6008 749 -6004
rect 753 -6008 765 -6004
rect 967 -6008 1014 -6004
rect 1050 -6008 1063 -6004
rect 1067 -6008 1098 -6004
rect 1134 -6008 1147 -6004
rect 1151 -6008 1163 -6004
rect 1325 -6008 1372 -6004
rect 1408 -6008 1421 -6004
rect 1425 -6008 1456 -6004
rect 1492 -6008 1505 -6004
rect 1509 -6008 1521 -6004
rect -1267 -6015 -1253 -6011
rect -1249 -6015 -1139 -6011
rect -1118 -6015 -1087 -6011
rect -936 -6015 -924 -6011
rect -920 -6015 -810 -6011
rect -789 -6015 -758 -6011
rect -580 -6015 -566 -6011
rect -562 -6015 -452 -6011
rect -431 -6015 -400 -6011
rect -223 -6015 -208 -6011
rect -204 -6015 -94 -6011
rect -73 -6015 -42 -6011
rect 205 -6015 220 -6011
rect 224 -6015 334 -6011
rect 355 -6015 386 -6011
rect 563 -6015 576 -6011
rect 580 -6015 690 -6011
rect 711 -6015 742 -6011
rect 961 -6015 974 -6011
rect 978 -6015 1088 -6011
rect 1109 -6015 1140 -6011
rect 1318 -6015 1332 -6011
rect 1336 -6015 1446 -6011
rect 1467 -6015 1498 -6011
rect -1218 -6022 -1195 -6018
rect -1176 -6022 -1157 -6018
rect -889 -6022 -866 -6018
rect -847 -6022 -828 -6018
rect -531 -6022 -508 -6018
rect -489 -6022 -470 -6018
rect -173 -6022 -150 -6018
rect -131 -6022 -112 -6018
rect 255 -6022 278 -6018
rect 297 -6022 316 -6018
rect 611 -6022 634 -6018
rect 653 -6022 672 -6018
rect 1009 -6022 1032 -6018
rect 1051 -6022 1070 -6018
rect 1367 -6022 1390 -6018
rect 1409 -6022 1428 -6018
rect 1633 -6033 1695 -5914
rect -1421 -6037 -1255 -6033
rect -1251 -6037 -1238 -6033
rect -1234 -6037 -1197 -6033
rect -1193 -6037 -1155 -6033
rect -1151 -6037 -1113 -6033
rect -1109 -6037 -1072 -6033
rect -1068 -6037 -926 -6033
rect -922 -6037 -909 -6033
rect -905 -6037 -868 -6033
rect -864 -6037 -826 -6033
rect -822 -6037 -784 -6033
rect -780 -6037 -743 -6033
rect -739 -6037 -568 -6033
rect -564 -6037 -551 -6033
rect -547 -6037 -510 -6033
rect -506 -6037 -468 -6033
rect -464 -6037 -426 -6033
rect -422 -6037 -385 -6033
rect -381 -6037 -210 -6033
rect -206 -6037 -193 -6033
rect -189 -6037 -152 -6033
rect -148 -6037 -110 -6033
rect -106 -6037 -68 -6033
rect -64 -6037 -27 -6033
rect -23 -6037 218 -6033
rect 222 -6037 235 -6033
rect 239 -6037 276 -6033
rect 280 -6037 318 -6033
rect 322 -6037 360 -6033
rect 364 -6037 401 -6033
rect 405 -6037 574 -6033
rect 578 -6037 591 -6033
rect 595 -6037 632 -6033
rect 636 -6037 674 -6033
rect 678 -6037 716 -6033
rect 720 -6037 757 -6033
rect 761 -6037 972 -6033
rect 976 -6037 989 -6033
rect 993 -6037 1030 -6033
rect 1034 -6037 1072 -6033
rect 1076 -6037 1114 -6033
rect 1118 -6037 1155 -6033
rect 1159 -6037 1330 -6033
rect 1334 -6037 1347 -6033
rect 1351 -6037 1388 -6033
rect 1392 -6037 1430 -6033
rect 1434 -6037 1472 -6033
rect 1476 -6037 1513 -6033
rect 1517 -6037 1695 -6033
rect 1319 -6044 1561 -6040
rect -1495 -6063 1330 -6059
rect 1334 -6063 1347 -6059
rect 1351 -6063 1367 -6059
rect 1371 -6063 1388 -6059
rect 1392 -6063 1409 -6059
rect 1413 -6063 1430 -6059
rect 1434 -6063 1451 -6059
rect 1455 -6063 1472 -6059
rect 1476 -6063 1493 -6059
rect 1497 -6063 1513 -6059
rect 1517 -6063 1617 -6059
rect -1495 -6155 -1433 -6063
rect 1352 -6111 1386 -6107
rect 1450 -6111 1470 -6107
rect 1485 -6111 1521 -6107
rect 1319 -6119 1328 -6115
rect 1332 -6119 1362 -6115
rect 1383 -6119 1414 -6115
rect 1443 -6119 1474 -6115
rect 1485 -6119 1512 -6115
rect 1325 -6126 1372 -6122
rect 1408 -6126 1421 -6122
rect 1425 -6126 1456 -6122
rect 1492 -6126 1505 -6122
rect 1509 -6126 1521 -6122
rect 1320 -6133 1332 -6129
rect 1336 -6133 1446 -6129
rect 1467 -6133 1498 -6129
rect 1367 -6140 1390 -6136
rect 1409 -6140 1428 -6136
rect 1633 -6151 1695 -6037
rect -1421 -6155 1330 -6151
rect 1334 -6155 1347 -6151
rect 1351 -6155 1388 -6151
rect 1392 -6155 1430 -6151
rect 1434 -6155 1472 -6151
rect 1476 -6155 1513 -6151
rect 1517 -6155 1695 -6151
<< metal3 >>
rect -1009 -1167 -989 -1161
rect -1275 -1214 -1269 -1213
rect -1275 -1218 -1274 -1214
rect -1270 -1218 -1269 -1214
rect -1275 -1257 -1269 -1218
rect -1009 -1241 -1003 -1167
rect -995 -1234 -989 -1167
rect -981 -1167 -962 -1161
rect -981 -1234 -975 -1167
rect -995 -1240 -975 -1234
rect -968 -1234 -962 -1167
rect -295 -1166 -273 -1160
rect -957 -1214 -951 -1212
rect -957 -1218 -956 -1214
rect -952 -1218 -951 -1214
rect -957 -1234 -951 -1218
rect -968 -1240 -951 -1234
rect -588 -1214 -582 -1213
rect -588 -1218 -587 -1214
rect -583 -1218 -582 -1214
rect -1254 -1247 -1230 -1241
rect -1254 -1257 -1248 -1247
rect -1275 -1263 -1248 -1257
rect -1236 -1257 -1230 -1247
rect -1221 -1247 -1003 -1241
rect -588 -1241 -582 -1218
rect -295 -1241 -289 -1166
rect -279 -1233 -273 -1166
rect -265 -1166 -246 -1160
rect -265 -1233 -259 -1166
rect -279 -1239 -259 -1233
rect -252 -1233 -246 -1166
rect 484 -1167 504 -1161
rect -241 -1214 -235 -1213
rect -241 -1218 -240 -1214
rect -236 -1218 -235 -1214
rect -241 -1233 -235 -1218
rect -252 -1239 -235 -1233
rect 197 -1214 203 -1213
rect 197 -1218 198 -1214
rect 202 -1218 203 -1214
rect -588 -1247 -530 -1241
rect -1221 -1257 -1215 -1247
rect -1236 -1263 -1215 -1257
rect -1056 -1563 -1036 -1557
rect -1271 -1567 -1260 -1566
rect -1271 -1571 -1265 -1567
rect -1261 -1571 -1260 -1567
rect -1271 -1572 -1260 -1571
rect -1271 -1644 -1265 -1572
rect -1056 -1644 -1050 -1563
rect -1271 -1650 -1050 -1644
rect -1271 -1688 -1265 -1650
rect -1271 -1692 -1270 -1688
rect -1266 -1692 -1265 -1688
rect -1271 -1809 -1265 -1692
rect -1042 -1708 -1036 -1563
rect -1030 -1563 -1013 -1557
rect -1030 -1708 -1024 -1563
rect -1019 -1670 -1013 -1563
rect -1009 -1670 -1003 -1247
rect -536 -1257 -530 -1247
rect -519 -1247 -495 -1241
rect -519 -1257 -513 -1247
rect -536 -1263 -513 -1257
rect -501 -1257 -495 -1247
rect -486 -1247 -289 -1241
rect 197 -1241 203 -1218
rect 484 -1241 490 -1167
rect 498 -1234 504 -1167
rect 512 -1167 531 -1161
rect 512 -1234 518 -1167
rect 498 -1240 518 -1234
rect 525 -1234 531 -1167
rect 535 -1214 542 -1213
rect 535 -1218 536 -1214
rect 540 -1218 542 -1214
rect 535 -1234 542 -1218
rect 525 -1240 542 -1234
rect 951 -1214 957 -1213
rect 951 -1218 952 -1214
rect 956 -1218 957 -1214
rect 197 -1247 254 -1241
rect -486 -1257 -480 -1247
rect -501 -1263 -480 -1257
rect -999 -1563 -982 -1557
rect -999 -1670 -993 -1563
rect -1019 -1676 -993 -1670
rect -1042 -1714 -1024 -1708
rect -1009 -1787 -1003 -1676
rect -988 -1709 -982 -1563
rect -977 -1563 -961 -1557
rect -977 -1709 -971 -1563
rect -988 -1715 -971 -1709
rect -967 -1709 -961 -1563
rect -346 -1563 -326 -1557
rect -947 -1567 -941 -1565
rect -947 -1571 -946 -1567
rect -942 -1571 -941 -1567
rect -947 -1687 -941 -1571
rect -589 -1567 -583 -1565
rect -589 -1571 -588 -1567
rect -584 -1571 -583 -1567
rect -589 -1644 -583 -1571
rect -346 -1644 -340 -1563
rect -589 -1650 -340 -1644
rect -957 -1688 -936 -1687
rect -957 -1692 -941 -1688
rect -937 -1692 -936 -1688
rect -957 -1693 -936 -1692
rect -589 -1688 -583 -1650
rect -589 -1692 -588 -1688
rect -584 -1692 -583 -1688
rect -957 -1709 -951 -1693
rect -967 -1715 -951 -1709
rect -1271 -1813 -1270 -1809
rect -1266 -1813 -1265 -1809
rect -1271 -1814 -1265 -1813
rect -1038 -1793 -1024 -1787
rect -1014 -1788 -1003 -1787
rect -1014 -1792 -1013 -1788
rect -1009 -1792 -1003 -1788
rect -1014 -1793 -1003 -1792
rect -1038 -1834 -1032 -1793
rect -947 -1809 -941 -1693
rect -947 -1813 -946 -1809
rect -942 -1813 -941 -1809
rect -947 -1815 -941 -1813
rect -589 -1809 -583 -1692
rect -332 -1708 -326 -1563
rect -320 -1563 -303 -1557
rect -320 -1708 -314 -1563
rect -309 -1670 -303 -1563
rect -295 -1670 -289 -1247
rect 248 -1257 254 -1247
rect 265 -1247 289 -1241
rect 265 -1257 271 -1247
rect 248 -1263 271 -1257
rect 283 -1257 289 -1247
rect 298 -1247 490 -1241
rect 951 -1241 957 -1218
rect 951 -1247 1011 -1241
rect 298 -1257 304 -1247
rect 283 -1263 304 -1257
rect -283 -1563 -266 -1557
rect -283 -1670 -277 -1563
rect -309 -1676 -277 -1670
rect -332 -1714 -314 -1708
rect -295 -1726 -289 -1676
rect -272 -1709 -266 -1563
rect -261 -1563 -245 -1557
rect -261 -1709 -255 -1563
rect -272 -1715 -255 -1709
rect -251 -1709 -245 -1563
rect 431 -1563 451 -1557
rect -231 -1567 -225 -1566
rect -231 -1571 -230 -1567
rect -226 -1571 -225 -1567
rect -231 -1687 -225 -1571
rect -241 -1688 -225 -1687
rect -241 -1692 -230 -1688
rect -226 -1692 -225 -1688
rect -241 -1693 -225 -1692
rect -241 -1709 -235 -1693
rect -251 -1715 -235 -1709
rect -315 -1732 -289 -1726
rect -315 -1787 -309 -1732
rect -589 -1813 -588 -1809
rect -584 -1813 -583 -1809
rect -589 -1814 -583 -1813
rect -341 -1793 -327 -1787
rect -317 -1788 -309 -1787
rect -317 -1792 -316 -1788
rect -312 -1792 -309 -1788
rect -317 -1793 -309 -1792
rect -341 -1815 -335 -1793
rect -231 -1809 -225 -1693
rect -231 -1813 -230 -1809
rect -226 -1813 -225 -1809
rect -231 -1814 -225 -1813
rect 198 -1567 204 -1565
rect 198 -1571 199 -1567
rect 203 -1571 204 -1567
rect 198 -1644 204 -1571
rect 431 -1644 437 -1563
rect 198 -1650 437 -1644
rect 198 -1688 204 -1650
rect 198 -1692 199 -1688
rect 203 -1692 204 -1688
rect 198 -1809 204 -1692
rect 445 -1708 451 -1563
rect 457 -1563 474 -1557
rect 457 -1708 463 -1563
rect 468 -1670 474 -1563
rect 484 -1670 490 -1247
rect 1005 -1257 1011 -1247
rect 1022 -1247 1046 -1241
rect 1022 -1257 1028 -1247
rect 1005 -1263 1028 -1257
rect 1040 -1257 1046 -1247
rect 1055 -1247 1244 -1241
rect 1055 -1257 1061 -1247
rect 1040 -1263 1061 -1257
rect 499 -1563 516 -1557
rect 499 -1670 505 -1563
rect 468 -1676 505 -1670
rect 445 -1714 463 -1708
rect 484 -1787 490 -1676
rect 510 -1709 516 -1563
rect 521 -1563 537 -1557
rect 521 -1709 527 -1563
rect 510 -1715 527 -1709
rect 531 -1709 537 -1563
rect 1183 -1563 1203 -1557
rect 552 -1567 558 -1566
rect 552 -1571 553 -1567
rect 557 -1571 558 -1567
rect 552 -1687 558 -1571
rect 950 -1567 956 -1565
rect 950 -1571 951 -1567
rect 955 -1571 956 -1567
rect 950 -1644 956 -1571
rect 1183 -1644 1189 -1563
rect 950 -1650 1189 -1644
rect 541 -1688 565 -1687
rect 541 -1692 560 -1688
rect 564 -1692 565 -1688
rect 541 -1693 565 -1692
rect 950 -1688 956 -1650
rect 950 -1692 951 -1688
rect 955 -1692 956 -1688
rect 541 -1709 547 -1693
rect 531 -1715 547 -1709
rect 198 -1813 199 -1809
rect 203 -1813 204 -1809
rect 198 -1815 204 -1813
rect 455 -1793 469 -1787
rect 479 -1788 490 -1787
rect 479 -1792 480 -1788
rect 484 -1792 490 -1788
rect 479 -1793 490 -1792
rect -700 -1824 -653 -1816
rect -1038 -1840 -1003 -1834
rect -700 -1840 -692 -1824
rect -1009 -1848 -692 -1840
rect -661 -1840 -653 -1824
rect -643 -1824 -596 -1816
rect -341 -1821 -287 -1815
rect -643 -1840 -635 -1824
rect -661 -1848 -635 -1840
rect -604 -1840 -596 -1824
rect -293 -1840 -287 -1821
rect 455 -1834 461 -1793
rect 552 -1809 558 -1693
rect 552 -1813 553 -1809
rect 557 -1813 558 -1809
rect 552 -1814 558 -1813
rect 950 -1809 956 -1692
rect 1197 -1708 1203 -1563
rect 1209 -1563 1226 -1557
rect 1209 -1708 1215 -1563
rect 1220 -1670 1226 -1563
rect 1238 -1670 1244 -1247
rect 1255 -1563 1272 -1557
rect 1255 -1670 1261 -1563
rect 1220 -1676 1261 -1670
rect 1197 -1714 1215 -1708
rect 1238 -1726 1244 -1676
rect 1266 -1709 1272 -1563
rect 1277 -1563 1293 -1557
rect 1277 -1709 1283 -1563
rect 1266 -1715 1283 -1709
rect 1287 -1709 1293 -1563
rect 1297 -1688 1316 -1687
rect 1297 -1692 1311 -1688
rect 1315 -1692 1316 -1688
rect 1297 -1693 1316 -1692
rect 1297 -1709 1303 -1693
rect 1287 -1715 1303 -1709
rect 1220 -1733 1244 -1726
rect 1220 -1787 1226 -1733
rect 950 -1813 951 -1809
rect 955 -1813 956 -1809
rect 950 -1815 956 -1813
rect 1194 -1793 1208 -1787
rect 1218 -1788 1226 -1787
rect 1218 -1792 1219 -1788
rect 1223 -1792 1226 -1788
rect 1218 -1793 1226 -1792
rect 1194 -1815 1200 -1793
rect 1308 -1809 1314 -1693
rect 1308 -1813 1309 -1809
rect 1313 -1813 1314 -1809
rect 1308 -1814 1314 -1813
rect 1194 -1821 1248 -1815
rect 828 -1834 861 -1826
rect 455 -1840 490 -1834
rect -604 -1848 -287 -1840
rect 484 -1842 490 -1840
rect 828 -1842 836 -1834
rect 484 -1848 836 -1842
rect -1038 -1854 -1003 -1848
rect -1038 -1902 -1032 -1854
rect -653 -1899 -643 -1848
rect -293 -1871 -287 -1848
rect -1038 -1908 -1024 -1902
rect -1014 -1903 -1003 -1902
rect -1014 -1907 -1013 -1903
rect -1009 -1907 -1003 -1903
rect -1014 -1908 -1003 -1907
rect -1274 -1924 -1268 -1923
rect -1274 -1928 -1273 -1924
rect -1269 -1928 -1268 -1924
rect -1274 -1962 -1268 -1928
rect -1274 -1968 -1242 -1962
rect -1248 -2007 -1242 -1968
rect -1233 -1968 -1212 -1962
rect -1233 -2007 -1227 -1968
rect -1248 -2013 -1227 -2007
rect -1218 -2007 -1212 -1968
rect -1203 -1968 -1181 -1962
rect -1203 -2007 -1197 -1968
rect -1218 -2013 -1197 -2007
rect -1187 -2007 -1181 -1968
rect -1172 -1968 -1150 -1962
rect -1172 -2007 -1166 -1968
rect -1187 -2013 -1166 -2007
rect -1156 -2007 -1150 -1968
rect -1140 -1967 -1119 -1961
rect -1140 -2007 -1134 -1967
rect -1156 -2013 -1134 -2007
rect -1125 -2007 -1119 -1967
rect -1110 -1967 -1089 -1961
rect -1110 -2007 -1104 -1967
rect -1125 -2013 -1104 -2007
rect -1095 -2007 -1089 -1967
rect -1009 -1981 -1003 -1908
rect -691 -1910 -668 -1900
rect -658 -1903 -643 -1899
rect -658 -1907 -657 -1903
rect -653 -1907 -643 -1903
rect -658 -1909 -643 -1907
rect -341 -1877 -287 -1871
rect 455 -1850 836 -1848
rect 853 -1842 861 -1834
rect 871 -1834 904 -1826
rect 871 -1842 879 -1834
rect 853 -1850 879 -1842
rect 896 -1842 904 -1834
rect 1242 -1842 1248 -1821
rect 896 -1850 1248 -1842
rect 455 -1854 490 -1850
rect -341 -1902 -335 -1877
rect 455 -1902 461 -1854
rect 861 -1899 871 -1850
rect 1242 -1871 1248 -1850
rect -341 -1908 -327 -1902
rect -317 -1903 -308 -1902
rect -317 -1907 -316 -1903
rect -312 -1907 -308 -1903
rect -317 -1908 -308 -1907
rect 455 -1908 469 -1902
rect 479 -1903 490 -1902
rect 479 -1907 480 -1903
rect 484 -1907 490 -1903
rect 479 -1908 490 -1907
rect -691 -1953 -681 -1910
rect -314 -1949 -308 -1908
rect -691 -1963 -655 -1953
rect -314 -1955 -287 -1949
rect -1080 -1987 -1003 -1981
rect -1080 -2007 -1074 -1987
rect -1095 -2013 -1074 -2007
rect -1285 -2299 -1279 -2297
rect -1285 -2303 -1284 -2299
rect -1280 -2303 -1279 -2299
rect -1285 -2353 -1279 -2303
rect -1259 -2332 -1227 -2326
rect -1259 -2353 -1253 -2332
rect -1285 -2359 -1253 -2353
rect -1233 -2353 -1227 -2332
rect -1209 -2332 -1175 -2326
rect -1209 -2353 -1203 -2332
rect -1233 -2359 -1203 -2353
rect -1181 -2353 -1175 -2332
rect -1152 -2332 -1121 -2326
rect -1152 -2353 -1146 -2332
rect -1181 -2359 -1146 -2353
rect -1127 -2353 -1121 -2332
rect -1099 -2332 -1068 -2326
rect -1099 -2353 -1093 -2332
rect -1127 -2359 -1093 -2353
rect -1074 -2353 -1068 -2332
rect -1049 -2332 -1015 -2326
rect -1049 -2353 -1043 -2332
rect -1074 -2359 -1043 -2353
rect -1021 -2353 -1015 -2332
rect -1009 -2353 -1003 -1987
rect -997 -2240 -980 -2234
rect -997 -2353 -991 -2240
rect -1021 -2359 -991 -2353
rect -1285 -2430 -1279 -2359
rect -986 -2386 -980 -2240
rect -975 -2240 -959 -2234
rect -975 -2386 -969 -2240
rect -986 -2392 -969 -2386
rect -965 -2386 -959 -2240
rect -955 -2299 -949 -2297
rect -955 -2303 -954 -2299
rect -950 -2303 -949 -2299
rect -955 -2386 -949 -2303
rect -965 -2392 -949 -2386
rect -1285 -2434 -1284 -2430
rect -1280 -2434 -1279 -2430
rect -1285 -2436 -1279 -2434
rect -955 -2430 -949 -2392
rect -955 -2434 -954 -2430
rect -950 -2434 -949 -2430
rect -955 -2435 -949 -2434
rect -665 -2470 -655 -1963
rect -596 -2299 -590 -2298
rect -596 -2303 -595 -2299
rect -591 -2303 -590 -2299
rect -596 -2353 -590 -2303
rect -570 -2332 -538 -2326
rect -570 -2353 -564 -2332
rect -596 -2359 -564 -2353
rect -544 -2353 -538 -2332
rect -520 -2332 -486 -2326
rect -520 -2353 -514 -2332
rect -544 -2359 -514 -2353
rect -492 -2353 -486 -2332
rect -463 -2332 -432 -2326
rect -463 -2353 -457 -2332
rect -492 -2359 -457 -2353
rect -438 -2353 -432 -2332
rect -410 -2332 -379 -2326
rect -410 -2353 -404 -2332
rect -438 -2359 -404 -2353
rect -385 -2353 -379 -2332
rect -360 -2332 -326 -2326
rect -360 -2353 -354 -2332
rect -385 -2359 -354 -2353
rect -332 -2353 -326 -2332
rect -293 -2353 -287 -1955
rect -282 -2240 -265 -2234
rect -282 -2353 -276 -2240
rect -332 -2359 -276 -2353
rect -596 -2430 -590 -2359
rect -271 -2386 -265 -2240
rect -260 -2240 -244 -2234
rect -260 -2386 -254 -2240
rect -271 -2392 -254 -2386
rect -250 -2386 -244 -2240
rect -240 -2299 -234 -2297
rect -240 -2303 -239 -2299
rect -235 -2303 -234 -2299
rect -240 -2386 -234 -2303
rect -250 -2392 -234 -2386
rect -596 -2434 -595 -2430
rect -591 -2434 -590 -2430
rect -596 -2436 -590 -2434
rect -240 -2430 -234 -2392
rect -240 -2434 -239 -2430
rect -235 -2434 -234 -2430
rect -240 -2435 -234 -2434
rect 191 -2299 197 -2298
rect 191 -2303 192 -2299
rect 196 -2303 197 -2299
rect 191 -2353 197 -2303
rect 215 -2332 247 -2326
rect 215 -2353 221 -2332
rect 191 -2359 221 -2353
rect 241 -2353 247 -2332
rect 265 -2332 299 -2326
rect 265 -2353 271 -2332
rect 241 -2359 271 -2353
rect 293 -2353 299 -2332
rect 322 -2332 353 -2326
rect 322 -2353 328 -2332
rect 293 -2359 328 -2353
rect 347 -2353 353 -2332
rect 375 -2332 406 -2326
rect 375 -2353 381 -2332
rect 347 -2359 381 -2353
rect 400 -2353 406 -2332
rect 425 -2332 459 -2326
rect 425 -2353 431 -2332
rect 400 -2359 431 -2353
rect 453 -2353 459 -2332
rect 484 -2353 490 -1908
rect 817 -1910 846 -1900
rect 856 -1903 871 -1899
rect 856 -1907 857 -1903
rect 861 -1907 871 -1903
rect 856 -1909 871 -1907
rect 1194 -1877 1248 -1871
rect 1194 -1902 1200 -1877
rect 1194 -1908 1208 -1902
rect 1218 -1903 1227 -1902
rect 1218 -1907 1219 -1903
rect 1223 -1907 1227 -1903
rect 1218 -1908 1227 -1907
rect 817 -1953 827 -1910
rect 1221 -1949 1227 -1908
rect 817 -1963 850 -1953
rect 1221 -1955 1248 -1949
rect 496 -2240 513 -2234
rect 496 -2353 502 -2240
rect 453 -2359 502 -2353
rect 191 -2430 197 -2359
rect 507 -2386 513 -2240
rect 518 -2240 534 -2234
rect 518 -2386 524 -2240
rect 507 -2392 524 -2386
rect 528 -2386 534 -2240
rect 542 -2299 548 -2298
rect 542 -2303 543 -2299
rect 547 -2303 548 -2299
rect 542 -2386 548 -2303
rect 528 -2392 548 -2386
rect 191 -2434 192 -2430
rect 196 -2434 197 -2430
rect 191 -2435 197 -2434
rect 542 -2430 548 -2392
rect 542 -2434 543 -2430
rect 547 -2434 548 -2430
rect 542 -2436 548 -2434
rect 78 -2470 106 -2457
rect 128 -2464 156 -2451
rect 128 -2470 140 -2464
rect -665 -2482 90 -2470
rect 94 -2482 140 -2470
rect -1059 -2552 -1036 -2546
rect -1276 -2561 -1270 -2560
rect -1276 -2565 -1275 -2561
rect -1271 -2565 -1270 -2561
rect -1276 -2593 -1270 -2565
rect -1059 -2593 -1053 -2552
rect -1276 -2599 -1053 -2593
rect -1276 -2673 -1270 -2599
rect -1042 -2611 -1036 -2552
rect -1024 -2552 -989 -2546
rect -1024 -2611 -1018 -2552
rect -1042 -2617 -1018 -2611
rect -1276 -2677 -1275 -2673
rect -1271 -2677 -1270 -2673
rect -1276 -2679 -1270 -2677
rect -1152 -2863 -1136 -2857
rect -1152 -2989 -1146 -2863
rect -1142 -2902 -1136 -2863
rect -1127 -2863 -1107 -2857
rect -1127 -2902 -1121 -2863
rect -1142 -2908 -1121 -2902
rect -1113 -2902 -1107 -2863
rect -1097 -2863 -1075 -2857
rect -1097 -2902 -1091 -2863
rect -1113 -2908 -1091 -2902
rect -1081 -2902 -1075 -2863
rect -1066 -2863 -1045 -2857
rect -1066 -2902 -1060 -2863
rect -1081 -2908 -1060 -2902
rect -1051 -2902 -1045 -2863
rect -1035 -2863 -1014 -2857
rect -1035 -2902 -1029 -2863
rect -1051 -2908 -1029 -2902
rect -1020 -2902 -1014 -2863
rect -1006 -2902 -1000 -2552
rect -995 -2636 -989 -2552
rect -985 -2552 -969 -2546
rect -985 -2636 -979 -2552
rect -995 -2642 -979 -2636
rect -975 -2636 -969 -2552
rect -965 -2552 -947 -2546
rect -965 -2636 -959 -2552
rect -953 -2595 -947 -2552
rect -943 -2561 -937 -2560
rect -943 -2565 -942 -2561
rect -938 -2565 -937 -2561
rect -943 -2595 -937 -2565
rect -953 -2601 -937 -2595
rect -975 -2642 -959 -2636
rect -943 -2673 -937 -2601
rect -943 -2677 -942 -2673
rect -938 -2677 -937 -2673
rect -943 -2678 -937 -2677
rect -996 -2794 -979 -2788
rect -996 -2902 -990 -2794
rect -1020 -2908 -990 -2902
rect -1268 -2995 -1146 -2989
rect -1268 -3024 -1262 -2995
rect -1006 -3003 -1000 -2908
rect -985 -2940 -979 -2794
rect -974 -2794 -958 -2788
rect -974 -2940 -968 -2794
rect -985 -2946 -968 -2940
rect -964 -2940 -958 -2794
rect -665 -2880 -655 -2482
rect 110 -2537 124 -2482
rect 144 -2488 156 -2464
rect 840 -2470 850 -1963
rect 973 -2332 1005 -2326
rect 973 -2353 979 -2332
rect 949 -2359 979 -2353
rect 999 -2353 1005 -2332
rect 1023 -2332 1057 -2326
rect 1023 -2353 1029 -2332
rect 999 -2359 1029 -2353
rect 1051 -2353 1057 -2332
rect 1080 -2332 1111 -2326
rect 1080 -2353 1086 -2332
rect 1051 -2359 1086 -2353
rect 1105 -2353 1111 -2332
rect 1133 -2332 1164 -2326
rect 1133 -2353 1139 -2332
rect 1105 -2359 1139 -2353
rect 1158 -2353 1164 -2332
rect 1183 -2332 1217 -2326
rect 1183 -2353 1189 -2332
rect 1158 -2359 1189 -2353
rect 1211 -2353 1217 -2332
rect 1242 -2353 1248 -1955
rect 1255 -2240 1272 -2234
rect 1255 -2353 1261 -2240
rect 1211 -2359 1261 -2353
rect 949 -2430 955 -2359
rect 1266 -2386 1272 -2240
rect 1277 -2240 1293 -2234
rect 1277 -2386 1283 -2240
rect 1266 -2392 1283 -2386
rect 1287 -2386 1293 -2240
rect 1287 -2392 1307 -2386
rect 949 -2434 950 -2430
rect 954 -2434 955 -2430
rect 949 -2435 955 -2434
rect 1301 -2430 1307 -2392
rect 1301 -2434 1302 -2430
rect 1306 -2434 1307 -2430
rect 1301 -2435 1307 -2434
rect 160 -2482 850 -2470
rect 160 -2488 172 -2482
rect 144 -2500 172 -2488
rect -371 -2551 -345 -2545
rect -587 -2561 -581 -2559
rect -587 -2565 -586 -2561
rect -582 -2565 -581 -2561
rect -587 -2592 -581 -2565
rect -371 -2592 -365 -2551
rect -587 -2598 -365 -2592
rect -351 -2610 -345 -2551
rect -333 -2551 -296 -2545
rect -333 -2610 -327 -2551
rect -351 -2616 -327 -2610
rect -433 -2783 -413 -2777
rect -433 -2870 -427 -2783
rect -419 -2822 -413 -2783
rect -403 -2783 -381 -2777
rect -403 -2822 -397 -2783
rect -419 -2828 -397 -2822
rect -387 -2822 -381 -2783
rect -372 -2783 -351 -2777
rect -372 -2822 -366 -2783
rect -387 -2828 -366 -2822
rect -357 -2822 -351 -2783
rect -341 -2783 -320 -2777
rect -341 -2822 -335 -2783
rect -357 -2828 -335 -2822
rect -326 -2822 -320 -2783
rect -312 -2822 -306 -2551
rect -302 -2635 -296 -2551
rect -292 -2551 -276 -2545
rect -292 -2635 -286 -2551
rect -302 -2641 -286 -2635
rect -282 -2635 -276 -2551
rect -272 -2551 -254 -2545
rect -272 -2635 -266 -2551
rect -260 -2594 -254 -2551
rect 70 -2551 93 -2537
rect 105 -2542 124 -2537
rect 105 -2546 106 -2542
rect 110 -2546 124 -2542
rect 105 -2551 124 -2546
rect 427 -2549 453 -2543
rect -229 -2561 -223 -2560
rect -229 -2565 -228 -2561
rect -224 -2565 -223 -2561
rect -229 -2594 -223 -2565
rect -260 -2600 -223 -2594
rect 70 -2596 84 -2551
rect 197 -2561 203 -2559
rect 197 -2565 198 -2561
rect 202 -2565 203 -2561
rect 197 -2590 203 -2565
rect 427 -2590 433 -2549
rect 197 -2596 433 -2590
rect 70 -2610 101 -2596
rect -282 -2641 -266 -2635
rect -326 -2828 -306 -2822
rect -466 -2876 -427 -2870
rect -665 -2890 -631 -2880
rect -954 -2915 -935 -2909
rect -641 -2911 -631 -2890
rect -954 -2940 -948 -2915
rect -964 -2946 -948 -2940
rect -1268 -3028 -1267 -3024
rect -1263 -3028 -1262 -3024
rect -1268 -3029 -1262 -3028
rect -1035 -3009 -1021 -3003
rect -1011 -3004 -1000 -3003
rect -1011 -3008 -1010 -3004
rect -1006 -3008 -1000 -3004
rect -1011 -3009 -1000 -3008
rect -1035 -3050 -1029 -3009
rect -941 -3024 -935 -2915
rect -665 -2921 -631 -2911
rect -665 -2941 -655 -2921
rect -690 -2951 -655 -2941
rect -466 -2944 -460 -2876
rect -591 -2950 -460 -2944
rect -312 -2891 -306 -2828
rect -299 -2783 -282 -2777
rect -299 -2891 -293 -2783
rect -312 -2897 -293 -2891
rect -690 -3000 -680 -2951
rect -690 -3010 -667 -3000
rect -657 -3003 -640 -3000
rect -657 -3007 -656 -3003
rect -652 -3007 -640 -3003
rect -657 -3010 -640 -3007
rect -941 -3028 -940 -3024
rect -936 -3028 -935 -3024
rect -941 -3029 -935 -3028
rect -1035 -3056 -1000 -3050
rect -1006 -3057 -1000 -3056
rect -650 -3057 -640 -3010
rect -591 -3024 -585 -2950
rect -312 -3004 -306 -2897
rect -288 -2929 -282 -2783
rect -277 -2783 -261 -2777
rect -277 -2929 -271 -2783
rect -288 -2935 -271 -2929
rect -267 -2929 -261 -2783
rect -257 -2904 -222 -2898
rect -257 -2929 -251 -2904
rect -267 -2935 -251 -2929
rect -591 -3028 -590 -3024
rect -586 -3028 -585 -3024
rect -591 -3031 -585 -3028
rect -338 -3010 -324 -3004
rect -314 -3005 -306 -3004
rect -314 -3009 -313 -3005
rect -309 -3009 -306 -3005
rect -314 -3010 -306 -3009
rect -338 -3032 -332 -3010
rect -228 -3024 -222 -2904
rect -228 -3028 -227 -3024
rect -223 -3028 -222 -3024
rect -228 -3029 -222 -3028
rect -338 -3038 -284 -3032
rect -290 -3057 -284 -3038
rect -1006 -3064 -689 -3057
rect -1035 -3065 -689 -3064
rect -1035 -3070 -1000 -3065
rect -1035 -3118 -1029 -3070
rect -697 -3081 -689 -3065
rect -658 -3065 -632 -3057
rect -658 -3081 -650 -3065
rect -697 -3089 -650 -3081
rect -640 -3081 -632 -3065
rect -601 -3065 -284 -3057
rect -601 -3081 -593 -3065
rect -640 -3089 -593 -3081
rect -290 -3088 -284 -3065
rect -338 -3094 -284 -3088
rect -1035 -3124 -1021 -3118
rect -1011 -3119 -1000 -3118
rect -1011 -3123 -1010 -3119
rect -1006 -3123 -1000 -3119
rect -1011 -3124 -1000 -3123
rect -1279 -3140 -1273 -3139
rect -1279 -3144 -1278 -3140
rect -1274 -3144 -1273 -3140
rect -1279 -3230 -1273 -3144
rect -1059 -3183 -1040 -3177
rect -1059 -3230 -1053 -3183
rect -1279 -3236 -1053 -3230
rect -1279 -3261 -1273 -3236
rect -1279 -3265 -1278 -3261
rect -1274 -3265 -1273 -3261
rect -1279 -3375 -1273 -3265
rect -1046 -3300 -1040 -3183
rect -1033 -3183 -1012 -3177
rect -1033 -3300 -1027 -3183
rect -1046 -3306 -1027 -3300
rect -1018 -3300 -1012 -3183
rect -1006 -3300 -1000 -3124
rect -338 -3119 -332 -3094
rect -338 -3125 -324 -3119
rect -314 -3120 -305 -3119
rect -314 -3124 -313 -3120
rect -309 -3124 -305 -3120
rect -314 -3125 -305 -3124
rect -941 -3140 -935 -3139
rect -941 -3144 -940 -3140
rect -936 -3144 -935 -3140
rect -995 -3183 -978 -3177
rect -995 -3300 -989 -3183
rect -1018 -3306 -989 -3300
rect -1279 -3379 -1278 -3375
rect -1274 -3379 -1273 -3375
rect -1279 -3380 -1273 -3379
rect -1006 -3701 -1000 -3306
rect -984 -3343 -978 -3183
rect -973 -3183 -956 -3177
rect -973 -3343 -967 -3183
rect -984 -3349 -967 -3343
rect -962 -3343 -956 -3183
rect -941 -3261 -935 -3144
rect -941 -3265 -940 -3261
rect -936 -3265 -935 -3261
rect -941 -3288 -935 -3265
rect -951 -3294 -935 -3288
rect -951 -3343 -945 -3294
rect -962 -3349 -945 -3343
rect -941 -3375 -935 -3294
rect -941 -3379 -940 -3375
rect -936 -3379 -935 -3375
rect -941 -3380 -935 -3379
rect -585 -3140 -579 -3139
rect -585 -3144 -584 -3140
rect -580 -3144 -579 -3140
rect -585 -3230 -579 -3144
rect -311 -3166 -305 -3125
rect -226 -3140 -220 -3139
rect -226 -3144 -225 -3140
rect -221 -3144 -220 -3140
rect -311 -3172 -284 -3166
rect -365 -3183 -346 -3177
rect -365 -3230 -359 -3183
rect -585 -3236 -359 -3230
rect -585 -3261 -579 -3236
rect -585 -3265 -584 -3261
rect -580 -3265 -579 -3261
rect -585 -3375 -579 -3265
rect -352 -3300 -346 -3183
rect -339 -3183 -318 -3177
rect -339 -3300 -333 -3183
rect -352 -3306 -333 -3300
rect -324 -3300 -318 -3183
rect -290 -3300 -284 -3172
rect -280 -3182 -263 -3176
rect -280 -3300 -274 -3182
rect -324 -3306 -274 -3300
rect -585 -3379 -584 -3375
rect -580 -3379 -579 -3375
rect -585 -3380 -579 -3379
rect -1282 -3707 -1000 -3701
rect -1282 -3746 -1276 -3707
rect -1282 -3750 -1281 -3746
rect -1277 -3750 -1276 -3746
rect -1282 -3751 -1276 -3750
rect -1006 -3747 -1000 -3707
rect -290 -3714 -284 -3306
rect -269 -3342 -263 -3182
rect -258 -3182 -241 -3176
rect -258 -3342 -252 -3182
rect -269 -3348 -252 -3342
rect -247 -3342 -241 -3182
rect -226 -3261 -220 -3144
rect -226 -3265 -225 -3261
rect -221 -3265 -220 -3261
rect -226 -3287 -220 -3265
rect -236 -3293 -220 -3287
rect -236 -3342 -230 -3293
rect -247 -3348 -230 -3342
rect -581 -3720 -284 -3714
rect -995 -3730 -978 -3724
rect -995 -3747 -989 -3730
rect -1006 -3753 -989 -3747
rect -984 -3747 -978 -3730
rect -974 -3730 -958 -3724
rect -974 -3747 -968 -3730
rect -984 -3753 -968 -3747
rect -964 -3745 -958 -3730
rect -964 -3746 -935 -3745
rect -964 -3750 -940 -3746
rect -936 -3750 -935 -3746
rect -964 -3751 -935 -3750
rect -581 -3746 -575 -3720
rect -581 -3750 -580 -3746
rect -576 -3750 -575 -3746
rect -581 -3751 -575 -3750
rect -290 -3747 -284 -3720
rect -275 -3730 -258 -3724
rect -275 -3747 -269 -3730
rect -290 -3753 -269 -3747
rect -264 -3747 -258 -3730
rect -254 -3730 -238 -3724
rect -254 -3747 -248 -3730
rect -264 -3753 -248 -3747
rect -244 -3745 -238 -3730
rect -244 -3746 -220 -3745
rect -244 -3750 -225 -3746
rect -221 -3750 -220 -3746
rect -244 -3751 -220 -3750
rect -1599 -3837 73 -3836
rect -1599 -3851 -1598 -3837
rect -1584 -3851 73 -3837
rect -1599 -3852 73 -3851
rect 87 -3842 101 -2610
rect 447 -2608 453 -2549
rect 465 -2549 509 -2543
rect 465 -2608 471 -2549
rect 447 -2614 471 -2608
rect 352 -2786 372 -2780
rect 352 -2873 358 -2786
rect 366 -2825 372 -2786
rect 382 -2786 404 -2780
rect 382 -2825 388 -2786
rect 366 -2831 388 -2825
rect 398 -2825 404 -2786
rect 413 -2786 434 -2780
rect 413 -2825 419 -2786
rect 398 -2831 419 -2825
rect 428 -2825 434 -2786
rect 444 -2786 465 -2780
rect 444 -2825 450 -2786
rect 428 -2831 450 -2825
rect 459 -2825 465 -2786
rect 492 -2825 498 -2549
rect 503 -2633 509 -2549
rect 513 -2549 529 -2543
rect 513 -2633 519 -2549
rect 503 -2639 519 -2633
rect 523 -2633 529 -2549
rect 533 -2549 551 -2543
rect 533 -2633 539 -2549
rect 545 -2592 551 -2549
rect 555 -2561 561 -2560
rect 555 -2565 556 -2561
rect 560 -2565 561 -2561
rect 555 -2592 561 -2565
rect 545 -2598 561 -2592
rect 523 -2639 539 -2633
rect 459 -2831 498 -2825
rect 319 -2879 358 -2873
rect 319 -2947 325 -2879
rect 194 -2953 325 -2947
rect 194 -3024 200 -2953
rect 492 -3002 498 -2831
rect 840 -2880 850 -2482
rect 1173 -2547 1199 -2541
rect 943 -2561 949 -2560
rect 943 -2565 944 -2561
rect 948 -2565 949 -2561
rect 943 -2588 949 -2565
rect 1173 -2588 1179 -2547
rect 943 -2594 1179 -2588
rect 1193 -2606 1199 -2547
rect 1211 -2547 1256 -2541
rect 1211 -2606 1217 -2547
rect 1193 -2612 1217 -2606
rect 840 -2890 874 -2880
rect 864 -2911 874 -2890
rect 840 -2921 874 -2911
rect 840 -2941 850 -2921
rect 194 -3028 195 -3024
rect 199 -3028 200 -3024
rect 194 -3031 200 -3028
rect 463 -3008 477 -3002
rect 487 -3003 498 -3002
rect 487 -3007 488 -3003
rect 492 -3007 498 -3003
rect 487 -3008 498 -3007
rect 820 -2951 850 -2941
rect 1238 -2947 1244 -2547
rect 1250 -2631 1256 -2547
rect 1260 -2547 1276 -2541
rect 1260 -2631 1266 -2547
rect 1250 -2637 1266 -2631
rect 1270 -2631 1276 -2547
rect 1280 -2547 1298 -2541
rect 1280 -2631 1286 -2547
rect 1292 -2590 1298 -2547
rect 1312 -2561 1318 -2560
rect 1312 -2565 1313 -2561
rect 1317 -2565 1318 -2561
rect 1312 -2590 1318 -2565
rect 1292 -2596 1318 -2590
rect 1270 -2637 1286 -2631
rect 820 -3000 830 -2951
rect 1216 -2953 1244 -2947
rect 463 -3049 469 -3008
rect 820 -3010 846 -3000
rect 856 -3003 873 -3000
rect 1216 -3003 1222 -2953
rect 856 -3007 857 -3003
rect 861 -3007 873 -3003
rect 856 -3010 873 -3007
rect 463 -3055 498 -3049
rect 492 -3058 498 -3055
rect 863 -3058 873 -3010
rect 1190 -3009 1204 -3003
rect 1214 -3004 1222 -3003
rect 1214 -3008 1215 -3004
rect 1219 -3008 1222 -3004
rect 1214 -3009 1222 -3008
rect 1190 -3031 1196 -3009
rect 1190 -3037 1244 -3031
rect 1238 -3058 1244 -3037
rect 492 -3064 838 -3058
rect 463 -3066 838 -3064
rect 463 -3070 498 -3066
rect 463 -3118 469 -3070
rect 830 -3074 838 -3066
rect 855 -3066 881 -3058
rect 855 -3074 863 -3066
rect 830 -3082 863 -3074
rect 873 -3074 881 -3066
rect 898 -3066 1244 -3058
rect 898 -3074 906 -3066
rect 873 -3082 906 -3074
rect 1238 -3087 1244 -3066
rect 1190 -3093 1244 -3087
rect 1190 -3118 1196 -3093
rect 463 -3124 477 -3118
rect 487 -3119 498 -3118
rect 487 -3123 488 -3119
rect 492 -3123 498 -3119
rect 487 -3124 498 -3123
rect 1190 -3124 1204 -3118
rect 1214 -3119 1223 -3118
rect 1214 -3123 1215 -3119
rect 1219 -3123 1223 -3119
rect 1214 -3124 1223 -3123
rect 200 -3140 206 -3139
rect 200 -3144 201 -3140
rect 205 -3144 206 -3140
rect 200 -3230 206 -3144
rect 420 -3183 439 -3177
rect 420 -3230 426 -3183
rect 200 -3236 426 -3230
rect 200 -3261 206 -3236
rect 200 -3265 201 -3261
rect 205 -3265 206 -3261
rect 200 -3266 206 -3265
rect 433 -3300 439 -3183
rect 446 -3183 467 -3177
rect 446 -3300 452 -3183
rect 433 -3306 452 -3300
rect 461 -3300 467 -3183
rect 492 -3300 498 -3124
rect 557 -3140 563 -3139
rect 557 -3144 558 -3140
rect 562 -3144 563 -3140
rect 503 -3183 520 -3177
rect 503 -3300 509 -3183
rect 461 -3306 509 -3300
rect 514 -3343 520 -3183
rect 525 -3183 542 -3177
rect 525 -3343 531 -3183
rect 514 -3349 531 -3343
rect 536 -3343 542 -3183
rect 557 -3261 563 -3144
rect 557 -3265 558 -3261
rect 562 -3265 563 -3261
rect 557 -3288 563 -3265
rect 953 -3140 959 -3139
rect 953 -3144 954 -3140
rect 958 -3144 959 -3140
rect 953 -3230 959 -3144
rect 1217 -3165 1223 -3124
rect 1313 -3140 1319 -3139
rect 1313 -3144 1314 -3140
rect 1318 -3144 1319 -3140
rect 1217 -3171 1244 -3165
rect 1173 -3183 1192 -3177
rect 1173 -3230 1179 -3183
rect 953 -3236 1179 -3230
rect 953 -3261 959 -3236
rect 953 -3265 954 -3261
rect 958 -3265 959 -3261
rect 953 -3267 959 -3265
rect 547 -3294 563 -3288
rect 547 -3343 553 -3294
rect 1186 -3300 1192 -3183
rect 1199 -3183 1220 -3177
rect 1199 -3300 1205 -3183
rect 1186 -3306 1205 -3300
rect 1214 -3300 1220 -3183
rect 1238 -3300 1244 -3171
rect 1248 -3183 1265 -3177
rect 1248 -3300 1254 -3183
rect 1214 -3306 1254 -3300
rect 536 -3349 553 -3343
rect 1259 -3343 1265 -3183
rect 1270 -3183 1287 -3177
rect 1270 -3343 1276 -3183
rect 1259 -3349 1276 -3343
rect 1281 -3343 1287 -3183
rect 1313 -3261 1319 -3144
rect 1313 -3265 1314 -3261
rect 1318 -3265 1319 -3261
rect 1313 -3288 1319 -3265
rect 1292 -3294 1319 -3288
rect 1292 -3343 1298 -3294
rect 1281 -3349 1298 -3343
rect 87 -3846 92 -3842
rect 96 -3846 101 -3842
rect 87 -3911 101 -3846
rect 87 -3925 189 -3911
rect 175 -3930 189 -3925
rect 2 -3944 189 -3930
rect 2 -3949 16 -3944
rect 2 -3963 101 -3949
rect -1273 -3977 -1267 -3976
rect -1273 -3981 -1272 -3977
rect -1268 -3981 -1267 -3977
rect -942 -3977 -936 -3976
rect -1273 -4067 -1267 -3981
rect -1058 -3986 -1038 -3980
rect -1058 -4067 -1052 -3986
rect -1273 -4073 -1052 -4067
rect -1273 -4102 -1267 -4073
rect -1273 -4106 -1272 -4102
rect -1268 -4106 -1267 -4102
rect -1273 -4226 -1267 -4106
rect -1044 -4131 -1038 -3986
rect -1032 -3986 -1015 -3980
rect -1032 -4131 -1026 -3986
rect -1021 -4093 -1015 -3986
rect -996 -3986 -979 -3980
rect -996 -4093 -990 -3986
rect -1021 -4099 -990 -4093
rect -1044 -4137 -1026 -4131
rect -1009 -4200 -1003 -4099
rect -985 -4132 -979 -3986
rect -974 -3986 -958 -3980
rect -974 -4132 -968 -3986
rect -985 -4138 -968 -4132
rect -964 -4132 -958 -3986
rect -942 -3981 -941 -3977
rect -937 -3981 -936 -3977
rect -942 -4101 -936 -3981
rect -954 -4102 -936 -4101
rect -954 -4106 -941 -4102
rect -937 -4106 -936 -4102
rect -954 -4107 -936 -4106
rect -954 -4132 -948 -4107
rect -964 -4138 -948 -4132
rect -1273 -4230 -1272 -4226
rect -1268 -4230 -1267 -4226
rect -1273 -4231 -1267 -4230
rect -1038 -4206 -1024 -4200
rect -1014 -4201 -1003 -4200
rect -1014 -4205 -1013 -4201
rect -1009 -4205 -1003 -4201
rect -1014 -4206 -1003 -4205
rect -1038 -4247 -1032 -4206
rect -942 -4226 -936 -4107
rect -942 -4230 -941 -4226
rect -937 -4230 -936 -4226
rect -942 -4231 -936 -4230
rect -584 -3977 -578 -3976
rect -227 -3977 -221 -3975
rect -584 -3981 -583 -3977
rect -579 -3981 -578 -3977
rect -584 -4064 -578 -3981
rect -364 -3983 -344 -3977
rect -364 -4064 -358 -3983
rect -584 -4070 -358 -4064
rect -584 -4102 -578 -4070
rect -584 -4106 -583 -4102
rect -579 -4106 -578 -4102
rect -584 -4226 -578 -4106
rect -350 -4128 -344 -3983
rect -338 -3983 -321 -3977
rect -338 -4128 -332 -3983
rect -327 -4090 -321 -3983
rect -301 -3983 -284 -3977
rect -301 -4090 -295 -3983
rect -327 -4096 -295 -4090
rect -350 -4134 -332 -4128
rect -315 -4202 -309 -4096
rect -290 -4129 -284 -3983
rect -279 -3983 -263 -3977
rect -279 -4129 -273 -3983
rect -290 -4135 -273 -4129
rect -269 -4129 -263 -3983
rect -227 -3981 -226 -3977
rect -222 -3981 -221 -3977
rect -227 -4101 -221 -3981
rect -259 -4102 -221 -4101
rect -259 -4106 -226 -4102
rect -222 -4106 -221 -4102
rect -259 -4107 -221 -4106
rect -259 -4129 -253 -4107
rect -269 -4135 -253 -4129
rect -584 -4230 -583 -4226
rect -579 -4230 -578 -4226
rect -700 -4239 -653 -4231
rect -1038 -4253 -1003 -4247
rect -1009 -4255 -1003 -4253
rect -700 -4255 -692 -4239
rect -1009 -4261 -692 -4255
rect -1038 -4263 -692 -4261
rect -661 -4255 -653 -4239
rect -643 -4239 -596 -4231
rect -584 -4232 -578 -4230
rect -341 -4208 -327 -4202
rect -317 -4203 -309 -4202
rect -317 -4207 -316 -4203
rect -312 -4207 -309 -4203
rect -317 -4208 -309 -4207
rect -341 -4230 -335 -4208
rect -227 -4226 -221 -4107
rect -227 -4230 -226 -4226
rect -222 -4230 -221 -4226
rect -341 -4236 -287 -4230
rect -227 -4231 -221 -4230
rect -643 -4255 -635 -4239
rect -661 -4263 -635 -4255
rect -604 -4255 -596 -4239
rect -295 -4255 -287 -4236
rect -604 -4263 -287 -4255
rect -1038 -4267 -1003 -4263
rect -1038 -4316 -1032 -4267
rect -653 -4313 -643 -4263
rect -293 -4286 -287 -4263
rect -1014 -4316 -1003 -4315
rect -1038 -4322 -1024 -4316
rect -1014 -4320 -1013 -4316
rect -1009 -4320 -1003 -4316
rect -1014 -4321 -1003 -4320
rect -1283 -4579 -1266 -4578
rect -1283 -4583 -1271 -4579
rect -1267 -4583 -1266 -4579
rect -1283 -4584 -1266 -4583
rect -1009 -4580 -1003 -4321
rect -693 -4324 -668 -4314
rect -658 -4317 -643 -4313
rect -658 -4321 -657 -4317
rect -653 -4321 -643 -4317
rect -658 -4323 -643 -4321
rect -341 -4292 -287 -4286
rect -341 -4317 -335 -4292
rect -341 -4323 -327 -4317
rect -317 -4318 -308 -4317
rect -317 -4322 -316 -4318
rect -312 -4322 -308 -4318
rect -317 -4323 -308 -4322
rect -693 -4372 -683 -4324
rect -693 -4382 -662 -4372
rect -672 -4390 -662 -4382
rect -672 -4400 -642 -4390
rect -652 -4416 -642 -4400
rect -672 -4426 -642 -4416
rect -997 -4501 -980 -4495
rect -997 -4580 -991 -4501
rect -1283 -4628 -1277 -4584
rect -1009 -4586 -991 -4580
rect -1262 -4607 -1240 -4601
rect -1262 -4628 -1256 -4607
rect -1283 -4634 -1256 -4628
rect -1246 -4628 -1240 -4607
rect -1226 -4607 -1200 -4601
rect -1226 -4628 -1220 -4607
rect -1246 -4634 -1220 -4628
rect -1206 -4628 -1200 -4607
rect -1184 -4607 -1158 -4601
rect -1184 -4628 -1178 -4607
rect -1206 -4634 -1178 -4628
rect -1164 -4628 -1158 -4607
rect -1141 -4607 -1114 -4601
rect -1141 -4628 -1135 -4607
rect -1164 -4634 -1135 -4628
rect -1120 -4628 -1114 -4607
rect -1094 -4607 -1066 -4601
rect -1094 -4628 -1088 -4607
rect -1120 -4634 -1088 -4628
rect -1072 -4628 -1066 -4607
rect -1050 -4607 -1023 -4601
rect -1050 -4628 -1044 -4607
rect -1072 -4634 -1044 -4628
rect -1029 -4628 -1023 -4607
rect -1009 -4628 -1003 -4586
rect -986 -4603 -980 -4501
rect -975 -4501 -958 -4495
rect -975 -4603 -969 -4501
rect -986 -4609 -969 -4603
rect -964 -4603 -958 -4501
rect -953 -4501 -937 -4495
rect -953 -4603 -947 -4501
rect -943 -4579 -937 -4501
rect -943 -4583 -942 -4579
rect -938 -4583 -937 -4579
rect -943 -4585 -937 -4583
rect -964 -4609 -947 -4603
rect -1029 -4634 -1003 -4628
rect -1273 -4700 -1267 -4699
rect -1273 -4704 -1272 -4700
rect -1268 -4704 -1267 -4700
rect -1273 -4749 -1267 -4704
rect -1257 -4728 -1225 -4722
rect -1257 -4749 -1251 -4728
rect -1273 -4755 -1251 -4749
rect -1231 -4749 -1225 -4728
rect -1207 -4728 -1173 -4722
rect -1207 -4749 -1201 -4728
rect -1231 -4755 -1201 -4749
rect -1179 -4749 -1173 -4728
rect -1150 -4728 -1119 -4722
rect -1150 -4749 -1144 -4728
rect -1179 -4755 -1144 -4749
rect -1125 -4749 -1119 -4728
rect -1097 -4728 -1066 -4722
rect -1097 -4749 -1091 -4728
rect -1125 -4755 -1091 -4749
rect -1072 -4749 -1066 -4728
rect -1047 -4728 -1013 -4722
rect -1047 -4749 -1041 -4728
rect -1072 -4755 -1041 -4749
rect -1019 -4749 -1013 -4728
rect -1009 -4749 -1003 -4634
rect -997 -4636 -980 -4630
rect -997 -4749 -991 -4636
rect -1019 -4755 -991 -4749
rect -1273 -4821 -1267 -4755
rect -986 -4782 -980 -4636
rect -975 -4636 -959 -4630
rect -975 -4782 -969 -4636
rect -986 -4788 -969 -4782
rect -965 -4782 -959 -4636
rect -942 -4700 -936 -4698
rect -942 -4704 -941 -4700
rect -937 -4704 -936 -4700
rect -942 -4782 -936 -4704
rect -965 -4788 -936 -4782
rect -1273 -4825 -1272 -4821
rect -1268 -4825 -1267 -4821
rect -1273 -4826 -1267 -4825
rect -942 -4821 -936 -4788
rect -942 -4825 -941 -4821
rect -937 -4825 -936 -4821
rect -942 -4826 -936 -4825
rect -672 -4849 -662 -4426
rect -588 -4579 -582 -4578
rect -588 -4583 -587 -4579
rect -583 -4583 -582 -4579
rect -588 -4628 -582 -4583
rect -567 -4607 -545 -4601
rect -567 -4628 -561 -4607
rect -588 -4634 -561 -4628
rect -551 -4628 -545 -4607
rect -531 -4607 -505 -4601
rect -531 -4628 -525 -4607
rect -551 -4634 -525 -4628
rect -511 -4628 -505 -4607
rect -489 -4607 -463 -4601
rect -489 -4628 -483 -4607
rect -511 -4634 -483 -4628
rect -469 -4628 -463 -4607
rect -446 -4607 -419 -4601
rect -446 -4628 -440 -4607
rect -469 -4634 -440 -4628
rect -425 -4628 -419 -4607
rect -399 -4607 -371 -4601
rect -399 -4628 -393 -4607
rect -425 -4634 -393 -4628
rect -377 -4628 -371 -4607
rect -355 -4607 -328 -4601
rect -355 -4628 -349 -4607
rect -377 -4634 -349 -4628
rect -334 -4628 -328 -4607
rect -314 -4628 -308 -4323
rect -334 -4634 -308 -4628
rect -588 -4700 -582 -4699
rect -588 -4704 -587 -4700
rect -583 -4704 -582 -4700
rect -588 -4749 -582 -4704
rect -562 -4728 -530 -4722
rect -562 -4749 -556 -4728
rect -588 -4755 -556 -4749
rect -536 -4749 -530 -4728
rect -512 -4728 -478 -4722
rect -512 -4749 -506 -4728
rect -536 -4755 -506 -4749
rect -484 -4749 -478 -4728
rect -455 -4728 -424 -4722
rect -455 -4749 -449 -4728
rect -484 -4755 -449 -4749
rect -430 -4749 -424 -4728
rect -402 -4728 -371 -4722
rect -402 -4749 -396 -4728
rect -430 -4755 -396 -4749
rect -377 -4749 -371 -4728
rect -352 -4728 -318 -4722
rect -352 -4749 -346 -4728
rect -377 -4755 -346 -4749
rect -324 -4749 -318 -4728
rect -314 -4749 -308 -4634
rect -299 -4636 -282 -4630
rect -299 -4749 -293 -4636
rect -324 -4755 -293 -4749
rect -588 -4821 -582 -4755
rect -288 -4782 -282 -4636
rect -277 -4636 -261 -4630
rect -277 -4782 -271 -4636
rect -288 -4788 -271 -4782
rect -267 -4782 -261 -4636
rect -227 -4700 -221 -4698
rect -227 -4704 -226 -4700
rect -222 -4704 -221 -4700
rect -227 -4782 -221 -4704
rect 87 -4732 101 -3963
rect 203 -3977 209 -3976
rect 559 -3977 565 -3975
rect 203 -3981 204 -3977
rect 208 -3981 209 -3977
rect 203 -4066 209 -3981
rect 427 -3985 447 -3979
rect 427 -4066 433 -3985
rect 203 -4072 433 -4066
rect 203 -4102 209 -4072
rect 203 -4106 204 -4102
rect 208 -4106 209 -4102
rect 203 -4108 209 -4106
rect 441 -4130 447 -3985
rect 453 -3985 470 -3979
rect 453 -4130 459 -3985
rect 464 -4092 470 -3985
rect 490 -3983 507 -3977
rect 490 -4092 496 -3983
rect 464 -4098 496 -4092
rect 441 -4136 459 -4130
rect 476 -4200 482 -4098
rect 501 -4129 507 -3983
rect 512 -3983 528 -3977
rect 512 -4129 518 -3983
rect 501 -4135 518 -4129
rect 522 -4129 528 -3983
rect 559 -3981 560 -3977
rect 564 -3981 565 -3977
rect 559 -4051 565 -3981
rect 532 -4057 565 -4051
rect 532 -4129 538 -4057
rect 559 -4102 565 -4057
rect 559 -4106 560 -4102
rect 564 -4106 565 -4102
rect 559 -4107 565 -4106
rect 944 -3977 950 -3975
rect 1314 -3977 1320 -3976
rect 944 -3981 945 -3977
rect 949 -3981 950 -3977
rect 944 -4064 950 -3981
rect 1168 -3983 1188 -3977
rect 1168 -4064 1174 -3983
rect 944 -4070 1174 -4064
rect 944 -4102 950 -4070
rect 944 -4106 945 -4102
rect 949 -4106 950 -4102
rect 944 -4108 950 -4106
rect 522 -4135 538 -4129
rect 1182 -4128 1188 -3983
rect 1194 -3983 1211 -3977
rect 1194 -4128 1200 -3983
rect 1205 -4090 1211 -3983
rect 1233 -3983 1250 -3977
rect 1233 -4090 1239 -3983
rect 1205 -4096 1239 -4090
rect 1182 -4134 1200 -4128
rect 1218 -4200 1224 -4096
rect 1244 -4129 1250 -3983
rect 1255 -3983 1271 -3977
rect 1255 -4129 1261 -3983
rect 1244 -4135 1261 -4129
rect 1265 -4129 1271 -3983
rect 1314 -3981 1315 -3977
rect 1319 -3981 1320 -3977
rect 1314 -4101 1320 -3981
rect 1275 -4102 1320 -4101
rect 1275 -4106 1315 -4102
rect 1319 -4106 1320 -4102
rect 1275 -4107 1320 -4106
rect 1275 -4129 1281 -4107
rect 1265 -4135 1281 -4129
rect 447 -4206 461 -4200
rect 471 -4201 482 -4200
rect 471 -4205 472 -4201
rect 476 -4205 482 -4201
rect 471 -4206 482 -4205
rect 1192 -4206 1206 -4200
rect 1216 -4201 1224 -4200
rect 1216 -4205 1217 -4201
rect 1221 -4205 1224 -4201
rect 1216 -4206 1224 -4205
rect 447 -4246 453 -4206
rect 890 -4239 937 -4231
rect 1192 -4233 1198 -4206
rect 1192 -4239 1246 -4233
rect 447 -4252 482 -4246
rect 476 -4255 482 -4252
rect 890 -4255 898 -4239
rect 476 -4261 898 -4255
rect 447 -4263 898 -4261
rect 929 -4255 937 -4239
rect 1240 -4255 1246 -4239
rect 929 -4263 1246 -4255
rect 447 -4267 482 -4263
rect 447 -4316 453 -4267
rect 880 -4313 890 -4263
rect 1240 -4284 1246 -4263
rect 471 -4316 482 -4315
rect 447 -4322 461 -4316
rect 471 -4320 472 -4316
rect 476 -4320 482 -4316
rect 471 -4321 482 -4320
rect -267 -4788 -221 -4782
rect -588 -4825 -587 -4821
rect -583 -4825 -582 -4821
rect -588 -4826 -582 -4825
rect -227 -4821 -221 -4788
rect 73 -4746 101 -4732
rect 201 -4700 207 -4699
rect 201 -4704 202 -4700
rect 206 -4704 207 -4700
rect 73 -4796 87 -4746
rect 201 -4749 207 -4704
rect 227 -4728 259 -4722
rect 227 -4749 233 -4728
rect 201 -4755 233 -4749
rect 253 -4749 259 -4728
rect 277 -4728 311 -4722
rect 277 -4749 283 -4728
rect 253 -4755 283 -4749
rect 305 -4749 311 -4728
rect 334 -4728 365 -4722
rect 334 -4749 340 -4728
rect 305 -4755 340 -4749
rect 359 -4749 365 -4728
rect 387 -4728 418 -4722
rect 387 -4749 393 -4728
rect 359 -4755 393 -4749
rect 412 -4749 418 -4728
rect 437 -4728 471 -4722
rect 437 -4749 443 -4728
rect 412 -4755 443 -4749
rect 465 -4749 471 -4728
rect 476 -4749 482 -4321
rect 843 -4324 865 -4314
rect 875 -4317 890 -4313
rect 875 -4321 876 -4317
rect 880 -4321 890 -4317
rect 875 -4323 890 -4321
rect 1192 -4290 1246 -4284
rect 1192 -4316 1198 -4290
rect 1216 -4316 1225 -4315
rect 1192 -4322 1206 -4316
rect 1216 -4320 1217 -4316
rect 1221 -4320 1225 -4316
rect 1216 -4321 1225 -4320
rect 843 -4372 853 -4324
rect 1219 -4357 1225 -4321
rect 1219 -4363 1246 -4357
rect 843 -4382 878 -4372
rect 868 -4390 878 -4382
rect 868 -4400 898 -4390
rect 888 -4416 898 -4400
rect 868 -4426 898 -4416
rect 486 -4636 503 -4630
rect 486 -4749 492 -4636
rect 465 -4755 492 -4749
rect 73 -4812 95 -4796
rect 105 -4802 141 -4797
rect 105 -4806 106 -4802
rect 110 -4806 141 -4802
rect 105 -4811 141 -4806
rect -227 -4825 -226 -4821
rect -222 -4825 -221 -4821
rect -227 -4826 -221 -4825
rect 127 -4849 141 -4811
rect 201 -4821 207 -4755
rect 497 -4782 503 -4636
rect 508 -4636 524 -4630
rect 508 -4782 514 -4636
rect 497 -4788 514 -4782
rect 518 -4782 524 -4636
rect 557 -4700 563 -4699
rect 557 -4704 558 -4700
rect 562 -4704 563 -4700
rect 557 -4782 563 -4704
rect 518 -4788 563 -4782
rect 201 -4825 202 -4821
rect 206 -4825 207 -4821
rect 201 -4826 207 -4825
rect 557 -4821 563 -4788
rect 557 -4825 558 -4821
rect 562 -4825 563 -4821
rect 557 -4826 563 -4825
rect 147 -4844 175 -4832
rect 147 -4849 159 -4844
rect -672 -4861 159 -4849
rect -1059 -4932 -1036 -4926
rect -1276 -4939 -1270 -4938
rect -1276 -4943 -1275 -4939
rect -1271 -4943 -1270 -4939
rect -1276 -4973 -1270 -4943
rect -1059 -4973 -1053 -4932
rect -1276 -4979 -1053 -4973
rect -1042 -4991 -1036 -4932
rect -1024 -4932 -989 -4926
rect -1024 -4991 -1018 -4932
rect -1042 -4997 -1018 -4991
rect -1056 -5182 -1036 -5176
rect -1271 -5294 -1265 -5293
rect -1271 -5298 -1270 -5294
rect -1266 -5298 -1265 -5294
rect -1271 -5336 -1265 -5298
rect -1056 -5336 -1050 -5182
rect -1042 -5327 -1036 -5182
rect -1030 -5182 -1013 -5176
rect -1030 -5327 -1024 -5182
rect -1019 -5289 -1013 -5182
rect -1006 -5289 -1000 -4932
rect -995 -5016 -989 -4932
rect -985 -4932 -969 -4926
rect -985 -5016 -979 -4932
rect -995 -5022 -979 -5016
rect -975 -5016 -969 -4932
rect -965 -4932 -947 -4926
rect -965 -5016 -959 -4932
rect -953 -4975 -947 -4932
rect -941 -4939 -935 -4938
rect -941 -4943 -940 -4939
rect -936 -4943 -935 -4939
rect -941 -4975 -935 -4943
rect -953 -4981 -935 -4975
rect -975 -5022 -959 -5016
rect -995 -5182 -978 -5176
rect -995 -5289 -989 -5182
rect -1019 -5295 -989 -5289
rect -1042 -5333 -1024 -5327
rect -1271 -5342 -1050 -5336
rect -1271 -5415 -1265 -5342
rect -1006 -5389 -1000 -5295
rect -984 -5328 -978 -5182
rect -973 -5182 -957 -5176
rect -973 -5328 -967 -5182
rect -984 -5334 -967 -5328
rect -963 -5328 -957 -5182
rect -672 -5279 -662 -4861
rect 163 -4863 175 -4844
rect 868 -4849 878 -4426
rect 954 -4700 960 -4699
rect 954 -4704 955 -4700
rect 959 -4704 960 -4700
rect 954 -4749 960 -4704
rect 980 -4728 1012 -4722
rect 980 -4749 986 -4728
rect 954 -4755 986 -4749
rect 1006 -4749 1012 -4728
rect 1030 -4728 1064 -4722
rect 1030 -4749 1036 -4728
rect 1006 -4755 1036 -4749
rect 1058 -4749 1064 -4728
rect 1087 -4728 1118 -4722
rect 1087 -4749 1093 -4728
rect 1058 -4755 1093 -4749
rect 1112 -4749 1118 -4728
rect 1140 -4728 1171 -4722
rect 1140 -4749 1146 -4728
rect 1112 -4755 1146 -4749
rect 1165 -4749 1171 -4728
rect 1190 -4728 1224 -4722
rect 1190 -4749 1196 -4728
rect 1165 -4755 1196 -4749
rect 1218 -4749 1224 -4728
rect 1240 -4749 1246 -4363
rect 1252 -4636 1269 -4630
rect 1252 -4749 1258 -4636
rect 1218 -4755 1258 -4749
rect 954 -4821 960 -4755
rect 1263 -4782 1269 -4636
rect 1274 -4636 1290 -4630
rect 1274 -4782 1280 -4636
rect 1263 -4788 1280 -4782
rect 1284 -4782 1290 -4636
rect 1314 -4700 1320 -4699
rect 1314 -4704 1315 -4700
rect 1319 -4704 1320 -4700
rect 1314 -4782 1320 -4704
rect 1284 -4788 1320 -4782
rect 954 -4825 955 -4821
rect 959 -4825 960 -4821
rect 954 -4826 960 -4825
rect 1314 -4821 1320 -4788
rect 1314 -4825 1315 -4821
rect 1319 -4825 1320 -4821
rect 1314 -4826 1320 -4825
rect 180 -4861 878 -4849
rect 180 -4863 192 -4861
rect 163 -4875 192 -4863
rect -363 -4931 -340 -4925
rect -584 -4939 -578 -4938
rect -584 -4943 -583 -4939
rect -579 -4943 -578 -4939
rect -584 -4972 -578 -4943
rect -363 -4972 -357 -4931
rect -584 -4978 -357 -4972
rect -346 -4990 -340 -4931
rect -328 -4931 -292 -4925
rect -328 -4990 -322 -4931
rect -346 -4996 -322 -4990
rect -360 -5182 -340 -5176
rect -672 -5289 -642 -5279
rect -943 -5294 -937 -5293
rect -943 -5298 -942 -5294
rect -938 -5298 -937 -5294
rect -943 -5306 -937 -5298
rect -652 -5305 -642 -5289
rect -953 -5312 -937 -5306
rect -953 -5328 -947 -5312
rect -963 -5334 -947 -5328
rect -1271 -5419 -1270 -5415
rect -1266 -5419 -1265 -5415
rect -1271 -5420 -1265 -5419
rect -1035 -5395 -1021 -5389
rect -1011 -5390 -1000 -5389
rect -1011 -5394 -1010 -5390
rect -1006 -5394 -1000 -5390
rect -1011 -5395 -1000 -5394
rect -1035 -5435 -1029 -5395
rect -943 -5415 -937 -5312
rect -672 -5315 -642 -5305
rect -672 -5329 -662 -5315
rect -692 -5339 -662 -5329
rect -360 -5336 -354 -5182
rect -346 -5327 -340 -5182
rect -334 -5182 -317 -5176
rect -334 -5327 -328 -5182
rect -323 -5289 -317 -5182
rect -310 -5289 -304 -4931
rect -298 -5015 -292 -4931
rect -288 -4931 -272 -4925
rect -288 -5015 -282 -4931
rect -298 -5021 -282 -5015
rect -278 -5015 -272 -4931
rect -268 -4931 -250 -4925
rect -268 -5015 -262 -4931
rect -256 -4974 -250 -4931
rect 434 -4930 457 -4924
rect -226 -4939 -220 -4938
rect -226 -4943 -225 -4939
rect -221 -4943 -220 -4939
rect -226 -4974 -220 -4943
rect -256 -4980 -220 -4974
rect 201 -4939 207 -4938
rect 201 -4943 202 -4939
rect 206 -4943 207 -4939
rect 201 -4971 207 -4943
rect 434 -4971 440 -4930
rect 201 -4977 440 -4971
rect 451 -4989 457 -4930
rect 469 -4930 493 -4924
rect 469 -4989 475 -4930
rect 451 -4995 475 -4989
rect -278 -5021 -262 -5015
rect -296 -5182 -279 -5176
rect -296 -5289 -290 -5182
rect -323 -5295 -290 -5289
rect -346 -5333 -328 -5327
rect -692 -5392 -682 -5339
rect -586 -5342 -354 -5336
rect -692 -5402 -668 -5392
rect -658 -5395 -640 -5391
rect -658 -5399 -657 -5395
rect -653 -5399 -640 -5395
rect -658 -5401 -640 -5399
rect -943 -5419 -942 -5415
rect -938 -5419 -937 -5415
rect -943 -5421 -937 -5419
rect -1035 -5441 -1000 -5435
rect -1006 -5448 -1000 -5441
rect -650 -5448 -640 -5401
rect -586 -5415 -580 -5342
rect -310 -5395 -304 -5295
rect -285 -5328 -279 -5182
rect -274 -5182 -258 -5176
rect -274 -5328 -268 -5182
rect -285 -5334 -268 -5328
rect -264 -5328 -258 -5182
rect 435 -5182 455 -5176
rect -254 -5312 -221 -5306
rect -254 -5328 -248 -5312
rect -264 -5334 -248 -5328
rect -586 -5419 -585 -5415
rect -581 -5419 -580 -5415
rect -586 -5421 -580 -5419
rect -336 -5401 -322 -5395
rect -312 -5396 -304 -5395
rect -312 -5400 -311 -5396
rect -307 -5400 -304 -5396
rect -312 -5401 -304 -5400
rect -336 -5423 -330 -5401
rect -227 -5415 -221 -5312
rect 435 -5336 441 -5182
rect 449 -5327 455 -5182
rect 461 -5182 478 -5176
rect 461 -5327 467 -5182
rect 472 -5289 478 -5182
rect 486 -5289 492 -4930
rect 500 -5182 517 -5176
rect 500 -5289 506 -5182
rect 472 -5295 506 -5289
rect 449 -5333 467 -5327
rect -227 -5419 -226 -5415
rect -222 -5419 -221 -5415
rect -227 -5420 -221 -5419
rect 204 -5342 441 -5336
rect 204 -5415 210 -5342
rect 486 -5389 492 -5295
rect 511 -5328 517 -5182
rect 522 -5182 538 -5176
rect 522 -5328 528 -5182
rect 511 -5334 528 -5328
rect 532 -5328 538 -5182
rect 868 -5279 878 -4861
rect 1177 -5183 1197 -5177
rect 868 -5289 898 -5279
rect 888 -5305 898 -5289
rect 542 -5312 562 -5306
rect 542 -5328 548 -5312
rect 532 -5334 548 -5328
rect 204 -5419 205 -5415
rect 209 -5419 210 -5415
rect 204 -5420 210 -5419
rect 457 -5395 471 -5389
rect 481 -5390 492 -5389
rect 481 -5394 482 -5390
rect 486 -5394 492 -5390
rect 481 -5395 492 -5394
rect -336 -5429 -282 -5423
rect -288 -5448 -282 -5429
rect 457 -5435 463 -5395
rect 556 -5415 562 -5312
rect 868 -5315 898 -5305
rect 868 -5328 878 -5315
rect 851 -5338 878 -5328
rect 1177 -5337 1183 -5183
rect 1191 -5328 1197 -5183
rect 1203 -5183 1220 -5177
rect 1203 -5328 1209 -5183
rect 1214 -5290 1220 -5183
rect 1242 -5183 1259 -5177
rect 1242 -5290 1248 -5183
rect 1214 -5296 1248 -5290
rect 1191 -5334 1209 -5328
rect 851 -5392 861 -5338
rect 951 -5343 1183 -5337
rect 851 -5402 872 -5392
rect 882 -5395 900 -5391
rect 882 -5399 883 -5395
rect 887 -5399 900 -5395
rect 882 -5401 900 -5399
rect 556 -5419 557 -5415
rect 561 -5419 562 -5415
rect 556 -5420 562 -5419
rect 457 -5441 492 -5435
rect -1006 -5456 -689 -5448
rect -1006 -5459 -1000 -5456
rect -1035 -5465 -1000 -5459
rect -1035 -5514 -1029 -5465
rect -697 -5472 -689 -5456
rect -658 -5456 -632 -5448
rect -658 -5472 -650 -5456
rect -697 -5480 -650 -5472
rect -640 -5472 -632 -5456
rect -601 -5456 -282 -5448
rect -601 -5472 -593 -5456
rect -640 -5480 -593 -5472
rect -288 -5479 -282 -5456
rect 486 -5452 492 -5441
rect 890 -5452 900 -5401
rect 951 -5415 957 -5343
rect 1227 -5398 1233 -5296
rect 1253 -5329 1259 -5183
rect 1264 -5183 1280 -5177
rect 1264 -5329 1270 -5183
rect 1253 -5335 1270 -5329
rect 1274 -5329 1280 -5183
rect 1284 -5313 1318 -5307
rect 1284 -5329 1290 -5313
rect 1274 -5335 1290 -5329
rect 951 -5419 952 -5415
rect 956 -5419 957 -5415
rect 951 -5420 957 -5419
rect 1201 -5404 1215 -5398
rect 1225 -5399 1233 -5398
rect 1225 -5403 1226 -5399
rect 1230 -5403 1233 -5399
rect 1225 -5404 1233 -5403
rect 1201 -5422 1207 -5404
rect 1312 -5415 1318 -5313
rect 1312 -5419 1313 -5415
rect 1317 -5419 1318 -5415
rect 1312 -5421 1318 -5419
rect 1201 -5428 1255 -5422
rect 1249 -5452 1255 -5428
rect 486 -5459 908 -5452
rect -336 -5485 -282 -5479
rect 457 -5460 908 -5459
rect 457 -5465 492 -5460
rect -336 -5510 -330 -5485
rect -1011 -5514 -1000 -5513
rect -1035 -5520 -1021 -5514
rect -1011 -5518 -1010 -5514
rect -1006 -5518 -1000 -5514
rect -336 -5516 -322 -5510
rect -312 -5511 -303 -5510
rect -312 -5515 -311 -5511
rect -307 -5515 -303 -5511
rect -312 -5516 -303 -5515
rect -1011 -5519 -1000 -5518
rect -1279 -5535 -1273 -5533
rect -1279 -5539 -1278 -5535
rect -1274 -5539 -1273 -5535
rect -1279 -5616 -1273 -5539
rect -1059 -5569 -1040 -5563
rect -1059 -5616 -1053 -5569
rect -1279 -5622 -1053 -5616
rect -1279 -5652 -1273 -5622
rect -1279 -5656 -1278 -5652
rect -1274 -5656 -1273 -5652
rect -1279 -5658 -1273 -5656
rect -1046 -5686 -1040 -5569
rect -1033 -5569 -1012 -5563
rect -1033 -5686 -1027 -5569
rect -1046 -5692 -1027 -5686
rect -1018 -5686 -1012 -5569
rect -1006 -5686 -1000 -5519
rect -942 -5535 -936 -5534
rect -942 -5539 -941 -5535
rect -937 -5539 -936 -5535
rect -996 -5569 -979 -5563
rect -996 -5686 -990 -5569
rect -1018 -5692 -990 -5686
rect -1256 -5917 -1224 -5911
rect -1256 -5938 -1250 -5917
rect -1272 -5944 -1250 -5938
rect -1230 -5938 -1224 -5917
rect -1206 -5917 -1172 -5911
rect -1206 -5938 -1200 -5917
rect -1230 -5944 -1200 -5938
rect -1178 -5938 -1172 -5917
rect -1149 -5917 -1118 -5911
rect -1149 -5938 -1143 -5917
rect -1178 -5944 -1143 -5938
rect -1124 -5938 -1118 -5917
rect -1096 -5917 -1065 -5911
rect -1096 -5938 -1090 -5917
rect -1124 -5944 -1090 -5938
rect -1071 -5938 -1065 -5917
rect -1046 -5917 -1012 -5911
rect -1046 -5938 -1040 -5917
rect -1071 -5944 -1040 -5938
rect -1018 -5938 -1012 -5917
rect -1006 -5938 -1000 -5692
rect -985 -5729 -979 -5569
rect -974 -5569 -957 -5563
rect -974 -5729 -968 -5569
rect -985 -5735 -968 -5729
rect -963 -5729 -957 -5569
rect -942 -5652 -936 -5539
rect -942 -5656 -941 -5652
rect -937 -5656 -936 -5652
rect -942 -5674 -936 -5656
rect -582 -5535 -576 -5533
rect -582 -5539 -581 -5535
rect -577 -5539 -576 -5535
rect -582 -5620 -576 -5539
rect -362 -5573 -343 -5567
rect -362 -5620 -356 -5573
rect -582 -5626 -356 -5620
rect -582 -5652 -576 -5626
rect -582 -5656 -581 -5652
rect -577 -5656 -576 -5652
rect -582 -5657 -576 -5656
rect -952 -5680 -936 -5674
rect -952 -5729 -946 -5680
rect -349 -5690 -343 -5573
rect -336 -5573 -315 -5567
rect -336 -5690 -330 -5573
rect -349 -5696 -330 -5690
rect -321 -5690 -315 -5573
rect -309 -5690 -303 -5516
rect 457 -5514 463 -5465
rect 900 -5476 908 -5460
rect 939 -5460 1255 -5452
rect 939 -5476 947 -5460
rect 900 -5484 947 -5476
rect 1249 -5482 1255 -5460
rect 1201 -5488 1255 -5482
rect 481 -5514 492 -5513
rect 457 -5520 471 -5514
rect 481 -5518 482 -5514
rect 486 -5518 492 -5514
rect 481 -5519 492 -5518
rect -228 -5535 -222 -5534
rect -228 -5539 -227 -5535
rect -223 -5539 -222 -5535
rect -297 -5573 -280 -5567
rect -297 -5690 -291 -5573
rect -321 -5696 -291 -5690
rect -963 -5735 -946 -5729
rect -996 -5825 -979 -5819
rect -996 -5938 -990 -5825
rect -1018 -5944 -990 -5938
rect -1272 -6011 -1266 -5944
rect -985 -5971 -979 -5825
rect -974 -5825 -958 -5819
rect -974 -5971 -968 -5825
rect -985 -5977 -968 -5971
rect -964 -5971 -958 -5825
rect -569 -5917 -537 -5911
rect -569 -5938 -563 -5917
rect -585 -5944 -563 -5938
rect -543 -5938 -537 -5917
rect -519 -5917 -485 -5911
rect -519 -5938 -513 -5917
rect -543 -5944 -513 -5938
rect -491 -5938 -485 -5917
rect -462 -5917 -431 -5911
rect -462 -5938 -456 -5917
rect -491 -5944 -456 -5938
rect -437 -5938 -431 -5917
rect -409 -5917 -378 -5911
rect -409 -5938 -403 -5917
rect -437 -5944 -403 -5938
rect -384 -5938 -378 -5917
rect -359 -5917 -325 -5911
rect -359 -5938 -353 -5917
rect -384 -5944 -353 -5938
rect -331 -5938 -325 -5917
rect -309 -5938 -303 -5696
rect -286 -5733 -280 -5573
rect -275 -5573 -258 -5567
rect -275 -5733 -269 -5573
rect -286 -5739 -269 -5733
rect -264 -5733 -258 -5573
rect -228 -5652 -222 -5539
rect -228 -5656 -227 -5652
rect -223 -5656 -222 -5652
rect -228 -5678 -222 -5656
rect 202 -5535 208 -5534
rect 202 -5539 203 -5535
rect 207 -5539 208 -5535
rect 202 -5618 208 -5539
rect 433 -5571 452 -5565
rect 433 -5618 439 -5571
rect 202 -5624 439 -5618
rect 202 -5652 208 -5624
rect 202 -5656 203 -5652
rect 207 -5656 208 -5652
rect 202 -5657 208 -5656
rect -253 -5684 -222 -5678
rect -253 -5733 -247 -5684
rect 446 -5688 452 -5571
rect 459 -5571 480 -5565
rect 459 -5688 465 -5571
rect 446 -5694 465 -5688
rect 474 -5688 480 -5571
rect 486 -5688 492 -5519
rect 1201 -5514 1207 -5488
rect 1225 -5514 1234 -5513
rect 1201 -5520 1215 -5514
rect 1225 -5518 1226 -5514
rect 1230 -5518 1234 -5514
rect 1225 -5519 1234 -5518
rect 560 -5535 566 -5534
rect 560 -5539 561 -5535
rect 565 -5539 566 -5535
rect 496 -5571 513 -5565
rect 496 -5688 502 -5571
rect 474 -5694 502 -5688
rect -264 -5739 -247 -5733
rect -296 -5825 -279 -5819
rect -296 -5938 -290 -5825
rect -331 -5944 -290 -5938
rect -964 -5977 -935 -5971
rect -1272 -6015 -1271 -6011
rect -1267 -6015 -1266 -6011
rect -1272 -6017 -1266 -6015
rect -941 -6011 -935 -5977
rect -941 -6015 -940 -6011
rect -936 -6015 -935 -6011
rect -941 -6016 -935 -6015
rect -585 -6011 -579 -5944
rect -285 -5971 -279 -5825
rect -274 -5825 -258 -5819
rect -274 -5971 -268 -5825
rect -285 -5977 -268 -5971
rect -264 -5971 -258 -5825
rect 216 -5917 248 -5911
rect 216 -5938 222 -5917
rect 200 -5944 222 -5938
rect 242 -5938 248 -5917
rect 266 -5917 300 -5911
rect 266 -5938 272 -5917
rect 242 -5944 272 -5938
rect 294 -5938 300 -5917
rect 323 -5917 354 -5911
rect 323 -5938 329 -5917
rect 294 -5944 329 -5938
rect 348 -5938 354 -5917
rect 376 -5917 407 -5911
rect 376 -5938 382 -5917
rect 348 -5944 382 -5938
rect 401 -5938 407 -5917
rect 426 -5917 460 -5911
rect 426 -5938 432 -5917
rect 401 -5944 432 -5938
rect 454 -5938 460 -5917
rect 486 -5938 492 -5694
rect 507 -5731 513 -5571
rect 518 -5571 535 -5565
rect 518 -5731 524 -5571
rect 507 -5737 524 -5731
rect 529 -5731 535 -5571
rect 560 -5652 566 -5539
rect 952 -5535 958 -5533
rect 952 -5539 953 -5535
rect 957 -5539 958 -5535
rect 952 -5618 958 -5539
rect 1228 -5555 1234 -5519
rect 1306 -5535 1321 -5534
rect 1306 -5539 1316 -5535
rect 1320 -5539 1321 -5535
rect 1306 -5540 1321 -5539
rect 1228 -5561 1255 -5555
rect 1196 -5571 1215 -5565
rect 1196 -5618 1202 -5571
rect 952 -5624 1202 -5618
rect 560 -5656 561 -5652
rect 565 -5656 566 -5652
rect 560 -5676 566 -5656
rect 540 -5682 566 -5676
rect 540 -5731 546 -5682
rect 1209 -5688 1215 -5571
rect 1222 -5571 1243 -5565
rect 1222 -5688 1228 -5571
rect 1209 -5694 1228 -5688
rect 1237 -5688 1243 -5571
rect 1249 -5688 1255 -5561
rect 1262 -5571 1279 -5565
rect 1262 -5688 1268 -5571
rect 1237 -5694 1268 -5688
rect 529 -5737 546 -5731
rect 498 -5825 515 -5819
rect 498 -5938 504 -5825
rect 454 -5944 504 -5938
rect -264 -5977 -222 -5971
rect -585 -6015 -584 -6011
rect -580 -6015 -579 -6011
rect -585 -6016 -579 -6015
rect -228 -6011 -222 -5977
rect -228 -6015 -227 -6011
rect -223 -6015 -222 -6011
rect -228 -6016 -222 -6015
rect 200 -6011 206 -5944
rect 509 -5971 515 -5825
rect 520 -5825 536 -5819
rect 520 -5971 526 -5825
rect 509 -5977 526 -5971
rect 530 -5971 536 -5825
rect 979 -5916 1011 -5910
rect 979 -5937 985 -5916
rect 956 -5943 985 -5937
rect 1005 -5937 1011 -5916
rect 1029 -5916 1063 -5910
rect 1029 -5937 1035 -5916
rect 1005 -5943 1035 -5937
rect 1057 -5937 1063 -5916
rect 1086 -5916 1117 -5910
rect 1086 -5937 1092 -5916
rect 1057 -5943 1092 -5937
rect 1111 -5937 1117 -5916
rect 1139 -5916 1170 -5910
rect 1139 -5937 1145 -5916
rect 1111 -5943 1145 -5937
rect 1164 -5937 1170 -5916
rect 1189 -5916 1223 -5910
rect 1189 -5937 1195 -5916
rect 1164 -5943 1195 -5937
rect 1217 -5937 1223 -5916
rect 1249 -5937 1255 -5694
rect 1273 -5731 1279 -5571
rect 1284 -5571 1301 -5565
rect 1284 -5731 1290 -5571
rect 1273 -5737 1290 -5731
rect 1295 -5731 1301 -5571
rect 1306 -5731 1312 -5540
rect 1295 -5737 1312 -5731
rect 1259 -5824 1276 -5818
rect 1259 -5937 1265 -5824
rect 1217 -5943 1265 -5937
rect 530 -5977 564 -5971
rect 200 -6015 201 -6011
rect 205 -6015 206 -6011
rect 200 -6017 206 -6015
rect 558 -6011 564 -5977
rect 558 -6015 559 -6011
rect 563 -6015 564 -6011
rect 558 -6016 564 -6015
rect 956 -6011 962 -5943
rect 1270 -5970 1276 -5824
rect 1281 -5824 1297 -5818
rect 1281 -5970 1287 -5824
rect 1270 -5976 1287 -5970
rect 956 -6015 957 -6011
rect 961 -6015 962 -6011
rect 956 -6016 962 -6015
rect 1291 -6061 1297 -5824
rect 1313 -6011 1319 -6010
rect 1313 -6015 1314 -6011
rect 1318 -6015 1319 -6011
rect 1313 -6061 1319 -6015
rect 1291 -6067 1319 -6061
rect 1313 -6128 1319 -6067
rect 1313 -6129 1321 -6128
rect 1313 -6133 1316 -6129
rect 1320 -6133 1321 -6129
rect 1313 -6134 1321 -6133
<< ntransistor >>
rect -1332 -1118 -1330 -1114
rect -1324 -1118 -1322 -1114
rect -1314 -1118 -1312 -1114
rect -931 -1118 -929 -1114
rect -923 -1118 -921 -1114
rect -913 -1118 -911 -1114
rect -572 -1118 -570 -1114
rect -564 -1118 -562 -1114
rect -554 -1118 -552 -1114
rect -214 -1118 -212 -1114
rect -206 -1118 -204 -1114
rect -196 -1118 -194 -1114
rect 214 -1118 216 -1114
rect 222 -1118 224 -1114
rect 232 -1118 234 -1114
rect 570 -1118 572 -1114
rect 578 -1118 580 -1114
rect 588 -1118 590 -1114
rect 968 -1118 970 -1114
rect 976 -1118 978 -1114
rect 986 -1118 988 -1114
rect 1326 -1118 1328 -1114
rect 1334 -1118 1336 -1114
rect 1344 -1118 1346 -1114
rect -1255 -1232 -1253 -1228
rect -1245 -1232 -1243 -1228
rect -1229 -1232 -1227 -1228
rect -1221 -1232 -1219 -1228
rect -1205 -1232 -1203 -1228
rect -1197 -1232 -1195 -1228
rect -1187 -1232 -1185 -1228
rect -1179 -1232 -1177 -1228
rect -1163 -1232 -1161 -1228
rect -1155 -1232 -1153 -1228
rect -1145 -1232 -1143 -1228
rect -1137 -1232 -1135 -1228
rect -1121 -1232 -1119 -1228
rect -1113 -1232 -1111 -1228
rect -1103 -1232 -1101 -1228
rect -1095 -1232 -1093 -1228
rect -1079 -1232 -1077 -1228
rect -1071 -1232 -1069 -1228
rect -930 -1232 -928 -1228
rect -920 -1232 -918 -1228
rect -904 -1232 -902 -1228
rect -896 -1232 -894 -1228
rect -880 -1232 -878 -1228
rect -872 -1232 -870 -1228
rect -862 -1232 -860 -1228
rect -854 -1232 -852 -1228
rect -838 -1232 -836 -1228
rect -830 -1232 -828 -1228
rect -820 -1232 -818 -1228
rect -812 -1232 -810 -1228
rect -796 -1232 -794 -1228
rect -788 -1232 -786 -1228
rect -778 -1232 -776 -1228
rect -770 -1232 -768 -1228
rect -754 -1232 -752 -1228
rect -746 -1232 -744 -1228
rect -572 -1232 -570 -1228
rect -562 -1232 -560 -1228
rect -546 -1232 -544 -1228
rect -538 -1232 -536 -1228
rect -522 -1232 -520 -1228
rect -514 -1232 -512 -1228
rect -504 -1232 -502 -1228
rect -496 -1232 -494 -1228
rect -480 -1232 -478 -1228
rect -472 -1232 -470 -1228
rect -462 -1232 -460 -1228
rect -454 -1232 -452 -1228
rect -438 -1232 -436 -1228
rect -430 -1232 -428 -1228
rect -420 -1232 -418 -1228
rect -412 -1232 -410 -1228
rect -396 -1232 -394 -1228
rect -388 -1232 -386 -1228
rect -214 -1232 -212 -1228
rect -204 -1232 -202 -1228
rect -188 -1232 -186 -1228
rect -180 -1232 -178 -1228
rect -164 -1232 -162 -1228
rect -156 -1232 -154 -1228
rect -146 -1232 -144 -1228
rect -138 -1232 -136 -1228
rect -122 -1232 -120 -1228
rect -114 -1232 -112 -1228
rect -104 -1232 -102 -1228
rect -96 -1232 -94 -1228
rect -80 -1232 -78 -1228
rect -72 -1232 -70 -1228
rect -62 -1232 -60 -1228
rect -54 -1232 -52 -1228
rect -38 -1232 -36 -1228
rect -30 -1232 -28 -1228
rect 214 -1232 216 -1228
rect 224 -1232 226 -1228
rect 240 -1232 242 -1228
rect 248 -1232 250 -1228
rect 264 -1232 266 -1228
rect 272 -1232 274 -1228
rect 282 -1232 284 -1228
rect 290 -1232 292 -1228
rect 306 -1232 308 -1228
rect 314 -1232 316 -1228
rect 324 -1232 326 -1228
rect 332 -1232 334 -1228
rect 348 -1232 350 -1228
rect 356 -1232 358 -1228
rect 366 -1232 368 -1228
rect 374 -1232 376 -1228
rect 390 -1232 392 -1228
rect 398 -1232 400 -1228
rect 570 -1232 572 -1228
rect 580 -1232 582 -1228
rect 596 -1232 598 -1228
rect 604 -1232 606 -1228
rect 620 -1232 622 -1228
rect 628 -1232 630 -1228
rect 638 -1232 640 -1228
rect 646 -1232 648 -1228
rect 662 -1232 664 -1228
rect 670 -1232 672 -1228
rect 680 -1232 682 -1228
rect 688 -1232 690 -1228
rect 704 -1232 706 -1228
rect 712 -1232 714 -1228
rect 722 -1232 724 -1228
rect 730 -1232 732 -1228
rect 746 -1232 748 -1228
rect 754 -1232 756 -1228
rect 968 -1232 970 -1228
rect 978 -1232 980 -1228
rect 994 -1232 996 -1228
rect 1002 -1232 1004 -1228
rect 1018 -1232 1020 -1228
rect 1026 -1232 1028 -1228
rect 1036 -1232 1038 -1228
rect 1044 -1232 1046 -1228
rect 1060 -1232 1062 -1228
rect 1068 -1232 1070 -1228
rect 1078 -1232 1080 -1228
rect 1086 -1232 1088 -1228
rect 1102 -1232 1104 -1228
rect 1110 -1232 1112 -1228
rect 1120 -1232 1122 -1228
rect 1128 -1232 1130 -1228
rect 1144 -1232 1146 -1228
rect 1152 -1232 1154 -1228
rect -1334 -1348 -1332 -1344
rect -1326 -1348 -1324 -1344
rect -1316 -1348 -1314 -1344
rect -930 -1348 -928 -1344
rect -922 -1348 -920 -1344
rect -912 -1348 -910 -1344
rect -572 -1348 -570 -1344
rect -564 -1348 -562 -1344
rect -554 -1348 -552 -1344
rect -214 -1348 -212 -1344
rect -206 -1348 -204 -1344
rect -196 -1348 -194 -1344
rect 214 -1348 216 -1344
rect 222 -1348 224 -1344
rect 232 -1348 234 -1344
rect 570 -1348 572 -1344
rect 578 -1348 580 -1344
rect 588 -1348 590 -1344
rect 968 -1348 970 -1344
rect 976 -1348 978 -1344
rect 986 -1348 988 -1344
rect 1326 -1348 1328 -1344
rect 1334 -1348 1336 -1344
rect 1344 -1348 1346 -1344
rect -1255 -1462 -1253 -1458
rect -1245 -1462 -1243 -1458
rect -1229 -1462 -1227 -1458
rect -1219 -1462 -1217 -1458
rect -1211 -1462 -1209 -1458
rect -1201 -1462 -1199 -1458
rect -1185 -1462 -1183 -1458
rect -1177 -1462 -1175 -1458
rect -1167 -1462 -1165 -1458
rect -930 -1462 -928 -1458
rect -920 -1462 -918 -1458
rect -904 -1462 -902 -1458
rect -894 -1462 -892 -1458
rect -878 -1462 -876 -1458
rect -868 -1462 -866 -1458
rect -860 -1462 -858 -1458
rect -850 -1462 -848 -1458
rect -834 -1462 -832 -1458
rect -826 -1462 -824 -1458
rect -816 -1462 -814 -1458
rect -800 -1462 -798 -1458
rect -790 -1462 -788 -1458
rect -782 -1462 -780 -1458
rect -772 -1462 -770 -1458
rect -756 -1462 -754 -1458
rect -748 -1462 -746 -1458
rect -732 -1462 -730 -1458
rect -716 -1462 -714 -1458
rect -708 -1462 -706 -1458
rect -698 -1462 -696 -1458
rect -572 -1462 -570 -1458
rect -562 -1462 -560 -1458
rect -546 -1462 -544 -1458
rect -536 -1462 -534 -1458
rect -520 -1462 -518 -1458
rect -510 -1462 -508 -1458
rect -502 -1462 -500 -1458
rect -492 -1462 -490 -1458
rect -476 -1462 -474 -1458
rect -468 -1462 -466 -1458
rect -458 -1462 -456 -1458
rect -442 -1462 -440 -1458
rect -432 -1462 -430 -1458
rect -424 -1462 -422 -1458
rect -414 -1462 -412 -1458
rect -398 -1462 -396 -1458
rect -390 -1462 -388 -1458
rect -374 -1462 -372 -1458
rect -358 -1462 -356 -1458
rect -350 -1462 -348 -1458
rect -340 -1462 -338 -1458
rect -214 -1462 -212 -1458
rect -204 -1462 -202 -1458
rect -188 -1462 -186 -1458
rect -178 -1462 -176 -1458
rect -162 -1462 -160 -1458
rect -152 -1462 -150 -1458
rect -144 -1462 -142 -1458
rect -134 -1462 -132 -1458
rect -118 -1462 -116 -1458
rect -110 -1462 -108 -1458
rect -100 -1462 -98 -1458
rect -84 -1462 -82 -1458
rect -74 -1462 -72 -1458
rect -66 -1462 -64 -1458
rect -56 -1462 -54 -1458
rect -40 -1462 -38 -1458
rect -32 -1462 -30 -1458
rect -16 -1462 -14 -1458
rect 0 -1462 2 -1458
rect 8 -1462 10 -1458
rect 18 -1462 20 -1458
rect 214 -1462 216 -1458
rect 224 -1462 226 -1458
rect 240 -1462 242 -1458
rect 250 -1462 252 -1458
rect 266 -1462 268 -1458
rect 276 -1462 278 -1458
rect 284 -1462 286 -1458
rect 294 -1462 296 -1458
rect 310 -1462 312 -1458
rect 318 -1462 320 -1458
rect 328 -1462 330 -1458
rect 344 -1462 346 -1458
rect 354 -1462 356 -1458
rect 362 -1462 364 -1458
rect 372 -1462 374 -1458
rect 388 -1462 390 -1458
rect 396 -1462 398 -1458
rect 412 -1462 414 -1458
rect 428 -1462 430 -1458
rect 436 -1462 438 -1458
rect 446 -1462 448 -1458
rect 570 -1462 572 -1458
rect 580 -1462 582 -1458
rect 596 -1462 598 -1458
rect 606 -1462 608 -1458
rect 622 -1462 624 -1458
rect 632 -1462 634 -1458
rect 640 -1462 642 -1458
rect 650 -1462 652 -1458
rect 666 -1462 668 -1458
rect 674 -1462 676 -1458
rect 684 -1462 686 -1458
rect 700 -1462 702 -1458
rect 710 -1462 712 -1458
rect 718 -1462 720 -1458
rect 728 -1462 730 -1458
rect 744 -1462 746 -1458
rect 752 -1462 754 -1458
rect 768 -1462 770 -1458
rect 784 -1462 786 -1458
rect 792 -1462 794 -1458
rect 802 -1462 804 -1458
rect 968 -1462 970 -1458
rect 978 -1462 980 -1458
rect 994 -1462 996 -1458
rect 1004 -1462 1006 -1458
rect 1020 -1462 1022 -1458
rect 1030 -1462 1032 -1458
rect 1038 -1462 1040 -1458
rect 1048 -1462 1050 -1458
rect 1064 -1462 1066 -1458
rect 1072 -1462 1074 -1458
rect 1082 -1462 1084 -1458
rect 1098 -1462 1100 -1458
rect 1108 -1462 1110 -1458
rect 1116 -1462 1118 -1458
rect 1126 -1462 1128 -1458
rect 1142 -1462 1144 -1458
rect 1150 -1462 1152 -1458
rect 1166 -1462 1168 -1458
rect 1182 -1462 1184 -1458
rect 1190 -1462 1192 -1458
rect 1200 -1462 1202 -1458
rect 1326 -1462 1328 -1458
rect 1336 -1462 1338 -1458
rect 1352 -1462 1354 -1458
rect 1362 -1462 1364 -1458
rect 1370 -1462 1372 -1458
rect 1380 -1462 1382 -1458
rect 1396 -1462 1398 -1458
rect 1404 -1462 1406 -1458
rect 1414 -1462 1416 -1458
rect -1255 -1585 -1253 -1581
rect -1245 -1585 -1243 -1581
rect -1229 -1585 -1227 -1581
rect -1221 -1585 -1219 -1581
rect -1205 -1585 -1203 -1581
rect -1197 -1585 -1195 -1581
rect -1187 -1585 -1185 -1581
rect -1179 -1585 -1177 -1581
rect -1163 -1585 -1161 -1581
rect -1155 -1585 -1153 -1581
rect -1145 -1585 -1143 -1581
rect -1137 -1585 -1135 -1581
rect -1121 -1585 -1119 -1581
rect -1113 -1585 -1111 -1581
rect -1103 -1585 -1101 -1581
rect -1095 -1585 -1093 -1581
rect -1079 -1585 -1077 -1581
rect -1071 -1585 -1069 -1581
rect -930 -1585 -928 -1581
rect -920 -1585 -918 -1581
rect -904 -1585 -902 -1581
rect -896 -1585 -894 -1581
rect -880 -1585 -878 -1581
rect -872 -1585 -870 -1581
rect -862 -1585 -860 -1581
rect -854 -1585 -852 -1581
rect -838 -1585 -836 -1581
rect -830 -1585 -828 -1581
rect -820 -1585 -818 -1581
rect -812 -1585 -810 -1581
rect -796 -1585 -794 -1581
rect -788 -1585 -786 -1581
rect -778 -1585 -776 -1581
rect -770 -1585 -768 -1581
rect -754 -1585 -752 -1581
rect -746 -1585 -744 -1581
rect -572 -1585 -570 -1581
rect -562 -1585 -560 -1581
rect -546 -1585 -544 -1581
rect -538 -1585 -536 -1581
rect -522 -1585 -520 -1581
rect -514 -1585 -512 -1581
rect -504 -1585 -502 -1581
rect -496 -1585 -494 -1581
rect -480 -1585 -478 -1581
rect -472 -1585 -470 -1581
rect -462 -1585 -460 -1581
rect -454 -1585 -452 -1581
rect -438 -1585 -436 -1581
rect -430 -1585 -428 -1581
rect -420 -1585 -418 -1581
rect -412 -1585 -410 -1581
rect -396 -1585 -394 -1581
rect -388 -1585 -386 -1581
rect -214 -1585 -212 -1581
rect -204 -1585 -202 -1581
rect -188 -1585 -186 -1581
rect -180 -1585 -178 -1581
rect -164 -1585 -162 -1581
rect -156 -1585 -154 -1581
rect -146 -1585 -144 -1581
rect -138 -1585 -136 -1581
rect -122 -1585 -120 -1581
rect -114 -1585 -112 -1581
rect -104 -1585 -102 -1581
rect -96 -1585 -94 -1581
rect -80 -1585 -78 -1581
rect -72 -1585 -70 -1581
rect -62 -1585 -60 -1581
rect -54 -1585 -52 -1581
rect -38 -1585 -36 -1581
rect -30 -1585 -28 -1581
rect 214 -1585 216 -1581
rect 224 -1585 226 -1581
rect 240 -1585 242 -1581
rect 248 -1585 250 -1581
rect 264 -1585 266 -1581
rect 272 -1585 274 -1581
rect 282 -1585 284 -1581
rect 290 -1585 292 -1581
rect 306 -1585 308 -1581
rect 314 -1585 316 -1581
rect 324 -1585 326 -1581
rect 332 -1585 334 -1581
rect 348 -1585 350 -1581
rect 356 -1585 358 -1581
rect 366 -1585 368 -1581
rect 374 -1585 376 -1581
rect 390 -1585 392 -1581
rect 398 -1585 400 -1581
rect 570 -1585 572 -1581
rect 580 -1585 582 -1581
rect 596 -1585 598 -1581
rect 604 -1585 606 -1581
rect 620 -1585 622 -1581
rect 628 -1585 630 -1581
rect 638 -1585 640 -1581
rect 646 -1585 648 -1581
rect 662 -1585 664 -1581
rect 670 -1585 672 -1581
rect 680 -1585 682 -1581
rect 688 -1585 690 -1581
rect 704 -1585 706 -1581
rect 712 -1585 714 -1581
rect 722 -1585 724 -1581
rect 730 -1585 732 -1581
rect 746 -1585 748 -1581
rect 754 -1585 756 -1581
rect 968 -1585 970 -1581
rect 978 -1585 980 -1581
rect 994 -1585 996 -1581
rect 1002 -1585 1004 -1581
rect 1018 -1585 1020 -1581
rect 1026 -1585 1028 -1581
rect 1036 -1585 1038 -1581
rect 1044 -1585 1046 -1581
rect 1060 -1585 1062 -1581
rect 1068 -1585 1070 -1581
rect 1078 -1585 1080 -1581
rect 1086 -1585 1088 -1581
rect 1102 -1585 1104 -1581
rect 1110 -1585 1112 -1581
rect 1120 -1585 1122 -1581
rect 1128 -1585 1130 -1581
rect 1144 -1585 1146 -1581
rect 1152 -1585 1154 -1581
rect -1255 -1706 -1253 -1702
rect -1245 -1706 -1243 -1702
rect -1229 -1706 -1227 -1702
rect -1221 -1706 -1219 -1702
rect -1205 -1706 -1203 -1702
rect -1197 -1706 -1195 -1702
rect -1187 -1706 -1185 -1702
rect -1179 -1706 -1177 -1702
rect -1163 -1706 -1161 -1702
rect -1155 -1706 -1153 -1702
rect -1145 -1706 -1143 -1702
rect -1137 -1706 -1135 -1702
rect -1121 -1706 -1119 -1702
rect -1113 -1706 -1111 -1702
rect -1103 -1706 -1101 -1702
rect -1095 -1706 -1093 -1702
rect -1079 -1706 -1077 -1702
rect -1071 -1706 -1069 -1702
rect -930 -1706 -928 -1702
rect -920 -1706 -918 -1702
rect -904 -1706 -902 -1702
rect -896 -1706 -894 -1702
rect -880 -1706 -878 -1702
rect -872 -1706 -870 -1702
rect -862 -1706 -860 -1702
rect -854 -1706 -852 -1702
rect -838 -1706 -836 -1702
rect -830 -1706 -828 -1702
rect -820 -1706 -818 -1702
rect -812 -1706 -810 -1702
rect -796 -1706 -794 -1702
rect -788 -1706 -786 -1702
rect -778 -1706 -776 -1702
rect -770 -1706 -768 -1702
rect -754 -1706 -752 -1702
rect -746 -1706 -744 -1702
rect -572 -1706 -570 -1702
rect -562 -1706 -560 -1702
rect -546 -1706 -544 -1702
rect -538 -1706 -536 -1702
rect -522 -1706 -520 -1702
rect -514 -1706 -512 -1702
rect -504 -1706 -502 -1702
rect -496 -1706 -494 -1702
rect -480 -1706 -478 -1702
rect -472 -1706 -470 -1702
rect -462 -1706 -460 -1702
rect -454 -1706 -452 -1702
rect -438 -1706 -436 -1702
rect -430 -1706 -428 -1702
rect -420 -1706 -418 -1702
rect -412 -1706 -410 -1702
rect -396 -1706 -394 -1702
rect -388 -1706 -386 -1702
rect -214 -1706 -212 -1702
rect -204 -1706 -202 -1702
rect -188 -1706 -186 -1702
rect -180 -1706 -178 -1702
rect -164 -1706 -162 -1702
rect -156 -1706 -154 -1702
rect -146 -1706 -144 -1702
rect -138 -1706 -136 -1702
rect -122 -1706 -120 -1702
rect -114 -1706 -112 -1702
rect -104 -1706 -102 -1702
rect -96 -1706 -94 -1702
rect -80 -1706 -78 -1702
rect -72 -1706 -70 -1702
rect -62 -1706 -60 -1702
rect -54 -1706 -52 -1702
rect -38 -1706 -36 -1702
rect -30 -1706 -28 -1702
rect 214 -1706 216 -1702
rect 224 -1706 226 -1702
rect 240 -1706 242 -1702
rect 248 -1706 250 -1702
rect 264 -1706 266 -1702
rect 272 -1706 274 -1702
rect 282 -1706 284 -1702
rect 290 -1706 292 -1702
rect 306 -1706 308 -1702
rect 314 -1706 316 -1702
rect 324 -1706 326 -1702
rect 332 -1706 334 -1702
rect 348 -1706 350 -1702
rect 356 -1706 358 -1702
rect 366 -1706 368 -1702
rect 374 -1706 376 -1702
rect 390 -1706 392 -1702
rect 398 -1706 400 -1702
rect 570 -1706 572 -1702
rect 580 -1706 582 -1702
rect 596 -1706 598 -1702
rect 604 -1706 606 -1702
rect 620 -1706 622 -1702
rect 628 -1706 630 -1702
rect 638 -1706 640 -1702
rect 646 -1706 648 -1702
rect 662 -1706 664 -1702
rect 670 -1706 672 -1702
rect 680 -1706 682 -1702
rect 688 -1706 690 -1702
rect 704 -1706 706 -1702
rect 712 -1706 714 -1702
rect 722 -1706 724 -1702
rect 730 -1706 732 -1702
rect 746 -1706 748 -1702
rect 754 -1706 756 -1702
rect 968 -1706 970 -1702
rect 978 -1706 980 -1702
rect 994 -1706 996 -1702
rect 1002 -1706 1004 -1702
rect 1018 -1706 1020 -1702
rect 1026 -1706 1028 -1702
rect 1036 -1706 1038 -1702
rect 1044 -1706 1046 -1702
rect 1060 -1706 1062 -1702
rect 1068 -1706 1070 -1702
rect 1078 -1706 1080 -1702
rect 1086 -1706 1088 -1702
rect 1102 -1706 1104 -1702
rect 1110 -1706 1112 -1702
rect 1120 -1706 1122 -1702
rect 1128 -1706 1130 -1702
rect 1144 -1706 1146 -1702
rect 1152 -1706 1154 -1702
rect 1326 -1706 1328 -1702
rect 1336 -1706 1338 -1702
rect 1352 -1706 1354 -1702
rect 1360 -1706 1362 -1702
rect 1376 -1706 1378 -1702
rect 1384 -1706 1386 -1702
rect 1394 -1706 1396 -1702
rect 1402 -1706 1404 -1702
rect 1418 -1706 1420 -1702
rect 1426 -1706 1428 -1702
rect 1436 -1706 1438 -1702
rect 1444 -1706 1446 -1702
rect 1460 -1706 1462 -1702
rect 1468 -1706 1470 -1702
rect 1478 -1706 1480 -1702
rect 1486 -1706 1488 -1702
rect 1502 -1706 1504 -1702
rect 1510 -1706 1512 -1702
rect -1255 -1827 -1253 -1823
rect -1245 -1827 -1243 -1823
rect -1229 -1827 -1227 -1823
rect -1221 -1827 -1219 -1823
rect -1205 -1827 -1203 -1823
rect -1197 -1827 -1195 -1823
rect -1187 -1827 -1185 -1823
rect -1179 -1827 -1177 -1823
rect -1163 -1827 -1161 -1823
rect -1155 -1827 -1153 -1823
rect -1145 -1827 -1143 -1823
rect -1137 -1827 -1135 -1823
rect -1121 -1827 -1119 -1823
rect -1113 -1827 -1111 -1823
rect -1103 -1827 -1101 -1823
rect -1095 -1827 -1093 -1823
rect -1079 -1827 -1077 -1823
rect -1071 -1827 -1069 -1823
rect -1024 -1827 -1022 -1823
rect -930 -1827 -928 -1823
rect -920 -1827 -918 -1823
rect -904 -1827 -902 -1823
rect -896 -1827 -894 -1823
rect -880 -1827 -878 -1823
rect -872 -1827 -870 -1823
rect -862 -1827 -860 -1823
rect -854 -1827 -852 -1823
rect -838 -1827 -836 -1823
rect -830 -1827 -828 -1823
rect -820 -1827 -818 -1823
rect -812 -1827 -810 -1823
rect -796 -1827 -794 -1823
rect -788 -1827 -786 -1823
rect -778 -1827 -776 -1823
rect -770 -1827 -768 -1823
rect -754 -1827 -752 -1823
rect -746 -1827 -744 -1823
rect -572 -1827 -570 -1823
rect -562 -1827 -560 -1823
rect -546 -1827 -544 -1823
rect -538 -1827 -536 -1823
rect -522 -1827 -520 -1823
rect -514 -1827 -512 -1823
rect -504 -1827 -502 -1823
rect -496 -1827 -494 -1823
rect -480 -1827 -478 -1823
rect -472 -1827 -470 -1823
rect -462 -1827 -460 -1823
rect -454 -1827 -452 -1823
rect -438 -1827 -436 -1823
rect -430 -1827 -428 -1823
rect -420 -1827 -418 -1823
rect -412 -1827 -410 -1823
rect -396 -1827 -394 -1823
rect -388 -1827 -386 -1823
rect -327 -1827 -325 -1823
rect -214 -1827 -212 -1823
rect -204 -1827 -202 -1823
rect -188 -1827 -186 -1823
rect -180 -1827 -178 -1823
rect -164 -1827 -162 -1823
rect -156 -1827 -154 -1823
rect -146 -1827 -144 -1823
rect -138 -1827 -136 -1823
rect -122 -1827 -120 -1823
rect -114 -1827 -112 -1823
rect -104 -1827 -102 -1823
rect -96 -1827 -94 -1823
rect -80 -1827 -78 -1823
rect -72 -1827 -70 -1823
rect -62 -1827 -60 -1823
rect -54 -1827 -52 -1823
rect -38 -1827 -36 -1823
rect -30 -1827 -28 -1823
rect 214 -1827 216 -1823
rect 224 -1827 226 -1823
rect 240 -1827 242 -1823
rect 248 -1827 250 -1823
rect 264 -1827 266 -1823
rect 272 -1827 274 -1823
rect 282 -1827 284 -1823
rect 290 -1827 292 -1823
rect 306 -1827 308 -1823
rect 314 -1827 316 -1823
rect 324 -1827 326 -1823
rect 332 -1827 334 -1823
rect 348 -1827 350 -1823
rect 356 -1827 358 -1823
rect 366 -1827 368 -1823
rect 374 -1827 376 -1823
rect 390 -1827 392 -1823
rect 398 -1827 400 -1823
rect 469 -1827 471 -1823
rect 570 -1827 572 -1823
rect 580 -1827 582 -1823
rect 596 -1827 598 -1823
rect 604 -1827 606 -1823
rect 620 -1827 622 -1823
rect 628 -1827 630 -1823
rect 638 -1827 640 -1823
rect 646 -1827 648 -1823
rect 662 -1827 664 -1823
rect 670 -1827 672 -1823
rect 680 -1827 682 -1823
rect 688 -1827 690 -1823
rect 704 -1827 706 -1823
rect 712 -1827 714 -1823
rect 722 -1827 724 -1823
rect 730 -1827 732 -1823
rect 746 -1827 748 -1823
rect 754 -1827 756 -1823
rect 968 -1827 970 -1823
rect 978 -1827 980 -1823
rect 994 -1827 996 -1823
rect 1002 -1827 1004 -1823
rect 1018 -1827 1020 -1823
rect 1026 -1827 1028 -1823
rect 1036 -1827 1038 -1823
rect 1044 -1827 1046 -1823
rect 1060 -1827 1062 -1823
rect 1068 -1827 1070 -1823
rect 1078 -1827 1080 -1823
rect 1086 -1827 1088 -1823
rect 1102 -1827 1104 -1823
rect 1110 -1827 1112 -1823
rect 1120 -1827 1122 -1823
rect 1128 -1827 1130 -1823
rect 1144 -1827 1146 -1823
rect 1152 -1827 1154 -1823
rect 1208 -1827 1210 -1823
rect 1326 -1827 1328 -1823
rect 1336 -1827 1338 -1823
rect 1352 -1827 1354 -1823
rect 1360 -1827 1362 -1823
rect 1376 -1827 1378 -1823
rect 1384 -1827 1386 -1823
rect 1394 -1827 1396 -1823
rect 1402 -1827 1404 -1823
rect 1418 -1827 1420 -1823
rect 1426 -1827 1428 -1823
rect 1436 -1827 1438 -1823
rect 1444 -1827 1446 -1823
rect 1460 -1827 1462 -1823
rect 1468 -1827 1470 -1823
rect 1478 -1827 1480 -1823
rect 1486 -1827 1488 -1823
rect 1502 -1827 1504 -1823
rect 1510 -1827 1512 -1823
rect -1255 -1942 -1253 -1938
rect -1245 -1942 -1243 -1938
rect -1229 -1942 -1227 -1938
rect -1221 -1942 -1219 -1938
rect -1205 -1942 -1203 -1938
rect -1197 -1942 -1195 -1938
rect -1187 -1942 -1185 -1938
rect -1179 -1942 -1177 -1938
rect -1163 -1942 -1161 -1938
rect -1155 -1942 -1153 -1938
rect -1145 -1942 -1143 -1938
rect -1137 -1942 -1135 -1938
rect -1121 -1942 -1119 -1938
rect -1113 -1942 -1111 -1938
rect -1103 -1942 -1101 -1938
rect -1095 -1942 -1093 -1938
rect -1079 -1942 -1077 -1938
rect -1071 -1942 -1069 -1938
rect -1024 -1942 -1022 -1938
rect -668 -1942 -666 -1934
rect -327 -1942 -325 -1938
rect 469 -1942 471 -1938
rect 846 -1942 848 -1934
rect 1208 -1942 1210 -1938
rect -1334 -2054 -1332 -2050
rect -1326 -2054 -1324 -2050
rect -1316 -2054 -1314 -2050
rect -930 -2054 -928 -2050
rect -922 -2054 -920 -2050
rect -912 -2054 -910 -2050
rect -572 -2054 -570 -2050
rect -564 -2054 -562 -2050
rect -554 -2054 -552 -2050
rect -214 -2054 -212 -2050
rect -206 -2054 -204 -2050
rect -196 -2054 -194 -2050
rect 214 -2054 216 -2050
rect 222 -2054 224 -2050
rect 232 -2054 234 -2050
rect 570 -2054 572 -2050
rect 578 -2054 580 -2050
rect 588 -2054 590 -2050
rect 968 -2054 970 -2050
rect 976 -2054 978 -2050
rect 986 -2054 988 -2050
rect 1326 -2054 1328 -2050
rect 1334 -2054 1336 -2050
rect 1344 -2054 1346 -2050
rect -1255 -2173 -1253 -2169
rect -1245 -2173 -1243 -2169
rect -1229 -2173 -1227 -2169
rect -1219 -2173 -1217 -2169
rect -1211 -2173 -1209 -2169
rect -1201 -2173 -1199 -2169
rect -1185 -2173 -1183 -2169
rect -1177 -2173 -1175 -2169
rect -1167 -2173 -1165 -2169
rect -930 -2173 -928 -2169
rect -920 -2173 -918 -2169
rect -904 -2173 -902 -2169
rect -894 -2173 -892 -2169
rect -878 -2173 -876 -2169
rect -868 -2173 -866 -2169
rect -860 -2173 -858 -2169
rect -850 -2173 -848 -2169
rect -834 -2173 -832 -2169
rect -826 -2173 -824 -2169
rect -816 -2173 -814 -2169
rect -800 -2173 -798 -2169
rect -790 -2173 -788 -2169
rect -782 -2173 -780 -2169
rect -772 -2173 -770 -2169
rect -756 -2173 -754 -2169
rect -748 -2173 -746 -2169
rect -732 -2173 -730 -2169
rect -716 -2173 -714 -2169
rect -708 -2173 -706 -2169
rect -698 -2173 -696 -2169
rect -572 -2173 -570 -2169
rect -562 -2173 -560 -2169
rect -546 -2173 -544 -2169
rect -536 -2173 -534 -2169
rect -520 -2173 -518 -2169
rect -510 -2173 -508 -2169
rect -502 -2173 -500 -2169
rect -492 -2173 -490 -2169
rect -476 -2173 -474 -2169
rect -468 -2173 -466 -2169
rect -458 -2173 -456 -2169
rect -442 -2173 -440 -2169
rect -432 -2173 -430 -2169
rect -424 -2173 -422 -2169
rect -414 -2173 -412 -2169
rect -398 -2173 -396 -2169
rect -390 -2173 -388 -2169
rect -374 -2173 -372 -2169
rect -358 -2173 -356 -2169
rect -350 -2173 -348 -2169
rect -340 -2173 -338 -2169
rect -214 -2173 -212 -2169
rect -204 -2173 -202 -2169
rect -188 -2173 -186 -2169
rect -178 -2173 -176 -2169
rect -162 -2173 -160 -2169
rect -152 -2173 -150 -2169
rect -144 -2173 -142 -2169
rect -134 -2173 -132 -2169
rect -118 -2173 -116 -2169
rect -110 -2173 -108 -2169
rect -100 -2173 -98 -2169
rect -84 -2173 -82 -2169
rect -74 -2173 -72 -2169
rect -66 -2173 -64 -2169
rect -56 -2173 -54 -2169
rect -40 -2173 -38 -2169
rect -32 -2173 -30 -2169
rect -16 -2173 -14 -2169
rect 0 -2173 2 -2169
rect 8 -2173 10 -2169
rect 18 -2173 20 -2169
rect 214 -2173 216 -2169
rect 224 -2173 226 -2169
rect 240 -2173 242 -2169
rect 250 -2173 252 -2169
rect 266 -2173 268 -2169
rect 276 -2173 278 -2169
rect 284 -2173 286 -2169
rect 294 -2173 296 -2169
rect 310 -2173 312 -2169
rect 318 -2173 320 -2169
rect 328 -2173 330 -2169
rect 344 -2173 346 -2169
rect 354 -2173 356 -2169
rect 362 -2173 364 -2169
rect 372 -2173 374 -2169
rect 388 -2173 390 -2169
rect 396 -2173 398 -2169
rect 412 -2173 414 -2169
rect 428 -2173 430 -2169
rect 436 -2173 438 -2169
rect 446 -2173 448 -2169
rect 570 -2173 572 -2169
rect 580 -2173 582 -2169
rect 596 -2173 598 -2169
rect 606 -2173 608 -2169
rect 622 -2173 624 -2169
rect 632 -2173 634 -2169
rect 640 -2173 642 -2169
rect 650 -2173 652 -2169
rect 666 -2173 668 -2169
rect 674 -2173 676 -2169
rect 684 -2173 686 -2169
rect 700 -2173 702 -2169
rect 710 -2173 712 -2169
rect 718 -2173 720 -2169
rect 728 -2173 730 -2169
rect 744 -2173 746 -2169
rect 752 -2173 754 -2169
rect 768 -2173 770 -2169
rect 784 -2173 786 -2169
rect 792 -2173 794 -2169
rect 802 -2173 804 -2169
rect 968 -2173 970 -2169
rect 978 -2173 980 -2169
rect 994 -2173 996 -2169
rect 1004 -2173 1006 -2169
rect 1020 -2173 1022 -2169
rect 1030 -2173 1032 -2169
rect 1038 -2173 1040 -2169
rect 1048 -2173 1050 -2169
rect 1064 -2173 1066 -2169
rect 1072 -2173 1074 -2169
rect 1082 -2173 1084 -2169
rect 1098 -2173 1100 -2169
rect 1108 -2173 1110 -2169
rect 1116 -2173 1118 -2169
rect 1126 -2173 1128 -2169
rect 1142 -2173 1144 -2169
rect 1150 -2173 1152 -2169
rect 1166 -2173 1168 -2169
rect 1182 -2173 1184 -2169
rect 1190 -2173 1192 -2169
rect 1200 -2173 1202 -2169
rect 1326 -2173 1328 -2169
rect 1336 -2173 1338 -2169
rect 1352 -2173 1354 -2169
rect 1362 -2173 1364 -2169
rect 1378 -2173 1380 -2169
rect 1388 -2173 1390 -2169
rect 1396 -2173 1398 -2169
rect 1406 -2173 1408 -2169
rect 1422 -2173 1424 -2169
rect 1430 -2173 1432 -2169
rect 1440 -2173 1442 -2169
rect 1456 -2173 1458 -2169
rect 1466 -2173 1468 -2169
rect 1474 -2173 1476 -2169
rect 1484 -2173 1486 -2169
rect 1500 -2173 1502 -2169
rect 1508 -2173 1510 -2169
rect 1524 -2173 1526 -2169
rect 1540 -2173 1542 -2169
rect 1548 -2173 1550 -2169
rect 1558 -2173 1560 -2169
rect -1259 -2317 -1257 -2313
rect -1249 -2317 -1247 -2313
rect -1233 -2317 -1231 -2313
rect -1225 -2317 -1223 -2313
rect -1209 -2317 -1207 -2313
rect -1201 -2317 -1199 -2313
rect -1191 -2317 -1189 -2313
rect -1183 -2317 -1181 -2313
rect -1167 -2317 -1165 -2313
rect -1159 -2317 -1157 -2313
rect -1149 -2317 -1147 -2313
rect -1141 -2317 -1139 -2313
rect -1125 -2317 -1123 -2313
rect -1117 -2317 -1115 -2313
rect -1107 -2317 -1105 -2313
rect -1099 -2317 -1097 -2313
rect -1083 -2317 -1081 -2313
rect -1075 -2317 -1073 -2313
rect -930 -2317 -928 -2313
rect -920 -2317 -918 -2313
rect -904 -2317 -902 -2313
rect -896 -2317 -894 -2313
rect -880 -2317 -878 -2313
rect -872 -2317 -870 -2313
rect -862 -2317 -860 -2313
rect -854 -2317 -852 -2313
rect -838 -2317 -836 -2313
rect -830 -2317 -828 -2313
rect -820 -2317 -818 -2313
rect -812 -2317 -810 -2313
rect -796 -2317 -794 -2313
rect -788 -2317 -786 -2313
rect -778 -2317 -776 -2313
rect -770 -2317 -768 -2313
rect -754 -2317 -752 -2313
rect -746 -2317 -744 -2313
rect -572 -2317 -570 -2313
rect -562 -2317 -560 -2313
rect -546 -2317 -544 -2313
rect -538 -2317 -536 -2313
rect -522 -2317 -520 -2313
rect -514 -2317 -512 -2313
rect -504 -2317 -502 -2313
rect -496 -2317 -494 -2313
rect -480 -2317 -478 -2313
rect -472 -2317 -470 -2313
rect -462 -2317 -460 -2313
rect -454 -2317 -452 -2313
rect -438 -2317 -436 -2313
rect -430 -2317 -428 -2313
rect -420 -2317 -418 -2313
rect -412 -2317 -410 -2313
rect -396 -2317 -394 -2313
rect -388 -2317 -386 -2313
rect -214 -2317 -212 -2313
rect -204 -2317 -202 -2313
rect -188 -2317 -186 -2313
rect -180 -2317 -178 -2313
rect -164 -2317 -162 -2313
rect -156 -2317 -154 -2313
rect -146 -2317 -144 -2313
rect -138 -2317 -136 -2313
rect -122 -2317 -120 -2313
rect -114 -2317 -112 -2313
rect -104 -2317 -102 -2313
rect -96 -2317 -94 -2313
rect -80 -2317 -78 -2313
rect -72 -2317 -70 -2313
rect -62 -2317 -60 -2313
rect -54 -2317 -52 -2313
rect -38 -2317 -36 -2313
rect -30 -2317 -28 -2313
rect 214 -2317 216 -2313
rect 224 -2317 226 -2313
rect 240 -2317 242 -2313
rect 248 -2317 250 -2313
rect 264 -2317 266 -2313
rect 272 -2317 274 -2313
rect 282 -2317 284 -2313
rect 290 -2317 292 -2313
rect 306 -2317 308 -2313
rect 314 -2317 316 -2313
rect 324 -2317 326 -2313
rect 332 -2317 334 -2313
rect 348 -2317 350 -2313
rect 356 -2317 358 -2313
rect 366 -2317 368 -2313
rect 374 -2317 376 -2313
rect 390 -2317 392 -2313
rect 398 -2317 400 -2313
rect 570 -2317 572 -2313
rect 580 -2317 582 -2313
rect 596 -2317 598 -2313
rect 604 -2317 606 -2313
rect 620 -2317 622 -2313
rect 628 -2317 630 -2313
rect 638 -2317 640 -2313
rect 646 -2317 648 -2313
rect 662 -2317 664 -2313
rect 670 -2317 672 -2313
rect 680 -2317 682 -2313
rect 688 -2317 690 -2313
rect 704 -2317 706 -2313
rect 712 -2317 714 -2313
rect 722 -2317 724 -2313
rect 730 -2317 732 -2313
rect 746 -2317 748 -2313
rect 754 -2317 756 -2313
rect -1259 -2448 -1257 -2444
rect -1249 -2448 -1247 -2444
rect -1233 -2448 -1231 -2444
rect -1225 -2448 -1223 -2444
rect -1209 -2448 -1207 -2444
rect -1201 -2448 -1199 -2444
rect -1191 -2448 -1189 -2444
rect -1183 -2448 -1181 -2444
rect -1167 -2448 -1165 -2444
rect -1159 -2448 -1157 -2444
rect -1149 -2448 -1147 -2444
rect -1141 -2448 -1139 -2444
rect -1125 -2448 -1123 -2444
rect -1117 -2448 -1115 -2444
rect -1107 -2448 -1105 -2444
rect -1099 -2448 -1097 -2444
rect -1083 -2448 -1081 -2444
rect -1075 -2448 -1073 -2444
rect -930 -2448 -928 -2444
rect -920 -2448 -918 -2444
rect -904 -2448 -902 -2444
rect -896 -2448 -894 -2444
rect -880 -2448 -878 -2444
rect -872 -2448 -870 -2444
rect -862 -2448 -860 -2444
rect -854 -2448 -852 -2444
rect -838 -2448 -836 -2444
rect -830 -2448 -828 -2444
rect -820 -2448 -818 -2444
rect -812 -2448 -810 -2444
rect -796 -2448 -794 -2444
rect -788 -2448 -786 -2444
rect -778 -2448 -776 -2444
rect -770 -2448 -768 -2444
rect -754 -2448 -752 -2444
rect -746 -2448 -744 -2444
rect -572 -2448 -570 -2444
rect -562 -2448 -560 -2444
rect -546 -2448 -544 -2444
rect -538 -2448 -536 -2444
rect -522 -2448 -520 -2444
rect -514 -2448 -512 -2444
rect -504 -2448 -502 -2444
rect -496 -2448 -494 -2444
rect -480 -2448 -478 -2444
rect -472 -2448 -470 -2444
rect -462 -2448 -460 -2444
rect -454 -2448 -452 -2444
rect -438 -2448 -436 -2444
rect -430 -2448 -428 -2444
rect -420 -2448 -418 -2444
rect -412 -2448 -410 -2444
rect -396 -2448 -394 -2444
rect -388 -2448 -386 -2444
rect -214 -2448 -212 -2444
rect -204 -2448 -202 -2444
rect -188 -2448 -186 -2444
rect -180 -2448 -178 -2444
rect -164 -2448 -162 -2444
rect -156 -2448 -154 -2444
rect -146 -2448 -144 -2444
rect -138 -2448 -136 -2444
rect -122 -2448 -120 -2444
rect -114 -2448 -112 -2444
rect -104 -2448 -102 -2444
rect -96 -2448 -94 -2444
rect -80 -2448 -78 -2444
rect -72 -2448 -70 -2444
rect -62 -2448 -60 -2444
rect -54 -2448 -52 -2444
rect -38 -2448 -36 -2444
rect -30 -2448 -28 -2444
rect 214 -2448 216 -2444
rect 224 -2448 226 -2444
rect 240 -2448 242 -2444
rect 248 -2448 250 -2444
rect 264 -2448 266 -2444
rect 272 -2448 274 -2444
rect 282 -2448 284 -2444
rect 290 -2448 292 -2444
rect 306 -2448 308 -2444
rect 314 -2448 316 -2444
rect 324 -2448 326 -2444
rect 332 -2448 334 -2444
rect 348 -2448 350 -2444
rect 356 -2448 358 -2444
rect 366 -2448 368 -2444
rect 374 -2448 376 -2444
rect 390 -2448 392 -2444
rect 398 -2448 400 -2444
rect 570 -2448 572 -2444
rect 580 -2448 582 -2444
rect 596 -2448 598 -2444
rect 604 -2448 606 -2444
rect 620 -2448 622 -2444
rect 628 -2448 630 -2444
rect 638 -2448 640 -2444
rect 646 -2448 648 -2444
rect 662 -2448 664 -2444
rect 670 -2448 672 -2444
rect 680 -2448 682 -2444
rect 688 -2448 690 -2444
rect 704 -2448 706 -2444
rect 712 -2448 714 -2444
rect 722 -2448 724 -2444
rect 730 -2448 732 -2444
rect 746 -2448 748 -2444
rect 754 -2448 756 -2444
rect 968 -2448 970 -2444
rect 978 -2448 980 -2444
rect 994 -2448 996 -2444
rect 1002 -2448 1004 -2444
rect 1018 -2448 1020 -2444
rect 1026 -2448 1028 -2444
rect 1036 -2448 1038 -2444
rect 1044 -2448 1046 -2444
rect 1060 -2448 1062 -2444
rect 1068 -2448 1070 -2444
rect 1078 -2448 1080 -2444
rect 1086 -2448 1088 -2444
rect 1102 -2448 1104 -2444
rect 1110 -2448 1112 -2444
rect 1120 -2448 1122 -2444
rect 1128 -2448 1130 -2444
rect 1144 -2448 1146 -2444
rect 1152 -2448 1154 -2444
rect 1326 -2448 1328 -2444
rect 1336 -2448 1338 -2444
rect 1352 -2448 1354 -2444
rect 1360 -2448 1362 -2444
rect 1376 -2448 1378 -2444
rect 1384 -2448 1386 -2444
rect 1394 -2448 1396 -2444
rect 1402 -2448 1404 -2444
rect 1418 -2448 1420 -2444
rect 1426 -2448 1428 -2444
rect 1436 -2448 1438 -2444
rect 1444 -2448 1446 -2444
rect 1460 -2448 1462 -2444
rect 1468 -2448 1470 -2444
rect 1478 -2448 1480 -2444
rect 1486 -2448 1488 -2444
rect 1502 -2448 1504 -2444
rect 1510 -2448 1512 -2444
rect -1259 -2579 -1257 -2575
rect -1249 -2579 -1247 -2575
rect -1233 -2579 -1231 -2575
rect -1225 -2579 -1223 -2575
rect -1209 -2579 -1207 -2575
rect -1201 -2579 -1199 -2575
rect -1191 -2579 -1189 -2575
rect -1183 -2579 -1181 -2575
rect -1167 -2579 -1165 -2575
rect -1159 -2579 -1157 -2575
rect -1149 -2579 -1147 -2575
rect -1141 -2579 -1139 -2575
rect -1125 -2579 -1123 -2575
rect -1117 -2579 -1115 -2575
rect -1107 -2579 -1105 -2575
rect -1099 -2579 -1097 -2575
rect -1083 -2579 -1081 -2575
rect -1075 -2579 -1073 -2575
rect -930 -2579 -928 -2575
rect -920 -2579 -918 -2575
rect -904 -2579 -902 -2575
rect -896 -2579 -894 -2575
rect -880 -2579 -878 -2575
rect -872 -2579 -870 -2575
rect -862 -2579 -860 -2575
rect -854 -2579 -852 -2575
rect -838 -2579 -836 -2575
rect -830 -2579 -828 -2575
rect -820 -2579 -818 -2575
rect -812 -2579 -810 -2575
rect -796 -2579 -794 -2575
rect -788 -2579 -786 -2575
rect -778 -2579 -776 -2575
rect -770 -2579 -768 -2575
rect -754 -2579 -752 -2575
rect -746 -2579 -744 -2575
rect -572 -2579 -570 -2575
rect -562 -2579 -560 -2575
rect -546 -2579 -544 -2575
rect -538 -2579 -536 -2575
rect -522 -2579 -520 -2575
rect -514 -2579 -512 -2575
rect -504 -2579 -502 -2575
rect -496 -2579 -494 -2575
rect -480 -2579 -478 -2575
rect -472 -2579 -470 -2575
rect -462 -2579 -460 -2575
rect -454 -2579 -452 -2575
rect -438 -2579 -436 -2575
rect -430 -2579 -428 -2575
rect -420 -2579 -418 -2575
rect -412 -2579 -410 -2575
rect -396 -2579 -394 -2575
rect -388 -2579 -386 -2575
rect -214 -2579 -212 -2575
rect -204 -2579 -202 -2575
rect -188 -2579 -186 -2575
rect -180 -2579 -178 -2575
rect -164 -2579 -162 -2575
rect -156 -2579 -154 -2575
rect -146 -2579 -144 -2575
rect -138 -2579 -136 -2575
rect -122 -2579 -120 -2575
rect -114 -2579 -112 -2575
rect -104 -2579 -102 -2575
rect -96 -2579 -94 -2575
rect -80 -2579 -78 -2575
rect -72 -2579 -70 -2575
rect -62 -2579 -60 -2575
rect -54 -2579 -52 -2575
rect -38 -2579 -36 -2575
rect -30 -2579 -28 -2575
rect 95 -2579 97 -2563
rect 214 -2579 216 -2575
rect 224 -2579 226 -2575
rect 240 -2579 242 -2575
rect 248 -2579 250 -2575
rect 264 -2579 266 -2575
rect 272 -2579 274 -2575
rect 282 -2579 284 -2575
rect 290 -2579 292 -2575
rect 306 -2579 308 -2575
rect 314 -2579 316 -2575
rect 324 -2579 326 -2575
rect 332 -2579 334 -2575
rect 348 -2579 350 -2575
rect 356 -2579 358 -2575
rect 366 -2579 368 -2575
rect 374 -2579 376 -2575
rect 390 -2579 392 -2575
rect 398 -2579 400 -2575
rect 570 -2579 572 -2575
rect 580 -2579 582 -2575
rect 596 -2579 598 -2575
rect 604 -2579 606 -2575
rect 620 -2579 622 -2575
rect 628 -2579 630 -2575
rect 638 -2579 640 -2575
rect 646 -2579 648 -2575
rect 662 -2579 664 -2575
rect 670 -2579 672 -2575
rect 680 -2579 682 -2575
rect 688 -2579 690 -2575
rect 704 -2579 706 -2575
rect 712 -2579 714 -2575
rect 722 -2579 724 -2575
rect 730 -2579 732 -2575
rect 746 -2579 748 -2575
rect 754 -2579 756 -2575
rect 968 -2579 970 -2575
rect 978 -2579 980 -2575
rect 994 -2579 996 -2575
rect 1002 -2579 1004 -2575
rect 1018 -2579 1020 -2575
rect 1026 -2579 1028 -2575
rect 1036 -2579 1038 -2575
rect 1044 -2579 1046 -2575
rect 1060 -2579 1062 -2575
rect 1068 -2579 1070 -2575
rect 1078 -2579 1080 -2575
rect 1086 -2579 1088 -2575
rect 1102 -2579 1104 -2575
rect 1110 -2579 1112 -2575
rect 1120 -2579 1122 -2575
rect 1128 -2579 1130 -2575
rect 1144 -2579 1146 -2575
rect 1152 -2579 1154 -2575
rect 1326 -2579 1328 -2575
rect 1336 -2579 1338 -2575
rect 1352 -2579 1354 -2575
rect 1360 -2579 1362 -2575
rect 1376 -2579 1378 -2575
rect 1384 -2579 1386 -2575
rect 1394 -2579 1396 -2575
rect 1402 -2579 1404 -2575
rect 1418 -2579 1420 -2575
rect 1426 -2579 1428 -2575
rect 1436 -2579 1438 -2575
rect 1444 -2579 1446 -2575
rect 1460 -2579 1462 -2575
rect 1468 -2579 1470 -2575
rect 1478 -2579 1480 -2575
rect 1486 -2579 1488 -2575
rect 1502 -2579 1504 -2575
rect 1510 -2579 1512 -2575
rect -1259 -2691 -1257 -2687
rect -1249 -2691 -1247 -2687
rect -1233 -2691 -1231 -2687
rect -1225 -2691 -1223 -2687
rect -1209 -2691 -1207 -2687
rect -1201 -2691 -1199 -2687
rect -1191 -2691 -1189 -2687
rect -1183 -2691 -1181 -2687
rect -1167 -2691 -1165 -2687
rect -1159 -2691 -1157 -2687
rect -1149 -2691 -1147 -2687
rect -1141 -2691 -1139 -2687
rect -1125 -2691 -1123 -2687
rect -1117 -2691 -1115 -2687
rect -1107 -2691 -1105 -2687
rect -1099 -2691 -1097 -2687
rect -1083 -2691 -1081 -2687
rect -1075 -2691 -1073 -2687
rect -930 -2691 -928 -2687
rect -920 -2691 -918 -2687
rect -904 -2691 -902 -2687
rect -896 -2691 -894 -2687
rect -880 -2691 -878 -2687
rect -872 -2691 -870 -2687
rect -862 -2691 -860 -2687
rect -854 -2691 -852 -2687
rect -838 -2691 -836 -2687
rect -830 -2691 -828 -2687
rect -820 -2691 -818 -2687
rect -812 -2691 -810 -2687
rect -796 -2691 -794 -2687
rect -788 -2691 -786 -2687
rect -778 -2691 -776 -2687
rect -770 -2691 -768 -2687
rect -754 -2691 -752 -2687
rect -746 -2691 -744 -2687
rect -1334 -2804 -1332 -2800
rect -1326 -2804 -1324 -2800
rect -1316 -2804 -1314 -2800
rect -930 -2804 -928 -2800
rect -922 -2804 -920 -2800
rect -912 -2804 -910 -2800
rect -572 -2804 -570 -2800
rect -564 -2804 -562 -2800
rect -554 -2804 -552 -2800
rect -214 -2804 -212 -2800
rect -206 -2804 -204 -2800
rect -196 -2804 -194 -2800
rect 214 -2804 216 -2800
rect 222 -2804 224 -2800
rect 232 -2804 234 -2800
rect 570 -2804 572 -2800
rect 578 -2804 580 -2800
rect 588 -2804 590 -2800
rect 968 -2804 970 -2800
rect 976 -2804 978 -2800
rect 986 -2804 988 -2800
rect 1326 -2804 1328 -2800
rect 1334 -2804 1336 -2800
rect 1344 -2804 1346 -2800
rect -1259 -2923 -1257 -2919
rect -1249 -2923 -1247 -2919
rect -1233 -2923 -1231 -2919
rect -1223 -2923 -1221 -2919
rect -1215 -2923 -1213 -2919
rect -1205 -2923 -1203 -2919
rect -1189 -2923 -1187 -2919
rect -1181 -2923 -1179 -2919
rect -1171 -2923 -1169 -2919
rect -930 -2923 -928 -2919
rect -920 -2923 -918 -2919
rect -904 -2923 -902 -2919
rect -894 -2923 -892 -2919
rect -878 -2923 -876 -2919
rect -868 -2923 -866 -2919
rect -860 -2923 -858 -2919
rect -850 -2923 -848 -2919
rect -834 -2923 -832 -2919
rect -826 -2923 -824 -2919
rect -816 -2923 -814 -2919
rect -800 -2923 -798 -2919
rect -790 -2923 -788 -2919
rect -782 -2923 -780 -2919
rect -772 -2923 -770 -2919
rect -756 -2923 -754 -2919
rect -748 -2923 -746 -2919
rect -732 -2923 -730 -2919
rect -716 -2923 -714 -2919
rect -708 -2923 -706 -2919
rect -698 -2923 -696 -2919
rect -572 -2923 -570 -2919
rect -562 -2923 -560 -2919
rect -546 -2923 -544 -2919
rect -536 -2923 -534 -2919
rect -520 -2923 -518 -2919
rect -510 -2923 -508 -2919
rect -502 -2923 -500 -2919
rect -492 -2923 -490 -2919
rect -476 -2923 -474 -2919
rect -468 -2923 -466 -2919
rect -458 -2923 -456 -2919
rect -442 -2923 -440 -2919
rect -432 -2923 -430 -2919
rect -424 -2923 -422 -2919
rect -414 -2923 -412 -2919
rect -398 -2923 -396 -2919
rect -390 -2923 -388 -2919
rect -374 -2923 -372 -2919
rect -358 -2923 -356 -2919
rect -350 -2923 -348 -2919
rect -340 -2923 -338 -2919
rect -214 -2923 -212 -2919
rect -204 -2923 -202 -2919
rect -188 -2923 -186 -2919
rect -178 -2923 -176 -2919
rect -162 -2923 -160 -2919
rect -152 -2923 -150 -2919
rect -144 -2923 -142 -2919
rect -134 -2923 -132 -2919
rect -118 -2923 -116 -2919
rect -110 -2923 -108 -2919
rect -100 -2923 -98 -2919
rect -84 -2923 -82 -2919
rect -74 -2923 -72 -2919
rect -66 -2923 -64 -2919
rect -56 -2923 -54 -2919
rect -40 -2923 -38 -2919
rect -32 -2923 -30 -2919
rect -16 -2923 -14 -2919
rect 0 -2923 2 -2919
rect 8 -2923 10 -2919
rect 18 -2923 20 -2919
rect 214 -2923 216 -2919
rect 224 -2923 226 -2919
rect 240 -2923 242 -2919
rect 250 -2923 252 -2919
rect 266 -2923 268 -2919
rect 276 -2923 278 -2919
rect 284 -2923 286 -2919
rect 294 -2923 296 -2919
rect 310 -2923 312 -2919
rect 318 -2923 320 -2919
rect 328 -2923 330 -2919
rect 344 -2923 346 -2919
rect 354 -2923 356 -2919
rect 362 -2923 364 -2919
rect 372 -2923 374 -2919
rect 388 -2923 390 -2919
rect 396 -2923 398 -2919
rect 412 -2923 414 -2919
rect 428 -2923 430 -2919
rect 436 -2923 438 -2919
rect 446 -2923 448 -2919
rect 570 -2923 572 -2919
rect 580 -2923 582 -2919
rect 596 -2923 598 -2919
rect 606 -2923 608 -2919
rect 622 -2923 624 -2919
rect 632 -2923 634 -2919
rect 640 -2923 642 -2919
rect 650 -2923 652 -2919
rect 666 -2923 668 -2919
rect 674 -2923 676 -2919
rect 684 -2923 686 -2919
rect 700 -2923 702 -2919
rect 710 -2923 712 -2919
rect 718 -2923 720 -2919
rect 728 -2923 730 -2919
rect 744 -2923 746 -2919
rect 752 -2923 754 -2919
rect 768 -2923 770 -2919
rect 784 -2923 786 -2919
rect 792 -2923 794 -2919
rect 802 -2923 804 -2919
rect 968 -2923 970 -2919
rect 978 -2923 980 -2919
rect 994 -2923 996 -2919
rect 1004 -2923 1006 -2919
rect 1020 -2923 1022 -2919
rect 1030 -2923 1032 -2919
rect 1038 -2923 1040 -2919
rect 1048 -2923 1050 -2919
rect 1064 -2923 1066 -2919
rect 1072 -2923 1074 -2919
rect 1082 -2923 1084 -2919
rect 1098 -2923 1100 -2919
rect 1108 -2923 1110 -2919
rect 1116 -2923 1118 -2919
rect 1126 -2923 1128 -2919
rect 1142 -2923 1144 -2919
rect 1150 -2923 1152 -2919
rect 1166 -2923 1168 -2919
rect 1182 -2923 1184 -2919
rect 1190 -2923 1192 -2919
rect 1200 -2923 1202 -2919
rect 1326 -2923 1328 -2919
rect 1336 -2923 1338 -2919
rect 1352 -2923 1354 -2919
rect 1362 -2923 1364 -2919
rect 1378 -2923 1380 -2919
rect 1388 -2923 1390 -2919
rect 1396 -2923 1398 -2919
rect 1406 -2923 1408 -2919
rect 1422 -2923 1424 -2919
rect 1430 -2923 1432 -2919
rect 1440 -2923 1442 -2919
rect 1456 -2923 1458 -2919
rect 1466 -2923 1468 -2919
rect 1474 -2923 1476 -2919
rect 1484 -2923 1486 -2919
rect 1500 -2923 1502 -2919
rect 1508 -2923 1510 -2919
rect 1524 -2923 1526 -2919
rect 1540 -2923 1542 -2919
rect 1548 -2923 1550 -2919
rect 1558 -2923 1560 -2919
rect -1259 -3042 -1257 -3038
rect -1249 -3042 -1247 -3038
rect -1233 -3042 -1231 -3038
rect -1225 -3042 -1223 -3038
rect -1209 -3042 -1207 -3038
rect -1201 -3042 -1199 -3038
rect -1191 -3042 -1189 -3038
rect -1183 -3042 -1181 -3038
rect -1167 -3042 -1165 -3038
rect -1159 -3042 -1157 -3038
rect -1149 -3042 -1147 -3038
rect -1141 -3042 -1139 -3038
rect -1125 -3042 -1123 -3038
rect -1117 -3042 -1115 -3038
rect -1107 -3042 -1105 -3038
rect -1099 -3042 -1097 -3038
rect -1083 -3042 -1081 -3038
rect -1075 -3042 -1073 -3038
rect -1021 -3042 -1019 -3038
rect -930 -3042 -928 -3038
rect -920 -3042 -918 -3038
rect -904 -3042 -902 -3038
rect -896 -3042 -894 -3038
rect -880 -3042 -878 -3038
rect -872 -3042 -870 -3038
rect -862 -3042 -860 -3038
rect -854 -3042 -852 -3038
rect -838 -3042 -836 -3038
rect -830 -3042 -828 -3038
rect -820 -3042 -818 -3038
rect -812 -3042 -810 -3038
rect -796 -3042 -794 -3038
rect -788 -3042 -786 -3038
rect -778 -3042 -776 -3038
rect -770 -3042 -768 -3038
rect -754 -3042 -752 -3038
rect -746 -3042 -744 -3038
rect -667 -3042 -665 -3034
rect -572 -3042 -570 -3038
rect -562 -3042 -560 -3038
rect -546 -3042 -544 -3038
rect -538 -3042 -536 -3038
rect -522 -3042 -520 -3038
rect -514 -3042 -512 -3038
rect -504 -3042 -502 -3038
rect -496 -3042 -494 -3038
rect -480 -3042 -478 -3038
rect -472 -3042 -470 -3038
rect -462 -3042 -460 -3038
rect -454 -3042 -452 -3038
rect -438 -3042 -436 -3038
rect -430 -3042 -428 -3038
rect -420 -3042 -418 -3038
rect -412 -3042 -410 -3038
rect -396 -3042 -394 -3038
rect -388 -3042 -386 -3038
rect -324 -3042 -322 -3038
rect -214 -3042 -212 -3038
rect -204 -3042 -202 -3038
rect -188 -3042 -186 -3038
rect -180 -3042 -178 -3038
rect -164 -3042 -162 -3038
rect -156 -3042 -154 -3038
rect -146 -3042 -144 -3038
rect -138 -3042 -136 -3038
rect -122 -3042 -120 -3038
rect -114 -3042 -112 -3038
rect -104 -3042 -102 -3038
rect -96 -3042 -94 -3038
rect -80 -3042 -78 -3038
rect -72 -3042 -70 -3038
rect -62 -3042 -60 -3038
rect -54 -3042 -52 -3038
rect -38 -3042 -36 -3038
rect -30 -3042 -28 -3038
rect 214 -3042 216 -3038
rect 224 -3042 226 -3038
rect 240 -3042 242 -3038
rect 248 -3042 250 -3038
rect 264 -3042 266 -3038
rect 272 -3042 274 -3038
rect 282 -3042 284 -3038
rect 290 -3042 292 -3038
rect 306 -3042 308 -3038
rect 314 -3042 316 -3038
rect 324 -3042 326 -3038
rect 332 -3042 334 -3038
rect 348 -3042 350 -3038
rect 356 -3042 358 -3038
rect 366 -3042 368 -3038
rect 374 -3042 376 -3038
rect 390 -3042 392 -3038
rect 398 -3042 400 -3038
rect 477 -3042 479 -3038
rect 846 -3042 848 -3034
rect 1204 -3042 1206 -3038
rect -1259 -3158 -1257 -3154
rect -1249 -3158 -1247 -3154
rect -1233 -3158 -1231 -3154
rect -1225 -3158 -1223 -3154
rect -1209 -3158 -1207 -3154
rect -1201 -3158 -1199 -3154
rect -1191 -3158 -1189 -3154
rect -1183 -3158 -1181 -3154
rect -1167 -3158 -1165 -3154
rect -1159 -3158 -1157 -3154
rect -1149 -3158 -1147 -3154
rect -1141 -3158 -1139 -3154
rect -1125 -3158 -1123 -3154
rect -1117 -3158 -1115 -3154
rect -1107 -3158 -1105 -3154
rect -1099 -3158 -1097 -3154
rect -1083 -3158 -1081 -3154
rect -1075 -3158 -1073 -3154
rect -1021 -3158 -1019 -3154
rect -930 -3158 -928 -3154
rect -920 -3158 -918 -3154
rect -904 -3158 -902 -3154
rect -896 -3158 -894 -3154
rect -880 -3158 -878 -3154
rect -872 -3158 -870 -3154
rect -862 -3158 -860 -3154
rect -854 -3158 -852 -3154
rect -838 -3158 -836 -3154
rect -830 -3158 -828 -3154
rect -820 -3158 -818 -3154
rect -812 -3158 -810 -3154
rect -796 -3158 -794 -3154
rect -788 -3158 -786 -3154
rect -778 -3158 -776 -3154
rect -770 -3158 -768 -3154
rect -754 -3158 -752 -3154
rect -746 -3158 -744 -3154
rect -572 -3158 -570 -3154
rect -562 -3158 -560 -3154
rect -546 -3158 -544 -3154
rect -538 -3158 -536 -3154
rect -522 -3158 -520 -3154
rect -514 -3158 -512 -3154
rect -504 -3158 -502 -3154
rect -496 -3158 -494 -3154
rect -480 -3158 -478 -3154
rect -472 -3158 -470 -3154
rect -462 -3158 -460 -3154
rect -454 -3158 -452 -3154
rect -438 -3158 -436 -3154
rect -430 -3158 -428 -3154
rect -420 -3158 -418 -3154
rect -412 -3158 -410 -3154
rect -396 -3158 -394 -3154
rect -388 -3158 -386 -3154
rect -324 -3158 -322 -3154
rect -214 -3158 -212 -3154
rect -204 -3158 -202 -3154
rect -188 -3158 -186 -3154
rect -180 -3158 -178 -3154
rect -164 -3158 -162 -3154
rect -156 -3158 -154 -3154
rect -146 -3158 -144 -3154
rect -138 -3158 -136 -3154
rect -122 -3158 -120 -3154
rect -114 -3158 -112 -3154
rect -104 -3158 -102 -3154
rect -96 -3158 -94 -3154
rect -80 -3158 -78 -3154
rect -72 -3158 -70 -3154
rect -62 -3158 -60 -3154
rect -54 -3158 -52 -3154
rect -38 -3158 -36 -3154
rect -30 -3158 -28 -3154
rect 214 -3158 216 -3154
rect 224 -3158 226 -3154
rect 240 -3158 242 -3154
rect 248 -3158 250 -3154
rect 264 -3158 266 -3154
rect 272 -3158 274 -3154
rect 282 -3158 284 -3154
rect 290 -3158 292 -3154
rect 306 -3158 308 -3154
rect 314 -3158 316 -3154
rect 324 -3158 326 -3154
rect 332 -3158 334 -3154
rect 348 -3158 350 -3154
rect 356 -3158 358 -3154
rect 366 -3158 368 -3154
rect 374 -3158 376 -3154
rect 390 -3158 392 -3154
rect 398 -3158 400 -3154
rect 477 -3158 479 -3154
rect 570 -3158 572 -3154
rect 580 -3158 582 -3154
rect 596 -3158 598 -3154
rect 604 -3158 606 -3154
rect 620 -3158 622 -3154
rect 628 -3158 630 -3154
rect 638 -3158 640 -3154
rect 646 -3158 648 -3154
rect 662 -3158 664 -3154
rect 670 -3158 672 -3154
rect 680 -3158 682 -3154
rect 688 -3158 690 -3154
rect 704 -3158 706 -3154
rect 712 -3158 714 -3154
rect 722 -3158 724 -3154
rect 730 -3158 732 -3154
rect 746 -3158 748 -3154
rect 754 -3158 756 -3154
rect 968 -3158 970 -3154
rect 978 -3158 980 -3154
rect 994 -3158 996 -3154
rect 1002 -3158 1004 -3154
rect 1018 -3158 1020 -3154
rect 1026 -3158 1028 -3154
rect 1036 -3158 1038 -3154
rect 1044 -3158 1046 -3154
rect 1060 -3158 1062 -3154
rect 1068 -3158 1070 -3154
rect 1078 -3158 1080 -3154
rect 1086 -3158 1088 -3154
rect 1102 -3158 1104 -3154
rect 1110 -3158 1112 -3154
rect 1120 -3158 1122 -3154
rect 1128 -3158 1130 -3154
rect 1144 -3158 1146 -3154
rect 1152 -3158 1154 -3154
rect 1204 -3158 1206 -3154
rect 1326 -3158 1328 -3154
rect 1336 -3158 1338 -3154
rect 1352 -3158 1354 -3154
rect 1360 -3158 1362 -3154
rect 1376 -3158 1378 -3154
rect 1384 -3158 1386 -3154
rect 1394 -3158 1396 -3154
rect 1402 -3158 1404 -3154
rect 1418 -3158 1420 -3154
rect 1426 -3158 1428 -3154
rect 1436 -3158 1438 -3154
rect 1444 -3158 1446 -3154
rect 1460 -3158 1462 -3154
rect 1468 -3158 1470 -3154
rect 1478 -3158 1480 -3154
rect 1486 -3158 1488 -3154
rect 1502 -3158 1504 -3154
rect 1510 -3158 1512 -3154
rect -1259 -3279 -1257 -3275
rect -1249 -3279 -1247 -3275
rect -1233 -3279 -1231 -3275
rect -1225 -3279 -1223 -3275
rect -1209 -3279 -1207 -3275
rect -1201 -3279 -1199 -3275
rect -1191 -3279 -1189 -3275
rect -1183 -3279 -1181 -3275
rect -1167 -3279 -1165 -3275
rect -1159 -3279 -1157 -3275
rect -1149 -3279 -1147 -3275
rect -1141 -3279 -1139 -3275
rect -1125 -3279 -1123 -3275
rect -1117 -3279 -1115 -3275
rect -1107 -3279 -1105 -3275
rect -1099 -3279 -1097 -3275
rect -1083 -3279 -1081 -3275
rect -1075 -3279 -1073 -3275
rect -930 -3279 -928 -3275
rect -920 -3279 -918 -3275
rect -904 -3279 -902 -3275
rect -896 -3279 -894 -3275
rect -880 -3279 -878 -3275
rect -872 -3279 -870 -3275
rect -862 -3279 -860 -3275
rect -854 -3279 -852 -3275
rect -838 -3279 -836 -3275
rect -830 -3279 -828 -3275
rect -820 -3279 -818 -3275
rect -812 -3279 -810 -3275
rect -796 -3279 -794 -3275
rect -788 -3279 -786 -3275
rect -778 -3279 -776 -3275
rect -770 -3279 -768 -3275
rect -754 -3279 -752 -3275
rect -746 -3279 -744 -3275
rect -572 -3279 -570 -3275
rect -562 -3279 -560 -3275
rect -546 -3279 -544 -3275
rect -538 -3279 -536 -3275
rect -522 -3279 -520 -3275
rect -514 -3279 -512 -3275
rect -504 -3279 -502 -3275
rect -496 -3279 -494 -3275
rect -480 -3279 -478 -3275
rect -472 -3279 -470 -3275
rect -462 -3279 -460 -3275
rect -454 -3279 -452 -3275
rect -438 -3279 -436 -3275
rect -430 -3279 -428 -3275
rect -420 -3279 -418 -3275
rect -412 -3279 -410 -3275
rect -396 -3279 -394 -3275
rect -388 -3279 -386 -3275
rect -214 -3279 -212 -3275
rect -204 -3279 -202 -3275
rect -188 -3279 -186 -3275
rect -180 -3279 -178 -3275
rect -164 -3279 -162 -3275
rect -156 -3279 -154 -3275
rect -146 -3279 -144 -3275
rect -138 -3279 -136 -3275
rect -122 -3279 -120 -3275
rect -114 -3279 -112 -3275
rect -104 -3279 -102 -3275
rect -96 -3279 -94 -3275
rect -80 -3279 -78 -3275
rect -72 -3279 -70 -3275
rect -62 -3279 -60 -3275
rect -54 -3279 -52 -3275
rect -38 -3279 -36 -3275
rect -30 -3279 -28 -3275
rect 214 -3279 216 -3275
rect 224 -3279 226 -3275
rect 240 -3279 242 -3275
rect 248 -3279 250 -3275
rect 264 -3279 266 -3275
rect 272 -3279 274 -3275
rect 282 -3279 284 -3275
rect 290 -3279 292 -3275
rect 306 -3279 308 -3275
rect 314 -3279 316 -3275
rect 324 -3279 326 -3275
rect 332 -3279 334 -3275
rect 348 -3279 350 -3275
rect 356 -3279 358 -3275
rect 366 -3279 368 -3275
rect 374 -3279 376 -3275
rect 390 -3279 392 -3275
rect 398 -3279 400 -3275
rect 570 -3279 572 -3275
rect 580 -3279 582 -3275
rect 596 -3279 598 -3275
rect 604 -3279 606 -3275
rect 620 -3279 622 -3275
rect 628 -3279 630 -3275
rect 638 -3279 640 -3275
rect 646 -3279 648 -3275
rect 662 -3279 664 -3275
rect 670 -3279 672 -3275
rect 680 -3279 682 -3275
rect 688 -3279 690 -3275
rect 704 -3279 706 -3275
rect 712 -3279 714 -3275
rect 722 -3279 724 -3275
rect 730 -3279 732 -3275
rect 746 -3279 748 -3275
rect 754 -3279 756 -3275
rect 968 -3279 970 -3275
rect 978 -3279 980 -3275
rect 994 -3279 996 -3275
rect 1002 -3279 1004 -3275
rect 1018 -3279 1020 -3275
rect 1026 -3279 1028 -3275
rect 1036 -3279 1038 -3275
rect 1044 -3279 1046 -3275
rect 1060 -3279 1062 -3275
rect 1068 -3279 1070 -3275
rect 1078 -3279 1080 -3275
rect 1086 -3279 1088 -3275
rect 1102 -3279 1104 -3275
rect 1110 -3279 1112 -3275
rect 1120 -3279 1122 -3275
rect 1128 -3279 1130 -3275
rect 1144 -3279 1146 -3275
rect 1152 -3279 1154 -3275
rect 1326 -3279 1328 -3275
rect 1336 -3279 1338 -3275
rect 1352 -3279 1354 -3275
rect 1360 -3279 1362 -3275
rect 1376 -3279 1378 -3275
rect 1384 -3279 1386 -3275
rect 1394 -3279 1396 -3275
rect 1402 -3279 1404 -3275
rect 1418 -3279 1420 -3275
rect 1426 -3279 1428 -3275
rect 1436 -3279 1438 -3275
rect 1444 -3279 1446 -3275
rect 1460 -3279 1462 -3275
rect 1468 -3279 1470 -3275
rect 1478 -3279 1480 -3275
rect 1486 -3279 1488 -3275
rect 1502 -3279 1504 -3275
rect 1510 -3279 1512 -3275
rect -1259 -3393 -1257 -3389
rect -1249 -3393 -1247 -3389
rect -1233 -3393 -1231 -3389
rect -1225 -3393 -1223 -3389
rect -1209 -3393 -1207 -3389
rect -1201 -3393 -1199 -3389
rect -1191 -3393 -1189 -3389
rect -1183 -3393 -1181 -3389
rect -1167 -3393 -1165 -3389
rect -1159 -3393 -1157 -3389
rect -1149 -3393 -1147 -3389
rect -1141 -3393 -1139 -3389
rect -1125 -3393 -1123 -3389
rect -1117 -3393 -1115 -3389
rect -1107 -3393 -1105 -3389
rect -1099 -3393 -1097 -3389
rect -1083 -3393 -1081 -3389
rect -1075 -3393 -1073 -3389
rect -930 -3393 -928 -3389
rect -920 -3393 -918 -3389
rect -904 -3393 -902 -3389
rect -896 -3393 -894 -3389
rect -880 -3393 -878 -3389
rect -872 -3393 -870 -3389
rect -862 -3393 -860 -3389
rect -854 -3393 -852 -3389
rect -838 -3393 -836 -3389
rect -830 -3393 -828 -3389
rect -820 -3393 -818 -3389
rect -812 -3393 -810 -3389
rect -796 -3393 -794 -3389
rect -788 -3393 -786 -3389
rect -778 -3393 -776 -3389
rect -770 -3393 -768 -3389
rect -754 -3393 -752 -3389
rect -746 -3393 -744 -3389
rect -572 -3393 -570 -3389
rect -562 -3393 -560 -3389
rect -546 -3393 -544 -3389
rect -538 -3393 -536 -3389
rect -522 -3393 -520 -3389
rect -514 -3393 -512 -3389
rect -504 -3393 -502 -3389
rect -496 -3393 -494 -3389
rect -480 -3393 -478 -3389
rect -472 -3393 -470 -3389
rect -462 -3393 -460 -3389
rect -454 -3393 -452 -3389
rect -438 -3393 -436 -3389
rect -430 -3393 -428 -3389
rect -420 -3393 -418 -3389
rect -412 -3393 -410 -3389
rect -396 -3393 -394 -3389
rect -388 -3393 -386 -3389
rect -1334 -3510 -1332 -3506
rect -1326 -3510 -1324 -3506
rect -1316 -3510 -1314 -3506
rect -930 -3510 -928 -3506
rect -922 -3510 -920 -3506
rect -912 -3510 -910 -3506
rect -572 -3510 -570 -3506
rect -564 -3510 -562 -3506
rect -554 -3510 -552 -3506
rect -214 -3510 -212 -3506
rect -206 -3510 -204 -3506
rect -196 -3510 -194 -3506
rect 214 -3510 216 -3506
rect 222 -3510 224 -3506
rect 232 -3510 234 -3506
rect 570 -3510 572 -3506
rect 578 -3510 580 -3506
rect 588 -3510 590 -3506
rect 968 -3510 970 -3506
rect 976 -3510 978 -3506
rect 986 -3510 988 -3506
rect 1326 -3510 1328 -3506
rect 1334 -3510 1336 -3506
rect 1344 -3510 1346 -3506
rect -1259 -3634 -1257 -3630
rect -1249 -3634 -1247 -3630
rect -1233 -3634 -1231 -3630
rect -1223 -3634 -1221 -3630
rect -1215 -3634 -1213 -3630
rect -1205 -3634 -1203 -3630
rect -1189 -3634 -1187 -3630
rect -1181 -3634 -1179 -3630
rect -1171 -3634 -1169 -3630
rect -930 -3634 -928 -3630
rect -920 -3634 -918 -3630
rect -904 -3634 -902 -3630
rect -894 -3634 -892 -3630
rect -878 -3634 -876 -3630
rect -868 -3634 -866 -3630
rect -860 -3634 -858 -3630
rect -850 -3634 -848 -3630
rect -834 -3634 -832 -3630
rect -826 -3634 -824 -3630
rect -816 -3634 -814 -3630
rect -800 -3634 -798 -3630
rect -790 -3634 -788 -3630
rect -782 -3634 -780 -3630
rect -772 -3634 -770 -3630
rect -756 -3634 -754 -3630
rect -748 -3634 -746 -3630
rect -732 -3634 -730 -3630
rect -716 -3634 -714 -3630
rect -708 -3634 -706 -3630
rect -698 -3634 -696 -3630
rect -572 -3634 -570 -3630
rect -562 -3634 -560 -3630
rect -546 -3634 -544 -3630
rect -536 -3634 -534 -3630
rect -520 -3634 -518 -3630
rect -510 -3634 -508 -3630
rect -502 -3634 -500 -3630
rect -492 -3634 -490 -3630
rect -476 -3634 -474 -3630
rect -468 -3634 -466 -3630
rect -458 -3634 -456 -3630
rect -442 -3634 -440 -3630
rect -432 -3634 -430 -3630
rect -424 -3634 -422 -3630
rect -414 -3634 -412 -3630
rect -398 -3634 -396 -3630
rect -390 -3634 -388 -3630
rect -374 -3634 -372 -3630
rect -358 -3634 -356 -3630
rect -350 -3634 -348 -3630
rect -340 -3634 -338 -3630
rect -214 -3634 -212 -3630
rect -204 -3634 -202 -3630
rect -188 -3634 -186 -3630
rect -178 -3634 -176 -3630
rect -162 -3634 -160 -3630
rect -152 -3634 -150 -3630
rect -144 -3634 -142 -3630
rect -134 -3634 -132 -3630
rect -118 -3634 -116 -3630
rect -110 -3634 -108 -3630
rect -100 -3634 -98 -3630
rect -84 -3634 -82 -3630
rect -74 -3634 -72 -3630
rect -66 -3634 -64 -3630
rect -56 -3634 -54 -3630
rect -40 -3634 -38 -3630
rect -32 -3634 -30 -3630
rect -16 -3634 -14 -3630
rect 0 -3634 2 -3630
rect 8 -3634 10 -3630
rect 18 -3634 20 -3630
rect 214 -3634 216 -3630
rect 224 -3634 226 -3630
rect 240 -3634 242 -3630
rect 250 -3634 252 -3630
rect 266 -3634 268 -3630
rect 276 -3634 278 -3630
rect 284 -3634 286 -3630
rect 294 -3634 296 -3630
rect 310 -3634 312 -3630
rect 318 -3634 320 -3630
rect 328 -3634 330 -3630
rect 344 -3634 346 -3630
rect 354 -3634 356 -3630
rect 362 -3634 364 -3630
rect 372 -3634 374 -3630
rect 388 -3634 390 -3630
rect 396 -3634 398 -3630
rect 412 -3634 414 -3630
rect 428 -3634 430 -3630
rect 436 -3634 438 -3630
rect 446 -3634 448 -3630
rect 570 -3634 572 -3630
rect 580 -3634 582 -3630
rect 596 -3634 598 -3630
rect 606 -3634 608 -3630
rect 622 -3634 624 -3630
rect 632 -3634 634 -3630
rect 640 -3634 642 -3630
rect 650 -3634 652 -3630
rect 666 -3634 668 -3630
rect 674 -3634 676 -3630
rect 684 -3634 686 -3630
rect 700 -3634 702 -3630
rect 710 -3634 712 -3630
rect 718 -3634 720 -3630
rect 728 -3634 730 -3630
rect 744 -3634 746 -3630
rect 752 -3634 754 -3630
rect 768 -3634 770 -3630
rect 784 -3634 786 -3630
rect 792 -3634 794 -3630
rect 802 -3634 804 -3630
rect 968 -3634 970 -3630
rect 978 -3634 980 -3630
rect 994 -3634 996 -3630
rect 1004 -3634 1006 -3630
rect 1020 -3634 1022 -3630
rect 1030 -3634 1032 -3630
rect 1038 -3634 1040 -3630
rect 1048 -3634 1050 -3630
rect 1064 -3634 1066 -3630
rect 1072 -3634 1074 -3630
rect 1082 -3634 1084 -3630
rect 1098 -3634 1100 -3630
rect 1108 -3634 1110 -3630
rect 1116 -3634 1118 -3630
rect 1126 -3634 1128 -3630
rect 1142 -3634 1144 -3630
rect 1150 -3634 1152 -3630
rect 1166 -3634 1168 -3630
rect 1182 -3634 1184 -3630
rect 1190 -3634 1192 -3630
rect 1200 -3634 1202 -3630
rect 1326 -3634 1328 -3630
rect 1336 -3634 1338 -3630
rect 1352 -3634 1354 -3630
rect 1362 -3634 1364 -3630
rect 1378 -3634 1380 -3630
rect 1388 -3634 1390 -3630
rect 1396 -3634 1398 -3630
rect 1406 -3634 1408 -3630
rect 1422 -3634 1424 -3630
rect 1430 -3634 1432 -3630
rect 1440 -3634 1442 -3630
rect 1456 -3634 1458 -3630
rect 1466 -3634 1468 -3630
rect 1474 -3634 1476 -3630
rect 1484 -3634 1486 -3630
rect 1500 -3634 1502 -3630
rect 1508 -3634 1510 -3630
rect 1524 -3634 1526 -3630
rect 1540 -3634 1542 -3630
rect 1548 -3634 1550 -3630
rect 1558 -3634 1560 -3630
rect -1259 -3764 -1257 -3760
rect -1249 -3764 -1247 -3760
rect -1233 -3764 -1231 -3760
rect -1225 -3764 -1223 -3760
rect -1209 -3764 -1207 -3760
rect -1201 -3764 -1199 -3760
rect -1191 -3764 -1189 -3760
rect -1183 -3764 -1181 -3760
rect -1167 -3764 -1165 -3760
rect -1159 -3764 -1157 -3760
rect -1149 -3764 -1147 -3760
rect -1141 -3764 -1139 -3760
rect -1125 -3764 -1123 -3760
rect -1117 -3764 -1115 -3760
rect -1107 -3764 -1105 -3760
rect -1099 -3764 -1097 -3760
rect -1083 -3764 -1081 -3760
rect -1075 -3764 -1073 -3760
rect -930 -3764 -928 -3760
rect -920 -3764 -918 -3760
rect -904 -3764 -902 -3760
rect -896 -3764 -894 -3760
rect -880 -3764 -878 -3760
rect -872 -3764 -870 -3760
rect -862 -3764 -860 -3760
rect -854 -3764 -852 -3760
rect -838 -3764 -836 -3760
rect -830 -3764 -828 -3760
rect -820 -3764 -818 -3760
rect -812 -3764 -810 -3760
rect -796 -3764 -794 -3760
rect -788 -3764 -786 -3760
rect -778 -3764 -776 -3760
rect -770 -3764 -768 -3760
rect -754 -3764 -752 -3760
rect -746 -3764 -744 -3760
rect -572 -3764 -570 -3760
rect -562 -3764 -560 -3760
rect -546 -3764 -544 -3760
rect -538 -3764 -536 -3760
rect -522 -3764 -520 -3760
rect -514 -3764 -512 -3760
rect -504 -3764 -502 -3760
rect -496 -3764 -494 -3760
rect -480 -3764 -478 -3760
rect -472 -3764 -470 -3760
rect -462 -3764 -460 -3760
rect -454 -3764 -452 -3760
rect -438 -3764 -436 -3760
rect -430 -3764 -428 -3760
rect -420 -3764 -418 -3760
rect -412 -3764 -410 -3760
rect -396 -3764 -394 -3760
rect -388 -3764 -386 -3760
rect -214 -3764 -212 -3760
rect -204 -3764 -202 -3760
rect -188 -3764 -186 -3760
rect -180 -3764 -178 -3760
rect -164 -3764 -162 -3760
rect -156 -3764 -154 -3760
rect -146 -3764 -144 -3760
rect -138 -3764 -136 -3760
rect -122 -3764 -120 -3760
rect -114 -3764 -112 -3760
rect -104 -3764 -102 -3760
rect -96 -3764 -94 -3760
rect -80 -3764 -78 -3760
rect -72 -3764 -70 -3760
rect -62 -3764 -60 -3760
rect -54 -3764 -52 -3760
rect -38 -3764 -36 -3760
rect -30 -3764 -28 -3760
rect 73 -3879 75 -3863
rect -1259 -3995 -1257 -3991
rect -1249 -3995 -1247 -3991
rect -1233 -3995 -1231 -3991
rect -1225 -3995 -1223 -3991
rect -1209 -3995 -1207 -3991
rect -1201 -3995 -1199 -3991
rect -1191 -3995 -1189 -3991
rect -1183 -3995 -1181 -3991
rect -1167 -3995 -1165 -3991
rect -1159 -3995 -1157 -3991
rect -1149 -3995 -1147 -3991
rect -1141 -3995 -1139 -3991
rect -1125 -3995 -1123 -3991
rect -1117 -3995 -1115 -3991
rect -1107 -3995 -1105 -3991
rect -1099 -3995 -1097 -3991
rect -1083 -3995 -1081 -3991
rect -1075 -3995 -1073 -3991
rect -930 -3995 -928 -3991
rect -920 -3995 -918 -3991
rect -904 -3995 -902 -3991
rect -896 -3995 -894 -3991
rect -880 -3995 -878 -3991
rect -872 -3995 -870 -3991
rect -862 -3995 -860 -3991
rect -854 -3995 -852 -3991
rect -838 -3995 -836 -3991
rect -830 -3995 -828 -3991
rect -820 -3995 -818 -3991
rect -812 -3995 -810 -3991
rect -796 -3995 -794 -3991
rect -788 -3995 -786 -3991
rect -778 -3995 -776 -3991
rect -770 -3995 -768 -3991
rect -754 -3995 -752 -3991
rect -746 -3995 -744 -3991
rect -572 -3995 -570 -3991
rect -562 -3995 -560 -3991
rect -546 -3995 -544 -3991
rect -538 -3995 -536 -3991
rect -522 -3995 -520 -3991
rect -514 -3995 -512 -3991
rect -504 -3995 -502 -3991
rect -496 -3995 -494 -3991
rect -480 -3995 -478 -3991
rect -472 -3995 -470 -3991
rect -462 -3995 -460 -3991
rect -454 -3995 -452 -3991
rect -438 -3995 -436 -3991
rect -430 -3995 -428 -3991
rect -420 -3995 -418 -3991
rect -412 -3995 -410 -3991
rect -396 -3995 -394 -3991
rect -388 -3995 -386 -3991
rect -214 -3995 -212 -3991
rect -204 -3995 -202 -3991
rect -188 -3995 -186 -3991
rect -180 -3995 -178 -3991
rect -164 -3995 -162 -3991
rect -156 -3995 -154 -3991
rect -146 -3995 -144 -3991
rect -138 -3995 -136 -3991
rect -122 -3995 -120 -3991
rect -114 -3995 -112 -3991
rect -104 -3995 -102 -3991
rect -96 -3995 -94 -3991
rect -80 -3995 -78 -3991
rect -72 -3995 -70 -3991
rect -62 -3995 -60 -3991
rect -54 -3995 -52 -3991
rect -38 -3995 -36 -3991
rect -30 -3995 -28 -3991
rect 214 -3995 216 -3991
rect 224 -3995 226 -3991
rect 240 -3995 242 -3991
rect 248 -3995 250 -3991
rect 264 -3995 266 -3991
rect 272 -3995 274 -3991
rect 282 -3995 284 -3991
rect 290 -3995 292 -3991
rect 306 -3995 308 -3991
rect 314 -3995 316 -3991
rect 324 -3995 326 -3991
rect 332 -3995 334 -3991
rect 348 -3995 350 -3991
rect 356 -3995 358 -3991
rect 366 -3995 368 -3991
rect 374 -3995 376 -3991
rect 390 -3995 392 -3991
rect 398 -3995 400 -3991
rect 570 -3995 572 -3991
rect 580 -3995 582 -3991
rect 596 -3995 598 -3991
rect 604 -3995 606 -3991
rect 620 -3995 622 -3991
rect 628 -3995 630 -3991
rect 638 -3995 640 -3991
rect 646 -3995 648 -3991
rect 662 -3995 664 -3991
rect 670 -3995 672 -3991
rect 680 -3995 682 -3991
rect 688 -3995 690 -3991
rect 704 -3995 706 -3991
rect 712 -3995 714 -3991
rect 722 -3995 724 -3991
rect 730 -3995 732 -3991
rect 746 -3995 748 -3991
rect 754 -3995 756 -3991
rect 968 -3995 970 -3991
rect 978 -3995 980 -3991
rect 994 -3995 996 -3991
rect 1002 -3995 1004 -3991
rect 1018 -3995 1020 -3991
rect 1026 -3995 1028 -3991
rect 1036 -3995 1038 -3991
rect 1044 -3995 1046 -3991
rect 1060 -3995 1062 -3991
rect 1068 -3995 1070 -3991
rect 1078 -3995 1080 -3991
rect 1086 -3995 1088 -3991
rect 1102 -3995 1104 -3991
rect 1110 -3995 1112 -3991
rect 1120 -3995 1122 -3991
rect 1128 -3995 1130 -3991
rect 1144 -3995 1146 -3991
rect 1152 -3995 1154 -3991
rect 1326 -3995 1328 -3991
rect 1336 -3995 1338 -3991
rect 1352 -3995 1354 -3991
rect 1360 -3995 1362 -3991
rect 1376 -3995 1378 -3991
rect 1384 -3995 1386 -3991
rect 1394 -3995 1396 -3991
rect 1402 -3995 1404 -3991
rect 1418 -3995 1420 -3991
rect 1426 -3995 1428 -3991
rect 1436 -3995 1438 -3991
rect 1444 -3995 1446 -3991
rect 1460 -3995 1462 -3991
rect 1468 -3995 1470 -3991
rect 1478 -3995 1480 -3991
rect 1486 -3995 1488 -3991
rect 1502 -3995 1504 -3991
rect 1510 -3995 1512 -3991
rect -1259 -4120 -1257 -4116
rect -1249 -4120 -1247 -4116
rect -1233 -4120 -1231 -4116
rect -1225 -4120 -1223 -4116
rect -1209 -4120 -1207 -4116
rect -1201 -4120 -1199 -4116
rect -1191 -4120 -1189 -4116
rect -1183 -4120 -1181 -4116
rect -1167 -4120 -1165 -4116
rect -1159 -4120 -1157 -4116
rect -1149 -4120 -1147 -4116
rect -1141 -4120 -1139 -4116
rect -1125 -4120 -1123 -4116
rect -1117 -4120 -1115 -4116
rect -1107 -4120 -1105 -4116
rect -1099 -4120 -1097 -4116
rect -1083 -4120 -1081 -4116
rect -1075 -4120 -1073 -4116
rect -930 -4120 -928 -4116
rect -920 -4120 -918 -4116
rect -904 -4120 -902 -4116
rect -896 -4120 -894 -4116
rect -880 -4120 -878 -4116
rect -872 -4120 -870 -4116
rect -862 -4120 -860 -4116
rect -854 -4120 -852 -4116
rect -838 -4120 -836 -4116
rect -830 -4120 -828 -4116
rect -820 -4120 -818 -4116
rect -812 -4120 -810 -4116
rect -796 -4120 -794 -4116
rect -788 -4120 -786 -4116
rect -778 -4120 -776 -4116
rect -770 -4120 -768 -4116
rect -754 -4120 -752 -4116
rect -746 -4120 -744 -4116
rect -572 -4120 -570 -4116
rect -562 -4120 -560 -4116
rect -546 -4120 -544 -4116
rect -538 -4120 -536 -4116
rect -522 -4120 -520 -4116
rect -514 -4120 -512 -4116
rect -504 -4120 -502 -4116
rect -496 -4120 -494 -4116
rect -480 -4120 -478 -4116
rect -472 -4120 -470 -4116
rect -462 -4120 -460 -4116
rect -454 -4120 -452 -4116
rect -438 -4120 -436 -4116
rect -430 -4120 -428 -4116
rect -420 -4120 -418 -4116
rect -412 -4120 -410 -4116
rect -396 -4120 -394 -4116
rect -388 -4120 -386 -4116
rect -214 -4120 -212 -4116
rect -204 -4120 -202 -4116
rect -188 -4120 -186 -4116
rect -180 -4120 -178 -4116
rect -164 -4120 -162 -4116
rect -156 -4120 -154 -4116
rect -146 -4120 -144 -4116
rect -138 -4120 -136 -4116
rect -122 -4120 -120 -4116
rect -114 -4120 -112 -4116
rect -104 -4120 -102 -4116
rect -96 -4120 -94 -4116
rect -80 -4120 -78 -4116
rect -72 -4120 -70 -4116
rect -62 -4120 -60 -4116
rect -54 -4120 -52 -4116
rect -38 -4120 -36 -4116
rect -30 -4120 -28 -4116
rect 214 -4120 216 -4116
rect 224 -4120 226 -4116
rect 240 -4120 242 -4116
rect 248 -4120 250 -4116
rect 264 -4120 266 -4116
rect 272 -4120 274 -4116
rect 282 -4120 284 -4116
rect 290 -4120 292 -4116
rect 306 -4120 308 -4116
rect 314 -4120 316 -4116
rect 324 -4120 326 -4116
rect 332 -4120 334 -4116
rect 348 -4120 350 -4116
rect 356 -4120 358 -4116
rect 366 -4120 368 -4116
rect 374 -4120 376 -4116
rect 390 -4120 392 -4116
rect 398 -4120 400 -4116
rect 570 -4120 572 -4116
rect 580 -4120 582 -4116
rect 596 -4120 598 -4116
rect 604 -4120 606 -4116
rect 620 -4120 622 -4116
rect 628 -4120 630 -4116
rect 638 -4120 640 -4116
rect 646 -4120 648 -4116
rect 662 -4120 664 -4116
rect 670 -4120 672 -4116
rect 680 -4120 682 -4116
rect 688 -4120 690 -4116
rect 704 -4120 706 -4116
rect 712 -4120 714 -4116
rect 722 -4120 724 -4116
rect 730 -4120 732 -4116
rect 746 -4120 748 -4116
rect 754 -4120 756 -4116
rect 968 -4120 970 -4116
rect 978 -4120 980 -4116
rect 994 -4120 996 -4116
rect 1002 -4120 1004 -4116
rect 1018 -4120 1020 -4116
rect 1026 -4120 1028 -4116
rect 1036 -4120 1038 -4116
rect 1044 -4120 1046 -4116
rect 1060 -4120 1062 -4116
rect 1068 -4120 1070 -4116
rect 1078 -4120 1080 -4116
rect 1086 -4120 1088 -4116
rect 1102 -4120 1104 -4116
rect 1110 -4120 1112 -4116
rect 1120 -4120 1122 -4116
rect 1128 -4120 1130 -4116
rect 1144 -4120 1146 -4116
rect 1152 -4120 1154 -4116
rect 1326 -4120 1328 -4116
rect 1336 -4120 1338 -4116
rect 1352 -4120 1354 -4116
rect 1360 -4120 1362 -4116
rect 1376 -4120 1378 -4116
rect 1384 -4120 1386 -4116
rect 1394 -4120 1396 -4116
rect 1402 -4120 1404 -4116
rect 1418 -4120 1420 -4116
rect 1426 -4120 1428 -4116
rect 1436 -4120 1438 -4116
rect 1444 -4120 1446 -4116
rect 1460 -4120 1462 -4116
rect 1468 -4120 1470 -4116
rect 1478 -4120 1480 -4116
rect 1486 -4120 1488 -4116
rect 1502 -4120 1504 -4116
rect 1510 -4120 1512 -4116
rect -1259 -4244 -1257 -4240
rect -1249 -4244 -1247 -4240
rect -1233 -4244 -1231 -4240
rect -1225 -4244 -1223 -4240
rect -1209 -4244 -1207 -4240
rect -1201 -4244 -1199 -4240
rect -1191 -4244 -1189 -4240
rect -1183 -4244 -1181 -4240
rect -1167 -4244 -1165 -4240
rect -1159 -4244 -1157 -4240
rect -1149 -4244 -1147 -4240
rect -1141 -4244 -1139 -4240
rect -1125 -4244 -1123 -4240
rect -1117 -4244 -1115 -4240
rect -1107 -4244 -1105 -4240
rect -1099 -4244 -1097 -4240
rect -1083 -4244 -1081 -4240
rect -1075 -4244 -1073 -4240
rect -1024 -4244 -1022 -4240
rect -930 -4244 -928 -4240
rect -920 -4244 -918 -4240
rect -904 -4244 -902 -4240
rect -896 -4244 -894 -4240
rect -880 -4244 -878 -4240
rect -872 -4244 -870 -4240
rect -862 -4244 -860 -4240
rect -854 -4244 -852 -4240
rect -838 -4244 -836 -4240
rect -830 -4244 -828 -4240
rect -820 -4244 -818 -4240
rect -812 -4244 -810 -4240
rect -796 -4244 -794 -4240
rect -788 -4244 -786 -4240
rect -778 -4244 -776 -4240
rect -770 -4244 -768 -4240
rect -754 -4244 -752 -4240
rect -746 -4244 -744 -4240
rect -572 -4244 -570 -4240
rect -562 -4244 -560 -4240
rect -546 -4244 -544 -4240
rect -538 -4244 -536 -4240
rect -522 -4244 -520 -4240
rect -514 -4244 -512 -4240
rect -504 -4244 -502 -4240
rect -496 -4244 -494 -4240
rect -480 -4244 -478 -4240
rect -472 -4244 -470 -4240
rect -462 -4244 -460 -4240
rect -454 -4244 -452 -4240
rect -438 -4244 -436 -4240
rect -430 -4244 -428 -4240
rect -420 -4244 -418 -4240
rect -412 -4244 -410 -4240
rect -396 -4244 -394 -4240
rect -388 -4244 -386 -4240
rect -327 -4244 -325 -4240
rect -214 -4244 -212 -4240
rect -204 -4244 -202 -4240
rect -188 -4244 -186 -4240
rect -180 -4244 -178 -4240
rect -164 -4244 -162 -4240
rect -156 -4244 -154 -4240
rect -146 -4244 -144 -4240
rect -138 -4244 -136 -4240
rect -122 -4244 -120 -4240
rect -114 -4244 -112 -4240
rect -104 -4244 -102 -4240
rect -96 -4244 -94 -4240
rect -80 -4244 -78 -4240
rect -72 -4244 -70 -4240
rect -62 -4244 -60 -4240
rect -54 -4244 -52 -4240
rect -38 -4244 -36 -4240
rect -30 -4244 -28 -4240
rect 461 -4244 463 -4240
rect 1206 -4244 1208 -4240
rect -1334 -4355 -1332 -4351
rect -1326 -4355 -1324 -4351
rect -1316 -4355 -1314 -4351
rect -1024 -4355 -1022 -4351
rect -930 -4355 -928 -4351
rect -922 -4355 -920 -4351
rect -912 -4355 -910 -4351
rect -668 -4355 -666 -4347
rect -572 -4355 -570 -4351
rect -564 -4355 -562 -4351
rect -554 -4355 -552 -4351
rect -327 -4355 -325 -4351
rect -214 -4355 -212 -4351
rect -206 -4355 -204 -4351
rect -196 -4355 -194 -4351
rect 214 -4355 216 -4351
rect 222 -4355 224 -4351
rect 232 -4355 234 -4351
rect 461 -4355 463 -4351
rect 570 -4355 572 -4351
rect 578 -4355 580 -4351
rect 588 -4355 590 -4351
rect 865 -4355 867 -4347
rect 968 -4355 970 -4351
rect 976 -4355 978 -4351
rect 986 -4355 988 -4351
rect 1206 -4355 1208 -4351
rect 1326 -4355 1328 -4351
rect 1334 -4355 1336 -4351
rect 1344 -4355 1346 -4351
rect -1259 -4474 -1257 -4470
rect -1249 -4474 -1247 -4470
rect -1233 -4474 -1231 -4470
rect -1223 -4474 -1221 -4470
rect -1215 -4474 -1213 -4470
rect -1205 -4474 -1203 -4470
rect -1189 -4474 -1187 -4470
rect -1181 -4474 -1179 -4470
rect -1171 -4474 -1169 -4470
rect -930 -4474 -928 -4470
rect -920 -4474 -918 -4470
rect -904 -4474 -902 -4470
rect -894 -4474 -892 -4470
rect -878 -4474 -876 -4470
rect -868 -4474 -866 -4470
rect -860 -4474 -858 -4470
rect -850 -4474 -848 -4470
rect -834 -4474 -832 -4470
rect -826 -4474 -824 -4470
rect -816 -4474 -814 -4470
rect -800 -4474 -798 -4470
rect -790 -4474 -788 -4470
rect -782 -4474 -780 -4470
rect -772 -4474 -770 -4470
rect -756 -4474 -754 -4470
rect -748 -4474 -746 -4470
rect -732 -4474 -730 -4470
rect -716 -4474 -714 -4470
rect -708 -4474 -706 -4470
rect -698 -4474 -696 -4470
rect -572 -4474 -570 -4470
rect -562 -4474 -560 -4470
rect -546 -4474 -544 -4470
rect -536 -4474 -534 -4470
rect -520 -4474 -518 -4470
rect -510 -4474 -508 -4470
rect -502 -4474 -500 -4470
rect -492 -4474 -490 -4470
rect -476 -4474 -474 -4470
rect -468 -4474 -466 -4470
rect -458 -4474 -456 -4470
rect -442 -4474 -440 -4470
rect -432 -4474 -430 -4470
rect -424 -4474 -422 -4470
rect -414 -4474 -412 -4470
rect -398 -4474 -396 -4470
rect -390 -4474 -388 -4470
rect -374 -4474 -372 -4470
rect -358 -4474 -356 -4470
rect -350 -4474 -348 -4470
rect -340 -4474 -338 -4470
rect -214 -4474 -212 -4470
rect -204 -4474 -202 -4470
rect -188 -4474 -186 -4470
rect -178 -4474 -176 -4470
rect -162 -4474 -160 -4470
rect -152 -4474 -150 -4470
rect -144 -4474 -142 -4470
rect -134 -4474 -132 -4470
rect -118 -4474 -116 -4470
rect -110 -4474 -108 -4470
rect -100 -4474 -98 -4470
rect -84 -4474 -82 -4470
rect -74 -4474 -72 -4470
rect -66 -4474 -64 -4470
rect -56 -4474 -54 -4470
rect -40 -4474 -38 -4470
rect -32 -4474 -30 -4470
rect -16 -4474 -14 -4470
rect 0 -4474 2 -4470
rect 8 -4474 10 -4470
rect 18 -4474 20 -4470
rect 214 -4474 216 -4470
rect 224 -4474 226 -4470
rect 240 -4474 242 -4470
rect 250 -4474 252 -4470
rect 266 -4474 268 -4470
rect 276 -4474 278 -4470
rect 284 -4474 286 -4470
rect 294 -4474 296 -4470
rect 310 -4474 312 -4470
rect 318 -4474 320 -4470
rect 328 -4474 330 -4470
rect 344 -4474 346 -4470
rect 354 -4474 356 -4470
rect 362 -4474 364 -4470
rect 372 -4474 374 -4470
rect 388 -4474 390 -4470
rect 396 -4474 398 -4470
rect 412 -4474 414 -4470
rect 428 -4474 430 -4470
rect 436 -4474 438 -4470
rect 446 -4474 448 -4470
rect 570 -4474 572 -4470
rect 580 -4474 582 -4470
rect 596 -4474 598 -4470
rect 606 -4474 608 -4470
rect 622 -4474 624 -4470
rect 632 -4474 634 -4470
rect 640 -4474 642 -4470
rect 650 -4474 652 -4470
rect 666 -4474 668 -4470
rect 674 -4474 676 -4470
rect 684 -4474 686 -4470
rect 700 -4474 702 -4470
rect 710 -4474 712 -4470
rect 718 -4474 720 -4470
rect 728 -4474 730 -4470
rect 744 -4474 746 -4470
rect 752 -4474 754 -4470
rect 768 -4474 770 -4470
rect 784 -4474 786 -4470
rect 792 -4474 794 -4470
rect 802 -4474 804 -4470
rect 968 -4474 970 -4470
rect 978 -4474 980 -4470
rect 994 -4474 996 -4470
rect 1004 -4474 1006 -4470
rect 1020 -4474 1022 -4470
rect 1030 -4474 1032 -4470
rect 1038 -4474 1040 -4470
rect 1048 -4474 1050 -4470
rect 1064 -4474 1066 -4470
rect 1072 -4474 1074 -4470
rect 1082 -4474 1084 -4470
rect 1098 -4474 1100 -4470
rect 1108 -4474 1110 -4470
rect 1116 -4474 1118 -4470
rect 1126 -4474 1128 -4470
rect 1142 -4474 1144 -4470
rect 1150 -4474 1152 -4470
rect 1166 -4474 1168 -4470
rect 1182 -4474 1184 -4470
rect 1190 -4474 1192 -4470
rect 1200 -4474 1202 -4470
rect 1326 -4474 1328 -4470
rect 1336 -4474 1338 -4470
rect 1352 -4474 1354 -4470
rect 1362 -4474 1364 -4470
rect 1378 -4474 1380 -4470
rect 1388 -4474 1390 -4470
rect 1396 -4474 1398 -4470
rect 1406 -4474 1408 -4470
rect 1422 -4474 1424 -4470
rect 1430 -4474 1432 -4470
rect 1440 -4474 1442 -4470
rect 1456 -4474 1458 -4470
rect 1466 -4474 1468 -4470
rect 1474 -4474 1476 -4470
rect 1484 -4474 1486 -4470
rect 1500 -4474 1502 -4470
rect 1508 -4474 1510 -4470
rect 1524 -4474 1526 -4470
rect 1540 -4474 1542 -4470
rect 1548 -4474 1550 -4470
rect 1558 -4474 1560 -4470
rect -1259 -4597 -1257 -4593
rect -1249 -4597 -1247 -4593
rect -1233 -4597 -1231 -4593
rect -1225 -4597 -1223 -4593
rect -1209 -4597 -1207 -4593
rect -1201 -4597 -1199 -4593
rect -1191 -4597 -1189 -4593
rect -1183 -4597 -1181 -4593
rect -1167 -4597 -1165 -4593
rect -1159 -4597 -1157 -4593
rect -1149 -4597 -1147 -4593
rect -1141 -4597 -1139 -4593
rect -1125 -4597 -1123 -4593
rect -1117 -4597 -1115 -4593
rect -1107 -4597 -1105 -4593
rect -1099 -4597 -1097 -4593
rect -1083 -4597 -1081 -4593
rect -1075 -4597 -1073 -4593
rect -930 -4597 -928 -4593
rect -920 -4597 -918 -4593
rect -904 -4597 -902 -4593
rect -896 -4597 -894 -4593
rect -880 -4597 -878 -4593
rect -872 -4597 -870 -4593
rect -862 -4597 -860 -4593
rect -854 -4597 -852 -4593
rect -838 -4597 -836 -4593
rect -830 -4597 -828 -4593
rect -820 -4597 -818 -4593
rect -812 -4597 -810 -4593
rect -796 -4597 -794 -4593
rect -788 -4597 -786 -4593
rect -778 -4597 -776 -4593
rect -770 -4597 -768 -4593
rect -754 -4597 -752 -4593
rect -746 -4597 -744 -4593
rect -572 -4597 -570 -4593
rect -562 -4597 -560 -4593
rect -546 -4597 -544 -4593
rect -538 -4597 -536 -4593
rect -522 -4597 -520 -4593
rect -514 -4597 -512 -4593
rect -504 -4597 -502 -4593
rect -496 -4597 -494 -4593
rect -480 -4597 -478 -4593
rect -472 -4597 -470 -4593
rect -462 -4597 -460 -4593
rect -454 -4597 -452 -4593
rect -438 -4597 -436 -4593
rect -430 -4597 -428 -4593
rect -420 -4597 -418 -4593
rect -412 -4597 -410 -4593
rect -396 -4597 -394 -4593
rect -388 -4597 -386 -4593
rect -1259 -4718 -1257 -4714
rect -1249 -4718 -1247 -4714
rect -1233 -4718 -1231 -4714
rect -1225 -4718 -1223 -4714
rect -1209 -4718 -1207 -4714
rect -1201 -4718 -1199 -4714
rect -1191 -4718 -1189 -4714
rect -1183 -4718 -1181 -4714
rect -1167 -4718 -1165 -4714
rect -1159 -4718 -1157 -4714
rect -1149 -4718 -1147 -4714
rect -1141 -4718 -1139 -4714
rect -1125 -4718 -1123 -4714
rect -1117 -4718 -1115 -4714
rect -1107 -4718 -1105 -4714
rect -1099 -4718 -1097 -4714
rect -1083 -4718 -1081 -4714
rect -1075 -4718 -1073 -4714
rect -930 -4718 -928 -4714
rect -920 -4718 -918 -4714
rect -904 -4718 -902 -4714
rect -896 -4718 -894 -4714
rect -880 -4718 -878 -4714
rect -872 -4718 -870 -4714
rect -862 -4718 -860 -4714
rect -854 -4718 -852 -4714
rect -838 -4718 -836 -4714
rect -830 -4718 -828 -4714
rect -820 -4718 -818 -4714
rect -812 -4718 -810 -4714
rect -796 -4718 -794 -4714
rect -788 -4718 -786 -4714
rect -778 -4718 -776 -4714
rect -770 -4718 -768 -4714
rect -754 -4718 -752 -4714
rect -746 -4718 -744 -4714
rect -572 -4718 -570 -4714
rect -562 -4718 -560 -4714
rect -546 -4718 -544 -4714
rect -538 -4718 -536 -4714
rect -522 -4718 -520 -4714
rect -514 -4718 -512 -4714
rect -504 -4718 -502 -4714
rect -496 -4718 -494 -4714
rect -480 -4718 -478 -4714
rect -472 -4718 -470 -4714
rect -462 -4718 -460 -4714
rect -454 -4718 -452 -4714
rect -438 -4718 -436 -4714
rect -430 -4718 -428 -4714
rect -420 -4718 -418 -4714
rect -412 -4718 -410 -4714
rect -396 -4718 -394 -4714
rect -388 -4718 -386 -4714
rect -214 -4718 -212 -4714
rect -204 -4718 -202 -4714
rect -188 -4718 -186 -4714
rect -180 -4718 -178 -4714
rect -164 -4718 -162 -4714
rect -156 -4718 -154 -4714
rect -146 -4718 -144 -4714
rect -138 -4718 -136 -4714
rect -122 -4718 -120 -4714
rect -114 -4718 -112 -4714
rect -104 -4718 -102 -4714
rect -96 -4718 -94 -4714
rect -80 -4718 -78 -4714
rect -72 -4718 -70 -4714
rect -62 -4718 -60 -4714
rect -54 -4718 -52 -4714
rect -38 -4718 -36 -4714
rect -30 -4718 -28 -4714
rect 214 -4718 216 -4714
rect 224 -4718 226 -4714
rect 240 -4718 242 -4714
rect 248 -4718 250 -4714
rect 264 -4718 266 -4714
rect 272 -4718 274 -4714
rect 282 -4718 284 -4714
rect 290 -4718 292 -4714
rect 306 -4718 308 -4714
rect 314 -4718 316 -4714
rect 324 -4718 326 -4714
rect 332 -4718 334 -4714
rect 348 -4718 350 -4714
rect 356 -4718 358 -4714
rect 366 -4718 368 -4714
rect 374 -4718 376 -4714
rect 390 -4718 392 -4714
rect 398 -4718 400 -4714
rect 570 -4718 572 -4714
rect 580 -4718 582 -4714
rect 596 -4718 598 -4714
rect 604 -4718 606 -4714
rect 620 -4718 622 -4714
rect 628 -4718 630 -4714
rect 638 -4718 640 -4714
rect 646 -4718 648 -4714
rect 662 -4718 664 -4714
rect 670 -4718 672 -4714
rect 680 -4718 682 -4714
rect 688 -4718 690 -4714
rect 704 -4718 706 -4714
rect 712 -4718 714 -4714
rect 722 -4718 724 -4714
rect 730 -4718 732 -4714
rect 746 -4718 748 -4714
rect 754 -4718 756 -4714
rect 968 -4718 970 -4714
rect 978 -4718 980 -4714
rect 994 -4718 996 -4714
rect 1002 -4718 1004 -4714
rect 1018 -4718 1020 -4714
rect 1026 -4718 1028 -4714
rect 1036 -4718 1038 -4714
rect 1044 -4718 1046 -4714
rect 1060 -4718 1062 -4714
rect 1068 -4718 1070 -4714
rect 1078 -4718 1080 -4714
rect 1086 -4718 1088 -4714
rect 1102 -4718 1104 -4714
rect 1110 -4718 1112 -4714
rect 1120 -4718 1122 -4714
rect 1128 -4718 1130 -4714
rect 1144 -4718 1146 -4714
rect 1152 -4718 1154 -4714
rect 1326 -4718 1328 -4714
rect 1336 -4718 1338 -4714
rect 1352 -4718 1354 -4714
rect 1360 -4718 1362 -4714
rect 1376 -4718 1378 -4714
rect 1384 -4718 1386 -4714
rect 1394 -4718 1396 -4714
rect 1402 -4718 1404 -4714
rect 1418 -4718 1420 -4714
rect 1426 -4718 1428 -4714
rect 1436 -4718 1438 -4714
rect 1444 -4718 1446 -4714
rect 1460 -4718 1462 -4714
rect 1468 -4718 1470 -4714
rect 1478 -4718 1480 -4714
rect 1486 -4718 1488 -4714
rect 1502 -4718 1504 -4714
rect 1510 -4718 1512 -4714
rect -1259 -4839 -1257 -4835
rect -1249 -4839 -1247 -4835
rect -1233 -4839 -1231 -4835
rect -1225 -4839 -1223 -4835
rect -1209 -4839 -1207 -4835
rect -1201 -4839 -1199 -4835
rect -1191 -4839 -1189 -4835
rect -1183 -4839 -1181 -4835
rect -1167 -4839 -1165 -4835
rect -1159 -4839 -1157 -4835
rect -1149 -4839 -1147 -4835
rect -1141 -4839 -1139 -4835
rect -1125 -4839 -1123 -4835
rect -1117 -4839 -1115 -4835
rect -1107 -4839 -1105 -4835
rect -1099 -4839 -1097 -4835
rect -1083 -4839 -1081 -4835
rect -1075 -4839 -1073 -4835
rect -930 -4839 -928 -4835
rect -920 -4839 -918 -4835
rect -904 -4839 -902 -4835
rect -896 -4839 -894 -4835
rect -880 -4839 -878 -4835
rect -872 -4839 -870 -4835
rect -862 -4839 -860 -4835
rect -854 -4839 -852 -4835
rect -838 -4839 -836 -4835
rect -830 -4839 -828 -4835
rect -820 -4839 -818 -4835
rect -812 -4839 -810 -4835
rect -796 -4839 -794 -4835
rect -788 -4839 -786 -4835
rect -778 -4839 -776 -4835
rect -770 -4839 -768 -4835
rect -754 -4839 -752 -4835
rect -746 -4839 -744 -4835
rect -572 -4839 -570 -4835
rect -562 -4839 -560 -4835
rect -546 -4839 -544 -4835
rect -538 -4839 -536 -4835
rect -522 -4839 -520 -4835
rect -514 -4839 -512 -4835
rect -504 -4839 -502 -4835
rect -496 -4839 -494 -4835
rect -480 -4839 -478 -4835
rect -472 -4839 -470 -4835
rect -462 -4839 -460 -4835
rect -454 -4839 -452 -4835
rect -438 -4839 -436 -4835
rect -430 -4839 -428 -4835
rect -420 -4839 -418 -4835
rect -412 -4839 -410 -4835
rect -396 -4839 -394 -4835
rect -388 -4839 -386 -4835
rect -214 -4839 -212 -4835
rect -204 -4839 -202 -4835
rect -188 -4839 -186 -4835
rect -180 -4839 -178 -4835
rect -164 -4839 -162 -4835
rect -156 -4839 -154 -4835
rect -146 -4839 -144 -4835
rect -138 -4839 -136 -4835
rect -122 -4839 -120 -4835
rect -114 -4839 -112 -4835
rect -104 -4839 -102 -4835
rect -96 -4839 -94 -4835
rect -80 -4839 -78 -4835
rect -72 -4839 -70 -4835
rect -62 -4839 -60 -4835
rect -54 -4839 -52 -4835
rect -38 -4839 -36 -4835
rect -30 -4839 -28 -4835
rect 95 -4839 97 -4823
rect 214 -4839 216 -4835
rect 224 -4839 226 -4835
rect 240 -4839 242 -4835
rect 248 -4839 250 -4835
rect 264 -4839 266 -4835
rect 272 -4839 274 -4835
rect 282 -4839 284 -4835
rect 290 -4839 292 -4835
rect 306 -4839 308 -4835
rect 314 -4839 316 -4835
rect 324 -4839 326 -4835
rect 332 -4839 334 -4835
rect 348 -4839 350 -4835
rect 356 -4839 358 -4835
rect 366 -4839 368 -4835
rect 374 -4839 376 -4835
rect 390 -4839 392 -4835
rect 398 -4839 400 -4835
rect 570 -4839 572 -4835
rect 580 -4839 582 -4835
rect 596 -4839 598 -4835
rect 604 -4839 606 -4835
rect 620 -4839 622 -4835
rect 628 -4839 630 -4835
rect 638 -4839 640 -4835
rect 646 -4839 648 -4835
rect 662 -4839 664 -4835
rect 670 -4839 672 -4835
rect 680 -4839 682 -4835
rect 688 -4839 690 -4835
rect 704 -4839 706 -4835
rect 712 -4839 714 -4835
rect 722 -4839 724 -4835
rect 730 -4839 732 -4835
rect 746 -4839 748 -4835
rect 754 -4839 756 -4835
rect 968 -4839 970 -4835
rect 978 -4839 980 -4835
rect 994 -4839 996 -4835
rect 1002 -4839 1004 -4835
rect 1018 -4839 1020 -4835
rect 1026 -4839 1028 -4835
rect 1036 -4839 1038 -4835
rect 1044 -4839 1046 -4835
rect 1060 -4839 1062 -4835
rect 1068 -4839 1070 -4835
rect 1078 -4839 1080 -4835
rect 1086 -4839 1088 -4835
rect 1102 -4839 1104 -4835
rect 1110 -4839 1112 -4835
rect 1120 -4839 1122 -4835
rect 1128 -4839 1130 -4835
rect 1144 -4839 1146 -4835
rect 1152 -4839 1154 -4835
rect 1326 -4839 1328 -4835
rect 1336 -4839 1338 -4835
rect 1352 -4839 1354 -4835
rect 1360 -4839 1362 -4835
rect 1376 -4839 1378 -4835
rect 1384 -4839 1386 -4835
rect 1394 -4839 1396 -4835
rect 1402 -4839 1404 -4835
rect 1418 -4839 1420 -4835
rect 1426 -4839 1428 -4835
rect 1436 -4839 1438 -4835
rect 1444 -4839 1446 -4835
rect 1460 -4839 1462 -4835
rect 1468 -4839 1470 -4835
rect 1478 -4839 1480 -4835
rect 1486 -4839 1488 -4835
rect 1502 -4839 1504 -4835
rect 1510 -4839 1512 -4835
rect -1259 -4957 -1257 -4953
rect -1249 -4957 -1247 -4953
rect -1233 -4957 -1231 -4953
rect -1225 -4957 -1223 -4953
rect -1209 -4957 -1207 -4953
rect -1201 -4957 -1199 -4953
rect -1191 -4957 -1189 -4953
rect -1183 -4957 -1181 -4953
rect -1167 -4957 -1165 -4953
rect -1159 -4957 -1157 -4953
rect -1149 -4957 -1147 -4953
rect -1141 -4957 -1139 -4953
rect -1125 -4957 -1123 -4953
rect -1117 -4957 -1115 -4953
rect -1107 -4957 -1105 -4953
rect -1099 -4957 -1097 -4953
rect -1083 -4957 -1081 -4953
rect -1075 -4957 -1073 -4953
rect -930 -4957 -928 -4953
rect -920 -4957 -918 -4953
rect -904 -4957 -902 -4953
rect -896 -4957 -894 -4953
rect -880 -4957 -878 -4953
rect -872 -4957 -870 -4953
rect -862 -4957 -860 -4953
rect -854 -4957 -852 -4953
rect -838 -4957 -836 -4953
rect -830 -4957 -828 -4953
rect -820 -4957 -818 -4953
rect -812 -4957 -810 -4953
rect -796 -4957 -794 -4953
rect -788 -4957 -786 -4953
rect -778 -4957 -776 -4953
rect -770 -4957 -768 -4953
rect -754 -4957 -752 -4953
rect -746 -4957 -744 -4953
rect -572 -4957 -570 -4953
rect -562 -4957 -560 -4953
rect -546 -4957 -544 -4953
rect -538 -4957 -536 -4953
rect -522 -4957 -520 -4953
rect -514 -4957 -512 -4953
rect -504 -4957 -502 -4953
rect -496 -4957 -494 -4953
rect -480 -4957 -478 -4953
rect -472 -4957 -470 -4953
rect -462 -4957 -460 -4953
rect -454 -4957 -452 -4953
rect -438 -4957 -436 -4953
rect -430 -4957 -428 -4953
rect -420 -4957 -418 -4953
rect -412 -4957 -410 -4953
rect -396 -4957 -394 -4953
rect -388 -4957 -386 -4953
rect -214 -4957 -212 -4953
rect -204 -4957 -202 -4953
rect -188 -4957 -186 -4953
rect -180 -4957 -178 -4953
rect -164 -4957 -162 -4953
rect -156 -4957 -154 -4953
rect -146 -4957 -144 -4953
rect -138 -4957 -136 -4953
rect -122 -4957 -120 -4953
rect -114 -4957 -112 -4953
rect -104 -4957 -102 -4953
rect -96 -4957 -94 -4953
rect -80 -4957 -78 -4953
rect -72 -4957 -70 -4953
rect -62 -4957 -60 -4953
rect -54 -4957 -52 -4953
rect -38 -4957 -36 -4953
rect -30 -4957 -28 -4953
rect 214 -4957 216 -4953
rect 224 -4957 226 -4953
rect 240 -4957 242 -4953
rect 248 -4957 250 -4953
rect 264 -4957 266 -4953
rect 272 -4957 274 -4953
rect 282 -4957 284 -4953
rect 290 -4957 292 -4953
rect 306 -4957 308 -4953
rect 314 -4957 316 -4953
rect 324 -4957 326 -4953
rect 332 -4957 334 -4953
rect 348 -4957 350 -4953
rect 356 -4957 358 -4953
rect 366 -4957 368 -4953
rect 374 -4957 376 -4953
rect 390 -4957 392 -4953
rect 398 -4957 400 -4953
rect -1334 -5074 -1332 -5070
rect -1326 -5074 -1324 -5070
rect -1316 -5074 -1314 -5070
rect -930 -5074 -928 -5070
rect -922 -5074 -920 -5070
rect -912 -5074 -910 -5070
rect -572 -5074 -570 -5070
rect -564 -5074 -562 -5070
rect -554 -5074 -552 -5070
rect -214 -5074 -212 -5070
rect -206 -5074 -204 -5070
rect -196 -5074 -194 -5070
rect 214 -5074 216 -5070
rect 222 -5074 224 -5070
rect 232 -5074 234 -5070
rect 570 -5074 572 -5070
rect 578 -5074 580 -5070
rect 588 -5074 590 -5070
rect 968 -5074 970 -5070
rect 976 -5074 978 -5070
rect 986 -5074 988 -5070
rect 1326 -5074 1328 -5070
rect 1334 -5074 1336 -5070
rect 1344 -5074 1346 -5070
rect -1259 -5193 -1257 -5189
rect -1249 -5193 -1247 -5189
rect -1233 -5193 -1231 -5189
rect -1223 -5193 -1221 -5189
rect -1215 -5193 -1213 -5189
rect -1205 -5193 -1203 -5189
rect -1189 -5193 -1187 -5189
rect -1181 -5193 -1179 -5189
rect -1171 -5193 -1169 -5189
rect -930 -5193 -928 -5189
rect -920 -5193 -918 -5189
rect -904 -5193 -902 -5189
rect -894 -5193 -892 -5189
rect -878 -5193 -876 -5189
rect -868 -5193 -866 -5189
rect -860 -5193 -858 -5189
rect -850 -5193 -848 -5189
rect -834 -5193 -832 -5189
rect -826 -5193 -824 -5189
rect -816 -5193 -814 -5189
rect -800 -5193 -798 -5189
rect -790 -5193 -788 -5189
rect -782 -5193 -780 -5189
rect -772 -5193 -770 -5189
rect -756 -5193 -754 -5189
rect -748 -5193 -746 -5189
rect -732 -5193 -730 -5189
rect -716 -5193 -714 -5189
rect -708 -5193 -706 -5189
rect -698 -5193 -696 -5189
rect -572 -5193 -570 -5189
rect -562 -5193 -560 -5189
rect -546 -5193 -544 -5189
rect -536 -5193 -534 -5189
rect -520 -5193 -518 -5189
rect -510 -5193 -508 -5189
rect -502 -5193 -500 -5189
rect -492 -5193 -490 -5189
rect -476 -5193 -474 -5189
rect -468 -5193 -466 -5189
rect -458 -5193 -456 -5189
rect -442 -5193 -440 -5189
rect -432 -5193 -430 -5189
rect -424 -5193 -422 -5189
rect -414 -5193 -412 -5189
rect -398 -5193 -396 -5189
rect -390 -5193 -388 -5189
rect -374 -5193 -372 -5189
rect -358 -5193 -356 -5189
rect -350 -5193 -348 -5189
rect -340 -5193 -338 -5189
rect -214 -5193 -212 -5189
rect -204 -5193 -202 -5189
rect -188 -5193 -186 -5189
rect -178 -5193 -176 -5189
rect -162 -5193 -160 -5189
rect -152 -5193 -150 -5189
rect -144 -5193 -142 -5189
rect -134 -5193 -132 -5189
rect -118 -5193 -116 -5189
rect -110 -5193 -108 -5189
rect -100 -5193 -98 -5189
rect -84 -5193 -82 -5189
rect -74 -5193 -72 -5189
rect -66 -5193 -64 -5189
rect -56 -5193 -54 -5189
rect -40 -5193 -38 -5189
rect -32 -5193 -30 -5189
rect -16 -5193 -14 -5189
rect 0 -5193 2 -5189
rect 8 -5193 10 -5189
rect 18 -5193 20 -5189
rect 214 -5193 216 -5189
rect 224 -5193 226 -5189
rect 240 -5193 242 -5189
rect 250 -5193 252 -5189
rect 266 -5193 268 -5189
rect 276 -5193 278 -5189
rect 284 -5193 286 -5189
rect 294 -5193 296 -5189
rect 310 -5193 312 -5189
rect 318 -5193 320 -5189
rect 328 -5193 330 -5189
rect 344 -5193 346 -5189
rect 354 -5193 356 -5189
rect 362 -5193 364 -5189
rect 372 -5193 374 -5189
rect 388 -5193 390 -5189
rect 396 -5193 398 -5189
rect 412 -5193 414 -5189
rect 428 -5193 430 -5189
rect 436 -5193 438 -5189
rect 446 -5193 448 -5189
rect 570 -5193 572 -5189
rect 580 -5193 582 -5189
rect 596 -5193 598 -5189
rect 606 -5193 608 -5189
rect 622 -5193 624 -5189
rect 632 -5193 634 -5189
rect 640 -5193 642 -5189
rect 650 -5193 652 -5189
rect 666 -5193 668 -5189
rect 674 -5193 676 -5189
rect 684 -5193 686 -5189
rect 700 -5193 702 -5189
rect 710 -5193 712 -5189
rect 718 -5193 720 -5189
rect 728 -5193 730 -5189
rect 744 -5193 746 -5189
rect 752 -5193 754 -5189
rect 768 -5193 770 -5189
rect 784 -5193 786 -5189
rect 792 -5193 794 -5189
rect 802 -5193 804 -5189
rect 968 -5193 970 -5189
rect 978 -5193 980 -5189
rect 994 -5193 996 -5189
rect 1004 -5193 1006 -5189
rect 1020 -5193 1022 -5189
rect 1030 -5193 1032 -5189
rect 1038 -5193 1040 -5189
rect 1048 -5193 1050 -5189
rect 1064 -5193 1066 -5189
rect 1072 -5193 1074 -5189
rect 1082 -5193 1084 -5189
rect 1098 -5193 1100 -5189
rect 1108 -5193 1110 -5189
rect 1116 -5193 1118 -5189
rect 1126 -5193 1128 -5189
rect 1142 -5193 1144 -5189
rect 1150 -5193 1152 -5189
rect 1166 -5193 1168 -5189
rect 1182 -5193 1184 -5189
rect 1190 -5193 1192 -5189
rect 1200 -5193 1202 -5189
rect 1326 -5193 1328 -5189
rect 1336 -5193 1338 -5189
rect 1352 -5193 1354 -5189
rect 1362 -5193 1364 -5189
rect 1378 -5193 1380 -5189
rect 1388 -5193 1390 -5189
rect 1396 -5193 1398 -5189
rect 1406 -5193 1408 -5189
rect 1422 -5193 1424 -5189
rect 1430 -5193 1432 -5189
rect 1440 -5193 1442 -5189
rect 1456 -5193 1458 -5189
rect 1466 -5193 1468 -5189
rect 1474 -5193 1476 -5189
rect 1484 -5193 1486 -5189
rect 1500 -5193 1502 -5189
rect 1508 -5193 1510 -5189
rect 1524 -5193 1526 -5189
rect 1540 -5193 1542 -5189
rect 1548 -5193 1550 -5189
rect 1558 -5193 1560 -5189
rect -1259 -5312 -1257 -5308
rect -1249 -5312 -1247 -5308
rect -1233 -5312 -1231 -5308
rect -1225 -5312 -1223 -5308
rect -1209 -5312 -1207 -5308
rect -1201 -5312 -1199 -5308
rect -1191 -5312 -1189 -5308
rect -1183 -5312 -1181 -5308
rect -1167 -5312 -1165 -5308
rect -1159 -5312 -1157 -5308
rect -1149 -5312 -1147 -5308
rect -1141 -5312 -1139 -5308
rect -1125 -5312 -1123 -5308
rect -1117 -5312 -1115 -5308
rect -1107 -5312 -1105 -5308
rect -1099 -5312 -1097 -5308
rect -1083 -5312 -1081 -5308
rect -1075 -5312 -1073 -5308
rect -930 -5312 -928 -5308
rect -920 -5312 -918 -5308
rect -904 -5312 -902 -5308
rect -896 -5312 -894 -5308
rect -880 -5312 -878 -5308
rect -872 -5312 -870 -5308
rect -862 -5312 -860 -5308
rect -854 -5312 -852 -5308
rect -838 -5312 -836 -5308
rect -830 -5312 -828 -5308
rect -820 -5312 -818 -5308
rect -812 -5312 -810 -5308
rect -796 -5312 -794 -5308
rect -788 -5312 -786 -5308
rect -778 -5312 -776 -5308
rect -770 -5312 -768 -5308
rect -754 -5312 -752 -5308
rect -746 -5312 -744 -5308
rect -1259 -5433 -1257 -5429
rect -1249 -5433 -1247 -5429
rect -1233 -5433 -1231 -5429
rect -1225 -5433 -1223 -5429
rect -1209 -5433 -1207 -5429
rect -1201 -5433 -1199 -5429
rect -1191 -5433 -1189 -5429
rect -1183 -5433 -1181 -5429
rect -1167 -5433 -1165 -5429
rect -1159 -5433 -1157 -5429
rect -1149 -5433 -1147 -5429
rect -1141 -5433 -1139 -5429
rect -1125 -5433 -1123 -5429
rect -1117 -5433 -1115 -5429
rect -1107 -5433 -1105 -5429
rect -1099 -5433 -1097 -5429
rect -1083 -5433 -1081 -5429
rect -1075 -5433 -1073 -5429
rect -1021 -5433 -1019 -5429
rect -930 -5433 -928 -5429
rect -920 -5433 -918 -5429
rect -904 -5433 -902 -5429
rect -896 -5433 -894 -5429
rect -880 -5433 -878 -5429
rect -872 -5433 -870 -5429
rect -862 -5433 -860 -5429
rect -854 -5433 -852 -5429
rect -838 -5433 -836 -5429
rect -830 -5433 -828 -5429
rect -820 -5433 -818 -5429
rect -812 -5433 -810 -5429
rect -796 -5433 -794 -5429
rect -788 -5433 -786 -5429
rect -778 -5433 -776 -5429
rect -770 -5433 -768 -5429
rect -754 -5433 -752 -5429
rect -746 -5433 -744 -5429
rect -668 -5433 -666 -5425
rect -572 -5433 -570 -5429
rect -562 -5433 -560 -5429
rect -546 -5433 -544 -5429
rect -538 -5433 -536 -5429
rect -522 -5433 -520 -5429
rect -514 -5433 -512 -5429
rect -504 -5433 -502 -5429
rect -496 -5433 -494 -5429
rect -480 -5433 -478 -5429
rect -472 -5433 -470 -5429
rect -462 -5433 -460 -5429
rect -454 -5433 -452 -5429
rect -438 -5433 -436 -5429
rect -430 -5433 -428 -5429
rect -420 -5433 -418 -5429
rect -412 -5433 -410 -5429
rect -396 -5433 -394 -5429
rect -388 -5433 -386 -5429
rect -322 -5433 -320 -5429
rect -214 -5433 -212 -5429
rect -204 -5433 -202 -5429
rect -188 -5433 -186 -5429
rect -180 -5433 -178 -5429
rect -164 -5433 -162 -5429
rect -156 -5433 -154 -5429
rect -146 -5433 -144 -5429
rect -138 -5433 -136 -5429
rect -122 -5433 -120 -5429
rect -114 -5433 -112 -5429
rect -104 -5433 -102 -5429
rect -96 -5433 -94 -5429
rect -80 -5433 -78 -5429
rect -72 -5433 -70 -5429
rect -62 -5433 -60 -5429
rect -54 -5433 -52 -5429
rect -38 -5433 -36 -5429
rect -30 -5433 -28 -5429
rect 214 -5433 216 -5429
rect 224 -5433 226 -5429
rect 240 -5433 242 -5429
rect 248 -5433 250 -5429
rect 264 -5433 266 -5429
rect 272 -5433 274 -5429
rect 282 -5433 284 -5429
rect 290 -5433 292 -5429
rect 306 -5433 308 -5429
rect 314 -5433 316 -5429
rect 324 -5433 326 -5429
rect 332 -5433 334 -5429
rect 348 -5433 350 -5429
rect 356 -5433 358 -5429
rect 366 -5433 368 -5429
rect 374 -5433 376 -5429
rect 390 -5433 392 -5429
rect 398 -5433 400 -5429
rect 471 -5433 473 -5429
rect 570 -5433 572 -5429
rect 580 -5433 582 -5429
rect 596 -5433 598 -5429
rect 604 -5433 606 -5429
rect 620 -5433 622 -5429
rect 628 -5433 630 -5429
rect 638 -5433 640 -5429
rect 646 -5433 648 -5429
rect 662 -5433 664 -5429
rect 670 -5433 672 -5429
rect 680 -5433 682 -5429
rect 688 -5433 690 -5429
rect 704 -5433 706 -5429
rect 712 -5433 714 -5429
rect 722 -5433 724 -5429
rect 730 -5433 732 -5429
rect 746 -5433 748 -5429
rect 754 -5433 756 -5429
rect 872 -5433 874 -5425
rect 968 -5433 970 -5429
rect 978 -5433 980 -5429
rect 994 -5433 996 -5429
rect 1002 -5433 1004 -5429
rect 1018 -5433 1020 -5429
rect 1026 -5433 1028 -5429
rect 1036 -5433 1038 -5429
rect 1044 -5433 1046 -5429
rect 1060 -5433 1062 -5429
rect 1068 -5433 1070 -5429
rect 1078 -5433 1080 -5429
rect 1086 -5433 1088 -5429
rect 1102 -5433 1104 -5429
rect 1110 -5433 1112 -5429
rect 1120 -5433 1122 -5429
rect 1128 -5433 1130 -5429
rect 1144 -5433 1146 -5429
rect 1152 -5433 1154 -5429
rect 1215 -5433 1217 -5429
rect 1326 -5433 1328 -5429
rect 1336 -5433 1338 -5429
rect 1352 -5433 1354 -5429
rect 1360 -5433 1362 -5429
rect 1376 -5433 1378 -5429
rect 1384 -5433 1386 -5429
rect 1394 -5433 1396 -5429
rect 1402 -5433 1404 -5429
rect 1418 -5433 1420 -5429
rect 1426 -5433 1428 -5429
rect 1436 -5433 1438 -5429
rect 1444 -5433 1446 -5429
rect 1460 -5433 1462 -5429
rect 1468 -5433 1470 -5429
rect 1478 -5433 1480 -5429
rect 1486 -5433 1488 -5429
rect 1502 -5433 1504 -5429
rect 1510 -5433 1512 -5429
rect -1259 -5553 -1257 -5549
rect -1249 -5553 -1247 -5549
rect -1233 -5553 -1231 -5549
rect -1225 -5553 -1223 -5549
rect -1209 -5553 -1207 -5549
rect -1201 -5553 -1199 -5549
rect -1191 -5553 -1189 -5549
rect -1183 -5553 -1181 -5549
rect -1167 -5553 -1165 -5549
rect -1159 -5553 -1157 -5549
rect -1149 -5553 -1147 -5549
rect -1141 -5553 -1139 -5549
rect -1125 -5553 -1123 -5549
rect -1117 -5553 -1115 -5549
rect -1107 -5553 -1105 -5549
rect -1099 -5553 -1097 -5549
rect -1083 -5553 -1081 -5549
rect -1075 -5553 -1073 -5549
rect -1021 -5553 -1019 -5549
rect -930 -5553 -928 -5549
rect -920 -5553 -918 -5549
rect -904 -5553 -902 -5549
rect -896 -5553 -894 -5549
rect -880 -5553 -878 -5549
rect -872 -5553 -870 -5549
rect -862 -5553 -860 -5549
rect -854 -5553 -852 -5549
rect -838 -5553 -836 -5549
rect -830 -5553 -828 -5549
rect -820 -5553 -818 -5549
rect -812 -5553 -810 -5549
rect -796 -5553 -794 -5549
rect -788 -5553 -786 -5549
rect -778 -5553 -776 -5549
rect -770 -5553 -768 -5549
rect -754 -5553 -752 -5549
rect -746 -5553 -744 -5549
rect -572 -5553 -570 -5549
rect -562 -5553 -560 -5549
rect -546 -5553 -544 -5549
rect -538 -5553 -536 -5549
rect -522 -5553 -520 -5549
rect -514 -5553 -512 -5549
rect -504 -5553 -502 -5549
rect -496 -5553 -494 -5549
rect -480 -5553 -478 -5549
rect -472 -5553 -470 -5549
rect -462 -5553 -460 -5549
rect -454 -5553 -452 -5549
rect -438 -5553 -436 -5549
rect -430 -5553 -428 -5549
rect -420 -5553 -418 -5549
rect -412 -5553 -410 -5549
rect -396 -5553 -394 -5549
rect -388 -5553 -386 -5549
rect -322 -5553 -320 -5549
rect -214 -5553 -212 -5549
rect -204 -5553 -202 -5549
rect -188 -5553 -186 -5549
rect -180 -5553 -178 -5549
rect -164 -5553 -162 -5549
rect -156 -5553 -154 -5549
rect -146 -5553 -144 -5549
rect -138 -5553 -136 -5549
rect -122 -5553 -120 -5549
rect -114 -5553 -112 -5549
rect -104 -5553 -102 -5549
rect -96 -5553 -94 -5549
rect -80 -5553 -78 -5549
rect -72 -5553 -70 -5549
rect -62 -5553 -60 -5549
rect -54 -5553 -52 -5549
rect -38 -5553 -36 -5549
rect -30 -5553 -28 -5549
rect 214 -5553 216 -5549
rect 224 -5553 226 -5549
rect 240 -5553 242 -5549
rect 248 -5553 250 -5549
rect 264 -5553 266 -5549
rect 272 -5553 274 -5549
rect 282 -5553 284 -5549
rect 290 -5553 292 -5549
rect 306 -5553 308 -5549
rect 314 -5553 316 -5549
rect 324 -5553 326 -5549
rect 332 -5553 334 -5549
rect 348 -5553 350 -5549
rect 356 -5553 358 -5549
rect 366 -5553 368 -5549
rect 374 -5553 376 -5549
rect 390 -5553 392 -5549
rect 398 -5553 400 -5549
rect 471 -5553 473 -5549
rect 570 -5553 572 -5549
rect 580 -5553 582 -5549
rect 596 -5553 598 -5549
rect 604 -5553 606 -5549
rect 620 -5553 622 -5549
rect 628 -5553 630 -5549
rect 638 -5553 640 -5549
rect 646 -5553 648 -5549
rect 662 -5553 664 -5549
rect 670 -5553 672 -5549
rect 680 -5553 682 -5549
rect 688 -5553 690 -5549
rect 704 -5553 706 -5549
rect 712 -5553 714 -5549
rect 722 -5553 724 -5549
rect 730 -5553 732 -5549
rect 746 -5553 748 -5549
rect 754 -5553 756 -5549
rect 968 -5553 970 -5549
rect 978 -5553 980 -5549
rect 994 -5553 996 -5549
rect 1002 -5553 1004 -5549
rect 1018 -5553 1020 -5549
rect 1026 -5553 1028 -5549
rect 1036 -5553 1038 -5549
rect 1044 -5553 1046 -5549
rect 1060 -5553 1062 -5549
rect 1068 -5553 1070 -5549
rect 1078 -5553 1080 -5549
rect 1086 -5553 1088 -5549
rect 1102 -5553 1104 -5549
rect 1110 -5553 1112 -5549
rect 1120 -5553 1122 -5549
rect 1128 -5553 1130 -5549
rect 1144 -5553 1146 -5549
rect 1152 -5553 1154 -5549
rect 1215 -5553 1217 -5549
rect 1326 -5553 1328 -5549
rect 1336 -5553 1338 -5549
rect 1352 -5553 1354 -5549
rect 1360 -5553 1362 -5549
rect 1376 -5553 1378 -5549
rect 1384 -5553 1386 -5549
rect 1394 -5553 1396 -5549
rect 1402 -5553 1404 -5549
rect 1418 -5553 1420 -5549
rect 1426 -5553 1428 -5549
rect 1436 -5553 1438 -5549
rect 1444 -5553 1446 -5549
rect 1460 -5553 1462 -5549
rect 1468 -5553 1470 -5549
rect 1478 -5553 1480 -5549
rect 1486 -5553 1488 -5549
rect 1502 -5553 1504 -5549
rect 1510 -5553 1512 -5549
rect -1259 -5670 -1257 -5666
rect -1249 -5670 -1247 -5666
rect -1233 -5670 -1231 -5666
rect -1225 -5670 -1223 -5666
rect -1209 -5670 -1207 -5666
rect -1201 -5670 -1199 -5666
rect -1191 -5670 -1189 -5666
rect -1183 -5670 -1181 -5666
rect -1167 -5670 -1165 -5666
rect -1159 -5670 -1157 -5666
rect -1149 -5670 -1147 -5666
rect -1141 -5670 -1139 -5666
rect -1125 -5670 -1123 -5666
rect -1117 -5670 -1115 -5666
rect -1107 -5670 -1105 -5666
rect -1099 -5670 -1097 -5666
rect -1083 -5670 -1081 -5666
rect -1075 -5670 -1073 -5666
rect -930 -5670 -928 -5666
rect -920 -5670 -918 -5666
rect -904 -5670 -902 -5666
rect -896 -5670 -894 -5666
rect -880 -5670 -878 -5666
rect -872 -5670 -870 -5666
rect -862 -5670 -860 -5666
rect -854 -5670 -852 -5666
rect -838 -5670 -836 -5666
rect -830 -5670 -828 -5666
rect -820 -5670 -818 -5666
rect -812 -5670 -810 -5666
rect -796 -5670 -794 -5666
rect -788 -5670 -786 -5666
rect -778 -5670 -776 -5666
rect -770 -5670 -768 -5666
rect -754 -5670 -752 -5666
rect -746 -5670 -744 -5666
rect -572 -5670 -570 -5666
rect -562 -5670 -560 -5666
rect -546 -5670 -544 -5666
rect -538 -5670 -536 -5666
rect -522 -5670 -520 -5666
rect -514 -5670 -512 -5666
rect -504 -5670 -502 -5666
rect -496 -5670 -494 -5666
rect -480 -5670 -478 -5666
rect -472 -5670 -470 -5666
rect -462 -5670 -460 -5666
rect -454 -5670 -452 -5666
rect -438 -5670 -436 -5666
rect -430 -5670 -428 -5666
rect -420 -5670 -418 -5666
rect -412 -5670 -410 -5666
rect -396 -5670 -394 -5666
rect -388 -5670 -386 -5666
rect -214 -5670 -212 -5666
rect -204 -5670 -202 -5666
rect -188 -5670 -186 -5666
rect -180 -5670 -178 -5666
rect -164 -5670 -162 -5666
rect -156 -5670 -154 -5666
rect -146 -5670 -144 -5666
rect -138 -5670 -136 -5666
rect -122 -5670 -120 -5666
rect -114 -5670 -112 -5666
rect -104 -5670 -102 -5666
rect -96 -5670 -94 -5666
rect -80 -5670 -78 -5666
rect -72 -5670 -70 -5666
rect -62 -5670 -60 -5666
rect -54 -5670 -52 -5666
rect -38 -5670 -36 -5666
rect -30 -5670 -28 -5666
rect 214 -5670 216 -5666
rect 224 -5670 226 -5666
rect 240 -5670 242 -5666
rect 248 -5670 250 -5666
rect 264 -5670 266 -5666
rect 272 -5670 274 -5666
rect 282 -5670 284 -5666
rect 290 -5670 292 -5666
rect 306 -5670 308 -5666
rect 314 -5670 316 -5666
rect 324 -5670 326 -5666
rect 332 -5670 334 -5666
rect 348 -5670 350 -5666
rect 356 -5670 358 -5666
rect 366 -5670 368 -5666
rect 374 -5670 376 -5666
rect 390 -5670 392 -5666
rect 398 -5670 400 -5666
rect 570 -5670 572 -5666
rect 580 -5670 582 -5666
rect 596 -5670 598 -5666
rect 604 -5670 606 -5666
rect 620 -5670 622 -5666
rect 628 -5670 630 -5666
rect 638 -5670 640 -5666
rect 646 -5670 648 -5666
rect 662 -5670 664 -5666
rect 670 -5670 672 -5666
rect 680 -5670 682 -5666
rect 688 -5670 690 -5666
rect 704 -5670 706 -5666
rect 712 -5670 714 -5666
rect 722 -5670 724 -5666
rect 730 -5670 732 -5666
rect 746 -5670 748 -5666
rect 754 -5670 756 -5666
rect -1334 -5787 -1332 -5783
rect -1326 -5787 -1324 -5783
rect -1316 -5787 -1314 -5783
rect -930 -5787 -928 -5783
rect -922 -5787 -920 -5783
rect -912 -5787 -910 -5783
rect -572 -5787 -570 -5783
rect -564 -5787 -562 -5783
rect -554 -5787 -552 -5783
rect -214 -5787 -212 -5783
rect -206 -5787 -204 -5783
rect -196 -5787 -194 -5783
rect 214 -5787 216 -5783
rect 222 -5787 224 -5783
rect 232 -5787 234 -5783
rect 570 -5787 572 -5783
rect 578 -5787 580 -5783
rect 588 -5787 590 -5783
rect 968 -5787 970 -5783
rect 976 -5787 978 -5783
rect 986 -5787 988 -5783
rect 1326 -5787 1328 -5783
rect 1334 -5787 1336 -5783
rect 1344 -5787 1346 -5783
rect -1259 -5906 -1257 -5902
rect -1249 -5906 -1247 -5902
rect -1233 -5906 -1231 -5902
rect -1223 -5906 -1221 -5902
rect -1215 -5906 -1213 -5902
rect -1205 -5906 -1203 -5902
rect -1189 -5906 -1187 -5902
rect -1181 -5906 -1179 -5902
rect -1171 -5906 -1169 -5902
rect -930 -5906 -928 -5902
rect -920 -5906 -918 -5902
rect -904 -5906 -902 -5902
rect -894 -5906 -892 -5902
rect -878 -5906 -876 -5902
rect -868 -5906 -866 -5902
rect -860 -5906 -858 -5902
rect -850 -5906 -848 -5902
rect -834 -5906 -832 -5902
rect -826 -5906 -824 -5902
rect -816 -5906 -814 -5902
rect -800 -5906 -798 -5902
rect -790 -5906 -788 -5902
rect -782 -5906 -780 -5902
rect -772 -5906 -770 -5902
rect -756 -5906 -754 -5902
rect -748 -5906 -746 -5902
rect -732 -5906 -730 -5902
rect -716 -5906 -714 -5902
rect -708 -5906 -706 -5902
rect -698 -5906 -696 -5902
rect -572 -5906 -570 -5902
rect -562 -5906 -560 -5902
rect -546 -5906 -544 -5902
rect -536 -5906 -534 -5902
rect -520 -5906 -518 -5902
rect -510 -5906 -508 -5902
rect -502 -5906 -500 -5902
rect -492 -5906 -490 -5902
rect -476 -5906 -474 -5902
rect -468 -5906 -466 -5902
rect -458 -5906 -456 -5902
rect -442 -5906 -440 -5902
rect -432 -5906 -430 -5902
rect -424 -5906 -422 -5902
rect -414 -5906 -412 -5902
rect -398 -5906 -396 -5902
rect -390 -5906 -388 -5902
rect -374 -5906 -372 -5902
rect -358 -5906 -356 -5902
rect -350 -5906 -348 -5902
rect -340 -5906 -338 -5902
rect -214 -5906 -212 -5902
rect -204 -5906 -202 -5902
rect -188 -5906 -186 -5902
rect -178 -5906 -176 -5902
rect -162 -5906 -160 -5902
rect -152 -5906 -150 -5902
rect -144 -5906 -142 -5902
rect -134 -5906 -132 -5902
rect -118 -5906 -116 -5902
rect -110 -5906 -108 -5902
rect -100 -5906 -98 -5902
rect -84 -5906 -82 -5902
rect -74 -5906 -72 -5902
rect -66 -5906 -64 -5902
rect -56 -5906 -54 -5902
rect -40 -5906 -38 -5902
rect -32 -5906 -30 -5902
rect -16 -5906 -14 -5902
rect 0 -5906 2 -5902
rect 8 -5906 10 -5902
rect 18 -5906 20 -5902
rect 214 -5906 216 -5902
rect 224 -5906 226 -5902
rect 240 -5906 242 -5902
rect 250 -5906 252 -5902
rect 266 -5906 268 -5902
rect 276 -5906 278 -5902
rect 284 -5906 286 -5902
rect 294 -5906 296 -5902
rect 310 -5906 312 -5902
rect 318 -5906 320 -5902
rect 328 -5906 330 -5902
rect 344 -5906 346 -5902
rect 354 -5906 356 -5902
rect 362 -5906 364 -5902
rect 372 -5906 374 -5902
rect 388 -5906 390 -5902
rect 396 -5906 398 -5902
rect 412 -5906 414 -5902
rect 428 -5906 430 -5902
rect 436 -5906 438 -5902
rect 446 -5906 448 -5902
rect 570 -5906 572 -5902
rect 580 -5906 582 -5902
rect 596 -5906 598 -5902
rect 606 -5906 608 -5902
rect 622 -5906 624 -5902
rect 632 -5906 634 -5902
rect 640 -5906 642 -5902
rect 650 -5906 652 -5902
rect 666 -5906 668 -5902
rect 674 -5906 676 -5902
rect 684 -5906 686 -5902
rect 700 -5906 702 -5902
rect 710 -5906 712 -5902
rect 718 -5906 720 -5902
rect 728 -5906 730 -5902
rect 744 -5906 746 -5902
rect 752 -5906 754 -5902
rect 768 -5906 770 -5902
rect 784 -5906 786 -5902
rect 792 -5906 794 -5902
rect 802 -5906 804 -5902
rect 968 -5906 970 -5902
rect 978 -5906 980 -5902
rect 994 -5906 996 -5902
rect 1004 -5906 1006 -5902
rect 1020 -5906 1022 -5902
rect 1030 -5906 1032 -5902
rect 1038 -5906 1040 -5902
rect 1048 -5906 1050 -5902
rect 1064 -5906 1066 -5902
rect 1072 -5906 1074 -5902
rect 1082 -5906 1084 -5902
rect 1098 -5906 1100 -5902
rect 1108 -5906 1110 -5902
rect 1116 -5906 1118 -5902
rect 1126 -5906 1128 -5902
rect 1142 -5906 1144 -5902
rect 1150 -5906 1152 -5902
rect 1166 -5906 1168 -5902
rect 1182 -5906 1184 -5902
rect 1190 -5906 1192 -5902
rect 1200 -5906 1202 -5902
rect 1326 -5906 1328 -5902
rect 1336 -5906 1338 -5902
rect 1352 -5906 1354 -5902
rect 1362 -5906 1364 -5902
rect 1378 -5906 1380 -5902
rect 1388 -5906 1390 -5902
rect 1396 -5906 1398 -5902
rect 1406 -5906 1408 -5902
rect 1422 -5906 1424 -5902
rect 1430 -5906 1432 -5902
rect 1440 -5906 1442 -5902
rect 1456 -5906 1458 -5902
rect 1466 -5906 1468 -5902
rect 1474 -5906 1476 -5902
rect 1484 -5906 1486 -5902
rect 1500 -5906 1502 -5902
rect 1508 -5906 1510 -5902
rect 1524 -5906 1526 -5902
rect 1540 -5906 1542 -5902
rect 1548 -5906 1550 -5902
rect 1558 -5906 1560 -5902
rect -1259 -6029 -1257 -6025
rect -1249 -6029 -1247 -6025
rect -1233 -6029 -1231 -6025
rect -1225 -6029 -1223 -6025
rect -1209 -6029 -1207 -6025
rect -1201 -6029 -1199 -6025
rect -1191 -6029 -1189 -6025
rect -1183 -6029 -1181 -6025
rect -1167 -6029 -1165 -6025
rect -1159 -6029 -1157 -6025
rect -1149 -6029 -1147 -6025
rect -1141 -6029 -1139 -6025
rect -1125 -6029 -1123 -6025
rect -1117 -6029 -1115 -6025
rect -1107 -6029 -1105 -6025
rect -1099 -6029 -1097 -6025
rect -1083 -6029 -1081 -6025
rect -1075 -6029 -1073 -6025
rect -930 -6029 -928 -6025
rect -920 -6029 -918 -6025
rect -904 -6029 -902 -6025
rect -896 -6029 -894 -6025
rect -880 -6029 -878 -6025
rect -872 -6029 -870 -6025
rect -862 -6029 -860 -6025
rect -854 -6029 -852 -6025
rect -838 -6029 -836 -6025
rect -830 -6029 -828 -6025
rect -820 -6029 -818 -6025
rect -812 -6029 -810 -6025
rect -796 -6029 -794 -6025
rect -788 -6029 -786 -6025
rect -778 -6029 -776 -6025
rect -770 -6029 -768 -6025
rect -754 -6029 -752 -6025
rect -746 -6029 -744 -6025
rect -572 -6029 -570 -6025
rect -562 -6029 -560 -6025
rect -546 -6029 -544 -6025
rect -538 -6029 -536 -6025
rect -522 -6029 -520 -6025
rect -514 -6029 -512 -6025
rect -504 -6029 -502 -6025
rect -496 -6029 -494 -6025
rect -480 -6029 -478 -6025
rect -472 -6029 -470 -6025
rect -462 -6029 -460 -6025
rect -454 -6029 -452 -6025
rect -438 -6029 -436 -6025
rect -430 -6029 -428 -6025
rect -420 -6029 -418 -6025
rect -412 -6029 -410 -6025
rect -396 -6029 -394 -6025
rect -388 -6029 -386 -6025
rect -214 -6029 -212 -6025
rect -204 -6029 -202 -6025
rect -188 -6029 -186 -6025
rect -180 -6029 -178 -6025
rect -164 -6029 -162 -6025
rect -156 -6029 -154 -6025
rect -146 -6029 -144 -6025
rect -138 -6029 -136 -6025
rect -122 -6029 -120 -6025
rect -114 -6029 -112 -6025
rect -104 -6029 -102 -6025
rect -96 -6029 -94 -6025
rect -80 -6029 -78 -6025
rect -72 -6029 -70 -6025
rect -62 -6029 -60 -6025
rect -54 -6029 -52 -6025
rect -38 -6029 -36 -6025
rect -30 -6029 -28 -6025
rect 214 -6029 216 -6025
rect 224 -6029 226 -6025
rect 240 -6029 242 -6025
rect 248 -6029 250 -6025
rect 264 -6029 266 -6025
rect 272 -6029 274 -6025
rect 282 -6029 284 -6025
rect 290 -6029 292 -6025
rect 306 -6029 308 -6025
rect 314 -6029 316 -6025
rect 324 -6029 326 -6025
rect 332 -6029 334 -6025
rect 348 -6029 350 -6025
rect 356 -6029 358 -6025
rect 366 -6029 368 -6025
rect 374 -6029 376 -6025
rect 390 -6029 392 -6025
rect 398 -6029 400 -6025
rect 570 -6029 572 -6025
rect 580 -6029 582 -6025
rect 596 -6029 598 -6025
rect 604 -6029 606 -6025
rect 620 -6029 622 -6025
rect 628 -6029 630 -6025
rect 638 -6029 640 -6025
rect 646 -6029 648 -6025
rect 662 -6029 664 -6025
rect 670 -6029 672 -6025
rect 680 -6029 682 -6025
rect 688 -6029 690 -6025
rect 704 -6029 706 -6025
rect 712 -6029 714 -6025
rect 722 -6029 724 -6025
rect 730 -6029 732 -6025
rect 746 -6029 748 -6025
rect 754 -6029 756 -6025
rect 968 -6029 970 -6025
rect 978 -6029 980 -6025
rect 994 -6029 996 -6025
rect 1002 -6029 1004 -6025
rect 1018 -6029 1020 -6025
rect 1026 -6029 1028 -6025
rect 1036 -6029 1038 -6025
rect 1044 -6029 1046 -6025
rect 1060 -6029 1062 -6025
rect 1068 -6029 1070 -6025
rect 1078 -6029 1080 -6025
rect 1086 -6029 1088 -6025
rect 1102 -6029 1104 -6025
rect 1110 -6029 1112 -6025
rect 1120 -6029 1122 -6025
rect 1128 -6029 1130 -6025
rect 1144 -6029 1146 -6025
rect 1152 -6029 1154 -6025
rect 1326 -6029 1328 -6025
rect 1336 -6029 1338 -6025
rect 1352 -6029 1354 -6025
rect 1360 -6029 1362 -6025
rect 1376 -6029 1378 -6025
rect 1384 -6029 1386 -6025
rect 1394 -6029 1396 -6025
rect 1402 -6029 1404 -6025
rect 1418 -6029 1420 -6025
rect 1426 -6029 1428 -6025
rect 1436 -6029 1438 -6025
rect 1444 -6029 1446 -6025
rect 1460 -6029 1462 -6025
rect 1468 -6029 1470 -6025
rect 1478 -6029 1480 -6025
rect 1486 -6029 1488 -6025
rect 1502 -6029 1504 -6025
rect 1510 -6029 1512 -6025
rect 1326 -6147 1328 -6143
rect 1336 -6147 1338 -6143
rect 1352 -6147 1354 -6143
rect 1360 -6147 1362 -6143
rect 1376 -6147 1378 -6143
rect 1384 -6147 1386 -6143
rect 1394 -6147 1396 -6143
rect 1402 -6147 1404 -6143
rect 1418 -6147 1420 -6143
rect 1426 -6147 1428 -6143
rect 1436 -6147 1438 -6143
rect 1444 -6147 1446 -6143
rect 1460 -6147 1462 -6143
rect 1468 -6147 1470 -6143
rect 1478 -6147 1480 -6143
rect 1486 -6147 1488 -6143
rect 1502 -6147 1504 -6143
rect 1510 -6147 1512 -6143
<< ptransistor >>
rect -1332 -1046 -1330 -1038
rect -1324 -1046 -1322 -1038
rect -1314 -1046 -1312 -1038
rect -931 -1046 -929 -1038
rect -923 -1046 -921 -1038
rect -913 -1046 -911 -1038
rect -572 -1046 -570 -1038
rect -564 -1046 -562 -1038
rect -554 -1046 -552 -1038
rect -214 -1046 -212 -1038
rect -206 -1046 -204 -1038
rect -196 -1046 -194 -1038
rect 214 -1046 216 -1038
rect 222 -1046 224 -1038
rect 232 -1046 234 -1038
rect 570 -1046 572 -1038
rect 578 -1046 580 -1038
rect 588 -1046 590 -1038
rect 968 -1046 970 -1038
rect 976 -1046 978 -1038
rect 986 -1046 988 -1038
rect 1326 -1046 1328 -1038
rect 1334 -1046 1336 -1038
rect 1344 -1046 1346 -1038
rect -1255 -1160 -1253 -1152
rect -1245 -1160 -1243 -1152
rect -1229 -1160 -1227 -1152
rect -1221 -1160 -1219 -1152
rect -1205 -1160 -1203 -1152
rect -1197 -1160 -1195 -1152
rect -1187 -1160 -1185 -1152
rect -1179 -1160 -1177 -1152
rect -1163 -1160 -1161 -1152
rect -1155 -1160 -1153 -1152
rect -1145 -1160 -1143 -1152
rect -1137 -1160 -1135 -1152
rect -1121 -1160 -1119 -1152
rect -1113 -1160 -1111 -1152
rect -1103 -1160 -1101 -1152
rect -1095 -1160 -1093 -1152
rect -1079 -1160 -1077 -1152
rect -1071 -1160 -1069 -1152
rect -930 -1160 -928 -1152
rect -920 -1160 -918 -1152
rect -904 -1160 -902 -1152
rect -896 -1160 -894 -1152
rect -880 -1160 -878 -1152
rect -872 -1160 -870 -1152
rect -862 -1160 -860 -1152
rect -854 -1160 -852 -1152
rect -838 -1160 -836 -1152
rect -830 -1160 -828 -1152
rect -820 -1160 -818 -1152
rect -812 -1160 -810 -1152
rect -796 -1160 -794 -1152
rect -788 -1160 -786 -1152
rect -778 -1160 -776 -1152
rect -770 -1160 -768 -1152
rect -754 -1160 -752 -1152
rect -746 -1160 -744 -1152
rect -572 -1160 -570 -1152
rect -562 -1160 -560 -1152
rect -546 -1160 -544 -1152
rect -538 -1160 -536 -1152
rect -522 -1160 -520 -1152
rect -514 -1160 -512 -1152
rect -504 -1160 -502 -1152
rect -496 -1160 -494 -1152
rect -480 -1160 -478 -1152
rect -472 -1160 -470 -1152
rect -462 -1160 -460 -1152
rect -454 -1160 -452 -1152
rect -438 -1160 -436 -1152
rect -430 -1160 -428 -1152
rect -420 -1160 -418 -1152
rect -412 -1160 -410 -1152
rect -396 -1160 -394 -1152
rect -388 -1160 -386 -1152
rect -214 -1160 -212 -1152
rect -204 -1160 -202 -1152
rect -188 -1160 -186 -1152
rect -180 -1160 -178 -1152
rect -164 -1160 -162 -1152
rect -156 -1160 -154 -1152
rect -146 -1160 -144 -1152
rect -138 -1160 -136 -1152
rect -122 -1160 -120 -1152
rect -114 -1160 -112 -1152
rect -104 -1160 -102 -1152
rect -96 -1160 -94 -1152
rect -80 -1160 -78 -1152
rect -72 -1160 -70 -1152
rect -62 -1160 -60 -1152
rect -54 -1160 -52 -1152
rect -38 -1160 -36 -1152
rect -30 -1160 -28 -1152
rect 214 -1160 216 -1152
rect 224 -1160 226 -1152
rect 240 -1160 242 -1152
rect 248 -1160 250 -1152
rect 264 -1160 266 -1152
rect 272 -1160 274 -1152
rect 282 -1160 284 -1152
rect 290 -1160 292 -1152
rect 306 -1160 308 -1152
rect 314 -1160 316 -1152
rect 324 -1160 326 -1152
rect 332 -1160 334 -1152
rect 348 -1160 350 -1152
rect 356 -1160 358 -1152
rect 366 -1160 368 -1152
rect 374 -1160 376 -1152
rect 390 -1160 392 -1152
rect 398 -1160 400 -1152
rect 570 -1160 572 -1152
rect 580 -1160 582 -1152
rect 596 -1160 598 -1152
rect 604 -1160 606 -1152
rect 620 -1160 622 -1152
rect 628 -1160 630 -1152
rect 638 -1160 640 -1152
rect 646 -1160 648 -1152
rect 662 -1160 664 -1152
rect 670 -1160 672 -1152
rect 680 -1160 682 -1152
rect 688 -1160 690 -1152
rect 704 -1160 706 -1152
rect 712 -1160 714 -1152
rect 722 -1160 724 -1152
rect 730 -1160 732 -1152
rect 746 -1160 748 -1152
rect 754 -1160 756 -1152
rect 968 -1160 970 -1152
rect 978 -1160 980 -1152
rect 994 -1160 996 -1152
rect 1002 -1160 1004 -1152
rect 1018 -1160 1020 -1152
rect 1026 -1160 1028 -1152
rect 1036 -1160 1038 -1152
rect 1044 -1160 1046 -1152
rect 1060 -1160 1062 -1152
rect 1068 -1160 1070 -1152
rect 1078 -1160 1080 -1152
rect 1086 -1160 1088 -1152
rect 1102 -1160 1104 -1152
rect 1110 -1160 1112 -1152
rect 1120 -1160 1122 -1152
rect 1128 -1160 1130 -1152
rect 1144 -1160 1146 -1152
rect 1152 -1160 1154 -1152
rect -1334 -1276 -1332 -1268
rect -1326 -1276 -1324 -1268
rect -1316 -1276 -1314 -1268
rect -930 -1276 -928 -1268
rect -922 -1276 -920 -1268
rect -912 -1276 -910 -1268
rect -572 -1276 -570 -1268
rect -564 -1276 -562 -1268
rect -554 -1276 -552 -1268
rect -214 -1276 -212 -1268
rect -206 -1276 -204 -1268
rect -196 -1276 -194 -1268
rect 214 -1276 216 -1268
rect 222 -1276 224 -1268
rect 232 -1276 234 -1268
rect 570 -1276 572 -1268
rect 578 -1276 580 -1268
rect 588 -1276 590 -1268
rect 968 -1276 970 -1268
rect 976 -1276 978 -1268
rect 986 -1276 988 -1268
rect 1326 -1276 1328 -1268
rect 1334 -1276 1336 -1268
rect 1344 -1276 1346 -1268
rect -1255 -1390 -1253 -1382
rect -1245 -1390 -1243 -1382
rect -1229 -1390 -1227 -1382
rect -1219 -1390 -1217 -1382
rect -1211 -1390 -1209 -1382
rect -1201 -1390 -1199 -1382
rect -1185 -1390 -1183 -1382
rect -1177 -1390 -1175 -1382
rect -1167 -1390 -1165 -1382
rect -930 -1390 -928 -1382
rect -920 -1390 -918 -1382
rect -904 -1390 -902 -1382
rect -894 -1390 -892 -1382
rect -878 -1390 -876 -1382
rect -868 -1390 -866 -1382
rect -860 -1390 -858 -1382
rect -850 -1390 -848 -1382
rect -834 -1390 -832 -1382
rect -826 -1390 -824 -1382
rect -816 -1390 -814 -1382
rect -800 -1390 -798 -1382
rect -790 -1390 -788 -1382
rect -782 -1390 -780 -1382
rect -772 -1390 -770 -1382
rect -756 -1390 -754 -1382
rect -748 -1390 -746 -1382
rect -732 -1390 -730 -1382
rect -716 -1390 -714 -1382
rect -708 -1390 -706 -1382
rect -698 -1390 -696 -1382
rect -572 -1390 -570 -1382
rect -562 -1390 -560 -1382
rect -546 -1390 -544 -1382
rect -536 -1390 -534 -1382
rect -520 -1390 -518 -1382
rect -510 -1390 -508 -1382
rect -502 -1390 -500 -1382
rect -492 -1390 -490 -1382
rect -476 -1390 -474 -1382
rect -468 -1390 -466 -1382
rect -458 -1390 -456 -1382
rect -442 -1390 -440 -1382
rect -432 -1390 -430 -1382
rect -424 -1390 -422 -1382
rect -414 -1390 -412 -1382
rect -398 -1390 -396 -1382
rect -390 -1390 -388 -1382
rect -374 -1390 -372 -1382
rect -358 -1390 -356 -1382
rect -350 -1390 -348 -1382
rect -340 -1390 -338 -1382
rect -214 -1390 -212 -1382
rect -204 -1390 -202 -1382
rect -188 -1390 -186 -1382
rect -178 -1390 -176 -1382
rect -162 -1390 -160 -1382
rect -152 -1390 -150 -1382
rect -144 -1390 -142 -1382
rect -134 -1390 -132 -1382
rect -118 -1390 -116 -1382
rect -110 -1390 -108 -1382
rect -100 -1390 -98 -1382
rect -84 -1390 -82 -1382
rect -74 -1390 -72 -1382
rect -66 -1390 -64 -1382
rect -56 -1390 -54 -1382
rect -40 -1390 -38 -1382
rect -32 -1390 -30 -1382
rect -16 -1390 -14 -1382
rect 0 -1390 2 -1382
rect 8 -1390 10 -1382
rect 18 -1390 20 -1382
rect 214 -1390 216 -1382
rect 224 -1390 226 -1382
rect 240 -1390 242 -1382
rect 250 -1390 252 -1382
rect 266 -1390 268 -1382
rect 276 -1390 278 -1382
rect 284 -1390 286 -1382
rect 294 -1390 296 -1382
rect 310 -1390 312 -1382
rect 318 -1390 320 -1382
rect 328 -1390 330 -1382
rect 344 -1390 346 -1382
rect 354 -1390 356 -1382
rect 362 -1390 364 -1382
rect 372 -1390 374 -1382
rect 388 -1390 390 -1382
rect 396 -1390 398 -1382
rect 412 -1390 414 -1382
rect 428 -1390 430 -1382
rect 436 -1390 438 -1382
rect 446 -1390 448 -1382
rect 570 -1390 572 -1382
rect 580 -1390 582 -1382
rect 596 -1390 598 -1382
rect 606 -1390 608 -1382
rect 622 -1390 624 -1382
rect 632 -1390 634 -1382
rect 640 -1390 642 -1382
rect 650 -1390 652 -1382
rect 666 -1390 668 -1382
rect 674 -1390 676 -1382
rect 684 -1390 686 -1382
rect 700 -1390 702 -1382
rect 710 -1390 712 -1382
rect 718 -1390 720 -1382
rect 728 -1390 730 -1382
rect 744 -1390 746 -1382
rect 752 -1390 754 -1382
rect 768 -1390 770 -1382
rect 784 -1390 786 -1382
rect 792 -1390 794 -1382
rect 802 -1390 804 -1382
rect 968 -1390 970 -1382
rect 978 -1390 980 -1382
rect 994 -1390 996 -1382
rect 1004 -1390 1006 -1382
rect 1020 -1390 1022 -1382
rect 1030 -1390 1032 -1382
rect 1038 -1390 1040 -1382
rect 1048 -1390 1050 -1382
rect 1064 -1390 1066 -1382
rect 1072 -1390 1074 -1382
rect 1082 -1390 1084 -1382
rect 1098 -1390 1100 -1382
rect 1108 -1390 1110 -1382
rect 1116 -1390 1118 -1382
rect 1126 -1390 1128 -1382
rect 1142 -1390 1144 -1382
rect 1150 -1390 1152 -1382
rect 1166 -1390 1168 -1382
rect 1182 -1390 1184 -1382
rect 1190 -1390 1192 -1382
rect 1200 -1390 1202 -1382
rect 1326 -1390 1328 -1382
rect 1336 -1390 1338 -1382
rect 1352 -1390 1354 -1382
rect 1362 -1390 1364 -1382
rect 1370 -1390 1372 -1382
rect 1380 -1390 1382 -1382
rect 1396 -1390 1398 -1382
rect 1404 -1390 1406 -1382
rect 1414 -1390 1416 -1382
rect -1255 -1513 -1253 -1505
rect -1245 -1513 -1243 -1505
rect -1229 -1513 -1227 -1505
rect -1221 -1513 -1219 -1505
rect -1205 -1513 -1203 -1505
rect -1197 -1513 -1195 -1505
rect -1187 -1513 -1185 -1505
rect -1179 -1513 -1177 -1505
rect -1163 -1513 -1161 -1505
rect -1155 -1513 -1153 -1505
rect -1145 -1513 -1143 -1505
rect -1137 -1513 -1135 -1505
rect -1121 -1513 -1119 -1505
rect -1113 -1513 -1111 -1505
rect -1103 -1513 -1101 -1505
rect -1095 -1513 -1093 -1505
rect -1079 -1513 -1077 -1505
rect -1071 -1513 -1069 -1505
rect -930 -1513 -928 -1505
rect -920 -1513 -918 -1505
rect -904 -1513 -902 -1505
rect -896 -1513 -894 -1505
rect -880 -1513 -878 -1505
rect -872 -1513 -870 -1505
rect -862 -1513 -860 -1505
rect -854 -1513 -852 -1505
rect -838 -1513 -836 -1505
rect -830 -1513 -828 -1505
rect -820 -1513 -818 -1505
rect -812 -1513 -810 -1505
rect -796 -1513 -794 -1505
rect -788 -1513 -786 -1505
rect -778 -1513 -776 -1505
rect -770 -1513 -768 -1505
rect -754 -1513 -752 -1505
rect -746 -1513 -744 -1505
rect -572 -1513 -570 -1505
rect -562 -1513 -560 -1505
rect -546 -1513 -544 -1505
rect -538 -1513 -536 -1505
rect -522 -1513 -520 -1505
rect -514 -1513 -512 -1505
rect -504 -1513 -502 -1505
rect -496 -1513 -494 -1505
rect -480 -1513 -478 -1505
rect -472 -1513 -470 -1505
rect -462 -1513 -460 -1505
rect -454 -1513 -452 -1505
rect -438 -1513 -436 -1505
rect -430 -1513 -428 -1505
rect -420 -1513 -418 -1505
rect -412 -1513 -410 -1505
rect -396 -1513 -394 -1505
rect -388 -1513 -386 -1505
rect -214 -1513 -212 -1505
rect -204 -1513 -202 -1505
rect -188 -1513 -186 -1505
rect -180 -1513 -178 -1505
rect -164 -1513 -162 -1505
rect -156 -1513 -154 -1505
rect -146 -1513 -144 -1505
rect -138 -1513 -136 -1505
rect -122 -1513 -120 -1505
rect -114 -1513 -112 -1505
rect -104 -1513 -102 -1505
rect -96 -1513 -94 -1505
rect -80 -1513 -78 -1505
rect -72 -1513 -70 -1505
rect -62 -1513 -60 -1505
rect -54 -1513 -52 -1505
rect -38 -1513 -36 -1505
rect -30 -1513 -28 -1505
rect 214 -1513 216 -1505
rect 224 -1513 226 -1505
rect 240 -1513 242 -1505
rect 248 -1513 250 -1505
rect 264 -1513 266 -1505
rect 272 -1513 274 -1505
rect 282 -1513 284 -1505
rect 290 -1513 292 -1505
rect 306 -1513 308 -1505
rect 314 -1513 316 -1505
rect 324 -1513 326 -1505
rect 332 -1513 334 -1505
rect 348 -1513 350 -1505
rect 356 -1513 358 -1505
rect 366 -1513 368 -1505
rect 374 -1513 376 -1505
rect 390 -1513 392 -1505
rect 398 -1513 400 -1505
rect 570 -1513 572 -1505
rect 580 -1513 582 -1505
rect 596 -1513 598 -1505
rect 604 -1513 606 -1505
rect 620 -1513 622 -1505
rect 628 -1513 630 -1505
rect 638 -1513 640 -1505
rect 646 -1513 648 -1505
rect 662 -1513 664 -1505
rect 670 -1513 672 -1505
rect 680 -1513 682 -1505
rect 688 -1513 690 -1505
rect 704 -1513 706 -1505
rect 712 -1513 714 -1505
rect 722 -1513 724 -1505
rect 730 -1513 732 -1505
rect 746 -1513 748 -1505
rect 754 -1513 756 -1505
rect 968 -1513 970 -1505
rect 978 -1513 980 -1505
rect 994 -1513 996 -1505
rect 1002 -1513 1004 -1505
rect 1018 -1513 1020 -1505
rect 1026 -1513 1028 -1505
rect 1036 -1513 1038 -1505
rect 1044 -1513 1046 -1505
rect 1060 -1513 1062 -1505
rect 1068 -1513 1070 -1505
rect 1078 -1513 1080 -1505
rect 1086 -1513 1088 -1505
rect 1102 -1513 1104 -1505
rect 1110 -1513 1112 -1505
rect 1120 -1513 1122 -1505
rect 1128 -1513 1130 -1505
rect 1144 -1513 1146 -1505
rect 1152 -1513 1154 -1505
rect -1255 -1634 -1253 -1626
rect -1245 -1634 -1243 -1626
rect -1229 -1634 -1227 -1626
rect -1221 -1634 -1219 -1626
rect -1205 -1634 -1203 -1626
rect -1197 -1634 -1195 -1626
rect -1187 -1634 -1185 -1626
rect -1179 -1634 -1177 -1626
rect -1163 -1634 -1161 -1626
rect -1155 -1634 -1153 -1626
rect -1145 -1634 -1143 -1626
rect -1137 -1634 -1135 -1626
rect -1121 -1634 -1119 -1626
rect -1113 -1634 -1111 -1626
rect -1103 -1634 -1101 -1626
rect -1095 -1634 -1093 -1626
rect -1079 -1634 -1077 -1626
rect -1071 -1634 -1069 -1626
rect -930 -1634 -928 -1626
rect -920 -1634 -918 -1626
rect -904 -1634 -902 -1626
rect -896 -1634 -894 -1626
rect -880 -1634 -878 -1626
rect -872 -1634 -870 -1626
rect -862 -1634 -860 -1626
rect -854 -1634 -852 -1626
rect -838 -1634 -836 -1626
rect -830 -1634 -828 -1626
rect -820 -1634 -818 -1626
rect -812 -1634 -810 -1626
rect -796 -1634 -794 -1626
rect -788 -1634 -786 -1626
rect -778 -1634 -776 -1626
rect -770 -1634 -768 -1626
rect -754 -1634 -752 -1626
rect -746 -1634 -744 -1626
rect -572 -1634 -570 -1626
rect -562 -1634 -560 -1626
rect -546 -1634 -544 -1626
rect -538 -1634 -536 -1626
rect -522 -1634 -520 -1626
rect -514 -1634 -512 -1626
rect -504 -1634 -502 -1626
rect -496 -1634 -494 -1626
rect -480 -1634 -478 -1626
rect -472 -1634 -470 -1626
rect -462 -1634 -460 -1626
rect -454 -1634 -452 -1626
rect -438 -1634 -436 -1626
rect -430 -1634 -428 -1626
rect -420 -1634 -418 -1626
rect -412 -1634 -410 -1626
rect -396 -1634 -394 -1626
rect -388 -1634 -386 -1626
rect -214 -1634 -212 -1626
rect -204 -1634 -202 -1626
rect -188 -1634 -186 -1626
rect -180 -1634 -178 -1626
rect -164 -1634 -162 -1626
rect -156 -1634 -154 -1626
rect -146 -1634 -144 -1626
rect -138 -1634 -136 -1626
rect -122 -1634 -120 -1626
rect -114 -1634 -112 -1626
rect -104 -1634 -102 -1626
rect -96 -1634 -94 -1626
rect -80 -1634 -78 -1626
rect -72 -1634 -70 -1626
rect -62 -1634 -60 -1626
rect -54 -1634 -52 -1626
rect -38 -1634 -36 -1626
rect -30 -1634 -28 -1626
rect 214 -1634 216 -1626
rect 224 -1634 226 -1626
rect 240 -1634 242 -1626
rect 248 -1634 250 -1626
rect 264 -1634 266 -1626
rect 272 -1634 274 -1626
rect 282 -1634 284 -1626
rect 290 -1634 292 -1626
rect 306 -1634 308 -1626
rect 314 -1634 316 -1626
rect 324 -1634 326 -1626
rect 332 -1634 334 -1626
rect 348 -1634 350 -1626
rect 356 -1634 358 -1626
rect 366 -1634 368 -1626
rect 374 -1634 376 -1626
rect 390 -1634 392 -1626
rect 398 -1634 400 -1626
rect 570 -1634 572 -1626
rect 580 -1634 582 -1626
rect 596 -1634 598 -1626
rect 604 -1634 606 -1626
rect 620 -1634 622 -1626
rect 628 -1634 630 -1626
rect 638 -1634 640 -1626
rect 646 -1634 648 -1626
rect 662 -1634 664 -1626
rect 670 -1634 672 -1626
rect 680 -1634 682 -1626
rect 688 -1634 690 -1626
rect 704 -1634 706 -1626
rect 712 -1634 714 -1626
rect 722 -1634 724 -1626
rect 730 -1634 732 -1626
rect 746 -1634 748 -1626
rect 754 -1634 756 -1626
rect 968 -1634 970 -1626
rect 978 -1634 980 -1626
rect 994 -1634 996 -1626
rect 1002 -1634 1004 -1626
rect 1018 -1634 1020 -1626
rect 1026 -1634 1028 -1626
rect 1036 -1634 1038 -1626
rect 1044 -1634 1046 -1626
rect 1060 -1634 1062 -1626
rect 1068 -1634 1070 -1626
rect 1078 -1634 1080 -1626
rect 1086 -1634 1088 -1626
rect 1102 -1634 1104 -1626
rect 1110 -1634 1112 -1626
rect 1120 -1634 1122 -1626
rect 1128 -1634 1130 -1626
rect 1144 -1634 1146 -1626
rect 1152 -1634 1154 -1626
rect 1326 -1634 1328 -1626
rect 1336 -1634 1338 -1626
rect 1352 -1634 1354 -1626
rect 1360 -1634 1362 -1626
rect 1376 -1634 1378 -1626
rect 1384 -1634 1386 -1626
rect 1394 -1634 1396 -1626
rect 1402 -1634 1404 -1626
rect 1418 -1634 1420 -1626
rect 1426 -1634 1428 -1626
rect 1436 -1634 1438 -1626
rect 1444 -1634 1446 -1626
rect 1460 -1634 1462 -1626
rect 1468 -1634 1470 -1626
rect 1478 -1634 1480 -1626
rect 1486 -1634 1488 -1626
rect 1502 -1634 1504 -1626
rect 1510 -1634 1512 -1626
rect -1255 -1755 -1253 -1747
rect -1245 -1755 -1243 -1747
rect -1229 -1755 -1227 -1747
rect -1221 -1755 -1219 -1747
rect -1205 -1755 -1203 -1747
rect -1197 -1755 -1195 -1747
rect -1187 -1755 -1185 -1747
rect -1179 -1755 -1177 -1747
rect -1163 -1755 -1161 -1747
rect -1155 -1755 -1153 -1747
rect -1145 -1755 -1143 -1747
rect -1137 -1755 -1135 -1747
rect -1121 -1755 -1119 -1747
rect -1113 -1755 -1111 -1747
rect -1103 -1755 -1101 -1747
rect -1095 -1755 -1093 -1747
rect -1079 -1755 -1077 -1747
rect -1071 -1755 -1069 -1747
rect -1024 -1755 -1022 -1747
rect -930 -1755 -928 -1747
rect -920 -1755 -918 -1747
rect -904 -1755 -902 -1747
rect -896 -1755 -894 -1747
rect -880 -1755 -878 -1747
rect -872 -1755 -870 -1747
rect -862 -1755 -860 -1747
rect -854 -1755 -852 -1747
rect -838 -1755 -836 -1747
rect -830 -1755 -828 -1747
rect -820 -1755 -818 -1747
rect -812 -1755 -810 -1747
rect -796 -1755 -794 -1747
rect -788 -1755 -786 -1747
rect -778 -1755 -776 -1747
rect -770 -1755 -768 -1747
rect -754 -1755 -752 -1747
rect -746 -1755 -744 -1747
rect -572 -1755 -570 -1747
rect -562 -1755 -560 -1747
rect -546 -1755 -544 -1747
rect -538 -1755 -536 -1747
rect -522 -1755 -520 -1747
rect -514 -1755 -512 -1747
rect -504 -1755 -502 -1747
rect -496 -1755 -494 -1747
rect -480 -1755 -478 -1747
rect -472 -1755 -470 -1747
rect -462 -1755 -460 -1747
rect -454 -1755 -452 -1747
rect -438 -1755 -436 -1747
rect -430 -1755 -428 -1747
rect -420 -1755 -418 -1747
rect -412 -1755 -410 -1747
rect -396 -1755 -394 -1747
rect -388 -1755 -386 -1747
rect -327 -1755 -325 -1747
rect -214 -1755 -212 -1747
rect -204 -1755 -202 -1747
rect -188 -1755 -186 -1747
rect -180 -1755 -178 -1747
rect -164 -1755 -162 -1747
rect -156 -1755 -154 -1747
rect -146 -1755 -144 -1747
rect -138 -1755 -136 -1747
rect -122 -1755 -120 -1747
rect -114 -1755 -112 -1747
rect -104 -1755 -102 -1747
rect -96 -1755 -94 -1747
rect -80 -1755 -78 -1747
rect -72 -1755 -70 -1747
rect -62 -1755 -60 -1747
rect -54 -1755 -52 -1747
rect -38 -1755 -36 -1747
rect -30 -1755 -28 -1747
rect 214 -1755 216 -1747
rect 224 -1755 226 -1747
rect 240 -1755 242 -1747
rect 248 -1755 250 -1747
rect 264 -1755 266 -1747
rect 272 -1755 274 -1747
rect 282 -1755 284 -1747
rect 290 -1755 292 -1747
rect 306 -1755 308 -1747
rect 314 -1755 316 -1747
rect 324 -1755 326 -1747
rect 332 -1755 334 -1747
rect 348 -1755 350 -1747
rect 356 -1755 358 -1747
rect 366 -1755 368 -1747
rect 374 -1755 376 -1747
rect 390 -1755 392 -1747
rect 398 -1755 400 -1747
rect 469 -1755 471 -1747
rect 570 -1755 572 -1747
rect 580 -1755 582 -1747
rect 596 -1755 598 -1747
rect 604 -1755 606 -1747
rect 620 -1755 622 -1747
rect 628 -1755 630 -1747
rect 638 -1755 640 -1747
rect 646 -1755 648 -1747
rect 662 -1755 664 -1747
rect 670 -1755 672 -1747
rect 680 -1755 682 -1747
rect 688 -1755 690 -1747
rect 704 -1755 706 -1747
rect 712 -1755 714 -1747
rect 722 -1755 724 -1747
rect 730 -1755 732 -1747
rect 746 -1755 748 -1747
rect 754 -1755 756 -1747
rect 968 -1755 970 -1747
rect 978 -1755 980 -1747
rect 994 -1755 996 -1747
rect 1002 -1755 1004 -1747
rect 1018 -1755 1020 -1747
rect 1026 -1755 1028 -1747
rect 1036 -1755 1038 -1747
rect 1044 -1755 1046 -1747
rect 1060 -1755 1062 -1747
rect 1068 -1755 1070 -1747
rect 1078 -1755 1080 -1747
rect 1086 -1755 1088 -1747
rect 1102 -1755 1104 -1747
rect 1110 -1755 1112 -1747
rect 1120 -1755 1122 -1747
rect 1128 -1755 1130 -1747
rect 1144 -1755 1146 -1747
rect 1152 -1755 1154 -1747
rect 1208 -1755 1210 -1747
rect 1326 -1755 1328 -1747
rect 1336 -1755 1338 -1747
rect 1352 -1755 1354 -1747
rect 1360 -1755 1362 -1747
rect 1376 -1755 1378 -1747
rect 1384 -1755 1386 -1747
rect 1394 -1755 1396 -1747
rect 1402 -1755 1404 -1747
rect 1418 -1755 1420 -1747
rect 1426 -1755 1428 -1747
rect 1436 -1755 1438 -1747
rect 1444 -1755 1446 -1747
rect 1460 -1755 1462 -1747
rect 1468 -1755 1470 -1747
rect 1478 -1755 1480 -1747
rect 1486 -1755 1488 -1747
rect 1502 -1755 1504 -1747
rect 1510 -1755 1512 -1747
rect -1255 -1870 -1253 -1862
rect -1245 -1870 -1243 -1862
rect -1229 -1870 -1227 -1862
rect -1221 -1870 -1219 -1862
rect -1205 -1870 -1203 -1862
rect -1197 -1870 -1195 -1862
rect -1187 -1870 -1185 -1862
rect -1179 -1870 -1177 -1862
rect -1163 -1870 -1161 -1862
rect -1155 -1870 -1153 -1862
rect -1145 -1870 -1143 -1862
rect -1137 -1870 -1135 -1862
rect -1121 -1870 -1119 -1862
rect -1113 -1870 -1111 -1862
rect -1103 -1870 -1101 -1862
rect -1095 -1870 -1093 -1862
rect -1079 -1870 -1077 -1862
rect -1071 -1870 -1069 -1862
rect -1024 -1870 -1022 -1862
rect -668 -1878 -666 -1862
rect -327 -1870 -325 -1862
rect 469 -1870 471 -1862
rect 846 -1878 848 -1862
rect 1208 -1870 1210 -1862
rect -1334 -1982 -1332 -1974
rect -1326 -1982 -1324 -1974
rect -1316 -1982 -1314 -1974
rect -930 -1982 -928 -1974
rect -922 -1982 -920 -1974
rect -912 -1982 -910 -1974
rect -572 -1982 -570 -1974
rect -564 -1982 -562 -1974
rect -554 -1982 -552 -1974
rect -214 -1982 -212 -1974
rect -206 -1982 -204 -1974
rect -196 -1982 -194 -1974
rect 214 -1982 216 -1974
rect 222 -1982 224 -1974
rect 232 -1982 234 -1974
rect 570 -1982 572 -1974
rect 578 -1982 580 -1974
rect 588 -1982 590 -1974
rect 968 -1982 970 -1974
rect 976 -1982 978 -1974
rect 986 -1982 988 -1974
rect 1326 -1982 1328 -1974
rect 1334 -1982 1336 -1974
rect 1344 -1982 1346 -1974
rect -1255 -2101 -1253 -2093
rect -1245 -2101 -1243 -2093
rect -1229 -2101 -1227 -2093
rect -1219 -2101 -1217 -2093
rect -1211 -2101 -1209 -2093
rect -1201 -2101 -1199 -2093
rect -1185 -2101 -1183 -2093
rect -1177 -2101 -1175 -2093
rect -1167 -2101 -1165 -2093
rect -930 -2101 -928 -2093
rect -920 -2101 -918 -2093
rect -904 -2101 -902 -2093
rect -894 -2101 -892 -2093
rect -878 -2101 -876 -2093
rect -868 -2101 -866 -2093
rect -860 -2101 -858 -2093
rect -850 -2101 -848 -2093
rect -834 -2101 -832 -2093
rect -826 -2101 -824 -2093
rect -816 -2101 -814 -2093
rect -800 -2101 -798 -2093
rect -790 -2101 -788 -2093
rect -782 -2101 -780 -2093
rect -772 -2101 -770 -2093
rect -756 -2101 -754 -2093
rect -748 -2101 -746 -2093
rect -732 -2101 -730 -2093
rect -716 -2101 -714 -2093
rect -708 -2101 -706 -2093
rect -698 -2101 -696 -2093
rect -572 -2101 -570 -2093
rect -562 -2101 -560 -2093
rect -546 -2101 -544 -2093
rect -536 -2101 -534 -2093
rect -520 -2101 -518 -2093
rect -510 -2101 -508 -2093
rect -502 -2101 -500 -2093
rect -492 -2101 -490 -2093
rect -476 -2101 -474 -2093
rect -468 -2101 -466 -2093
rect -458 -2101 -456 -2093
rect -442 -2101 -440 -2093
rect -432 -2101 -430 -2093
rect -424 -2101 -422 -2093
rect -414 -2101 -412 -2093
rect -398 -2101 -396 -2093
rect -390 -2101 -388 -2093
rect -374 -2101 -372 -2093
rect -358 -2101 -356 -2093
rect -350 -2101 -348 -2093
rect -340 -2101 -338 -2093
rect -214 -2101 -212 -2093
rect -204 -2101 -202 -2093
rect -188 -2101 -186 -2093
rect -178 -2101 -176 -2093
rect -162 -2101 -160 -2093
rect -152 -2101 -150 -2093
rect -144 -2101 -142 -2093
rect -134 -2101 -132 -2093
rect -118 -2101 -116 -2093
rect -110 -2101 -108 -2093
rect -100 -2101 -98 -2093
rect -84 -2101 -82 -2093
rect -74 -2101 -72 -2093
rect -66 -2101 -64 -2093
rect -56 -2101 -54 -2093
rect -40 -2101 -38 -2093
rect -32 -2101 -30 -2093
rect -16 -2101 -14 -2093
rect 0 -2101 2 -2093
rect 8 -2101 10 -2093
rect 18 -2101 20 -2093
rect 214 -2101 216 -2093
rect 224 -2101 226 -2093
rect 240 -2101 242 -2093
rect 250 -2101 252 -2093
rect 266 -2101 268 -2093
rect 276 -2101 278 -2093
rect 284 -2101 286 -2093
rect 294 -2101 296 -2093
rect 310 -2101 312 -2093
rect 318 -2101 320 -2093
rect 328 -2101 330 -2093
rect 344 -2101 346 -2093
rect 354 -2101 356 -2093
rect 362 -2101 364 -2093
rect 372 -2101 374 -2093
rect 388 -2101 390 -2093
rect 396 -2101 398 -2093
rect 412 -2101 414 -2093
rect 428 -2101 430 -2093
rect 436 -2101 438 -2093
rect 446 -2101 448 -2093
rect 570 -2101 572 -2093
rect 580 -2101 582 -2093
rect 596 -2101 598 -2093
rect 606 -2101 608 -2093
rect 622 -2101 624 -2093
rect 632 -2101 634 -2093
rect 640 -2101 642 -2093
rect 650 -2101 652 -2093
rect 666 -2101 668 -2093
rect 674 -2101 676 -2093
rect 684 -2101 686 -2093
rect 700 -2101 702 -2093
rect 710 -2101 712 -2093
rect 718 -2101 720 -2093
rect 728 -2101 730 -2093
rect 744 -2101 746 -2093
rect 752 -2101 754 -2093
rect 768 -2101 770 -2093
rect 784 -2101 786 -2093
rect 792 -2101 794 -2093
rect 802 -2101 804 -2093
rect 968 -2101 970 -2093
rect 978 -2101 980 -2093
rect 994 -2101 996 -2093
rect 1004 -2101 1006 -2093
rect 1020 -2101 1022 -2093
rect 1030 -2101 1032 -2093
rect 1038 -2101 1040 -2093
rect 1048 -2101 1050 -2093
rect 1064 -2101 1066 -2093
rect 1072 -2101 1074 -2093
rect 1082 -2101 1084 -2093
rect 1098 -2101 1100 -2093
rect 1108 -2101 1110 -2093
rect 1116 -2101 1118 -2093
rect 1126 -2101 1128 -2093
rect 1142 -2101 1144 -2093
rect 1150 -2101 1152 -2093
rect 1166 -2101 1168 -2093
rect 1182 -2101 1184 -2093
rect 1190 -2101 1192 -2093
rect 1200 -2101 1202 -2093
rect 1326 -2101 1328 -2093
rect 1336 -2101 1338 -2093
rect 1352 -2101 1354 -2093
rect 1362 -2101 1364 -2093
rect 1378 -2101 1380 -2093
rect 1388 -2101 1390 -2093
rect 1396 -2101 1398 -2093
rect 1406 -2101 1408 -2093
rect 1422 -2101 1424 -2093
rect 1430 -2101 1432 -2093
rect 1440 -2101 1442 -2093
rect 1456 -2101 1458 -2093
rect 1466 -2101 1468 -2093
rect 1474 -2101 1476 -2093
rect 1484 -2101 1486 -2093
rect 1500 -2101 1502 -2093
rect 1508 -2101 1510 -2093
rect 1524 -2101 1526 -2093
rect 1540 -2101 1542 -2093
rect 1548 -2101 1550 -2093
rect 1558 -2101 1560 -2093
rect -1259 -2245 -1257 -2237
rect -1249 -2245 -1247 -2237
rect -1233 -2245 -1231 -2237
rect -1225 -2245 -1223 -2237
rect -1209 -2245 -1207 -2237
rect -1201 -2245 -1199 -2237
rect -1191 -2245 -1189 -2237
rect -1183 -2245 -1181 -2237
rect -1167 -2245 -1165 -2237
rect -1159 -2245 -1157 -2237
rect -1149 -2245 -1147 -2237
rect -1141 -2245 -1139 -2237
rect -1125 -2245 -1123 -2237
rect -1117 -2245 -1115 -2237
rect -1107 -2245 -1105 -2237
rect -1099 -2245 -1097 -2237
rect -1083 -2245 -1081 -2237
rect -1075 -2245 -1073 -2237
rect -930 -2245 -928 -2237
rect -920 -2245 -918 -2237
rect -904 -2245 -902 -2237
rect -896 -2245 -894 -2237
rect -880 -2245 -878 -2237
rect -872 -2245 -870 -2237
rect -862 -2245 -860 -2237
rect -854 -2245 -852 -2237
rect -838 -2245 -836 -2237
rect -830 -2245 -828 -2237
rect -820 -2245 -818 -2237
rect -812 -2245 -810 -2237
rect -796 -2245 -794 -2237
rect -788 -2245 -786 -2237
rect -778 -2245 -776 -2237
rect -770 -2245 -768 -2237
rect -754 -2245 -752 -2237
rect -746 -2245 -744 -2237
rect -572 -2245 -570 -2237
rect -562 -2245 -560 -2237
rect -546 -2245 -544 -2237
rect -538 -2245 -536 -2237
rect -522 -2245 -520 -2237
rect -514 -2245 -512 -2237
rect -504 -2245 -502 -2237
rect -496 -2245 -494 -2237
rect -480 -2245 -478 -2237
rect -472 -2245 -470 -2237
rect -462 -2245 -460 -2237
rect -454 -2245 -452 -2237
rect -438 -2245 -436 -2237
rect -430 -2245 -428 -2237
rect -420 -2245 -418 -2237
rect -412 -2245 -410 -2237
rect -396 -2245 -394 -2237
rect -388 -2245 -386 -2237
rect -214 -2245 -212 -2237
rect -204 -2245 -202 -2237
rect -188 -2245 -186 -2237
rect -180 -2245 -178 -2237
rect -164 -2245 -162 -2237
rect -156 -2245 -154 -2237
rect -146 -2245 -144 -2237
rect -138 -2245 -136 -2237
rect -122 -2245 -120 -2237
rect -114 -2245 -112 -2237
rect -104 -2245 -102 -2237
rect -96 -2245 -94 -2237
rect -80 -2245 -78 -2237
rect -72 -2245 -70 -2237
rect -62 -2245 -60 -2237
rect -54 -2245 -52 -2237
rect -38 -2245 -36 -2237
rect -30 -2245 -28 -2237
rect 214 -2245 216 -2237
rect 224 -2245 226 -2237
rect 240 -2245 242 -2237
rect 248 -2245 250 -2237
rect 264 -2245 266 -2237
rect 272 -2245 274 -2237
rect 282 -2245 284 -2237
rect 290 -2245 292 -2237
rect 306 -2245 308 -2237
rect 314 -2245 316 -2237
rect 324 -2245 326 -2237
rect 332 -2245 334 -2237
rect 348 -2245 350 -2237
rect 356 -2245 358 -2237
rect 366 -2245 368 -2237
rect 374 -2245 376 -2237
rect 390 -2245 392 -2237
rect 398 -2245 400 -2237
rect 570 -2245 572 -2237
rect 580 -2245 582 -2237
rect 596 -2245 598 -2237
rect 604 -2245 606 -2237
rect 620 -2245 622 -2237
rect 628 -2245 630 -2237
rect 638 -2245 640 -2237
rect 646 -2245 648 -2237
rect 662 -2245 664 -2237
rect 670 -2245 672 -2237
rect 680 -2245 682 -2237
rect 688 -2245 690 -2237
rect 704 -2245 706 -2237
rect 712 -2245 714 -2237
rect 722 -2245 724 -2237
rect 730 -2245 732 -2237
rect 746 -2245 748 -2237
rect 754 -2245 756 -2237
rect -1259 -2376 -1257 -2368
rect -1249 -2376 -1247 -2368
rect -1233 -2376 -1231 -2368
rect -1225 -2376 -1223 -2368
rect -1209 -2376 -1207 -2368
rect -1201 -2376 -1199 -2368
rect -1191 -2376 -1189 -2368
rect -1183 -2376 -1181 -2368
rect -1167 -2376 -1165 -2368
rect -1159 -2376 -1157 -2368
rect -1149 -2376 -1147 -2368
rect -1141 -2376 -1139 -2368
rect -1125 -2376 -1123 -2368
rect -1117 -2376 -1115 -2368
rect -1107 -2376 -1105 -2368
rect -1099 -2376 -1097 -2368
rect -1083 -2376 -1081 -2368
rect -1075 -2376 -1073 -2368
rect -930 -2376 -928 -2368
rect -920 -2376 -918 -2368
rect -904 -2376 -902 -2368
rect -896 -2376 -894 -2368
rect -880 -2376 -878 -2368
rect -872 -2376 -870 -2368
rect -862 -2376 -860 -2368
rect -854 -2376 -852 -2368
rect -838 -2376 -836 -2368
rect -830 -2376 -828 -2368
rect -820 -2376 -818 -2368
rect -812 -2376 -810 -2368
rect -796 -2376 -794 -2368
rect -788 -2376 -786 -2368
rect -778 -2376 -776 -2368
rect -770 -2376 -768 -2368
rect -754 -2376 -752 -2368
rect -746 -2376 -744 -2368
rect -572 -2376 -570 -2368
rect -562 -2376 -560 -2368
rect -546 -2376 -544 -2368
rect -538 -2376 -536 -2368
rect -522 -2376 -520 -2368
rect -514 -2376 -512 -2368
rect -504 -2376 -502 -2368
rect -496 -2376 -494 -2368
rect -480 -2376 -478 -2368
rect -472 -2376 -470 -2368
rect -462 -2376 -460 -2368
rect -454 -2376 -452 -2368
rect -438 -2376 -436 -2368
rect -430 -2376 -428 -2368
rect -420 -2376 -418 -2368
rect -412 -2376 -410 -2368
rect -396 -2376 -394 -2368
rect -388 -2376 -386 -2368
rect -214 -2376 -212 -2368
rect -204 -2376 -202 -2368
rect -188 -2376 -186 -2368
rect -180 -2376 -178 -2368
rect -164 -2376 -162 -2368
rect -156 -2376 -154 -2368
rect -146 -2376 -144 -2368
rect -138 -2376 -136 -2368
rect -122 -2376 -120 -2368
rect -114 -2376 -112 -2368
rect -104 -2376 -102 -2368
rect -96 -2376 -94 -2368
rect -80 -2376 -78 -2368
rect -72 -2376 -70 -2368
rect -62 -2376 -60 -2368
rect -54 -2376 -52 -2368
rect -38 -2376 -36 -2368
rect -30 -2376 -28 -2368
rect 214 -2376 216 -2368
rect 224 -2376 226 -2368
rect 240 -2376 242 -2368
rect 248 -2376 250 -2368
rect 264 -2376 266 -2368
rect 272 -2376 274 -2368
rect 282 -2376 284 -2368
rect 290 -2376 292 -2368
rect 306 -2376 308 -2368
rect 314 -2376 316 -2368
rect 324 -2376 326 -2368
rect 332 -2376 334 -2368
rect 348 -2376 350 -2368
rect 356 -2376 358 -2368
rect 366 -2376 368 -2368
rect 374 -2376 376 -2368
rect 390 -2376 392 -2368
rect 398 -2376 400 -2368
rect 570 -2376 572 -2368
rect 580 -2376 582 -2368
rect 596 -2376 598 -2368
rect 604 -2376 606 -2368
rect 620 -2376 622 -2368
rect 628 -2376 630 -2368
rect 638 -2376 640 -2368
rect 646 -2376 648 -2368
rect 662 -2376 664 -2368
rect 670 -2376 672 -2368
rect 680 -2376 682 -2368
rect 688 -2376 690 -2368
rect 704 -2376 706 -2368
rect 712 -2376 714 -2368
rect 722 -2376 724 -2368
rect 730 -2376 732 -2368
rect 746 -2376 748 -2368
rect 754 -2376 756 -2368
rect 968 -2376 970 -2368
rect 978 -2376 980 -2368
rect 994 -2376 996 -2368
rect 1002 -2376 1004 -2368
rect 1018 -2376 1020 -2368
rect 1026 -2376 1028 -2368
rect 1036 -2376 1038 -2368
rect 1044 -2376 1046 -2368
rect 1060 -2376 1062 -2368
rect 1068 -2376 1070 -2368
rect 1078 -2376 1080 -2368
rect 1086 -2376 1088 -2368
rect 1102 -2376 1104 -2368
rect 1110 -2376 1112 -2368
rect 1120 -2376 1122 -2368
rect 1128 -2376 1130 -2368
rect 1144 -2376 1146 -2368
rect 1152 -2376 1154 -2368
rect 1326 -2376 1328 -2368
rect 1336 -2376 1338 -2368
rect 1352 -2376 1354 -2368
rect 1360 -2376 1362 -2368
rect 1376 -2376 1378 -2368
rect 1384 -2376 1386 -2368
rect 1394 -2376 1396 -2368
rect 1402 -2376 1404 -2368
rect 1418 -2376 1420 -2368
rect 1426 -2376 1428 -2368
rect 1436 -2376 1438 -2368
rect 1444 -2376 1446 -2368
rect 1460 -2376 1462 -2368
rect 1468 -2376 1470 -2368
rect 1478 -2376 1480 -2368
rect 1486 -2376 1488 -2368
rect 1502 -2376 1504 -2368
rect 1510 -2376 1512 -2368
rect -1259 -2507 -1257 -2499
rect -1249 -2507 -1247 -2499
rect -1233 -2507 -1231 -2499
rect -1225 -2507 -1223 -2499
rect -1209 -2507 -1207 -2499
rect -1201 -2507 -1199 -2499
rect -1191 -2507 -1189 -2499
rect -1183 -2507 -1181 -2499
rect -1167 -2507 -1165 -2499
rect -1159 -2507 -1157 -2499
rect -1149 -2507 -1147 -2499
rect -1141 -2507 -1139 -2499
rect -1125 -2507 -1123 -2499
rect -1117 -2507 -1115 -2499
rect -1107 -2507 -1105 -2499
rect -1099 -2507 -1097 -2499
rect -1083 -2507 -1081 -2499
rect -1075 -2507 -1073 -2499
rect -930 -2507 -928 -2499
rect -920 -2507 -918 -2499
rect -904 -2507 -902 -2499
rect -896 -2507 -894 -2499
rect -880 -2507 -878 -2499
rect -872 -2507 -870 -2499
rect -862 -2507 -860 -2499
rect -854 -2507 -852 -2499
rect -838 -2507 -836 -2499
rect -830 -2507 -828 -2499
rect -820 -2507 -818 -2499
rect -812 -2507 -810 -2499
rect -796 -2507 -794 -2499
rect -788 -2507 -786 -2499
rect -778 -2507 -776 -2499
rect -770 -2507 -768 -2499
rect -754 -2507 -752 -2499
rect -746 -2507 -744 -2499
rect -572 -2507 -570 -2499
rect -562 -2507 -560 -2499
rect -546 -2507 -544 -2499
rect -538 -2507 -536 -2499
rect -522 -2507 -520 -2499
rect -514 -2507 -512 -2499
rect -504 -2507 -502 -2499
rect -496 -2507 -494 -2499
rect -480 -2507 -478 -2499
rect -472 -2507 -470 -2499
rect -462 -2507 -460 -2499
rect -454 -2507 -452 -2499
rect -438 -2507 -436 -2499
rect -430 -2507 -428 -2499
rect -420 -2507 -418 -2499
rect -412 -2507 -410 -2499
rect -396 -2507 -394 -2499
rect -388 -2507 -386 -2499
rect -214 -2507 -212 -2499
rect -204 -2507 -202 -2499
rect -188 -2507 -186 -2499
rect -180 -2507 -178 -2499
rect -164 -2507 -162 -2499
rect -156 -2507 -154 -2499
rect -146 -2507 -144 -2499
rect -138 -2507 -136 -2499
rect -122 -2507 -120 -2499
rect -114 -2507 -112 -2499
rect -104 -2507 -102 -2499
rect -96 -2507 -94 -2499
rect -80 -2507 -78 -2499
rect -72 -2507 -70 -2499
rect -62 -2507 -60 -2499
rect -54 -2507 -52 -2499
rect -38 -2507 -36 -2499
rect -30 -2507 -28 -2499
rect 95 -2531 97 -2499
rect 214 -2507 216 -2499
rect 224 -2507 226 -2499
rect 240 -2507 242 -2499
rect 248 -2507 250 -2499
rect 264 -2507 266 -2499
rect 272 -2507 274 -2499
rect 282 -2507 284 -2499
rect 290 -2507 292 -2499
rect 306 -2507 308 -2499
rect 314 -2507 316 -2499
rect 324 -2507 326 -2499
rect 332 -2507 334 -2499
rect 348 -2507 350 -2499
rect 356 -2507 358 -2499
rect 366 -2507 368 -2499
rect 374 -2507 376 -2499
rect 390 -2507 392 -2499
rect 398 -2507 400 -2499
rect 570 -2507 572 -2499
rect 580 -2507 582 -2499
rect 596 -2507 598 -2499
rect 604 -2507 606 -2499
rect 620 -2507 622 -2499
rect 628 -2507 630 -2499
rect 638 -2507 640 -2499
rect 646 -2507 648 -2499
rect 662 -2507 664 -2499
rect 670 -2507 672 -2499
rect 680 -2507 682 -2499
rect 688 -2507 690 -2499
rect 704 -2507 706 -2499
rect 712 -2507 714 -2499
rect 722 -2507 724 -2499
rect 730 -2507 732 -2499
rect 746 -2507 748 -2499
rect 754 -2507 756 -2499
rect 968 -2507 970 -2499
rect 978 -2507 980 -2499
rect 994 -2507 996 -2499
rect 1002 -2507 1004 -2499
rect 1018 -2507 1020 -2499
rect 1026 -2507 1028 -2499
rect 1036 -2507 1038 -2499
rect 1044 -2507 1046 -2499
rect 1060 -2507 1062 -2499
rect 1068 -2507 1070 -2499
rect 1078 -2507 1080 -2499
rect 1086 -2507 1088 -2499
rect 1102 -2507 1104 -2499
rect 1110 -2507 1112 -2499
rect 1120 -2507 1122 -2499
rect 1128 -2507 1130 -2499
rect 1144 -2507 1146 -2499
rect 1152 -2507 1154 -2499
rect 1326 -2507 1328 -2499
rect 1336 -2507 1338 -2499
rect 1352 -2507 1354 -2499
rect 1360 -2507 1362 -2499
rect 1376 -2507 1378 -2499
rect 1384 -2507 1386 -2499
rect 1394 -2507 1396 -2499
rect 1402 -2507 1404 -2499
rect 1418 -2507 1420 -2499
rect 1426 -2507 1428 -2499
rect 1436 -2507 1438 -2499
rect 1444 -2507 1446 -2499
rect 1460 -2507 1462 -2499
rect 1468 -2507 1470 -2499
rect 1478 -2507 1480 -2499
rect 1486 -2507 1488 -2499
rect 1502 -2507 1504 -2499
rect 1510 -2507 1512 -2499
rect -1259 -2619 -1257 -2611
rect -1249 -2619 -1247 -2611
rect -1233 -2619 -1231 -2611
rect -1225 -2619 -1223 -2611
rect -1209 -2619 -1207 -2611
rect -1201 -2619 -1199 -2611
rect -1191 -2619 -1189 -2611
rect -1183 -2619 -1181 -2611
rect -1167 -2619 -1165 -2611
rect -1159 -2619 -1157 -2611
rect -1149 -2619 -1147 -2611
rect -1141 -2619 -1139 -2611
rect -1125 -2619 -1123 -2611
rect -1117 -2619 -1115 -2611
rect -1107 -2619 -1105 -2611
rect -1099 -2619 -1097 -2611
rect -1083 -2619 -1081 -2611
rect -1075 -2619 -1073 -2611
rect -930 -2619 -928 -2611
rect -920 -2619 -918 -2611
rect -904 -2619 -902 -2611
rect -896 -2619 -894 -2611
rect -880 -2619 -878 -2611
rect -872 -2619 -870 -2611
rect -862 -2619 -860 -2611
rect -854 -2619 -852 -2611
rect -838 -2619 -836 -2611
rect -830 -2619 -828 -2611
rect -820 -2619 -818 -2611
rect -812 -2619 -810 -2611
rect -796 -2619 -794 -2611
rect -788 -2619 -786 -2611
rect -778 -2619 -776 -2611
rect -770 -2619 -768 -2611
rect -754 -2619 -752 -2611
rect -746 -2619 -744 -2611
rect -1334 -2732 -1332 -2724
rect -1326 -2732 -1324 -2724
rect -1316 -2732 -1314 -2724
rect -930 -2732 -928 -2724
rect -922 -2732 -920 -2724
rect -912 -2732 -910 -2724
rect -572 -2732 -570 -2724
rect -564 -2732 -562 -2724
rect -554 -2732 -552 -2724
rect -214 -2732 -212 -2724
rect -206 -2732 -204 -2724
rect -196 -2732 -194 -2724
rect 214 -2732 216 -2724
rect 222 -2732 224 -2724
rect 232 -2732 234 -2724
rect 570 -2732 572 -2724
rect 578 -2732 580 -2724
rect 588 -2732 590 -2724
rect 968 -2732 970 -2724
rect 976 -2732 978 -2724
rect 986 -2732 988 -2724
rect 1326 -2732 1328 -2724
rect 1334 -2732 1336 -2724
rect 1344 -2732 1346 -2724
rect -1259 -2851 -1257 -2843
rect -1249 -2851 -1247 -2843
rect -1233 -2851 -1231 -2843
rect -1223 -2851 -1221 -2843
rect -1215 -2851 -1213 -2843
rect -1205 -2851 -1203 -2843
rect -1189 -2851 -1187 -2843
rect -1181 -2851 -1179 -2843
rect -1171 -2851 -1169 -2843
rect -930 -2851 -928 -2843
rect -920 -2851 -918 -2843
rect -904 -2851 -902 -2843
rect -894 -2851 -892 -2843
rect -878 -2851 -876 -2843
rect -868 -2851 -866 -2843
rect -860 -2851 -858 -2843
rect -850 -2851 -848 -2843
rect -834 -2851 -832 -2843
rect -826 -2851 -824 -2843
rect -816 -2851 -814 -2843
rect -800 -2851 -798 -2843
rect -790 -2851 -788 -2843
rect -782 -2851 -780 -2843
rect -772 -2851 -770 -2843
rect -756 -2851 -754 -2843
rect -748 -2851 -746 -2843
rect -732 -2851 -730 -2843
rect -716 -2851 -714 -2843
rect -708 -2851 -706 -2843
rect -698 -2851 -696 -2843
rect -572 -2851 -570 -2843
rect -562 -2851 -560 -2843
rect -546 -2851 -544 -2843
rect -536 -2851 -534 -2843
rect -520 -2851 -518 -2843
rect -510 -2851 -508 -2843
rect -502 -2851 -500 -2843
rect -492 -2851 -490 -2843
rect -476 -2851 -474 -2843
rect -468 -2851 -466 -2843
rect -458 -2851 -456 -2843
rect -442 -2851 -440 -2843
rect -432 -2851 -430 -2843
rect -424 -2851 -422 -2843
rect -414 -2851 -412 -2843
rect -398 -2851 -396 -2843
rect -390 -2851 -388 -2843
rect -374 -2851 -372 -2843
rect -358 -2851 -356 -2843
rect -350 -2851 -348 -2843
rect -340 -2851 -338 -2843
rect -214 -2851 -212 -2843
rect -204 -2851 -202 -2843
rect -188 -2851 -186 -2843
rect -178 -2851 -176 -2843
rect -162 -2851 -160 -2843
rect -152 -2851 -150 -2843
rect -144 -2851 -142 -2843
rect -134 -2851 -132 -2843
rect -118 -2851 -116 -2843
rect -110 -2851 -108 -2843
rect -100 -2851 -98 -2843
rect -84 -2851 -82 -2843
rect -74 -2851 -72 -2843
rect -66 -2851 -64 -2843
rect -56 -2851 -54 -2843
rect -40 -2851 -38 -2843
rect -32 -2851 -30 -2843
rect -16 -2851 -14 -2843
rect 0 -2851 2 -2843
rect 8 -2851 10 -2843
rect 18 -2851 20 -2843
rect 214 -2851 216 -2843
rect 224 -2851 226 -2843
rect 240 -2851 242 -2843
rect 250 -2851 252 -2843
rect 266 -2851 268 -2843
rect 276 -2851 278 -2843
rect 284 -2851 286 -2843
rect 294 -2851 296 -2843
rect 310 -2851 312 -2843
rect 318 -2851 320 -2843
rect 328 -2851 330 -2843
rect 344 -2851 346 -2843
rect 354 -2851 356 -2843
rect 362 -2851 364 -2843
rect 372 -2851 374 -2843
rect 388 -2851 390 -2843
rect 396 -2851 398 -2843
rect 412 -2851 414 -2843
rect 428 -2851 430 -2843
rect 436 -2851 438 -2843
rect 446 -2851 448 -2843
rect 570 -2851 572 -2843
rect 580 -2851 582 -2843
rect 596 -2851 598 -2843
rect 606 -2851 608 -2843
rect 622 -2851 624 -2843
rect 632 -2851 634 -2843
rect 640 -2851 642 -2843
rect 650 -2851 652 -2843
rect 666 -2851 668 -2843
rect 674 -2851 676 -2843
rect 684 -2851 686 -2843
rect 700 -2851 702 -2843
rect 710 -2851 712 -2843
rect 718 -2851 720 -2843
rect 728 -2851 730 -2843
rect 744 -2851 746 -2843
rect 752 -2851 754 -2843
rect 768 -2851 770 -2843
rect 784 -2851 786 -2843
rect 792 -2851 794 -2843
rect 802 -2851 804 -2843
rect 968 -2851 970 -2843
rect 978 -2851 980 -2843
rect 994 -2851 996 -2843
rect 1004 -2851 1006 -2843
rect 1020 -2851 1022 -2843
rect 1030 -2851 1032 -2843
rect 1038 -2851 1040 -2843
rect 1048 -2851 1050 -2843
rect 1064 -2851 1066 -2843
rect 1072 -2851 1074 -2843
rect 1082 -2851 1084 -2843
rect 1098 -2851 1100 -2843
rect 1108 -2851 1110 -2843
rect 1116 -2851 1118 -2843
rect 1126 -2851 1128 -2843
rect 1142 -2851 1144 -2843
rect 1150 -2851 1152 -2843
rect 1166 -2851 1168 -2843
rect 1182 -2851 1184 -2843
rect 1190 -2851 1192 -2843
rect 1200 -2851 1202 -2843
rect 1326 -2851 1328 -2843
rect 1336 -2851 1338 -2843
rect 1352 -2851 1354 -2843
rect 1362 -2851 1364 -2843
rect 1378 -2851 1380 -2843
rect 1388 -2851 1390 -2843
rect 1396 -2851 1398 -2843
rect 1406 -2851 1408 -2843
rect 1422 -2851 1424 -2843
rect 1430 -2851 1432 -2843
rect 1440 -2851 1442 -2843
rect 1456 -2851 1458 -2843
rect 1466 -2851 1468 -2843
rect 1474 -2851 1476 -2843
rect 1484 -2851 1486 -2843
rect 1500 -2851 1502 -2843
rect 1508 -2851 1510 -2843
rect 1524 -2851 1526 -2843
rect 1540 -2851 1542 -2843
rect 1548 -2851 1550 -2843
rect 1558 -2851 1560 -2843
rect -1259 -2970 -1257 -2962
rect -1249 -2970 -1247 -2962
rect -1233 -2970 -1231 -2962
rect -1225 -2970 -1223 -2962
rect -1209 -2970 -1207 -2962
rect -1201 -2970 -1199 -2962
rect -1191 -2970 -1189 -2962
rect -1183 -2970 -1181 -2962
rect -1167 -2970 -1165 -2962
rect -1159 -2970 -1157 -2962
rect -1149 -2970 -1147 -2962
rect -1141 -2970 -1139 -2962
rect -1125 -2970 -1123 -2962
rect -1117 -2970 -1115 -2962
rect -1107 -2970 -1105 -2962
rect -1099 -2970 -1097 -2962
rect -1083 -2970 -1081 -2962
rect -1075 -2970 -1073 -2962
rect -1021 -2970 -1019 -2962
rect -930 -2970 -928 -2962
rect -920 -2970 -918 -2962
rect -904 -2970 -902 -2962
rect -896 -2970 -894 -2962
rect -880 -2970 -878 -2962
rect -872 -2970 -870 -2962
rect -862 -2970 -860 -2962
rect -854 -2970 -852 -2962
rect -838 -2970 -836 -2962
rect -830 -2970 -828 -2962
rect -820 -2970 -818 -2962
rect -812 -2970 -810 -2962
rect -796 -2970 -794 -2962
rect -788 -2970 -786 -2962
rect -778 -2970 -776 -2962
rect -770 -2970 -768 -2962
rect -754 -2970 -752 -2962
rect -746 -2970 -744 -2962
rect -667 -2978 -665 -2962
rect -572 -2970 -570 -2962
rect -562 -2970 -560 -2962
rect -546 -2970 -544 -2962
rect -538 -2970 -536 -2962
rect -522 -2970 -520 -2962
rect -514 -2970 -512 -2962
rect -504 -2970 -502 -2962
rect -496 -2970 -494 -2962
rect -480 -2970 -478 -2962
rect -472 -2970 -470 -2962
rect -462 -2970 -460 -2962
rect -454 -2970 -452 -2962
rect -438 -2970 -436 -2962
rect -430 -2970 -428 -2962
rect -420 -2970 -418 -2962
rect -412 -2970 -410 -2962
rect -396 -2970 -394 -2962
rect -388 -2970 -386 -2962
rect -324 -2970 -322 -2962
rect -214 -2970 -212 -2962
rect -204 -2970 -202 -2962
rect -188 -2970 -186 -2962
rect -180 -2970 -178 -2962
rect -164 -2970 -162 -2962
rect -156 -2970 -154 -2962
rect -146 -2970 -144 -2962
rect -138 -2970 -136 -2962
rect -122 -2970 -120 -2962
rect -114 -2970 -112 -2962
rect -104 -2970 -102 -2962
rect -96 -2970 -94 -2962
rect -80 -2970 -78 -2962
rect -72 -2970 -70 -2962
rect -62 -2970 -60 -2962
rect -54 -2970 -52 -2962
rect -38 -2970 -36 -2962
rect -30 -2970 -28 -2962
rect 214 -2970 216 -2962
rect 224 -2970 226 -2962
rect 240 -2970 242 -2962
rect 248 -2970 250 -2962
rect 264 -2970 266 -2962
rect 272 -2970 274 -2962
rect 282 -2970 284 -2962
rect 290 -2970 292 -2962
rect 306 -2970 308 -2962
rect 314 -2970 316 -2962
rect 324 -2970 326 -2962
rect 332 -2970 334 -2962
rect 348 -2970 350 -2962
rect 356 -2970 358 -2962
rect 366 -2970 368 -2962
rect 374 -2970 376 -2962
rect 390 -2970 392 -2962
rect 398 -2970 400 -2962
rect 477 -2970 479 -2962
rect 846 -2978 848 -2962
rect 1204 -2970 1206 -2962
rect -1259 -3086 -1257 -3078
rect -1249 -3086 -1247 -3078
rect -1233 -3086 -1231 -3078
rect -1225 -3086 -1223 -3078
rect -1209 -3086 -1207 -3078
rect -1201 -3086 -1199 -3078
rect -1191 -3086 -1189 -3078
rect -1183 -3086 -1181 -3078
rect -1167 -3086 -1165 -3078
rect -1159 -3086 -1157 -3078
rect -1149 -3086 -1147 -3078
rect -1141 -3086 -1139 -3078
rect -1125 -3086 -1123 -3078
rect -1117 -3086 -1115 -3078
rect -1107 -3086 -1105 -3078
rect -1099 -3086 -1097 -3078
rect -1083 -3086 -1081 -3078
rect -1075 -3086 -1073 -3078
rect -1021 -3086 -1019 -3078
rect -930 -3086 -928 -3078
rect -920 -3086 -918 -3078
rect -904 -3086 -902 -3078
rect -896 -3086 -894 -3078
rect -880 -3086 -878 -3078
rect -872 -3086 -870 -3078
rect -862 -3086 -860 -3078
rect -854 -3086 -852 -3078
rect -838 -3086 -836 -3078
rect -830 -3086 -828 -3078
rect -820 -3086 -818 -3078
rect -812 -3086 -810 -3078
rect -796 -3086 -794 -3078
rect -788 -3086 -786 -3078
rect -778 -3086 -776 -3078
rect -770 -3086 -768 -3078
rect -754 -3086 -752 -3078
rect -746 -3086 -744 -3078
rect -572 -3086 -570 -3078
rect -562 -3086 -560 -3078
rect -546 -3086 -544 -3078
rect -538 -3086 -536 -3078
rect -522 -3086 -520 -3078
rect -514 -3086 -512 -3078
rect -504 -3086 -502 -3078
rect -496 -3086 -494 -3078
rect -480 -3086 -478 -3078
rect -472 -3086 -470 -3078
rect -462 -3086 -460 -3078
rect -454 -3086 -452 -3078
rect -438 -3086 -436 -3078
rect -430 -3086 -428 -3078
rect -420 -3086 -418 -3078
rect -412 -3086 -410 -3078
rect -396 -3086 -394 -3078
rect -388 -3086 -386 -3078
rect -324 -3086 -322 -3078
rect -214 -3086 -212 -3078
rect -204 -3086 -202 -3078
rect -188 -3086 -186 -3078
rect -180 -3086 -178 -3078
rect -164 -3086 -162 -3078
rect -156 -3086 -154 -3078
rect -146 -3086 -144 -3078
rect -138 -3086 -136 -3078
rect -122 -3086 -120 -3078
rect -114 -3086 -112 -3078
rect -104 -3086 -102 -3078
rect -96 -3086 -94 -3078
rect -80 -3086 -78 -3078
rect -72 -3086 -70 -3078
rect -62 -3086 -60 -3078
rect -54 -3086 -52 -3078
rect -38 -3086 -36 -3078
rect -30 -3086 -28 -3078
rect 214 -3086 216 -3078
rect 224 -3086 226 -3078
rect 240 -3086 242 -3078
rect 248 -3086 250 -3078
rect 264 -3086 266 -3078
rect 272 -3086 274 -3078
rect 282 -3086 284 -3078
rect 290 -3086 292 -3078
rect 306 -3086 308 -3078
rect 314 -3086 316 -3078
rect 324 -3086 326 -3078
rect 332 -3086 334 -3078
rect 348 -3086 350 -3078
rect 356 -3086 358 -3078
rect 366 -3086 368 -3078
rect 374 -3086 376 -3078
rect 390 -3086 392 -3078
rect 398 -3086 400 -3078
rect 477 -3086 479 -3078
rect 570 -3086 572 -3078
rect 580 -3086 582 -3078
rect 596 -3086 598 -3078
rect 604 -3086 606 -3078
rect 620 -3086 622 -3078
rect 628 -3086 630 -3078
rect 638 -3086 640 -3078
rect 646 -3086 648 -3078
rect 662 -3086 664 -3078
rect 670 -3086 672 -3078
rect 680 -3086 682 -3078
rect 688 -3086 690 -3078
rect 704 -3086 706 -3078
rect 712 -3086 714 -3078
rect 722 -3086 724 -3078
rect 730 -3086 732 -3078
rect 746 -3086 748 -3078
rect 754 -3086 756 -3078
rect 968 -3086 970 -3078
rect 978 -3086 980 -3078
rect 994 -3086 996 -3078
rect 1002 -3086 1004 -3078
rect 1018 -3086 1020 -3078
rect 1026 -3086 1028 -3078
rect 1036 -3086 1038 -3078
rect 1044 -3086 1046 -3078
rect 1060 -3086 1062 -3078
rect 1068 -3086 1070 -3078
rect 1078 -3086 1080 -3078
rect 1086 -3086 1088 -3078
rect 1102 -3086 1104 -3078
rect 1110 -3086 1112 -3078
rect 1120 -3086 1122 -3078
rect 1128 -3086 1130 -3078
rect 1144 -3086 1146 -3078
rect 1152 -3086 1154 -3078
rect 1204 -3086 1206 -3078
rect 1326 -3086 1328 -3078
rect 1336 -3086 1338 -3078
rect 1352 -3086 1354 -3078
rect 1360 -3086 1362 -3078
rect 1376 -3086 1378 -3078
rect 1384 -3086 1386 -3078
rect 1394 -3086 1396 -3078
rect 1402 -3086 1404 -3078
rect 1418 -3086 1420 -3078
rect 1426 -3086 1428 -3078
rect 1436 -3086 1438 -3078
rect 1444 -3086 1446 -3078
rect 1460 -3086 1462 -3078
rect 1468 -3086 1470 -3078
rect 1478 -3086 1480 -3078
rect 1486 -3086 1488 -3078
rect 1502 -3086 1504 -3078
rect 1510 -3086 1512 -3078
rect -1259 -3207 -1257 -3199
rect -1249 -3207 -1247 -3199
rect -1233 -3207 -1231 -3199
rect -1225 -3207 -1223 -3199
rect -1209 -3207 -1207 -3199
rect -1201 -3207 -1199 -3199
rect -1191 -3207 -1189 -3199
rect -1183 -3207 -1181 -3199
rect -1167 -3207 -1165 -3199
rect -1159 -3207 -1157 -3199
rect -1149 -3207 -1147 -3199
rect -1141 -3207 -1139 -3199
rect -1125 -3207 -1123 -3199
rect -1117 -3207 -1115 -3199
rect -1107 -3207 -1105 -3199
rect -1099 -3207 -1097 -3199
rect -1083 -3207 -1081 -3199
rect -1075 -3207 -1073 -3199
rect -930 -3207 -928 -3199
rect -920 -3207 -918 -3199
rect -904 -3207 -902 -3199
rect -896 -3207 -894 -3199
rect -880 -3207 -878 -3199
rect -872 -3207 -870 -3199
rect -862 -3207 -860 -3199
rect -854 -3207 -852 -3199
rect -838 -3207 -836 -3199
rect -830 -3207 -828 -3199
rect -820 -3207 -818 -3199
rect -812 -3207 -810 -3199
rect -796 -3207 -794 -3199
rect -788 -3207 -786 -3199
rect -778 -3207 -776 -3199
rect -770 -3207 -768 -3199
rect -754 -3207 -752 -3199
rect -746 -3207 -744 -3199
rect -572 -3207 -570 -3199
rect -562 -3207 -560 -3199
rect -546 -3207 -544 -3199
rect -538 -3207 -536 -3199
rect -522 -3207 -520 -3199
rect -514 -3207 -512 -3199
rect -504 -3207 -502 -3199
rect -496 -3207 -494 -3199
rect -480 -3207 -478 -3199
rect -472 -3207 -470 -3199
rect -462 -3207 -460 -3199
rect -454 -3207 -452 -3199
rect -438 -3207 -436 -3199
rect -430 -3207 -428 -3199
rect -420 -3207 -418 -3199
rect -412 -3207 -410 -3199
rect -396 -3207 -394 -3199
rect -388 -3207 -386 -3199
rect -214 -3207 -212 -3199
rect -204 -3207 -202 -3199
rect -188 -3207 -186 -3199
rect -180 -3207 -178 -3199
rect -164 -3207 -162 -3199
rect -156 -3207 -154 -3199
rect -146 -3207 -144 -3199
rect -138 -3207 -136 -3199
rect -122 -3207 -120 -3199
rect -114 -3207 -112 -3199
rect -104 -3207 -102 -3199
rect -96 -3207 -94 -3199
rect -80 -3207 -78 -3199
rect -72 -3207 -70 -3199
rect -62 -3207 -60 -3199
rect -54 -3207 -52 -3199
rect -38 -3207 -36 -3199
rect -30 -3207 -28 -3199
rect 214 -3207 216 -3199
rect 224 -3207 226 -3199
rect 240 -3207 242 -3199
rect 248 -3207 250 -3199
rect 264 -3207 266 -3199
rect 272 -3207 274 -3199
rect 282 -3207 284 -3199
rect 290 -3207 292 -3199
rect 306 -3207 308 -3199
rect 314 -3207 316 -3199
rect 324 -3207 326 -3199
rect 332 -3207 334 -3199
rect 348 -3207 350 -3199
rect 356 -3207 358 -3199
rect 366 -3207 368 -3199
rect 374 -3207 376 -3199
rect 390 -3207 392 -3199
rect 398 -3207 400 -3199
rect 570 -3207 572 -3199
rect 580 -3207 582 -3199
rect 596 -3207 598 -3199
rect 604 -3207 606 -3199
rect 620 -3207 622 -3199
rect 628 -3207 630 -3199
rect 638 -3207 640 -3199
rect 646 -3207 648 -3199
rect 662 -3207 664 -3199
rect 670 -3207 672 -3199
rect 680 -3207 682 -3199
rect 688 -3207 690 -3199
rect 704 -3207 706 -3199
rect 712 -3207 714 -3199
rect 722 -3207 724 -3199
rect 730 -3207 732 -3199
rect 746 -3207 748 -3199
rect 754 -3207 756 -3199
rect 968 -3207 970 -3199
rect 978 -3207 980 -3199
rect 994 -3207 996 -3199
rect 1002 -3207 1004 -3199
rect 1018 -3207 1020 -3199
rect 1026 -3207 1028 -3199
rect 1036 -3207 1038 -3199
rect 1044 -3207 1046 -3199
rect 1060 -3207 1062 -3199
rect 1068 -3207 1070 -3199
rect 1078 -3207 1080 -3199
rect 1086 -3207 1088 -3199
rect 1102 -3207 1104 -3199
rect 1110 -3207 1112 -3199
rect 1120 -3207 1122 -3199
rect 1128 -3207 1130 -3199
rect 1144 -3207 1146 -3199
rect 1152 -3207 1154 -3199
rect 1326 -3207 1328 -3199
rect 1336 -3207 1338 -3199
rect 1352 -3207 1354 -3199
rect 1360 -3207 1362 -3199
rect 1376 -3207 1378 -3199
rect 1384 -3207 1386 -3199
rect 1394 -3207 1396 -3199
rect 1402 -3207 1404 -3199
rect 1418 -3207 1420 -3199
rect 1426 -3207 1428 -3199
rect 1436 -3207 1438 -3199
rect 1444 -3207 1446 -3199
rect 1460 -3207 1462 -3199
rect 1468 -3207 1470 -3199
rect 1478 -3207 1480 -3199
rect 1486 -3207 1488 -3199
rect 1502 -3207 1504 -3199
rect 1510 -3207 1512 -3199
rect -1259 -3321 -1257 -3313
rect -1249 -3321 -1247 -3313
rect -1233 -3321 -1231 -3313
rect -1225 -3321 -1223 -3313
rect -1209 -3321 -1207 -3313
rect -1201 -3321 -1199 -3313
rect -1191 -3321 -1189 -3313
rect -1183 -3321 -1181 -3313
rect -1167 -3321 -1165 -3313
rect -1159 -3321 -1157 -3313
rect -1149 -3321 -1147 -3313
rect -1141 -3321 -1139 -3313
rect -1125 -3321 -1123 -3313
rect -1117 -3321 -1115 -3313
rect -1107 -3321 -1105 -3313
rect -1099 -3321 -1097 -3313
rect -1083 -3321 -1081 -3313
rect -1075 -3321 -1073 -3313
rect -930 -3321 -928 -3313
rect -920 -3321 -918 -3313
rect -904 -3321 -902 -3313
rect -896 -3321 -894 -3313
rect -880 -3321 -878 -3313
rect -872 -3321 -870 -3313
rect -862 -3321 -860 -3313
rect -854 -3321 -852 -3313
rect -838 -3321 -836 -3313
rect -830 -3321 -828 -3313
rect -820 -3321 -818 -3313
rect -812 -3321 -810 -3313
rect -796 -3321 -794 -3313
rect -788 -3321 -786 -3313
rect -778 -3321 -776 -3313
rect -770 -3321 -768 -3313
rect -754 -3321 -752 -3313
rect -746 -3321 -744 -3313
rect -572 -3321 -570 -3313
rect -562 -3321 -560 -3313
rect -546 -3321 -544 -3313
rect -538 -3321 -536 -3313
rect -522 -3321 -520 -3313
rect -514 -3321 -512 -3313
rect -504 -3321 -502 -3313
rect -496 -3321 -494 -3313
rect -480 -3321 -478 -3313
rect -472 -3321 -470 -3313
rect -462 -3321 -460 -3313
rect -454 -3321 -452 -3313
rect -438 -3321 -436 -3313
rect -430 -3321 -428 -3313
rect -420 -3321 -418 -3313
rect -412 -3321 -410 -3313
rect -396 -3321 -394 -3313
rect -388 -3321 -386 -3313
rect -1334 -3438 -1332 -3430
rect -1326 -3438 -1324 -3430
rect -1316 -3438 -1314 -3430
rect -930 -3438 -928 -3430
rect -922 -3438 -920 -3430
rect -912 -3438 -910 -3430
rect -572 -3438 -570 -3430
rect -564 -3438 -562 -3430
rect -554 -3438 -552 -3430
rect -214 -3438 -212 -3430
rect -206 -3438 -204 -3430
rect -196 -3438 -194 -3430
rect 214 -3438 216 -3430
rect 222 -3438 224 -3430
rect 232 -3438 234 -3430
rect 570 -3438 572 -3430
rect 578 -3438 580 -3430
rect 588 -3438 590 -3430
rect 968 -3438 970 -3430
rect 976 -3438 978 -3430
rect 986 -3438 988 -3430
rect 1326 -3438 1328 -3430
rect 1334 -3438 1336 -3430
rect 1344 -3438 1346 -3430
rect -1259 -3562 -1257 -3554
rect -1249 -3562 -1247 -3554
rect -1233 -3562 -1231 -3554
rect -1223 -3562 -1221 -3554
rect -1215 -3562 -1213 -3554
rect -1205 -3562 -1203 -3554
rect -1189 -3562 -1187 -3554
rect -1181 -3562 -1179 -3554
rect -1171 -3562 -1169 -3554
rect -930 -3562 -928 -3554
rect -920 -3562 -918 -3554
rect -904 -3562 -902 -3554
rect -894 -3562 -892 -3554
rect -878 -3562 -876 -3554
rect -868 -3562 -866 -3554
rect -860 -3562 -858 -3554
rect -850 -3562 -848 -3554
rect -834 -3562 -832 -3554
rect -826 -3562 -824 -3554
rect -816 -3562 -814 -3554
rect -800 -3562 -798 -3554
rect -790 -3562 -788 -3554
rect -782 -3562 -780 -3554
rect -772 -3562 -770 -3554
rect -756 -3562 -754 -3554
rect -748 -3562 -746 -3554
rect -732 -3562 -730 -3554
rect -716 -3562 -714 -3554
rect -708 -3562 -706 -3554
rect -698 -3562 -696 -3554
rect -572 -3562 -570 -3554
rect -562 -3562 -560 -3554
rect -546 -3562 -544 -3554
rect -536 -3562 -534 -3554
rect -520 -3562 -518 -3554
rect -510 -3562 -508 -3554
rect -502 -3562 -500 -3554
rect -492 -3562 -490 -3554
rect -476 -3562 -474 -3554
rect -468 -3562 -466 -3554
rect -458 -3562 -456 -3554
rect -442 -3562 -440 -3554
rect -432 -3562 -430 -3554
rect -424 -3562 -422 -3554
rect -414 -3562 -412 -3554
rect -398 -3562 -396 -3554
rect -390 -3562 -388 -3554
rect -374 -3562 -372 -3554
rect -358 -3562 -356 -3554
rect -350 -3562 -348 -3554
rect -340 -3562 -338 -3554
rect -214 -3562 -212 -3554
rect -204 -3562 -202 -3554
rect -188 -3562 -186 -3554
rect -178 -3562 -176 -3554
rect -162 -3562 -160 -3554
rect -152 -3562 -150 -3554
rect -144 -3562 -142 -3554
rect -134 -3562 -132 -3554
rect -118 -3562 -116 -3554
rect -110 -3562 -108 -3554
rect -100 -3562 -98 -3554
rect -84 -3562 -82 -3554
rect -74 -3562 -72 -3554
rect -66 -3562 -64 -3554
rect -56 -3562 -54 -3554
rect -40 -3562 -38 -3554
rect -32 -3562 -30 -3554
rect -16 -3562 -14 -3554
rect 0 -3562 2 -3554
rect 8 -3562 10 -3554
rect 18 -3562 20 -3554
rect 214 -3562 216 -3554
rect 224 -3562 226 -3554
rect 240 -3562 242 -3554
rect 250 -3562 252 -3554
rect 266 -3562 268 -3554
rect 276 -3562 278 -3554
rect 284 -3562 286 -3554
rect 294 -3562 296 -3554
rect 310 -3562 312 -3554
rect 318 -3562 320 -3554
rect 328 -3562 330 -3554
rect 344 -3562 346 -3554
rect 354 -3562 356 -3554
rect 362 -3562 364 -3554
rect 372 -3562 374 -3554
rect 388 -3562 390 -3554
rect 396 -3562 398 -3554
rect 412 -3562 414 -3554
rect 428 -3562 430 -3554
rect 436 -3562 438 -3554
rect 446 -3562 448 -3554
rect 570 -3562 572 -3554
rect 580 -3562 582 -3554
rect 596 -3562 598 -3554
rect 606 -3562 608 -3554
rect 622 -3562 624 -3554
rect 632 -3562 634 -3554
rect 640 -3562 642 -3554
rect 650 -3562 652 -3554
rect 666 -3562 668 -3554
rect 674 -3562 676 -3554
rect 684 -3562 686 -3554
rect 700 -3562 702 -3554
rect 710 -3562 712 -3554
rect 718 -3562 720 -3554
rect 728 -3562 730 -3554
rect 744 -3562 746 -3554
rect 752 -3562 754 -3554
rect 768 -3562 770 -3554
rect 784 -3562 786 -3554
rect 792 -3562 794 -3554
rect 802 -3562 804 -3554
rect 968 -3562 970 -3554
rect 978 -3562 980 -3554
rect 994 -3562 996 -3554
rect 1004 -3562 1006 -3554
rect 1020 -3562 1022 -3554
rect 1030 -3562 1032 -3554
rect 1038 -3562 1040 -3554
rect 1048 -3562 1050 -3554
rect 1064 -3562 1066 -3554
rect 1072 -3562 1074 -3554
rect 1082 -3562 1084 -3554
rect 1098 -3562 1100 -3554
rect 1108 -3562 1110 -3554
rect 1116 -3562 1118 -3554
rect 1126 -3562 1128 -3554
rect 1142 -3562 1144 -3554
rect 1150 -3562 1152 -3554
rect 1166 -3562 1168 -3554
rect 1182 -3562 1184 -3554
rect 1190 -3562 1192 -3554
rect 1200 -3562 1202 -3554
rect 1326 -3562 1328 -3554
rect 1336 -3562 1338 -3554
rect 1352 -3562 1354 -3554
rect 1362 -3562 1364 -3554
rect 1378 -3562 1380 -3554
rect 1388 -3562 1390 -3554
rect 1396 -3562 1398 -3554
rect 1406 -3562 1408 -3554
rect 1422 -3562 1424 -3554
rect 1430 -3562 1432 -3554
rect 1440 -3562 1442 -3554
rect 1456 -3562 1458 -3554
rect 1466 -3562 1468 -3554
rect 1474 -3562 1476 -3554
rect 1484 -3562 1486 -3554
rect 1500 -3562 1502 -3554
rect 1508 -3562 1510 -3554
rect 1524 -3562 1526 -3554
rect 1540 -3562 1542 -3554
rect 1548 -3562 1550 -3554
rect 1558 -3562 1560 -3554
rect -1259 -3692 -1257 -3684
rect -1249 -3692 -1247 -3684
rect -1233 -3692 -1231 -3684
rect -1225 -3692 -1223 -3684
rect -1209 -3692 -1207 -3684
rect -1201 -3692 -1199 -3684
rect -1191 -3692 -1189 -3684
rect -1183 -3692 -1181 -3684
rect -1167 -3692 -1165 -3684
rect -1159 -3692 -1157 -3684
rect -1149 -3692 -1147 -3684
rect -1141 -3692 -1139 -3684
rect -1125 -3692 -1123 -3684
rect -1117 -3692 -1115 -3684
rect -1107 -3692 -1105 -3684
rect -1099 -3692 -1097 -3684
rect -1083 -3692 -1081 -3684
rect -1075 -3692 -1073 -3684
rect -930 -3692 -928 -3684
rect -920 -3692 -918 -3684
rect -904 -3692 -902 -3684
rect -896 -3692 -894 -3684
rect -880 -3692 -878 -3684
rect -872 -3692 -870 -3684
rect -862 -3692 -860 -3684
rect -854 -3692 -852 -3684
rect -838 -3692 -836 -3684
rect -830 -3692 -828 -3684
rect -820 -3692 -818 -3684
rect -812 -3692 -810 -3684
rect -796 -3692 -794 -3684
rect -788 -3692 -786 -3684
rect -778 -3692 -776 -3684
rect -770 -3692 -768 -3684
rect -754 -3692 -752 -3684
rect -746 -3692 -744 -3684
rect -572 -3692 -570 -3684
rect -562 -3692 -560 -3684
rect -546 -3692 -544 -3684
rect -538 -3692 -536 -3684
rect -522 -3692 -520 -3684
rect -514 -3692 -512 -3684
rect -504 -3692 -502 -3684
rect -496 -3692 -494 -3684
rect -480 -3692 -478 -3684
rect -472 -3692 -470 -3684
rect -462 -3692 -460 -3684
rect -454 -3692 -452 -3684
rect -438 -3692 -436 -3684
rect -430 -3692 -428 -3684
rect -420 -3692 -418 -3684
rect -412 -3692 -410 -3684
rect -396 -3692 -394 -3684
rect -388 -3692 -386 -3684
rect -214 -3692 -212 -3684
rect -204 -3692 -202 -3684
rect -188 -3692 -186 -3684
rect -180 -3692 -178 -3684
rect -164 -3692 -162 -3684
rect -156 -3692 -154 -3684
rect -146 -3692 -144 -3684
rect -138 -3692 -136 -3684
rect -122 -3692 -120 -3684
rect -114 -3692 -112 -3684
rect -104 -3692 -102 -3684
rect -96 -3692 -94 -3684
rect -80 -3692 -78 -3684
rect -72 -3692 -70 -3684
rect -62 -3692 -60 -3684
rect -54 -3692 -52 -3684
rect -38 -3692 -36 -3684
rect -30 -3692 -28 -3684
rect 73 -3831 75 -3799
rect -1259 -3923 -1257 -3915
rect -1249 -3923 -1247 -3915
rect -1233 -3923 -1231 -3915
rect -1225 -3923 -1223 -3915
rect -1209 -3923 -1207 -3915
rect -1201 -3923 -1199 -3915
rect -1191 -3923 -1189 -3915
rect -1183 -3923 -1181 -3915
rect -1167 -3923 -1165 -3915
rect -1159 -3923 -1157 -3915
rect -1149 -3923 -1147 -3915
rect -1141 -3923 -1139 -3915
rect -1125 -3923 -1123 -3915
rect -1117 -3923 -1115 -3915
rect -1107 -3923 -1105 -3915
rect -1099 -3923 -1097 -3915
rect -1083 -3923 -1081 -3915
rect -1075 -3923 -1073 -3915
rect -930 -3923 -928 -3915
rect -920 -3923 -918 -3915
rect -904 -3923 -902 -3915
rect -896 -3923 -894 -3915
rect -880 -3923 -878 -3915
rect -872 -3923 -870 -3915
rect -862 -3923 -860 -3915
rect -854 -3923 -852 -3915
rect -838 -3923 -836 -3915
rect -830 -3923 -828 -3915
rect -820 -3923 -818 -3915
rect -812 -3923 -810 -3915
rect -796 -3923 -794 -3915
rect -788 -3923 -786 -3915
rect -778 -3923 -776 -3915
rect -770 -3923 -768 -3915
rect -754 -3923 -752 -3915
rect -746 -3923 -744 -3915
rect -572 -3923 -570 -3915
rect -562 -3923 -560 -3915
rect -546 -3923 -544 -3915
rect -538 -3923 -536 -3915
rect -522 -3923 -520 -3915
rect -514 -3923 -512 -3915
rect -504 -3923 -502 -3915
rect -496 -3923 -494 -3915
rect -480 -3923 -478 -3915
rect -472 -3923 -470 -3915
rect -462 -3923 -460 -3915
rect -454 -3923 -452 -3915
rect -438 -3923 -436 -3915
rect -430 -3923 -428 -3915
rect -420 -3923 -418 -3915
rect -412 -3923 -410 -3915
rect -396 -3923 -394 -3915
rect -388 -3923 -386 -3915
rect -214 -3923 -212 -3915
rect -204 -3923 -202 -3915
rect -188 -3923 -186 -3915
rect -180 -3923 -178 -3915
rect -164 -3923 -162 -3915
rect -156 -3923 -154 -3915
rect -146 -3923 -144 -3915
rect -138 -3923 -136 -3915
rect -122 -3923 -120 -3915
rect -114 -3923 -112 -3915
rect -104 -3923 -102 -3915
rect -96 -3923 -94 -3915
rect -80 -3923 -78 -3915
rect -72 -3923 -70 -3915
rect -62 -3923 -60 -3915
rect -54 -3923 -52 -3915
rect -38 -3923 -36 -3915
rect -30 -3923 -28 -3915
rect 214 -3923 216 -3915
rect 224 -3923 226 -3915
rect 240 -3923 242 -3915
rect 248 -3923 250 -3915
rect 264 -3923 266 -3915
rect 272 -3923 274 -3915
rect 282 -3923 284 -3915
rect 290 -3923 292 -3915
rect 306 -3923 308 -3915
rect 314 -3923 316 -3915
rect 324 -3923 326 -3915
rect 332 -3923 334 -3915
rect 348 -3923 350 -3915
rect 356 -3923 358 -3915
rect 366 -3923 368 -3915
rect 374 -3923 376 -3915
rect 390 -3923 392 -3915
rect 398 -3923 400 -3915
rect 570 -3923 572 -3915
rect 580 -3923 582 -3915
rect 596 -3923 598 -3915
rect 604 -3923 606 -3915
rect 620 -3923 622 -3915
rect 628 -3923 630 -3915
rect 638 -3923 640 -3915
rect 646 -3923 648 -3915
rect 662 -3923 664 -3915
rect 670 -3923 672 -3915
rect 680 -3923 682 -3915
rect 688 -3923 690 -3915
rect 704 -3923 706 -3915
rect 712 -3923 714 -3915
rect 722 -3923 724 -3915
rect 730 -3923 732 -3915
rect 746 -3923 748 -3915
rect 754 -3923 756 -3915
rect 968 -3923 970 -3915
rect 978 -3923 980 -3915
rect 994 -3923 996 -3915
rect 1002 -3923 1004 -3915
rect 1018 -3923 1020 -3915
rect 1026 -3923 1028 -3915
rect 1036 -3923 1038 -3915
rect 1044 -3923 1046 -3915
rect 1060 -3923 1062 -3915
rect 1068 -3923 1070 -3915
rect 1078 -3923 1080 -3915
rect 1086 -3923 1088 -3915
rect 1102 -3923 1104 -3915
rect 1110 -3923 1112 -3915
rect 1120 -3923 1122 -3915
rect 1128 -3923 1130 -3915
rect 1144 -3923 1146 -3915
rect 1152 -3923 1154 -3915
rect 1326 -3923 1328 -3915
rect 1336 -3923 1338 -3915
rect 1352 -3923 1354 -3915
rect 1360 -3923 1362 -3915
rect 1376 -3923 1378 -3915
rect 1384 -3923 1386 -3915
rect 1394 -3923 1396 -3915
rect 1402 -3923 1404 -3915
rect 1418 -3923 1420 -3915
rect 1426 -3923 1428 -3915
rect 1436 -3923 1438 -3915
rect 1444 -3923 1446 -3915
rect 1460 -3923 1462 -3915
rect 1468 -3923 1470 -3915
rect 1478 -3923 1480 -3915
rect 1486 -3923 1488 -3915
rect 1502 -3923 1504 -3915
rect 1510 -3923 1512 -3915
rect -1259 -4048 -1257 -4040
rect -1249 -4048 -1247 -4040
rect -1233 -4048 -1231 -4040
rect -1225 -4048 -1223 -4040
rect -1209 -4048 -1207 -4040
rect -1201 -4048 -1199 -4040
rect -1191 -4048 -1189 -4040
rect -1183 -4048 -1181 -4040
rect -1167 -4048 -1165 -4040
rect -1159 -4048 -1157 -4040
rect -1149 -4048 -1147 -4040
rect -1141 -4048 -1139 -4040
rect -1125 -4048 -1123 -4040
rect -1117 -4048 -1115 -4040
rect -1107 -4048 -1105 -4040
rect -1099 -4048 -1097 -4040
rect -1083 -4048 -1081 -4040
rect -1075 -4048 -1073 -4040
rect -930 -4048 -928 -4040
rect -920 -4048 -918 -4040
rect -904 -4048 -902 -4040
rect -896 -4048 -894 -4040
rect -880 -4048 -878 -4040
rect -872 -4048 -870 -4040
rect -862 -4048 -860 -4040
rect -854 -4048 -852 -4040
rect -838 -4048 -836 -4040
rect -830 -4048 -828 -4040
rect -820 -4048 -818 -4040
rect -812 -4048 -810 -4040
rect -796 -4048 -794 -4040
rect -788 -4048 -786 -4040
rect -778 -4048 -776 -4040
rect -770 -4048 -768 -4040
rect -754 -4048 -752 -4040
rect -746 -4048 -744 -4040
rect -572 -4048 -570 -4040
rect -562 -4048 -560 -4040
rect -546 -4048 -544 -4040
rect -538 -4048 -536 -4040
rect -522 -4048 -520 -4040
rect -514 -4048 -512 -4040
rect -504 -4048 -502 -4040
rect -496 -4048 -494 -4040
rect -480 -4048 -478 -4040
rect -472 -4048 -470 -4040
rect -462 -4048 -460 -4040
rect -454 -4048 -452 -4040
rect -438 -4048 -436 -4040
rect -430 -4048 -428 -4040
rect -420 -4048 -418 -4040
rect -412 -4048 -410 -4040
rect -396 -4048 -394 -4040
rect -388 -4048 -386 -4040
rect -214 -4048 -212 -4040
rect -204 -4048 -202 -4040
rect -188 -4048 -186 -4040
rect -180 -4048 -178 -4040
rect -164 -4048 -162 -4040
rect -156 -4048 -154 -4040
rect -146 -4048 -144 -4040
rect -138 -4048 -136 -4040
rect -122 -4048 -120 -4040
rect -114 -4048 -112 -4040
rect -104 -4048 -102 -4040
rect -96 -4048 -94 -4040
rect -80 -4048 -78 -4040
rect -72 -4048 -70 -4040
rect -62 -4048 -60 -4040
rect -54 -4048 -52 -4040
rect -38 -4048 -36 -4040
rect -30 -4048 -28 -4040
rect 214 -4048 216 -4040
rect 224 -4048 226 -4040
rect 240 -4048 242 -4040
rect 248 -4048 250 -4040
rect 264 -4048 266 -4040
rect 272 -4048 274 -4040
rect 282 -4048 284 -4040
rect 290 -4048 292 -4040
rect 306 -4048 308 -4040
rect 314 -4048 316 -4040
rect 324 -4048 326 -4040
rect 332 -4048 334 -4040
rect 348 -4048 350 -4040
rect 356 -4048 358 -4040
rect 366 -4048 368 -4040
rect 374 -4048 376 -4040
rect 390 -4048 392 -4040
rect 398 -4048 400 -4040
rect 570 -4048 572 -4040
rect 580 -4048 582 -4040
rect 596 -4048 598 -4040
rect 604 -4048 606 -4040
rect 620 -4048 622 -4040
rect 628 -4048 630 -4040
rect 638 -4048 640 -4040
rect 646 -4048 648 -4040
rect 662 -4048 664 -4040
rect 670 -4048 672 -4040
rect 680 -4048 682 -4040
rect 688 -4048 690 -4040
rect 704 -4048 706 -4040
rect 712 -4048 714 -4040
rect 722 -4048 724 -4040
rect 730 -4048 732 -4040
rect 746 -4048 748 -4040
rect 754 -4048 756 -4040
rect 968 -4048 970 -4040
rect 978 -4048 980 -4040
rect 994 -4048 996 -4040
rect 1002 -4048 1004 -4040
rect 1018 -4048 1020 -4040
rect 1026 -4048 1028 -4040
rect 1036 -4048 1038 -4040
rect 1044 -4048 1046 -4040
rect 1060 -4048 1062 -4040
rect 1068 -4048 1070 -4040
rect 1078 -4048 1080 -4040
rect 1086 -4048 1088 -4040
rect 1102 -4048 1104 -4040
rect 1110 -4048 1112 -4040
rect 1120 -4048 1122 -4040
rect 1128 -4048 1130 -4040
rect 1144 -4048 1146 -4040
rect 1152 -4048 1154 -4040
rect 1326 -4048 1328 -4040
rect 1336 -4048 1338 -4040
rect 1352 -4048 1354 -4040
rect 1360 -4048 1362 -4040
rect 1376 -4048 1378 -4040
rect 1384 -4048 1386 -4040
rect 1394 -4048 1396 -4040
rect 1402 -4048 1404 -4040
rect 1418 -4048 1420 -4040
rect 1426 -4048 1428 -4040
rect 1436 -4048 1438 -4040
rect 1444 -4048 1446 -4040
rect 1460 -4048 1462 -4040
rect 1468 -4048 1470 -4040
rect 1478 -4048 1480 -4040
rect 1486 -4048 1488 -4040
rect 1502 -4048 1504 -4040
rect 1510 -4048 1512 -4040
rect -1259 -4172 -1257 -4164
rect -1249 -4172 -1247 -4164
rect -1233 -4172 -1231 -4164
rect -1225 -4172 -1223 -4164
rect -1209 -4172 -1207 -4164
rect -1201 -4172 -1199 -4164
rect -1191 -4172 -1189 -4164
rect -1183 -4172 -1181 -4164
rect -1167 -4172 -1165 -4164
rect -1159 -4172 -1157 -4164
rect -1149 -4172 -1147 -4164
rect -1141 -4172 -1139 -4164
rect -1125 -4172 -1123 -4164
rect -1117 -4172 -1115 -4164
rect -1107 -4172 -1105 -4164
rect -1099 -4172 -1097 -4164
rect -1083 -4172 -1081 -4164
rect -1075 -4172 -1073 -4164
rect -1024 -4172 -1022 -4164
rect -930 -4172 -928 -4164
rect -920 -4172 -918 -4164
rect -904 -4172 -902 -4164
rect -896 -4172 -894 -4164
rect -880 -4172 -878 -4164
rect -872 -4172 -870 -4164
rect -862 -4172 -860 -4164
rect -854 -4172 -852 -4164
rect -838 -4172 -836 -4164
rect -830 -4172 -828 -4164
rect -820 -4172 -818 -4164
rect -812 -4172 -810 -4164
rect -796 -4172 -794 -4164
rect -788 -4172 -786 -4164
rect -778 -4172 -776 -4164
rect -770 -4172 -768 -4164
rect -754 -4172 -752 -4164
rect -746 -4172 -744 -4164
rect -572 -4172 -570 -4164
rect -562 -4172 -560 -4164
rect -546 -4172 -544 -4164
rect -538 -4172 -536 -4164
rect -522 -4172 -520 -4164
rect -514 -4172 -512 -4164
rect -504 -4172 -502 -4164
rect -496 -4172 -494 -4164
rect -480 -4172 -478 -4164
rect -472 -4172 -470 -4164
rect -462 -4172 -460 -4164
rect -454 -4172 -452 -4164
rect -438 -4172 -436 -4164
rect -430 -4172 -428 -4164
rect -420 -4172 -418 -4164
rect -412 -4172 -410 -4164
rect -396 -4172 -394 -4164
rect -388 -4172 -386 -4164
rect -327 -4172 -325 -4164
rect -214 -4172 -212 -4164
rect -204 -4172 -202 -4164
rect -188 -4172 -186 -4164
rect -180 -4172 -178 -4164
rect -164 -4172 -162 -4164
rect -156 -4172 -154 -4164
rect -146 -4172 -144 -4164
rect -138 -4172 -136 -4164
rect -122 -4172 -120 -4164
rect -114 -4172 -112 -4164
rect -104 -4172 -102 -4164
rect -96 -4172 -94 -4164
rect -80 -4172 -78 -4164
rect -72 -4172 -70 -4164
rect -62 -4172 -60 -4164
rect -54 -4172 -52 -4164
rect -38 -4172 -36 -4164
rect -30 -4172 -28 -4164
rect 461 -4172 463 -4164
rect 1206 -4172 1208 -4164
rect -1334 -4283 -1332 -4275
rect -1326 -4283 -1324 -4275
rect -1316 -4283 -1314 -4275
rect -1024 -4283 -1022 -4275
rect -930 -4283 -928 -4275
rect -922 -4283 -920 -4275
rect -912 -4283 -910 -4275
rect -668 -4291 -666 -4275
rect -572 -4283 -570 -4275
rect -564 -4283 -562 -4275
rect -554 -4283 -552 -4275
rect -327 -4283 -325 -4275
rect -214 -4283 -212 -4275
rect -206 -4283 -204 -4275
rect -196 -4283 -194 -4275
rect 214 -4283 216 -4275
rect 222 -4283 224 -4275
rect 232 -4283 234 -4275
rect 461 -4283 463 -4275
rect 570 -4283 572 -4275
rect 578 -4283 580 -4275
rect 588 -4283 590 -4275
rect 865 -4291 867 -4275
rect 968 -4283 970 -4275
rect 976 -4283 978 -4275
rect 986 -4283 988 -4275
rect 1206 -4283 1208 -4275
rect 1326 -4283 1328 -4275
rect 1334 -4283 1336 -4275
rect 1344 -4283 1346 -4275
rect -1259 -4402 -1257 -4394
rect -1249 -4402 -1247 -4394
rect -1233 -4402 -1231 -4394
rect -1223 -4402 -1221 -4394
rect -1215 -4402 -1213 -4394
rect -1205 -4402 -1203 -4394
rect -1189 -4402 -1187 -4394
rect -1181 -4402 -1179 -4394
rect -1171 -4402 -1169 -4394
rect -930 -4402 -928 -4394
rect -920 -4402 -918 -4394
rect -904 -4402 -902 -4394
rect -894 -4402 -892 -4394
rect -878 -4402 -876 -4394
rect -868 -4402 -866 -4394
rect -860 -4402 -858 -4394
rect -850 -4402 -848 -4394
rect -834 -4402 -832 -4394
rect -826 -4402 -824 -4394
rect -816 -4402 -814 -4394
rect -800 -4402 -798 -4394
rect -790 -4402 -788 -4394
rect -782 -4402 -780 -4394
rect -772 -4402 -770 -4394
rect -756 -4402 -754 -4394
rect -748 -4402 -746 -4394
rect -732 -4402 -730 -4394
rect -716 -4402 -714 -4394
rect -708 -4402 -706 -4394
rect -698 -4402 -696 -4394
rect -572 -4402 -570 -4394
rect -562 -4402 -560 -4394
rect -546 -4402 -544 -4394
rect -536 -4402 -534 -4394
rect -520 -4402 -518 -4394
rect -510 -4402 -508 -4394
rect -502 -4402 -500 -4394
rect -492 -4402 -490 -4394
rect -476 -4402 -474 -4394
rect -468 -4402 -466 -4394
rect -458 -4402 -456 -4394
rect -442 -4402 -440 -4394
rect -432 -4402 -430 -4394
rect -424 -4402 -422 -4394
rect -414 -4402 -412 -4394
rect -398 -4402 -396 -4394
rect -390 -4402 -388 -4394
rect -374 -4402 -372 -4394
rect -358 -4402 -356 -4394
rect -350 -4402 -348 -4394
rect -340 -4402 -338 -4394
rect -214 -4402 -212 -4394
rect -204 -4402 -202 -4394
rect -188 -4402 -186 -4394
rect -178 -4402 -176 -4394
rect -162 -4402 -160 -4394
rect -152 -4402 -150 -4394
rect -144 -4402 -142 -4394
rect -134 -4402 -132 -4394
rect -118 -4402 -116 -4394
rect -110 -4402 -108 -4394
rect -100 -4402 -98 -4394
rect -84 -4402 -82 -4394
rect -74 -4402 -72 -4394
rect -66 -4402 -64 -4394
rect -56 -4402 -54 -4394
rect -40 -4402 -38 -4394
rect -32 -4402 -30 -4394
rect -16 -4402 -14 -4394
rect 0 -4402 2 -4394
rect 8 -4402 10 -4394
rect 18 -4402 20 -4394
rect 214 -4402 216 -4394
rect 224 -4402 226 -4394
rect 240 -4402 242 -4394
rect 250 -4402 252 -4394
rect 266 -4402 268 -4394
rect 276 -4402 278 -4394
rect 284 -4402 286 -4394
rect 294 -4402 296 -4394
rect 310 -4402 312 -4394
rect 318 -4402 320 -4394
rect 328 -4402 330 -4394
rect 344 -4402 346 -4394
rect 354 -4402 356 -4394
rect 362 -4402 364 -4394
rect 372 -4402 374 -4394
rect 388 -4402 390 -4394
rect 396 -4402 398 -4394
rect 412 -4402 414 -4394
rect 428 -4402 430 -4394
rect 436 -4402 438 -4394
rect 446 -4402 448 -4394
rect 570 -4402 572 -4394
rect 580 -4402 582 -4394
rect 596 -4402 598 -4394
rect 606 -4402 608 -4394
rect 622 -4402 624 -4394
rect 632 -4402 634 -4394
rect 640 -4402 642 -4394
rect 650 -4402 652 -4394
rect 666 -4402 668 -4394
rect 674 -4402 676 -4394
rect 684 -4402 686 -4394
rect 700 -4402 702 -4394
rect 710 -4402 712 -4394
rect 718 -4402 720 -4394
rect 728 -4402 730 -4394
rect 744 -4402 746 -4394
rect 752 -4402 754 -4394
rect 768 -4402 770 -4394
rect 784 -4402 786 -4394
rect 792 -4402 794 -4394
rect 802 -4402 804 -4394
rect 968 -4402 970 -4394
rect 978 -4402 980 -4394
rect 994 -4402 996 -4394
rect 1004 -4402 1006 -4394
rect 1020 -4402 1022 -4394
rect 1030 -4402 1032 -4394
rect 1038 -4402 1040 -4394
rect 1048 -4402 1050 -4394
rect 1064 -4402 1066 -4394
rect 1072 -4402 1074 -4394
rect 1082 -4402 1084 -4394
rect 1098 -4402 1100 -4394
rect 1108 -4402 1110 -4394
rect 1116 -4402 1118 -4394
rect 1126 -4402 1128 -4394
rect 1142 -4402 1144 -4394
rect 1150 -4402 1152 -4394
rect 1166 -4402 1168 -4394
rect 1182 -4402 1184 -4394
rect 1190 -4402 1192 -4394
rect 1200 -4402 1202 -4394
rect 1326 -4402 1328 -4394
rect 1336 -4402 1338 -4394
rect 1352 -4402 1354 -4394
rect 1362 -4402 1364 -4394
rect 1378 -4402 1380 -4394
rect 1388 -4402 1390 -4394
rect 1396 -4402 1398 -4394
rect 1406 -4402 1408 -4394
rect 1422 -4402 1424 -4394
rect 1430 -4402 1432 -4394
rect 1440 -4402 1442 -4394
rect 1456 -4402 1458 -4394
rect 1466 -4402 1468 -4394
rect 1474 -4402 1476 -4394
rect 1484 -4402 1486 -4394
rect 1500 -4402 1502 -4394
rect 1508 -4402 1510 -4394
rect 1524 -4402 1526 -4394
rect 1540 -4402 1542 -4394
rect 1548 -4402 1550 -4394
rect 1558 -4402 1560 -4394
rect -1259 -4525 -1257 -4517
rect -1249 -4525 -1247 -4517
rect -1233 -4525 -1231 -4517
rect -1225 -4525 -1223 -4517
rect -1209 -4525 -1207 -4517
rect -1201 -4525 -1199 -4517
rect -1191 -4525 -1189 -4517
rect -1183 -4525 -1181 -4517
rect -1167 -4525 -1165 -4517
rect -1159 -4525 -1157 -4517
rect -1149 -4525 -1147 -4517
rect -1141 -4525 -1139 -4517
rect -1125 -4525 -1123 -4517
rect -1117 -4525 -1115 -4517
rect -1107 -4525 -1105 -4517
rect -1099 -4525 -1097 -4517
rect -1083 -4525 -1081 -4517
rect -1075 -4525 -1073 -4517
rect -930 -4525 -928 -4517
rect -920 -4525 -918 -4517
rect -904 -4525 -902 -4517
rect -896 -4525 -894 -4517
rect -880 -4525 -878 -4517
rect -872 -4525 -870 -4517
rect -862 -4525 -860 -4517
rect -854 -4525 -852 -4517
rect -838 -4525 -836 -4517
rect -830 -4525 -828 -4517
rect -820 -4525 -818 -4517
rect -812 -4525 -810 -4517
rect -796 -4525 -794 -4517
rect -788 -4525 -786 -4517
rect -778 -4525 -776 -4517
rect -770 -4525 -768 -4517
rect -754 -4525 -752 -4517
rect -746 -4525 -744 -4517
rect -572 -4525 -570 -4517
rect -562 -4525 -560 -4517
rect -546 -4525 -544 -4517
rect -538 -4525 -536 -4517
rect -522 -4525 -520 -4517
rect -514 -4525 -512 -4517
rect -504 -4525 -502 -4517
rect -496 -4525 -494 -4517
rect -480 -4525 -478 -4517
rect -472 -4525 -470 -4517
rect -462 -4525 -460 -4517
rect -454 -4525 -452 -4517
rect -438 -4525 -436 -4517
rect -430 -4525 -428 -4517
rect -420 -4525 -418 -4517
rect -412 -4525 -410 -4517
rect -396 -4525 -394 -4517
rect -388 -4525 -386 -4517
rect -1259 -4646 -1257 -4638
rect -1249 -4646 -1247 -4638
rect -1233 -4646 -1231 -4638
rect -1225 -4646 -1223 -4638
rect -1209 -4646 -1207 -4638
rect -1201 -4646 -1199 -4638
rect -1191 -4646 -1189 -4638
rect -1183 -4646 -1181 -4638
rect -1167 -4646 -1165 -4638
rect -1159 -4646 -1157 -4638
rect -1149 -4646 -1147 -4638
rect -1141 -4646 -1139 -4638
rect -1125 -4646 -1123 -4638
rect -1117 -4646 -1115 -4638
rect -1107 -4646 -1105 -4638
rect -1099 -4646 -1097 -4638
rect -1083 -4646 -1081 -4638
rect -1075 -4646 -1073 -4638
rect -930 -4646 -928 -4638
rect -920 -4646 -918 -4638
rect -904 -4646 -902 -4638
rect -896 -4646 -894 -4638
rect -880 -4646 -878 -4638
rect -872 -4646 -870 -4638
rect -862 -4646 -860 -4638
rect -854 -4646 -852 -4638
rect -838 -4646 -836 -4638
rect -830 -4646 -828 -4638
rect -820 -4646 -818 -4638
rect -812 -4646 -810 -4638
rect -796 -4646 -794 -4638
rect -788 -4646 -786 -4638
rect -778 -4646 -776 -4638
rect -770 -4646 -768 -4638
rect -754 -4646 -752 -4638
rect -746 -4646 -744 -4638
rect -572 -4646 -570 -4638
rect -562 -4646 -560 -4638
rect -546 -4646 -544 -4638
rect -538 -4646 -536 -4638
rect -522 -4646 -520 -4638
rect -514 -4646 -512 -4638
rect -504 -4646 -502 -4638
rect -496 -4646 -494 -4638
rect -480 -4646 -478 -4638
rect -472 -4646 -470 -4638
rect -462 -4646 -460 -4638
rect -454 -4646 -452 -4638
rect -438 -4646 -436 -4638
rect -430 -4646 -428 -4638
rect -420 -4646 -418 -4638
rect -412 -4646 -410 -4638
rect -396 -4646 -394 -4638
rect -388 -4646 -386 -4638
rect -214 -4646 -212 -4638
rect -204 -4646 -202 -4638
rect -188 -4646 -186 -4638
rect -180 -4646 -178 -4638
rect -164 -4646 -162 -4638
rect -156 -4646 -154 -4638
rect -146 -4646 -144 -4638
rect -138 -4646 -136 -4638
rect -122 -4646 -120 -4638
rect -114 -4646 -112 -4638
rect -104 -4646 -102 -4638
rect -96 -4646 -94 -4638
rect -80 -4646 -78 -4638
rect -72 -4646 -70 -4638
rect -62 -4646 -60 -4638
rect -54 -4646 -52 -4638
rect -38 -4646 -36 -4638
rect -30 -4646 -28 -4638
rect 214 -4646 216 -4638
rect 224 -4646 226 -4638
rect 240 -4646 242 -4638
rect 248 -4646 250 -4638
rect 264 -4646 266 -4638
rect 272 -4646 274 -4638
rect 282 -4646 284 -4638
rect 290 -4646 292 -4638
rect 306 -4646 308 -4638
rect 314 -4646 316 -4638
rect 324 -4646 326 -4638
rect 332 -4646 334 -4638
rect 348 -4646 350 -4638
rect 356 -4646 358 -4638
rect 366 -4646 368 -4638
rect 374 -4646 376 -4638
rect 390 -4646 392 -4638
rect 398 -4646 400 -4638
rect 570 -4646 572 -4638
rect 580 -4646 582 -4638
rect 596 -4646 598 -4638
rect 604 -4646 606 -4638
rect 620 -4646 622 -4638
rect 628 -4646 630 -4638
rect 638 -4646 640 -4638
rect 646 -4646 648 -4638
rect 662 -4646 664 -4638
rect 670 -4646 672 -4638
rect 680 -4646 682 -4638
rect 688 -4646 690 -4638
rect 704 -4646 706 -4638
rect 712 -4646 714 -4638
rect 722 -4646 724 -4638
rect 730 -4646 732 -4638
rect 746 -4646 748 -4638
rect 754 -4646 756 -4638
rect 968 -4646 970 -4638
rect 978 -4646 980 -4638
rect 994 -4646 996 -4638
rect 1002 -4646 1004 -4638
rect 1018 -4646 1020 -4638
rect 1026 -4646 1028 -4638
rect 1036 -4646 1038 -4638
rect 1044 -4646 1046 -4638
rect 1060 -4646 1062 -4638
rect 1068 -4646 1070 -4638
rect 1078 -4646 1080 -4638
rect 1086 -4646 1088 -4638
rect 1102 -4646 1104 -4638
rect 1110 -4646 1112 -4638
rect 1120 -4646 1122 -4638
rect 1128 -4646 1130 -4638
rect 1144 -4646 1146 -4638
rect 1152 -4646 1154 -4638
rect 1326 -4646 1328 -4638
rect 1336 -4646 1338 -4638
rect 1352 -4646 1354 -4638
rect 1360 -4646 1362 -4638
rect 1376 -4646 1378 -4638
rect 1384 -4646 1386 -4638
rect 1394 -4646 1396 -4638
rect 1402 -4646 1404 -4638
rect 1418 -4646 1420 -4638
rect 1426 -4646 1428 -4638
rect 1436 -4646 1438 -4638
rect 1444 -4646 1446 -4638
rect 1460 -4646 1462 -4638
rect 1468 -4646 1470 -4638
rect 1478 -4646 1480 -4638
rect 1486 -4646 1488 -4638
rect 1502 -4646 1504 -4638
rect 1510 -4646 1512 -4638
rect -1259 -4767 -1257 -4759
rect -1249 -4767 -1247 -4759
rect -1233 -4767 -1231 -4759
rect -1225 -4767 -1223 -4759
rect -1209 -4767 -1207 -4759
rect -1201 -4767 -1199 -4759
rect -1191 -4767 -1189 -4759
rect -1183 -4767 -1181 -4759
rect -1167 -4767 -1165 -4759
rect -1159 -4767 -1157 -4759
rect -1149 -4767 -1147 -4759
rect -1141 -4767 -1139 -4759
rect -1125 -4767 -1123 -4759
rect -1117 -4767 -1115 -4759
rect -1107 -4767 -1105 -4759
rect -1099 -4767 -1097 -4759
rect -1083 -4767 -1081 -4759
rect -1075 -4767 -1073 -4759
rect -930 -4767 -928 -4759
rect -920 -4767 -918 -4759
rect -904 -4767 -902 -4759
rect -896 -4767 -894 -4759
rect -880 -4767 -878 -4759
rect -872 -4767 -870 -4759
rect -862 -4767 -860 -4759
rect -854 -4767 -852 -4759
rect -838 -4767 -836 -4759
rect -830 -4767 -828 -4759
rect -820 -4767 -818 -4759
rect -812 -4767 -810 -4759
rect -796 -4767 -794 -4759
rect -788 -4767 -786 -4759
rect -778 -4767 -776 -4759
rect -770 -4767 -768 -4759
rect -754 -4767 -752 -4759
rect -746 -4767 -744 -4759
rect -572 -4767 -570 -4759
rect -562 -4767 -560 -4759
rect -546 -4767 -544 -4759
rect -538 -4767 -536 -4759
rect -522 -4767 -520 -4759
rect -514 -4767 -512 -4759
rect -504 -4767 -502 -4759
rect -496 -4767 -494 -4759
rect -480 -4767 -478 -4759
rect -472 -4767 -470 -4759
rect -462 -4767 -460 -4759
rect -454 -4767 -452 -4759
rect -438 -4767 -436 -4759
rect -430 -4767 -428 -4759
rect -420 -4767 -418 -4759
rect -412 -4767 -410 -4759
rect -396 -4767 -394 -4759
rect -388 -4767 -386 -4759
rect -214 -4767 -212 -4759
rect -204 -4767 -202 -4759
rect -188 -4767 -186 -4759
rect -180 -4767 -178 -4759
rect -164 -4767 -162 -4759
rect -156 -4767 -154 -4759
rect -146 -4767 -144 -4759
rect -138 -4767 -136 -4759
rect -122 -4767 -120 -4759
rect -114 -4767 -112 -4759
rect -104 -4767 -102 -4759
rect -96 -4767 -94 -4759
rect -80 -4767 -78 -4759
rect -72 -4767 -70 -4759
rect -62 -4767 -60 -4759
rect -54 -4767 -52 -4759
rect -38 -4767 -36 -4759
rect -30 -4767 -28 -4759
rect 95 -4791 97 -4759
rect 214 -4767 216 -4759
rect 224 -4767 226 -4759
rect 240 -4767 242 -4759
rect 248 -4767 250 -4759
rect 264 -4767 266 -4759
rect 272 -4767 274 -4759
rect 282 -4767 284 -4759
rect 290 -4767 292 -4759
rect 306 -4767 308 -4759
rect 314 -4767 316 -4759
rect 324 -4767 326 -4759
rect 332 -4767 334 -4759
rect 348 -4767 350 -4759
rect 356 -4767 358 -4759
rect 366 -4767 368 -4759
rect 374 -4767 376 -4759
rect 390 -4767 392 -4759
rect 398 -4767 400 -4759
rect 570 -4767 572 -4759
rect 580 -4767 582 -4759
rect 596 -4767 598 -4759
rect 604 -4767 606 -4759
rect 620 -4767 622 -4759
rect 628 -4767 630 -4759
rect 638 -4767 640 -4759
rect 646 -4767 648 -4759
rect 662 -4767 664 -4759
rect 670 -4767 672 -4759
rect 680 -4767 682 -4759
rect 688 -4767 690 -4759
rect 704 -4767 706 -4759
rect 712 -4767 714 -4759
rect 722 -4767 724 -4759
rect 730 -4767 732 -4759
rect 746 -4767 748 -4759
rect 754 -4767 756 -4759
rect 968 -4767 970 -4759
rect 978 -4767 980 -4759
rect 994 -4767 996 -4759
rect 1002 -4767 1004 -4759
rect 1018 -4767 1020 -4759
rect 1026 -4767 1028 -4759
rect 1036 -4767 1038 -4759
rect 1044 -4767 1046 -4759
rect 1060 -4767 1062 -4759
rect 1068 -4767 1070 -4759
rect 1078 -4767 1080 -4759
rect 1086 -4767 1088 -4759
rect 1102 -4767 1104 -4759
rect 1110 -4767 1112 -4759
rect 1120 -4767 1122 -4759
rect 1128 -4767 1130 -4759
rect 1144 -4767 1146 -4759
rect 1152 -4767 1154 -4759
rect 1326 -4767 1328 -4759
rect 1336 -4767 1338 -4759
rect 1352 -4767 1354 -4759
rect 1360 -4767 1362 -4759
rect 1376 -4767 1378 -4759
rect 1384 -4767 1386 -4759
rect 1394 -4767 1396 -4759
rect 1402 -4767 1404 -4759
rect 1418 -4767 1420 -4759
rect 1426 -4767 1428 -4759
rect 1436 -4767 1438 -4759
rect 1444 -4767 1446 -4759
rect 1460 -4767 1462 -4759
rect 1468 -4767 1470 -4759
rect 1478 -4767 1480 -4759
rect 1486 -4767 1488 -4759
rect 1502 -4767 1504 -4759
rect 1510 -4767 1512 -4759
rect -1259 -4885 -1257 -4877
rect -1249 -4885 -1247 -4877
rect -1233 -4885 -1231 -4877
rect -1225 -4885 -1223 -4877
rect -1209 -4885 -1207 -4877
rect -1201 -4885 -1199 -4877
rect -1191 -4885 -1189 -4877
rect -1183 -4885 -1181 -4877
rect -1167 -4885 -1165 -4877
rect -1159 -4885 -1157 -4877
rect -1149 -4885 -1147 -4877
rect -1141 -4885 -1139 -4877
rect -1125 -4885 -1123 -4877
rect -1117 -4885 -1115 -4877
rect -1107 -4885 -1105 -4877
rect -1099 -4885 -1097 -4877
rect -1083 -4885 -1081 -4877
rect -1075 -4885 -1073 -4877
rect -930 -4885 -928 -4877
rect -920 -4885 -918 -4877
rect -904 -4885 -902 -4877
rect -896 -4885 -894 -4877
rect -880 -4885 -878 -4877
rect -872 -4885 -870 -4877
rect -862 -4885 -860 -4877
rect -854 -4885 -852 -4877
rect -838 -4885 -836 -4877
rect -830 -4885 -828 -4877
rect -820 -4885 -818 -4877
rect -812 -4885 -810 -4877
rect -796 -4885 -794 -4877
rect -788 -4885 -786 -4877
rect -778 -4885 -776 -4877
rect -770 -4885 -768 -4877
rect -754 -4885 -752 -4877
rect -746 -4885 -744 -4877
rect -572 -4885 -570 -4877
rect -562 -4885 -560 -4877
rect -546 -4885 -544 -4877
rect -538 -4885 -536 -4877
rect -522 -4885 -520 -4877
rect -514 -4885 -512 -4877
rect -504 -4885 -502 -4877
rect -496 -4885 -494 -4877
rect -480 -4885 -478 -4877
rect -472 -4885 -470 -4877
rect -462 -4885 -460 -4877
rect -454 -4885 -452 -4877
rect -438 -4885 -436 -4877
rect -430 -4885 -428 -4877
rect -420 -4885 -418 -4877
rect -412 -4885 -410 -4877
rect -396 -4885 -394 -4877
rect -388 -4885 -386 -4877
rect -214 -4885 -212 -4877
rect -204 -4885 -202 -4877
rect -188 -4885 -186 -4877
rect -180 -4885 -178 -4877
rect -164 -4885 -162 -4877
rect -156 -4885 -154 -4877
rect -146 -4885 -144 -4877
rect -138 -4885 -136 -4877
rect -122 -4885 -120 -4877
rect -114 -4885 -112 -4877
rect -104 -4885 -102 -4877
rect -96 -4885 -94 -4877
rect -80 -4885 -78 -4877
rect -72 -4885 -70 -4877
rect -62 -4885 -60 -4877
rect -54 -4885 -52 -4877
rect -38 -4885 -36 -4877
rect -30 -4885 -28 -4877
rect 214 -4885 216 -4877
rect 224 -4885 226 -4877
rect 240 -4885 242 -4877
rect 248 -4885 250 -4877
rect 264 -4885 266 -4877
rect 272 -4885 274 -4877
rect 282 -4885 284 -4877
rect 290 -4885 292 -4877
rect 306 -4885 308 -4877
rect 314 -4885 316 -4877
rect 324 -4885 326 -4877
rect 332 -4885 334 -4877
rect 348 -4885 350 -4877
rect 356 -4885 358 -4877
rect 366 -4885 368 -4877
rect 374 -4885 376 -4877
rect 390 -4885 392 -4877
rect 398 -4885 400 -4877
rect -1334 -5002 -1332 -4994
rect -1326 -5002 -1324 -4994
rect -1316 -5002 -1314 -4994
rect -930 -5002 -928 -4994
rect -922 -5002 -920 -4994
rect -912 -5002 -910 -4994
rect -572 -5002 -570 -4994
rect -564 -5002 -562 -4994
rect -554 -5002 -552 -4994
rect -214 -5002 -212 -4994
rect -206 -5002 -204 -4994
rect -196 -5002 -194 -4994
rect 214 -5002 216 -4994
rect 222 -5002 224 -4994
rect 232 -5002 234 -4994
rect 570 -5002 572 -4994
rect 578 -5002 580 -4994
rect 588 -5002 590 -4994
rect 968 -5002 970 -4994
rect 976 -5002 978 -4994
rect 986 -5002 988 -4994
rect 1326 -5002 1328 -4994
rect 1334 -5002 1336 -4994
rect 1344 -5002 1346 -4994
rect -1259 -5121 -1257 -5113
rect -1249 -5121 -1247 -5113
rect -1233 -5121 -1231 -5113
rect -1223 -5121 -1221 -5113
rect -1215 -5121 -1213 -5113
rect -1205 -5121 -1203 -5113
rect -1189 -5121 -1187 -5113
rect -1181 -5121 -1179 -5113
rect -1171 -5121 -1169 -5113
rect -930 -5121 -928 -5113
rect -920 -5121 -918 -5113
rect -904 -5121 -902 -5113
rect -894 -5121 -892 -5113
rect -878 -5121 -876 -5113
rect -868 -5121 -866 -5113
rect -860 -5121 -858 -5113
rect -850 -5121 -848 -5113
rect -834 -5121 -832 -5113
rect -826 -5121 -824 -5113
rect -816 -5121 -814 -5113
rect -800 -5121 -798 -5113
rect -790 -5121 -788 -5113
rect -782 -5121 -780 -5113
rect -772 -5121 -770 -5113
rect -756 -5121 -754 -5113
rect -748 -5121 -746 -5113
rect -732 -5121 -730 -5113
rect -716 -5121 -714 -5113
rect -708 -5121 -706 -5113
rect -698 -5121 -696 -5113
rect -572 -5121 -570 -5113
rect -562 -5121 -560 -5113
rect -546 -5121 -544 -5113
rect -536 -5121 -534 -5113
rect -520 -5121 -518 -5113
rect -510 -5121 -508 -5113
rect -502 -5121 -500 -5113
rect -492 -5121 -490 -5113
rect -476 -5121 -474 -5113
rect -468 -5121 -466 -5113
rect -458 -5121 -456 -5113
rect -442 -5121 -440 -5113
rect -432 -5121 -430 -5113
rect -424 -5121 -422 -5113
rect -414 -5121 -412 -5113
rect -398 -5121 -396 -5113
rect -390 -5121 -388 -5113
rect -374 -5121 -372 -5113
rect -358 -5121 -356 -5113
rect -350 -5121 -348 -5113
rect -340 -5121 -338 -5113
rect -214 -5121 -212 -5113
rect -204 -5121 -202 -5113
rect -188 -5121 -186 -5113
rect -178 -5121 -176 -5113
rect -162 -5121 -160 -5113
rect -152 -5121 -150 -5113
rect -144 -5121 -142 -5113
rect -134 -5121 -132 -5113
rect -118 -5121 -116 -5113
rect -110 -5121 -108 -5113
rect -100 -5121 -98 -5113
rect -84 -5121 -82 -5113
rect -74 -5121 -72 -5113
rect -66 -5121 -64 -5113
rect -56 -5121 -54 -5113
rect -40 -5121 -38 -5113
rect -32 -5121 -30 -5113
rect -16 -5121 -14 -5113
rect 0 -5121 2 -5113
rect 8 -5121 10 -5113
rect 18 -5121 20 -5113
rect 214 -5121 216 -5113
rect 224 -5121 226 -5113
rect 240 -5121 242 -5113
rect 250 -5121 252 -5113
rect 266 -5121 268 -5113
rect 276 -5121 278 -5113
rect 284 -5121 286 -5113
rect 294 -5121 296 -5113
rect 310 -5121 312 -5113
rect 318 -5121 320 -5113
rect 328 -5121 330 -5113
rect 344 -5121 346 -5113
rect 354 -5121 356 -5113
rect 362 -5121 364 -5113
rect 372 -5121 374 -5113
rect 388 -5121 390 -5113
rect 396 -5121 398 -5113
rect 412 -5121 414 -5113
rect 428 -5121 430 -5113
rect 436 -5121 438 -5113
rect 446 -5121 448 -5113
rect 570 -5121 572 -5113
rect 580 -5121 582 -5113
rect 596 -5121 598 -5113
rect 606 -5121 608 -5113
rect 622 -5121 624 -5113
rect 632 -5121 634 -5113
rect 640 -5121 642 -5113
rect 650 -5121 652 -5113
rect 666 -5121 668 -5113
rect 674 -5121 676 -5113
rect 684 -5121 686 -5113
rect 700 -5121 702 -5113
rect 710 -5121 712 -5113
rect 718 -5121 720 -5113
rect 728 -5121 730 -5113
rect 744 -5121 746 -5113
rect 752 -5121 754 -5113
rect 768 -5121 770 -5113
rect 784 -5121 786 -5113
rect 792 -5121 794 -5113
rect 802 -5121 804 -5113
rect 968 -5121 970 -5113
rect 978 -5121 980 -5113
rect 994 -5121 996 -5113
rect 1004 -5121 1006 -5113
rect 1020 -5121 1022 -5113
rect 1030 -5121 1032 -5113
rect 1038 -5121 1040 -5113
rect 1048 -5121 1050 -5113
rect 1064 -5121 1066 -5113
rect 1072 -5121 1074 -5113
rect 1082 -5121 1084 -5113
rect 1098 -5121 1100 -5113
rect 1108 -5121 1110 -5113
rect 1116 -5121 1118 -5113
rect 1126 -5121 1128 -5113
rect 1142 -5121 1144 -5113
rect 1150 -5121 1152 -5113
rect 1166 -5121 1168 -5113
rect 1182 -5121 1184 -5113
rect 1190 -5121 1192 -5113
rect 1200 -5121 1202 -5113
rect 1326 -5121 1328 -5113
rect 1336 -5121 1338 -5113
rect 1352 -5121 1354 -5113
rect 1362 -5121 1364 -5113
rect 1378 -5121 1380 -5113
rect 1388 -5121 1390 -5113
rect 1396 -5121 1398 -5113
rect 1406 -5121 1408 -5113
rect 1422 -5121 1424 -5113
rect 1430 -5121 1432 -5113
rect 1440 -5121 1442 -5113
rect 1456 -5121 1458 -5113
rect 1466 -5121 1468 -5113
rect 1474 -5121 1476 -5113
rect 1484 -5121 1486 -5113
rect 1500 -5121 1502 -5113
rect 1508 -5121 1510 -5113
rect 1524 -5121 1526 -5113
rect 1540 -5121 1542 -5113
rect 1548 -5121 1550 -5113
rect 1558 -5121 1560 -5113
rect -1259 -5240 -1257 -5232
rect -1249 -5240 -1247 -5232
rect -1233 -5240 -1231 -5232
rect -1225 -5240 -1223 -5232
rect -1209 -5240 -1207 -5232
rect -1201 -5240 -1199 -5232
rect -1191 -5240 -1189 -5232
rect -1183 -5240 -1181 -5232
rect -1167 -5240 -1165 -5232
rect -1159 -5240 -1157 -5232
rect -1149 -5240 -1147 -5232
rect -1141 -5240 -1139 -5232
rect -1125 -5240 -1123 -5232
rect -1117 -5240 -1115 -5232
rect -1107 -5240 -1105 -5232
rect -1099 -5240 -1097 -5232
rect -1083 -5240 -1081 -5232
rect -1075 -5240 -1073 -5232
rect -930 -5240 -928 -5232
rect -920 -5240 -918 -5232
rect -904 -5240 -902 -5232
rect -896 -5240 -894 -5232
rect -880 -5240 -878 -5232
rect -872 -5240 -870 -5232
rect -862 -5240 -860 -5232
rect -854 -5240 -852 -5232
rect -838 -5240 -836 -5232
rect -830 -5240 -828 -5232
rect -820 -5240 -818 -5232
rect -812 -5240 -810 -5232
rect -796 -5240 -794 -5232
rect -788 -5240 -786 -5232
rect -778 -5240 -776 -5232
rect -770 -5240 -768 -5232
rect -754 -5240 -752 -5232
rect -746 -5240 -744 -5232
rect -1259 -5361 -1257 -5353
rect -1249 -5361 -1247 -5353
rect -1233 -5361 -1231 -5353
rect -1225 -5361 -1223 -5353
rect -1209 -5361 -1207 -5353
rect -1201 -5361 -1199 -5353
rect -1191 -5361 -1189 -5353
rect -1183 -5361 -1181 -5353
rect -1167 -5361 -1165 -5353
rect -1159 -5361 -1157 -5353
rect -1149 -5361 -1147 -5353
rect -1141 -5361 -1139 -5353
rect -1125 -5361 -1123 -5353
rect -1117 -5361 -1115 -5353
rect -1107 -5361 -1105 -5353
rect -1099 -5361 -1097 -5353
rect -1083 -5361 -1081 -5353
rect -1075 -5361 -1073 -5353
rect -1021 -5361 -1019 -5353
rect -930 -5361 -928 -5353
rect -920 -5361 -918 -5353
rect -904 -5361 -902 -5353
rect -896 -5361 -894 -5353
rect -880 -5361 -878 -5353
rect -872 -5361 -870 -5353
rect -862 -5361 -860 -5353
rect -854 -5361 -852 -5353
rect -838 -5361 -836 -5353
rect -830 -5361 -828 -5353
rect -820 -5361 -818 -5353
rect -812 -5361 -810 -5353
rect -796 -5361 -794 -5353
rect -788 -5361 -786 -5353
rect -778 -5361 -776 -5353
rect -770 -5361 -768 -5353
rect -754 -5361 -752 -5353
rect -746 -5361 -744 -5353
rect -668 -5369 -666 -5353
rect -572 -5361 -570 -5353
rect -562 -5361 -560 -5353
rect -546 -5361 -544 -5353
rect -538 -5361 -536 -5353
rect -522 -5361 -520 -5353
rect -514 -5361 -512 -5353
rect -504 -5361 -502 -5353
rect -496 -5361 -494 -5353
rect -480 -5361 -478 -5353
rect -472 -5361 -470 -5353
rect -462 -5361 -460 -5353
rect -454 -5361 -452 -5353
rect -438 -5361 -436 -5353
rect -430 -5361 -428 -5353
rect -420 -5361 -418 -5353
rect -412 -5361 -410 -5353
rect -396 -5361 -394 -5353
rect -388 -5361 -386 -5353
rect -322 -5361 -320 -5353
rect -214 -5361 -212 -5353
rect -204 -5361 -202 -5353
rect -188 -5361 -186 -5353
rect -180 -5361 -178 -5353
rect -164 -5361 -162 -5353
rect -156 -5361 -154 -5353
rect -146 -5361 -144 -5353
rect -138 -5361 -136 -5353
rect -122 -5361 -120 -5353
rect -114 -5361 -112 -5353
rect -104 -5361 -102 -5353
rect -96 -5361 -94 -5353
rect -80 -5361 -78 -5353
rect -72 -5361 -70 -5353
rect -62 -5361 -60 -5353
rect -54 -5361 -52 -5353
rect -38 -5361 -36 -5353
rect -30 -5361 -28 -5353
rect 214 -5361 216 -5353
rect 224 -5361 226 -5353
rect 240 -5361 242 -5353
rect 248 -5361 250 -5353
rect 264 -5361 266 -5353
rect 272 -5361 274 -5353
rect 282 -5361 284 -5353
rect 290 -5361 292 -5353
rect 306 -5361 308 -5353
rect 314 -5361 316 -5353
rect 324 -5361 326 -5353
rect 332 -5361 334 -5353
rect 348 -5361 350 -5353
rect 356 -5361 358 -5353
rect 366 -5361 368 -5353
rect 374 -5361 376 -5353
rect 390 -5361 392 -5353
rect 398 -5361 400 -5353
rect 471 -5361 473 -5353
rect 570 -5361 572 -5353
rect 580 -5361 582 -5353
rect 596 -5361 598 -5353
rect 604 -5361 606 -5353
rect 620 -5361 622 -5353
rect 628 -5361 630 -5353
rect 638 -5361 640 -5353
rect 646 -5361 648 -5353
rect 662 -5361 664 -5353
rect 670 -5361 672 -5353
rect 680 -5361 682 -5353
rect 688 -5361 690 -5353
rect 704 -5361 706 -5353
rect 712 -5361 714 -5353
rect 722 -5361 724 -5353
rect 730 -5361 732 -5353
rect 746 -5361 748 -5353
rect 754 -5361 756 -5353
rect 872 -5369 874 -5353
rect 968 -5361 970 -5353
rect 978 -5361 980 -5353
rect 994 -5361 996 -5353
rect 1002 -5361 1004 -5353
rect 1018 -5361 1020 -5353
rect 1026 -5361 1028 -5353
rect 1036 -5361 1038 -5353
rect 1044 -5361 1046 -5353
rect 1060 -5361 1062 -5353
rect 1068 -5361 1070 -5353
rect 1078 -5361 1080 -5353
rect 1086 -5361 1088 -5353
rect 1102 -5361 1104 -5353
rect 1110 -5361 1112 -5353
rect 1120 -5361 1122 -5353
rect 1128 -5361 1130 -5353
rect 1144 -5361 1146 -5353
rect 1152 -5361 1154 -5353
rect 1215 -5361 1217 -5353
rect 1326 -5361 1328 -5353
rect 1336 -5361 1338 -5353
rect 1352 -5361 1354 -5353
rect 1360 -5361 1362 -5353
rect 1376 -5361 1378 -5353
rect 1384 -5361 1386 -5353
rect 1394 -5361 1396 -5353
rect 1402 -5361 1404 -5353
rect 1418 -5361 1420 -5353
rect 1426 -5361 1428 -5353
rect 1436 -5361 1438 -5353
rect 1444 -5361 1446 -5353
rect 1460 -5361 1462 -5353
rect 1468 -5361 1470 -5353
rect 1478 -5361 1480 -5353
rect 1486 -5361 1488 -5353
rect 1502 -5361 1504 -5353
rect 1510 -5361 1512 -5353
rect -1259 -5481 -1257 -5473
rect -1249 -5481 -1247 -5473
rect -1233 -5481 -1231 -5473
rect -1225 -5481 -1223 -5473
rect -1209 -5481 -1207 -5473
rect -1201 -5481 -1199 -5473
rect -1191 -5481 -1189 -5473
rect -1183 -5481 -1181 -5473
rect -1167 -5481 -1165 -5473
rect -1159 -5481 -1157 -5473
rect -1149 -5481 -1147 -5473
rect -1141 -5481 -1139 -5473
rect -1125 -5481 -1123 -5473
rect -1117 -5481 -1115 -5473
rect -1107 -5481 -1105 -5473
rect -1099 -5481 -1097 -5473
rect -1083 -5481 -1081 -5473
rect -1075 -5481 -1073 -5473
rect -1021 -5481 -1019 -5473
rect -930 -5481 -928 -5473
rect -920 -5481 -918 -5473
rect -904 -5481 -902 -5473
rect -896 -5481 -894 -5473
rect -880 -5481 -878 -5473
rect -872 -5481 -870 -5473
rect -862 -5481 -860 -5473
rect -854 -5481 -852 -5473
rect -838 -5481 -836 -5473
rect -830 -5481 -828 -5473
rect -820 -5481 -818 -5473
rect -812 -5481 -810 -5473
rect -796 -5481 -794 -5473
rect -788 -5481 -786 -5473
rect -778 -5481 -776 -5473
rect -770 -5481 -768 -5473
rect -754 -5481 -752 -5473
rect -746 -5481 -744 -5473
rect -572 -5481 -570 -5473
rect -562 -5481 -560 -5473
rect -546 -5481 -544 -5473
rect -538 -5481 -536 -5473
rect -522 -5481 -520 -5473
rect -514 -5481 -512 -5473
rect -504 -5481 -502 -5473
rect -496 -5481 -494 -5473
rect -480 -5481 -478 -5473
rect -472 -5481 -470 -5473
rect -462 -5481 -460 -5473
rect -454 -5481 -452 -5473
rect -438 -5481 -436 -5473
rect -430 -5481 -428 -5473
rect -420 -5481 -418 -5473
rect -412 -5481 -410 -5473
rect -396 -5481 -394 -5473
rect -388 -5481 -386 -5473
rect -322 -5481 -320 -5473
rect -214 -5481 -212 -5473
rect -204 -5481 -202 -5473
rect -188 -5481 -186 -5473
rect -180 -5481 -178 -5473
rect -164 -5481 -162 -5473
rect -156 -5481 -154 -5473
rect -146 -5481 -144 -5473
rect -138 -5481 -136 -5473
rect -122 -5481 -120 -5473
rect -114 -5481 -112 -5473
rect -104 -5481 -102 -5473
rect -96 -5481 -94 -5473
rect -80 -5481 -78 -5473
rect -72 -5481 -70 -5473
rect -62 -5481 -60 -5473
rect -54 -5481 -52 -5473
rect -38 -5481 -36 -5473
rect -30 -5481 -28 -5473
rect 214 -5481 216 -5473
rect 224 -5481 226 -5473
rect 240 -5481 242 -5473
rect 248 -5481 250 -5473
rect 264 -5481 266 -5473
rect 272 -5481 274 -5473
rect 282 -5481 284 -5473
rect 290 -5481 292 -5473
rect 306 -5481 308 -5473
rect 314 -5481 316 -5473
rect 324 -5481 326 -5473
rect 332 -5481 334 -5473
rect 348 -5481 350 -5473
rect 356 -5481 358 -5473
rect 366 -5481 368 -5473
rect 374 -5481 376 -5473
rect 390 -5481 392 -5473
rect 398 -5481 400 -5473
rect 471 -5481 473 -5473
rect 570 -5481 572 -5473
rect 580 -5481 582 -5473
rect 596 -5481 598 -5473
rect 604 -5481 606 -5473
rect 620 -5481 622 -5473
rect 628 -5481 630 -5473
rect 638 -5481 640 -5473
rect 646 -5481 648 -5473
rect 662 -5481 664 -5473
rect 670 -5481 672 -5473
rect 680 -5481 682 -5473
rect 688 -5481 690 -5473
rect 704 -5481 706 -5473
rect 712 -5481 714 -5473
rect 722 -5481 724 -5473
rect 730 -5481 732 -5473
rect 746 -5481 748 -5473
rect 754 -5481 756 -5473
rect 968 -5481 970 -5473
rect 978 -5481 980 -5473
rect 994 -5481 996 -5473
rect 1002 -5481 1004 -5473
rect 1018 -5481 1020 -5473
rect 1026 -5481 1028 -5473
rect 1036 -5481 1038 -5473
rect 1044 -5481 1046 -5473
rect 1060 -5481 1062 -5473
rect 1068 -5481 1070 -5473
rect 1078 -5481 1080 -5473
rect 1086 -5481 1088 -5473
rect 1102 -5481 1104 -5473
rect 1110 -5481 1112 -5473
rect 1120 -5481 1122 -5473
rect 1128 -5481 1130 -5473
rect 1144 -5481 1146 -5473
rect 1152 -5481 1154 -5473
rect 1215 -5481 1217 -5473
rect 1326 -5481 1328 -5473
rect 1336 -5481 1338 -5473
rect 1352 -5481 1354 -5473
rect 1360 -5481 1362 -5473
rect 1376 -5481 1378 -5473
rect 1384 -5481 1386 -5473
rect 1394 -5481 1396 -5473
rect 1402 -5481 1404 -5473
rect 1418 -5481 1420 -5473
rect 1426 -5481 1428 -5473
rect 1436 -5481 1438 -5473
rect 1444 -5481 1446 -5473
rect 1460 -5481 1462 -5473
rect 1468 -5481 1470 -5473
rect 1478 -5481 1480 -5473
rect 1486 -5481 1488 -5473
rect 1502 -5481 1504 -5473
rect 1510 -5481 1512 -5473
rect -1259 -5598 -1257 -5590
rect -1249 -5598 -1247 -5590
rect -1233 -5598 -1231 -5590
rect -1225 -5598 -1223 -5590
rect -1209 -5598 -1207 -5590
rect -1201 -5598 -1199 -5590
rect -1191 -5598 -1189 -5590
rect -1183 -5598 -1181 -5590
rect -1167 -5598 -1165 -5590
rect -1159 -5598 -1157 -5590
rect -1149 -5598 -1147 -5590
rect -1141 -5598 -1139 -5590
rect -1125 -5598 -1123 -5590
rect -1117 -5598 -1115 -5590
rect -1107 -5598 -1105 -5590
rect -1099 -5598 -1097 -5590
rect -1083 -5598 -1081 -5590
rect -1075 -5598 -1073 -5590
rect -930 -5598 -928 -5590
rect -920 -5598 -918 -5590
rect -904 -5598 -902 -5590
rect -896 -5598 -894 -5590
rect -880 -5598 -878 -5590
rect -872 -5598 -870 -5590
rect -862 -5598 -860 -5590
rect -854 -5598 -852 -5590
rect -838 -5598 -836 -5590
rect -830 -5598 -828 -5590
rect -820 -5598 -818 -5590
rect -812 -5598 -810 -5590
rect -796 -5598 -794 -5590
rect -788 -5598 -786 -5590
rect -778 -5598 -776 -5590
rect -770 -5598 -768 -5590
rect -754 -5598 -752 -5590
rect -746 -5598 -744 -5590
rect -572 -5598 -570 -5590
rect -562 -5598 -560 -5590
rect -546 -5598 -544 -5590
rect -538 -5598 -536 -5590
rect -522 -5598 -520 -5590
rect -514 -5598 -512 -5590
rect -504 -5598 -502 -5590
rect -496 -5598 -494 -5590
rect -480 -5598 -478 -5590
rect -472 -5598 -470 -5590
rect -462 -5598 -460 -5590
rect -454 -5598 -452 -5590
rect -438 -5598 -436 -5590
rect -430 -5598 -428 -5590
rect -420 -5598 -418 -5590
rect -412 -5598 -410 -5590
rect -396 -5598 -394 -5590
rect -388 -5598 -386 -5590
rect -214 -5598 -212 -5590
rect -204 -5598 -202 -5590
rect -188 -5598 -186 -5590
rect -180 -5598 -178 -5590
rect -164 -5598 -162 -5590
rect -156 -5598 -154 -5590
rect -146 -5598 -144 -5590
rect -138 -5598 -136 -5590
rect -122 -5598 -120 -5590
rect -114 -5598 -112 -5590
rect -104 -5598 -102 -5590
rect -96 -5598 -94 -5590
rect -80 -5598 -78 -5590
rect -72 -5598 -70 -5590
rect -62 -5598 -60 -5590
rect -54 -5598 -52 -5590
rect -38 -5598 -36 -5590
rect -30 -5598 -28 -5590
rect 214 -5598 216 -5590
rect 224 -5598 226 -5590
rect 240 -5598 242 -5590
rect 248 -5598 250 -5590
rect 264 -5598 266 -5590
rect 272 -5598 274 -5590
rect 282 -5598 284 -5590
rect 290 -5598 292 -5590
rect 306 -5598 308 -5590
rect 314 -5598 316 -5590
rect 324 -5598 326 -5590
rect 332 -5598 334 -5590
rect 348 -5598 350 -5590
rect 356 -5598 358 -5590
rect 366 -5598 368 -5590
rect 374 -5598 376 -5590
rect 390 -5598 392 -5590
rect 398 -5598 400 -5590
rect 570 -5598 572 -5590
rect 580 -5598 582 -5590
rect 596 -5598 598 -5590
rect 604 -5598 606 -5590
rect 620 -5598 622 -5590
rect 628 -5598 630 -5590
rect 638 -5598 640 -5590
rect 646 -5598 648 -5590
rect 662 -5598 664 -5590
rect 670 -5598 672 -5590
rect 680 -5598 682 -5590
rect 688 -5598 690 -5590
rect 704 -5598 706 -5590
rect 712 -5598 714 -5590
rect 722 -5598 724 -5590
rect 730 -5598 732 -5590
rect 746 -5598 748 -5590
rect 754 -5598 756 -5590
rect -1334 -5715 -1332 -5707
rect -1326 -5715 -1324 -5707
rect -1316 -5715 -1314 -5707
rect -930 -5715 -928 -5707
rect -922 -5715 -920 -5707
rect -912 -5715 -910 -5707
rect -572 -5715 -570 -5707
rect -564 -5715 -562 -5707
rect -554 -5715 -552 -5707
rect -214 -5715 -212 -5707
rect -206 -5715 -204 -5707
rect -196 -5715 -194 -5707
rect 214 -5715 216 -5707
rect 222 -5715 224 -5707
rect 232 -5715 234 -5707
rect 570 -5715 572 -5707
rect 578 -5715 580 -5707
rect 588 -5715 590 -5707
rect 968 -5715 970 -5707
rect 976 -5715 978 -5707
rect 986 -5715 988 -5707
rect 1326 -5715 1328 -5707
rect 1334 -5715 1336 -5707
rect 1344 -5715 1346 -5707
rect -1259 -5834 -1257 -5826
rect -1249 -5834 -1247 -5826
rect -1233 -5834 -1231 -5826
rect -1223 -5834 -1221 -5826
rect -1215 -5834 -1213 -5826
rect -1205 -5834 -1203 -5826
rect -1189 -5834 -1187 -5826
rect -1181 -5834 -1179 -5826
rect -1171 -5834 -1169 -5826
rect -930 -5834 -928 -5826
rect -920 -5834 -918 -5826
rect -904 -5834 -902 -5826
rect -894 -5834 -892 -5826
rect -878 -5834 -876 -5826
rect -868 -5834 -866 -5826
rect -860 -5834 -858 -5826
rect -850 -5834 -848 -5826
rect -834 -5834 -832 -5826
rect -826 -5834 -824 -5826
rect -816 -5834 -814 -5826
rect -800 -5834 -798 -5826
rect -790 -5834 -788 -5826
rect -782 -5834 -780 -5826
rect -772 -5834 -770 -5826
rect -756 -5834 -754 -5826
rect -748 -5834 -746 -5826
rect -732 -5834 -730 -5826
rect -716 -5834 -714 -5826
rect -708 -5834 -706 -5826
rect -698 -5834 -696 -5826
rect -572 -5834 -570 -5826
rect -562 -5834 -560 -5826
rect -546 -5834 -544 -5826
rect -536 -5834 -534 -5826
rect -520 -5834 -518 -5826
rect -510 -5834 -508 -5826
rect -502 -5834 -500 -5826
rect -492 -5834 -490 -5826
rect -476 -5834 -474 -5826
rect -468 -5834 -466 -5826
rect -458 -5834 -456 -5826
rect -442 -5834 -440 -5826
rect -432 -5834 -430 -5826
rect -424 -5834 -422 -5826
rect -414 -5834 -412 -5826
rect -398 -5834 -396 -5826
rect -390 -5834 -388 -5826
rect -374 -5834 -372 -5826
rect -358 -5834 -356 -5826
rect -350 -5834 -348 -5826
rect -340 -5834 -338 -5826
rect -214 -5834 -212 -5826
rect -204 -5834 -202 -5826
rect -188 -5834 -186 -5826
rect -178 -5834 -176 -5826
rect -162 -5834 -160 -5826
rect -152 -5834 -150 -5826
rect -144 -5834 -142 -5826
rect -134 -5834 -132 -5826
rect -118 -5834 -116 -5826
rect -110 -5834 -108 -5826
rect -100 -5834 -98 -5826
rect -84 -5834 -82 -5826
rect -74 -5834 -72 -5826
rect -66 -5834 -64 -5826
rect -56 -5834 -54 -5826
rect -40 -5834 -38 -5826
rect -32 -5834 -30 -5826
rect -16 -5834 -14 -5826
rect 0 -5834 2 -5826
rect 8 -5834 10 -5826
rect 18 -5834 20 -5826
rect 214 -5834 216 -5826
rect 224 -5834 226 -5826
rect 240 -5834 242 -5826
rect 250 -5834 252 -5826
rect 266 -5834 268 -5826
rect 276 -5834 278 -5826
rect 284 -5834 286 -5826
rect 294 -5834 296 -5826
rect 310 -5834 312 -5826
rect 318 -5834 320 -5826
rect 328 -5834 330 -5826
rect 344 -5834 346 -5826
rect 354 -5834 356 -5826
rect 362 -5834 364 -5826
rect 372 -5834 374 -5826
rect 388 -5834 390 -5826
rect 396 -5834 398 -5826
rect 412 -5834 414 -5826
rect 428 -5834 430 -5826
rect 436 -5834 438 -5826
rect 446 -5834 448 -5826
rect 570 -5834 572 -5826
rect 580 -5834 582 -5826
rect 596 -5834 598 -5826
rect 606 -5834 608 -5826
rect 622 -5834 624 -5826
rect 632 -5834 634 -5826
rect 640 -5834 642 -5826
rect 650 -5834 652 -5826
rect 666 -5834 668 -5826
rect 674 -5834 676 -5826
rect 684 -5834 686 -5826
rect 700 -5834 702 -5826
rect 710 -5834 712 -5826
rect 718 -5834 720 -5826
rect 728 -5834 730 -5826
rect 744 -5834 746 -5826
rect 752 -5834 754 -5826
rect 768 -5834 770 -5826
rect 784 -5834 786 -5826
rect 792 -5834 794 -5826
rect 802 -5834 804 -5826
rect 968 -5834 970 -5826
rect 978 -5834 980 -5826
rect 994 -5834 996 -5826
rect 1004 -5834 1006 -5826
rect 1020 -5834 1022 -5826
rect 1030 -5834 1032 -5826
rect 1038 -5834 1040 -5826
rect 1048 -5834 1050 -5826
rect 1064 -5834 1066 -5826
rect 1072 -5834 1074 -5826
rect 1082 -5834 1084 -5826
rect 1098 -5834 1100 -5826
rect 1108 -5834 1110 -5826
rect 1116 -5834 1118 -5826
rect 1126 -5834 1128 -5826
rect 1142 -5834 1144 -5826
rect 1150 -5834 1152 -5826
rect 1166 -5834 1168 -5826
rect 1182 -5834 1184 -5826
rect 1190 -5834 1192 -5826
rect 1200 -5834 1202 -5826
rect 1326 -5834 1328 -5826
rect 1336 -5834 1338 -5826
rect 1352 -5834 1354 -5826
rect 1362 -5834 1364 -5826
rect 1378 -5834 1380 -5826
rect 1388 -5834 1390 -5826
rect 1396 -5834 1398 -5826
rect 1406 -5834 1408 -5826
rect 1422 -5834 1424 -5826
rect 1430 -5834 1432 -5826
rect 1440 -5834 1442 -5826
rect 1456 -5834 1458 -5826
rect 1466 -5834 1468 -5826
rect 1474 -5834 1476 -5826
rect 1484 -5834 1486 -5826
rect 1500 -5834 1502 -5826
rect 1508 -5834 1510 -5826
rect 1524 -5834 1526 -5826
rect 1540 -5834 1542 -5826
rect 1548 -5834 1550 -5826
rect 1558 -5834 1560 -5826
rect -1259 -5957 -1257 -5949
rect -1249 -5957 -1247 -5949
rect -1233 -5957 -1231 -5949
rect -1225 -5957 -1223 -5949
rect -1209 -5957 -1207 -5949
rect -1201 -5957 -1199 -5949
rect -1191 -5957 -1189 -5949
rect -1183 -5957 -1181 -5949
rect -1167 -5957 -1165 -5949
rect -1159 -5957 -1157 -5949
rect -1149 -5957 -1147 -5949
rect -1141 -5957 -1139 -5949
rect -1125 -5957 -1123 -5949
rect -1117 -5957 -1115 -5949
rect -1107 -5957 -1105 -5949
rect -1099 -5957 -1097 -5949
rect -1083 -5957 -1081 -5949
rect -1075 -5957 -1073 -5949
rect -930 -5957 -928 -5949
rect -920 -5957 -918 -5949
rect -904 -5957 -902 -5949
rect -896 -5957 -894 -5949
rect -880 -5957 -878 -5949
rect -872 -5957 -870 -5949
rect -862 -5957 -860 -5949
rect -854 -5957 -852 -5949
rect -838 -5957 -836 -5949
rect -830 -5957 -828 -5949
rect -820 -5957 -818 -5949
rect -812 -5957 -810 -5949
rect -796 -5957 -794 -5949
rect -788 -5957 -786 -5949
rect -778 -5957 -776 -5949
rect -770 -5957 -768 -5949
rect -754 -5957 -752 -5949
rect -746 -5957 -744 -5949
rect -572 -5957 -570 -5949
rect -562 -5957 -560 -5949
rect -546 -5957 -544 -5949
rect -538 -5957 -536 -5949
rect -522 -5957 -520 -5949
rect -514 -5957 -512 -5949
rect -504 -5957 -502 -5949
rect -496 -5957 -494 -5949
rect -480 -5957 -478 -5949
rect -472 -5957 -470 -5949
rect -462 -5957 -460 -5949
rect -454 -5957 -452 -5949
rect -438 -5957 -436 -5949
rect -430 -5957 -428 -5949
rect -420 -5957 -418 -5949
rect -412 -5957 -410 -5949
rect -396 -5957 -394 -5949
rect -388 -5957 -386 -5949
rect -214 -5957 -212 -5949
rect -204 -5957 -202 -5949
rect -188 -5957 -186 -5949
rect -180 -5957 -178 -5949
rect -164 -5957 -162 -5949
rect -156 -5957 -154 -5949
rect -146 -5957 -144 -5949
rect -138 -5957 -136 -5949
rect -122 -5957 -120 -5949
rect -114 -5957 -112 -5949
rect -104 -5957 -102 -5949
rect -96 -5957 -94 -5949
rect -80 -5957 -78 -5949
rect -72 -5957 -70 -5949
rect -62 -5957 -60 -5949
rect -54 -5957 -52 -5949
rect -38 -5957 -36 -5949
rect -30 -5957 -28 -5949
rect 214 -5957 216 -5949
rect 224 -5957 226 -5949
rect 240 -5957 242 -5949
rect 248 -5957 250 -5949
rect 264 -5957 266 -5949
rect 272 -5957 274 -5949
rect 282 -5957 284 -5949
rect 290 -5957 292 -5949
rect 306 -5957 308 -5949
rect 314 -5957 316 -5949
rect 324 -5957 326 -5949
rect 332 -5957 334 -5949
rect 348 -5957 350 -5949
rect 356 -5957 358 -5949
rect 366 -5957 368 -5949
rect 374 -5957 376 -5949
rect 390 -5957 392 -5949
rect 398 -5957 400 -5949
rect 570 -5957 572 -5949
rect 580 -5957 582 -5949
rect 596 -5957 598 -5949
rect 604 -5957 606 -5949
rect 620 -5957 622 -5949
rect 628 -5957 630 -5949
rect 638 -5957 640 -5949
rect 646 -5957 648 -5949
rect 662 -5957 664 -5949
rect 670 -5957 672 -5949
rect 680 -5957 682 -5949
rect 688 -5957 690 -5949
rect 704 -5957 706 -5949
rect 712 -5957 714 -5949
rect 722 -5957 724 -5949
rect 730 -5957 732 -5949
rect 746 -5957 748 -5949
rect 754 -5957 756 -5949
rect 968 -5957 970 -5949
rect 978 -5957 980 -5949
rect 994 -5957 996 -5949
rect 1002 -5957 1004 -5949
rect 1018 -5957 1020 -5949
rect 1026 -5957 1028 -5949
rect 1036 -5957 1038 -5949
rect 1044 -5957 1046 -5949
rect 1060 -5957 1062 -5949
rect 1068 -5957 1070 -5949
rect 1078 -5957 1080 -5949
rect 1086 -5957 1088 -5949
rect 1102 -5957 1104 -5949
rect 1110 -5957 1112 -5949
rect 1120 -5957 1122 -5949
rect 1128 -5957 1130 -5949
rect 1144 -5957 1146 -5949
rect 1152 -5957 1154 -5949
rect 1326 -5957 1328 -5949
rect 1336 -5957 1338 -5949
rect 1352 -5957 1354 -5949
rect 1360 -5957 1362 -5949
rect 1376 -5957 1378 -5949
rect 1384 -5957 1386 -5949
rect 1394 -5957 1396 -5949
rect 1402 -5957 1404 -5949
rect 1418 -5957 1420 -5949
rect 1426 -5957 1428 -5949
rect 1436 -5957 1438 -5949
rect 1444 -5957 1446 -5949
rect 1460 -5957 1462 -5949
rect 1468 -5957 1470 -5949
rect 1478 -5957 1480 -5949
rect 1486 -5957 1488 -5949
rect 1502 -5957 1504 -5949
rect 1510 -5957 1512 -5949
rect 1326 -6075 1328 -6067
rect 1336 -6075 1338 -6067
rect 1352 -6075 1354 -6067
rect 1360 -6075 1362 -6067
rect 1376 -6075 1378 -6067
rect 1384 -6075 1386 -6067
rect 1394 -6075 1396 -6067
rect 1402 -6075 1404 -6067
rect 1418 -6075 1420 -6067
rect 1426 -6075 1428 -6067
rect 1436 -6075 1438 -6067
rect 1444 -6075 1446 -6067
rect 1460 -6075 1462 -6067
rect 1468 -6075 1470 -6067
rect 1478 -6075 1480 -6067
rect 1486 -6075 1488 -6067
rect 1502 -6075 1504 -6067
rect 1510 -6075 1512 -6067
<< polycontact >>
rect -1336 -1066 -1332 -1062
rect -1325 -1074 -1321 -1070
rect -1318 -1096 -1314 -1092
rect -935 -1066 -931 -1062
rect -924 -1074 -920 -1070
rect -917 -1098 -913 -1094
rect -576 -1066 -572 -1062
rect -565 -1074 -561 -1070
rect -558 -1098 -554 -1094
rect -218 -1066 -214 -1062
rect -207 -1074 -203 -1070
rect -200 -1098 -196 -1094
rect 210 -1066 214 -1062
rect 221 -1074 225 -1070
rect 228 -1111 232 -1107
rect 566 -1066 570 -1062
rect 577 -1074 581 -1070
rect 584 -1111 588 -1107
rect 964 -1066 968 -1062
rect 975 -1074 979 -1070
rect 982 -1111 986 -1107
rect 1322 -1066 1326 -1062
rect 1333 -1074 1337 -1070
rect 1340 -1111 1344 -1107
rect -1253 -1204 -1249 -1200
rect -1249 -1218 -1245 -1214
rect -1233 -1196 -1229 -1192
rect -1233 -1225 -1229 -1221
rect -1219 -1204 -1215 -1200
rect -1209 -1211 -1205 -1207
rect -1195 -1196 -1191 -1192
rect -1191 -1225 -1187 -1221
rect -1167 -1204 -1163 -1200
rect -1177 -1211 -1173 -1207
rect -1153 -1225 -1149 -1221
rect -1135 -1196 -1131 -1192
rect -1125 -1211 -1121 -1207
rect -1135 -1218 -1131 -1214
rect -1111 -1196 -1107 -1192
rect -1107 -1204 -1103 -1200
rect -1093 -1211 -1089 -1207
rect -1083 -1218 -1079 -1214
rect -1069 -1204 -1065 -1200
rect -928 -1204 -924 -1200
rect -924 -1218 -920 -1214
rect -908 -1196 -904 -1192
rect -908 -1225 -904 -1221
rect -894 -1204 -890 -1200
rect -884 -1211 -880 -1207
rect -870 -1196 -866 -1192
rect -866 -1225 -862 -1221
rect -842 -1204 -838 -1200
rect -852 -1211 -848 -1207
rect -828 -1225 -824 -1221
rect -810 -1196 -806 -1192
rect -800 -1211 -796 -1207
rect -810 -1218 -806 -1214
rect -786 -1196 -782 -1192
rect -782 -1204 -778 -1200
rect -768 -1211 -764 -1207
rect -758 -1218 -754 -1214
rect -744 -1204 -740 -1200
rect -570 -1204 -566 -1200
rect -566 -1218 -562 -1214
rect -550 -1196 -546 -1192
rect -550 -1225 -546 -1221
rect -536 -1204 -532 -1200
rect -526 -1211 -522 -1207
rect -512 -1196 -508 -1192
rect -508 -1225 -504 -1221
rect -484 -1204 -480 -1200
rect -494 -1211 -490 -1207
rect -470 -1225 -466 -1221
rect -452 -1196 -448 -1192
rect -442 -1211 -438 -1207
rect -452 -1218 -448 -1214
rect -428 -1196 -424 -1192
rect -424 -1204 -420 -1200
rect -410 -1211 -406 -1207
rect -400 -1218 -396 -1214
rect -386 -1204 -382 -1200
rect -212 -1204 -208 -1200
rect -208 -1218 -204 -1214
rect -192 -1196 -188 -1192
rect -192 -1225 -188 -1221
rect -178 -1204 -174 -1200
rect -168 -1211 -164 -1207
rect -154 -1196 -150 -1192
rect -150 -1225 -146 -1221
rect -126 -1204 -122 -1200
rect -136 -1211 -132 -1207
rect -112 -1225 -108 -1221
rect -94 -1196 -90 -1192
rect -84 -1211 -80 -1207
rect -94 -1218 -90 -1214
rect -70 -1196 -66 -1192
rect -66 -1204 -62 -1200
rect -52 -1211 -48 -1207
rect -42 -1218 -38 -1214
rect -28 -1204 -24 -1200
rect 216 -1204 220 -1200
rect 220 -1218 224 -1214
rect 236 -1196 240 -1192
rect 236 -1225 240 -1221
rect 250 -1204 254 -1200
rect 260 -1211 264 -1207
rect 274 -1196 278 -1192
rect 278 -1225 282 -1221
rect 302 -1204 306 -1200
rect 292 -1211 296 -1207
rect 316 -1225 320 -1221
rect 334 -1196 338 -1192
rect 344 -1211 348 -1207
rect 334 -1218 338 -1214
rect 358 -1196 362 -1192
rect 362 -1204 366 -1200
rect 376 -1211 380 -1207
rect 386 -1218 390 -1214
rect 400 -1204 404 -1200
rect 572 -1204 576 -1200
rect 576 -1218 580 -1214
rect 592 -1196 596 -1192
rect 592 -1225 596 -1221
rect 606 -1204 610 -1200
rect 616 -1211 620 -1207
rect 630 -1196 634 -1192
rect 634 -1225 638 -1221
rect 658 -1204 662 -1200
rect 648 -1211 652 -1207
rect 672 -1225 676 -1221
rect 690 -1196 694 -1192
rect 700 -1211 704 -1207
rect 690 -1218 694 -1214
rect 714 -1196 718 -1192
rect 718 -1204 722 -1200
rect 732 -1211 736 -1207
rect 742 -1218 746 -1214
rect 756 -1204 760 -1200
rect 970 -1204 974 -1200
rect 974 -1218 978 -1214
rect 990 -1196 994 -1192
rect 990 -1225 994 -1221
rect 1004 -1204 1008 -1200
rect 1014 -1211 1018 -1207
rect 1028 -1196 1032 -1192
rect 1032 -1225 1036 -1221
rect 1056 -1204 1060 -1200
rect 1046 -1211 1050 -1207
rect 1070 -1225 1074 -1221
rect 1088 -1196 1092 -1192
rect 1098 -1211 1102 -1207
rect 1088 -1218 1092 -1214
rect 1112 -1196 1116 -1192
rect 1116 -1204 1120 -1200
rect 1130 -1211 1134 -1207
rect 1140 -1218 1144 -1214
rect 1154 -1204 1158 -1200
rect -1338 -1296 -1334 -1292
rect -1327 -1304 -1323 -1300
rect -1320 -1326 -1316 -1322
rect -934 -1296 -930 -1292
rect -923 -1304 -919 -1300
rect -916 -1326 -912 -1322
rect -576 -1296 -572 -1292
rect -565 -1304 -561 -1300
rect -558 -1326 -554 -1322
rect -218 -1296 -214 -1292
rect -207 -1304 -203 -1300
rect -200 -1326 -196 -1322
rect 210 -1296 214 -1292
rect 221 -1304 225 -1300
rect 228 -1326 232 -1322
rect 566 -1296 570 -1292
rect 577 -1304 581 -1300
rect 584 -1326 588 -1322
rect 964 -1296 968 -1292
rect 975 -1304 979 -1300
rect 982 -1326 986 -1322
rect 1322 -1296 1326 -1292
rect 1333 -1304 1337 -1300
rect 1340 -1326 1344 -1322
rect -1249 -1434 -1245 -1430
rect -1253 -1441 -1249 -1437
rect -1233 -1421 -1229 -1417
rect -1223 -1441 -1219 -1437
rect -1209 -1434 -1205 -1430
rect -1199 -1427 -1195 -1423
rect -1189 -1434 -1185 -1430
rect -1175 -1441 -1171 -1437
rect -1171 -1455 -1167 -1451
rect -924 -1397 -920 -1393
rect -928 -1418 -924 -1414
rect -924 -1433 -920 -1429
rect -928 -1447 -924 -1443
rect -898 -1418 -894 -1414
rect -902 -1426 -898 -1422
rect -902 -1440 -898 -1436
rect -882 -1404 -878 -1400
rect -872 -1447 -868 -1443
rect -858 -1397 -854 -1393
rect -848 -1411 -844 -1407
rect -838 -1447 -834 -1443
rect -824 -1397 -820 -1393
rect -820 -1455 -816 -1451
rect -804 -1426 -800 -1422
rect -794 -1440 -790 -1436
rect -780 -1397 -776 -1393
rect -780 -1418 -776 -1414
rect -776 -1433 -772 -1429
rect -760 -1440 -756 -1436
rect -746 -1397 -742 -1393
rect -736 -1448 -732 -1444
rect -720 -1455 -716 -1451
rect -706 -1411 -702 -1407
rect -702 -1448 -698 -1444
rect -566 -1397 -562 -1393
rect -570 -1418 -566 -1414
rect -566 -1433 -562 -1429
rect -570 -1447 -566 -1443
rect -540 -1418 -536 -1414
rect -544 -1426 -540 -1422
rect -544 -1440 -540 -1436
rect -524 -1404 -520 -1400
rect -514 -1447 -510 -1443
rect -500 -1397 -496 -1393
rect -490 -1411 -486 -1407
rect -480 -1447 -476 -1443
rect -466 -1397 -462 -1393
rect -462 -1455 -458 -1451
rect -446 -1426 -442 -1422
rect -436 -1440 -432 -1436
rect -422 -1397 -418 -1393
rect -422 -1418 -418 -1414
rect -418 -1433 -414 -1429
rect -402 -1440 -398 -1436
rect -388 -1397 -384 -1393
rect -378 -1448 -374 -1444
rect -362 -1455 -358 -1451
rect -348 -1411 -344 -1407
rect -344 -1448 -340 -1444
rect -208 -1397 -204 -1393
rect -212 -1418 -208 -1414
rect -208 -1433 -204 -1429
rect -212 -1447 -208 -1443
rect -182 -1418 -178 -1414
rect -186 -1426 -182 -1422
rect -186 -1440 -182 -1436
rect -166 -1404 -162 -1400
rect -156 -1447 -152 -1443
rect -142 -1397 -138 -1393
rect -132 -1411 -128 -1407
rect -122 -1447 -118 -1443
rect -108 -1397 -104 -1393
rect -104 -1455 -100 -1451
rect -88 -1426 -84 -1422
rect -78 -1440 -74 -1436
rect -64 -1397 -60 -1393
rect -64 -1418 -60 -1414
rect -60 -1433 -56 -1429
rect -44 -1440 -40 -1436
rect -30 -1397 -26 -1393
rect -20 -1448 -16 -1444
rect -4 -1455 0 -1451
rect 10 -1411 14 -1407
rect 14 -1448 18 -1444
rect 220 -1397 224 -1393
rect 216 -1418 220 -1414
rect 220 -1433 224 -1429
rect 216 -1447 220 -1443
rect 246 -1418 250 -1414
rect 242 -1426 246 -1422
rect 242 -1440 246 -1436
rect 262 -1404 266 -1400
rect 272 -1447 276 -1443
rect 286 -1397 290 -1393
rect 296 -1411 300 -1407
rect 306 -1447 310 -1443
rect 320 -1397 324 -1393
rect 324 -1455 328 -1451
rect 340 -1426 344 -1422
rect 350 -1440 354 -1436
rect 364 -1397 368 -1393
rect 364 -1418 368 -1414
rect 368 -1433 372 -1429
rect 384 -1440 388 -1436
rect 398 -1397 402 -1393
rect 408 -1448 412 -1444
rect 424 -1455 428 -1451
rect 438 -1411 442 -1407
rect 442 -1448 446 -1444
rect 576 -1397 580 -1393
rect 572 -1418 576 -1414
rect 576 -1433 580 -1429
rect 572 -1447 576 -1443
rect 602 -1418 606 -1414
rect 598 -1426 602 -1422
rect 598 -1440 602 -1436
rect 618 -1404 622 -1400
rect 628 -1447 632 -1443
rect 642 -1397 646 -1393
rect 652 -1411 656 -1407
rect 662 -1447 666 -1443
rect 676 -1397 680 -1393
rect 680 -1455 684 -1451
rect 696 -1426 700 -1422
rect 706 -1440 710 -1436
rect 720 -1397 724 -1393
rect 720 -1418 724 -1414
rect 724 -1433 728 -1429
rect 740 -1440 744 -1436
rect 754 -1397 758 -1393
rect 764 -1448 768 -1444
rect 780 -1455 784 -1451
rect 794 -1411 798 -1407
rect 798 -1448 802 -1444
rect 974 -1397 978 -1393
rect 970 -1418 974 -1414
rect 974 -1433 978 -1429
rect 970 -1447 974 -1443
rect 1000 -1418 1004 -1414
rect 996 -1426 1000 -1422
rect 996 -1440 1000 -1436
rect 1016 -1404 1020 -1400
rect 1026 -1447 1030 -1443
rect 1040 -1397 1044 -1393
rect 1050 -1411 1054 -1407
rect 1060 -1447 1064 -1443
rect 1074 -1397 1078 -1393
rect 1078 -1455 1082 -1451
rect 1094 -1426 1098 -1422
rect 1104 -1440 1108 -1436
rect 1118 -1397 1122 -1393
rect 1118 -1418 1122 -1414
rect 1122 -1433 1126 -1429
rect 1138 -1440 1142 -1436
rect 1152 -1397 1156 -1393
rect 1162 -1448 1166 -1444
rect 1178 -1455 1182 -1451
rect 1192 -1411 1196 -1407
rect 1196 -1448 1200 -1444
rect 1332 -1434 1336 -1430
rect 1328 -1441 1332 -1437
rect 1348 -1421 1352 -1417
rect 1358 -1441 1362 -1437
rect 1372 -1434 1376 -1430
rect 1382 -1427 1386 -1423
rect 1392 -1434 1396 -1430
rect 1406 -1441 1410 -1437
rect 1410 -1455 1414 -1451
rect -1253 -1557 -1249 -1553
rect -1249 -1571 -1245 -1567
rect -1233 -1549 -1229 -1545
rect -1233 -1578 -1229 -1574
rect -1219 -1557 -1215 -1553
rect -1209 -1564 -1205 -1560
rect -1195 -1549 -1191 -1545
rect -1191 -1578 -1187 -1574
rect -1167 -1557 -1163 -1553
rect -1177 -1564 -1173 -1560
rect -1153 -1578 -1149 -1574
rect -1135 -1549 -1131 -1545
rect -1125 -1564 -1121 -1560
rect -1135 -1571 -1131 -1567
rect -1111 -1549 -1107 -1545
rect -1107 -1557 -1103 -1553
rect -1093 -1564 -1089 -1560
rect -1083 -1571 -1079 -1567
rect -1069 -1557 -1065 -1553
rect -928 -1557 -924 -1553
rect -924 -1571 -920 -1567
rect -908 -1549 -904 -1545
rect -908 -1578 -904 -1574
rect -894 -1557 -890 -1553
rect -884 -1564 -880 -1560
rect -870 -1549 -866 -1545
rect -866 -1578 -862 -1574
rect -842 -1557 -838 -1553
rect -852 -1564 -848 -1560
rect -828 -1578 -824 -1574
rect -810 -1549 -806 -1545
rect -800 -1564 -796 -1560
rect -810 -1571 -806 -1567
rect -786 -1549 -782 -1545
rect -782 -1557 -778 -1553
rect -768 -1564 -764 -1560
rect -758 -1571 -754 -1567
rect -744 -1557 -740 -1553
rect -570 -1557 -566 -1553
rect -566 -1571 -562 -1567
rect -550 -1549 -546 -1545
rect -550 -1578 -546 -1574
rect -536 -1557 -532 -1553
rect -526 -1564 -522 -1560
rect -512 -1549 -508 -1545
rect -508 -1578 -504 -1574
rect -484 -1557 -480 -1553
rect -494 -1564 -490 -1560
rect -470 -1578 -466 -1574
rect -452 -1549 -448 -1545
rect -442 -1564 -438 -1560
rect -452 -1571 -448 -1567
rect -428 -1549 -424 -1545
rect -424 -1557 -420 -1553
rect -410 -1564 -406 -1560
rect -400 -1571 -396 -1567
rect -386 -1557 -382 -1553
rect -212 -1557 -208 -1553
rect -208 -1571 -204 -1567
rect -192 -1549 -188 -1545
rect -192 -1578 -188 -1574
rect -178 -1557 -174 -1553
rect -168 -1564 -164 -1560
rect -154 -1549 -150 -1545
rect -150 -1578 -146 -1574
rect -126 -1557 -122 -1553
rect -136 -1564 -132 -1560
rect -112 -1578 -108 -1574
rect -94 -1549 -90 -1545
rect -84 -1564 -80 -1560
rect -94 -1571 -90 -1567
rect -70 -1549 -66 -1545
rect -66 -1557 -62 -1553
rect -52 -1564 -48 -1560
rect -42 -1571 -38 -1567
rect -28 -1557 -24 -1553
rect 216 -1557 220 -1553
rect 220 -1571 224 -1567
rect 236 -1549 240 -1545
rect 236 -1578 240 -1574
rect 250 -1557 254 -1553
rect 260 -1564 264 -1560
rect 274 -1549 278 -1545
rect 278 -1578 282 -1574
rect 302 -1557 306 -1553
rect 292 -1564 296 -1560
rect 316 -1578 320 -1574
rect 334 -1549 338 -1545
rect 344 -1564 348 -1560
rect 334 -1571 338 -1567
rect 358 -1549 362 -1545
rect 362 -1557 366 -1553
rect 376 -1564 380 -1560
rect 386 -1571 390 -1567
rect 400 -1557 404 -1553
rect 572 -1557 576 -1553
rect 576 -1571 580 -1567
rect 592 -1549 596 -1545
rect 592 -1578 596 -1574
rect 606 -1557 610 -1553
rect 616 -1564 620 -1560
rect 630 -1549 634 -1545
rect 634 -1578 638 -1574
rect 658 -1557 662 -1553
rect 648 -1564 652 -1560
rect 672 -1578 676 -1574
rect 690 -1549 694 -1545
rect 700 -1564 704 -1560
rect 690 -1571 694 -1567
rect 714 -1549 718 -1545
rect 718 -1557 722 -1553
rect 732 -1564 736 -1560
rect 742 -1571 746 -1567
rect 756 -1557 760 -1553
rect 970 -1557 974 -1553
rect 974 -1571 978 -1567
rect 990 -1549 994 -1545
rect 990 -1578 994 -1574
rect 1004 -1557 1008 -1553
rect 1014 -1564 1018 -1560
rect 1028 -1549 1032 -1545
rect 1032 -1578 1036 -1574
rect 1056 -1557 1060 -1553
rect 1046 -1564 1050 -1560
rect 1070 -1578 1074 -1574
rect 1088 -1549 1092 -1545
rect 1098 -1564 1102 -1560
rect 1088 -1571 1092 -1567
rect 1112 -1549 1116 -1545
rect 1116 -1557 1120 -1553
rect 1130 -1564 1134 -1560
rect 1140 -1571 1144 -1567
rect 1154 -1557 1158 -1553
rect -1253 -1678 -1249 -1674
rect -1249 -1692 -1245 -1688
rect -1233 -1670 -1229 -1666
rect -1233 -1699 -1229 -1695
rect -1219 -1678 -1215 -1674
rect -1209 -1685 -1205 -1681
rect -1195 -1670 -1191 -1666
rect -1191 -1699 -1187 -1695
rect -1167 -1678 -1163 -1674
rect -1177 -1685 -1173 -1681
rect -1153 -1699 -1149 -1695
rect -1135 -1670 -1131 -1666
rect -1125 -1685 -1121 -1681
rect -1135 -1692 -1131 -1688
rect -1111 -1670 -1107 -1666
rect -1107 -1678 -1103 -1674
rect -1093 -1685 -1089 -1681
rect -1083 -1692 -1079 -1688
rect -1069 -1678 -1065 -1674
rect -928 -1678 -924 -1674
rect -924 -1692 -920 -1688
rect -908 -1670 -904 -1666
rect -908 -1699 -904 -1695
rect -894 -1678 -890 -1674
rect -884 -1685 -880 -1681
rect -870 -1670 -866 -1666
rect -866 -1699 -862 -1695
rect -842 -1678 -838 -1674
rect -852 -1685 -848 -1681
rect -828 -1699 -824 -1695
rect -810 -1670 -806 -1666
rect -800 -1685 -796 -1681
rect -810 -1692 -806 -1688
rect -786 -1670 -782 -1666
rect -782 -1678 -778 -1674
rect -768 -1685 -764 -1681
rect -758 -1692 -754 -1688
rect -744 -1678 -740 -1674
rect -570 -1678 -566 -1674
rect -566 -1692 -562 -1688
rect -550 -1670 -546 -1666
rect -550 -1699 -546 -1695
rect -536 -1678 -532 -1674
rect -526 -1685 -522 -1681
rect -512 -1670 -508 -1666
rect -508 -1699 -504 -1695
rect -484 -1678 -480 -1674
rect -494 -1685 -490 -1681
rect -470 -1699 -466 -1695
rect -452 -1670 -448 -1666
rect -442 -1685 -438 -1681
rect -452 -1692 -448 -1688
rect -428 -1670 -424 -1666
rect -424 -1678 -420 -1674
rect -410 -1685 -406 -1681
rect -400 -1692 -396 -1688
rect -386 -1678 -382 -1674
rect -212 -1678 -208 -1674
rect -208 -1692 -204 -1688
rect -192 -1670 -188 -1666
rect -192 -1699 -188 -1695
rect -178 -1678 -174 -1674
rect -168 -1685 -164 -1681
rect -154 -1670 -150 -1666
rect -150 -1699 -146 -1695
rect -126 -1678 -122 -1674
rect -136 -1685 -132 -1681
rect -112 -1699 -108 -1695
rect -94 -1670 -90 -1666
rect -84 -1685 -80 -1681
rect -94 -1692 -90 -1688
rect -70 -1670 -66 -1666
rect -66 -1678 -62 -1674
rect -52 -1685 -48 -1681
rect -42 -1692 -38 -1688
rect -28 -1678 -24 -1674
rect 216 -1678 220 -1674
rect 220 -1692 224 -1688
rect 236 -1670 240 -1666
rect 236 -1699 240 -1695
rect 250 -1678 254 -1674
rect 260 -1685 264 -1681
rect 274 -1670 278 -1666
rect 278 -1699 282 -1695
rect 302 -1678 306 -1674
rect 292 -1685 296 -1681
rect 316 -1699 320 -1695
rect 334 -1670 338 -1666
rect 344 -1685 348 -1681
rect 334 -1692 338 -1688
rect 358 -1670 362 -1666
rect 362 -1678 366 -1674
rect 376 -1685 380 -1681
rect 386 -1692 390 -1688
rect 400 -1678 404 -1674
rect 572 -1678 576 -1674
rect 576 -1692 580 -1688
rect 592 -1670 596 -1666
rect 592 -1699 596 -1695
rect 606 -1678 610 -1674
rect 616 -1685 620 -1681
rect 630 -1670 634 -1666
rect 634 -1699 638 -1695
rect 658 -1678 662 -1674
rect 648 -1685 652 -1681
rect 672 -1699 676 -1695
rect 690 -1670 694 -1666
rect 700 -1685 704 -1681
rect 690 -1692 694 -1688
rect 714 -1670 718 -1666
rect 718 -1678 722 -1674
rect 732 -1685 736 -1681
rect 742 -1692 746 -1688
rect 756 -1678 760 -1674
rect 970 -1678 974 -1674
rect 974 -1692 978 -1688
rect 990 -1670 994 -1666
rect 990 -1699 994 -1695
rect 1004 -1678 1008 -1674
rect 1014 -1685 1018 -1681
rect 1028 -1670 1032 -1666
rect 1032 -1699 1036 -1695
rect 1056 -1678 1060 -1674
rect 1046 -1685 1050 -1681
rect 1070 -1699 1074 -1695
rect 1088 -1670 1092 -1666
rect 1098 -1685 1102 -1681
rect 1088 -1692 1092 -1688
rect 1112 -1670 1116 -1666
rect 1116 -1678 1120 -1674
rect 1130 -1685 1134 -1681
rect 1140 -1692 1144 -1688
rect 1154 -1678 1158 -1674
rect 1328 -1678 1332 -1674
rect 1332 -1692 1336 -1688
rect 1348 -1670 1352 -1666
rect 1348 -1699 1352 -1695
rect 1362 -1678 1366 -1674
rect 1372 -1685 1376 -1681
rect 1386 -1670 1390 -1666
rect 1390 -1699 1394 -1695
rect 1414 -1678 1418 -1674
rect 1404 -1685 1408 -1681
rect 1428 -1699 1432 -1695
rect 1446 -1670 1450 -1666
rect 1456 -1685 1460 -1681
rect 1446 -1692 1450 -1688
rect 1470 -1670 1474 -1666
rect 1474 -1678 1478 -1674
rect 1488 -1685 1492 -1681
rect 1498 -1692 1502 -1688
rect 1512 -1678 1516 -1674
rect -1253 -1799 -1249 -1795
rect -1249 -1813 -1245 -1809
rect -1233 -1791 -1229 -1787
rect -1233 -1820 -1229 -1816
rect -1219 -1799 -1215 -1795
rect -1209 -1806 -1205 -1802
rect -1195 -1791 -1191 -1787
rect -1191 -1820 -1187 -1816
rect -1167 -1799 -1163 -1795
rect -1177 -1806 -1173 -1802
rect -1153 -1820 -1149 -1816
rect -1135 -1791 -1131 -1787
rect -1125 -1806 -1121 -1802
rect -1135 -1813 -1131 -1809
rect -1111 -1791 -1107 -1787
rect -1107 -1799 -1103 -1795
rect -1093 -1806 -1089 -1802
rect -1083 -1813 -1079 -1809
rect -1028 -1795 -1024 -1785
rect -1069 -1799 -1065 -1795
rect -928 -1799 -924 -1795
rect -924 -1813 -920 -1809
rect -908 -1791 -904 -1787
rect -908 -1820 -904 -1816
rect -894 -1799 -890 -1795
rect -884 -1806 -880 -1802
rect -870 -1791 -866 -1787
rect -866 -1820 -862 -1816
rect -842 -1799 -838 -1795
rect -852 -1806 -848 -1802
rect -828 -1820 -824 -1816
rect -810 -1791 -806 -1787
rect -800 -1806 -796 -1802
rect -810 -1813 -806 -1809
rect -786 -1791 -782 -1787
rect -782 -1799 -778 -1795
rect -768 -1806 -764 -1802
rect -758 -1813 -754 -1809
rect -744 -1799 -740 -1795
rect -570 -1799 -566 -1795
rect -566 -1813 -562 -1809
rect -550 -1791 -546 -1787
rect -550 -1820 -546 -1816
rect -536 -1799 -532 -1795
rect -526 -1806 -522 -1802
rect -512 -1791 -508 -1787
rect -508 -1820 -504 -1816
rect -484 -1799 -480 -1795
rect -494 -1806 -490 -1802
rect -470 -1820 -466 -1816
rect -452 -1791 -448 -1787
rect -442 -1806 -438 -1802
rect -452 -1813 -448 -1809
rect -428 -1791 -424 -1787
rect -424 -1799 -420 -1795
rect -410 -1806 -406 -1802
rect -400 -1813 -396 -1809
rect -331 -1795 -327 -1785
rect -386 -1799 -382 -1795
rect -212 -1799 -208 -1795
rect -208 -1813 -204 -1809
rect -192 -1791 -188 -1787
rect -192 -1820 -188 -1816
rect -178 -1799 -174 -1795
rect -168 -1806 -164 -1802
rect -154 -1791 -150 -1787
rect -150 -1820 -146 -1816
rect -126 -1799 -122 -1795
rect -136 -1806 -132 -1802
rect -112 -1820 -108 -1816
rect -94 -1791 -90 -1787
rect -84 -1806 -80 -1802
rect -94 -1813 -90 -1809
rect -70 -1791 -66 -1787
rect -66 -1799 -62 -1795
rect -52 -1806 -48 -1802
rect -42 -1813 -38 -1809
rect -28 -1799 -24 -1795
rect 216 -1799 220 -1795
rect 220 -1813 224 -1809
rect 236 -1791 240 -1787
rect 236 -1820 240 -1816
rect 250 -1799 254 -1795
rect 260 -1806 264 -1802
rect 274 -1791 278 -1787
rect 278 -1820 282 -1816
rect 302 -1799 306 -1795
rect 292 -1806 296 -1802
rect 316 -1820 320 -1816
rect 334 -1791 338 -1787
rect 344 -1806 348 -1802
rect 334 -1813 338 -1809
rect 358 -1791 362 -1787
rect 362 -1799 366 -1795
rect 376 -1806 380 -1802
rect 386 -1813 390 -1809
rect 465 -1795 469 -1785
rect 400 -1799 404 -1795
rect 572 -1799 576 -1795
rect 576 -1813 580 -1809
rect 592 -1791 596 -1787
rect 592 -1820 596 -1816
rect 606 -1799 610 -1795
rect 616 -1806 620 -1802
rect 630 -1791 634 -1787
rect 634 -1820 638 -1816
rect 658 -1799 662 -1795
rect 648 -1806 652 -1802
rect 672 -1820 676 -1816
rect 690 -1791 694 -1787
rect 700 -1806 704 -1802
rect 690 -1813 694 -1809
rect 714 -1791 718 -1787
rect 718 -1799 722 -1795
rect 732 -1806 736 -1802
rect 742 -1813 746 -1809
rect 756 -1799 760 -1795
rect 970 -1799 974 -1795
rect 974 -1813 978 -1809
rect 990 -1791 994 -1787
rect 990 -1820 994 -1816
rect 1004 -1799 1008 -1795
rect 1014 -1806 1018 -1802
rect 1028 -1791 1032 -1787
rect 1032 -1820 1036 -1816
rect 1056 -1799 1060 -1795
rect 1046 -1806 1050 -1802
rect 1070 -1820 1074 -1816
rect 1088 -1791 1092 -1787
rect 1098 -1806 1102 -1802
rect 1088 -1813 1092 -1809
rect 1112 -1791 1116 -1787
rect 1116 -1799 1120 -1795
rect 1130 -1806 1134 -1802
rect 1140 -1813 1144 -1809
rect 1204 -1795 1208 -1785
rect 1154 -1799 1158 -1795
rect 1328 -1799 1332 -1795
rect 1332 -1813 1336 -1809
rect 1348 -1791 1352 -1787
rect 1348 -1820 1352 -1816
rect 1362 -1799 1366 -1795
rect 1372 -1806 1376 -1802
rect 1386 -1791 1390 -1787
rect 1390 -1820 1394 -1816
rect 1414 -1799 1418 -1795
rect 1404 -1806 1408 -1802
rect 1428 -1820 1432 -1816
rect 1446 -1791 1450 -1787
rect 1456 -1806 1460 -1802
rect 1446 -1813 1450 -1809
rect 1470 -1791 1474 -1787
rect 1474 -1799 1478 -1795
rect 1488 -1806 1492 -1802
rect 1498 -1813 1502 -1809
rect 1512 -1799 1516 -1795
rect -1253 -1914 -1249 -1910
rect -1249 -1928 -1245 -1924
rect -1233 -1906 -1229 -1902
rect -1233 -1935 -1229 -1931
rect -1219 -1914 -1215 -1910
rect -1209 -1921 -1205 -1917
rect -1195 -1906 -1191 -1902
rect -1191 -1935 -1187 -1931
rect -1167 -1914 -1163 -1910
rect -1177 -1921 -1173 -1917
rect -1153 -1935 -1149 -1931
rect -1135 -1906 -1131 -1902
rect -1125 -1921 -1121 -1917
rect -1135 -1928 -1131 -1924
rect -1111 -1906 -1107 -1902
rect -1107 -1914 -1103 -1910
rect -1093 -1921 -1089 -1917
rect -1083 -1928 -1079 -1924
rect -1028 -1910 -1024 -1900
rect -1069 -1914 -1065 -1910
rect -672 -1910 -668 -1900
rect -331 -1910 -327 -1900
rect 465 -1910 469 -1900
rect 842 -1910 846 -1900
rect 1204 -1910 1208 -1900
rect -1338 -2002 -1334 -1998
rect -1327 -2010 -1323 -2006
rect -1320 -2032 -1316 -2028
rect -934 -2002 -930 -1998
rect -923 -2010 -919 -2006
rect -916 -2032 -912 -2028
rect -576 -2002 -572 -1998
rect -565 -2010 -561 -2006
rect -558 -2032 -554 -2028
rect -218 -2002 -214 -1998
rect -207 -2010 -203 -2006
rect -200 -2032 -196 -2028
rect 210 -2002 214 -1998
rect 221 -2010 225 -2006
rect 228 -2032 232 -2028
rect 566 -2002 570 -1998
rect 577 -2010 581 -2006
rect 584 -2032 588 -2028
rect 964 -2002 968 -1998
rect 975 -2010 979 -2006
rect 982 -2032 986 -2028
rect 1322 -2002 1326 -1998
rect 1333 -2010 1337 -2006
rect 1340 -2032 1344 -2028
rect -1249 -2145 -1245 -2141
rect -1253 -2152 -1249 -2148
rect -1233 -2132 -1229 -2128
rect -1223 -2152 -1219 -2148
rect -1209 -2145 -1205 -2141
rect -1199 -2138 -1195 -2134
rect -1189 -2145 -1185 -2141
rect -1175 -2152 -1171 -2148
rect -1171 -2166 -1167 -2162
rect -924 -2108 -920 -2104
rect -928 -2129 -924 -2125
rect -924 -2144 -920 -2140
rect -928 -2158 -924 -2154
rect -898 -2129 -894 -2125
rect -902 -2137 -898 -2133
rect -902 -2151 -898 -2147
rect -882 -2115 -878 -2111
rect -872 -2158 -868 -2154
rect -858 -2108 -854 -2104
rect -848 -2122 -844 -2118
rect -838 -2158 -834 -2154
rect -824 -2108 -820 -2104
rect -820 -2166 -816 -2162
rect -804 -2137 -800 -2133
rect -794 -2151 -790 -2147
rect -780 -2108 -776 -2104
rect -780 -2129 -776 -2125
rect -776 -2144 -772 -2140
rect -760 -2151 -756 -2147
rect -746 -2108 -742 -2104
rect -736 -2159 -732 -2155
rect -720 -2166 -716 -2162
rect -706 -2122 -702 -2118
rect -702 -2159 -698 -2155
rect -566 -2108 -562 -2104
rect -570 -2129 -566 -2125
rect -566 -2144 -562 -2140
rect -570 -2158 -566 -2154
rect -540 -2129 -536 -2125
rect -544 -2137 -540 -2133
rect -544 -2151 -540 -2147
rect -524 -2115 -520 -2111
rect -514 -2158 -510 -2154
rect -500 -2108 -496 -2104
rect -490 -2122 -486 -2118
rect -480 -2158 -476 -2154
rect -466 -2108 -462 -2104
rect -462 -2166 -458 -2162
rect -446 -2137 -442 -2133
rect -436 -2151 -432 -2147
rect -422 -2108 -418 -2104
rect -422 -2129 -418 -2125
rect -418 -2144 -414 -2140
rect -402 -2151 -398 -2147
rect -388 -2108 -384 -2104
rect -378 -2159 -374 -2155
rect -362 -2166 -358 -2162
rect -348 -2122 -344 -2118
rect -344 -2159 -340 -2155
rect -208 -2108 -204 -2104
rect -212 -2129 -208 -2125
rect -208 -2144 -204 -2140
rect -212 -2158 -208 -2154
rect -182 -2129 -178 -2125
rect -186 -2137 -182 -2133
rect -186 -2151 -182 -2147
rect -166 -2115 -162 -2111
rect -156 -2158 -152 -2154
rect -142 -2108 -138 -2104
rect -132 -2122 -128 -2118
rect -122 -2158 -118 -2154
rect -108 -2108 -104 -2104
rect -104 -2166 -100 -2162
rect -88 -2137 -84 -2133
rect -78 -2151 -74 -2147
rect -64 -2108 -60 -2104
rect -64 -2129 -60 -2125
rect -60 -2144 -56 -2140
rect -44 -2151 -40 -2147
rect -30 -2108 -26 -2104
rect -20 -2159 -16 -2155
rect -4 -2166 0 -2162
rect 10 -2122 14 -2118
rect 14 -2159 18 -2155
rect 220 -2108 224 -2104
rect 216 -2129 220 -2125
rect 220 -2144 224 -2140
rect 216 -2158 220 -2154
rect 246 -2129 250 -2125
rect 242 -2137 246 -2133
rect 242 -2151 246 -2147
rect 262 -2115 266 -2111
rect 272 -2158 276 -2154
rect 286 -2108 290 -2104
rect 296 -2122 300 -2118
rect 306 -2158 310 -2154
rect 320 -2108 324 -2104
rect 324 -2166 328 -2162
rect 340 -2137 344 -2133
rect 350 -2151 354 -2147
rect 364 -2108 368 -2104
rect 364 -2129 368 -2125
rect 368 -2144 372 -2140
rect 384 -2151 388 -2147
rect 398 -2108 402 -2104
rect 408 -2159 412 -2155
rect 424 -2166 428 -2162
rect 438 -2122 442 -2118
rect 442 -2159 446 -2155
rect 576 -2108 580 -2104
rect 572 -2129 576 -2125
rect 576 -2144 580 -2140
rect 572 -2158 576 -2154
rect 602 -2129 606 -2125
rect 598 -2137 602 -2133
rect 598 -2151 602 -2147
rect 618 -2115 622 -2111
rect 628 -2158 632 -2154
rect 642 -2108 646 -2104
rect 652 -2122 656 -2118
rect 662 -2158 666 -2154
rect 676 -2108 680 -2104
rect 680 -2166 684 -2162
rect 696 -2137 700 -2133
rect 706 -2151 710 -2147
rect 720 -2108 724 -2104
rect 720 -2129 724 -2125
rect 724 -2144 728 -2140
rect 740 -2151 744 -2147
rect 754 -2108 758 -2104
rect 764 -2159 768 -2155
rect 780 -2166 784 -2162
rect 794 -2122 798 -2118
rect 798 -2159 802 -2155
rect 974 -2108 978 -2104
rect 970 -2129 974 -2125
rect 974 -2144 978 -2140
rect 970 -2158 974 -2154
rect 1000 -2129 1004 -2125
rect 996 -2137 1000 -2133
rect 996 -2151 1000 -2147
rect 1016 -2115 1020 -2111
rect 1026 -2158 1030 -2154
rect 1040 -2108 1044 -2104
rect 1050 -2122 1054 -2118
rect 1060 -2158 1064 -2154
rect 1074 -2108 1078 -2104
rect 1078 -2166 1082 -2162
rect 1094 -2137 1098 -2133
rect 1104 -2151 1108 -2147
rect 1118 -2108 1122 -2104
rect 1118 -2129 1122 -2125
rect 1122 -2144 1126 -2140
rect 1138 -2151 1142 -2147
rect 1152 -2108 1156 -2104
rect 1162 -2159 1166 -2155
rect 1178 -2166 1182 -2162
rect 1192 -2122 1196 -2118
rect 1196 -2159 1200 -2155
rect 1332 -2108 1336 -2104
rect 1328 -2129 1332 -2125
rect 1332 -2144 1336 -2140
rect 1328 -2158 1332 -2154
rect 1358 -2129 1362 -2125
rect 1354 -2137 1358 -2133
rect 1354 -2151 1358 -2147
rect 1374 -2115 1378 -2111
rect 1384 -2158 1388 -2154
rect 1398 -2108 1402 -2104
rect 1408 -2122 1412 -2118
rect 1418 -2158 1422 -2154
rect 1432 -2108 1436 -2104
rect 1436 -2166 1440 -2162
rect 1452 -2137 1456 -2133
rect 1462 -2151 1466 -2147
rect 1476 -2108 1480 -2104
rect 1476 -2129 1480 -2125
rect 1480 -2144 1484 -2140
rect 1496 -2151 1500 -2147
rect 1510 -2108 1514 -2104
rect 1520 -2159 1524 -2155
rect 1536 -2166 1540 -2162
rect 1550 -2122 1554 -2118
rect 1554 -2159 1558 -2155
rect -1257 -2289 -1253 -2285
rect -1253 -2303 -1249 -2299
rect -1237 -2281 -1233 -2277
rect -1237 -2310 -1233 -2306
rect -1223 -2289 -1219 -2285
rect -1213 -2296 -1209 -2292
rect -1199 -2281 -1195 -2277
rect -1195 -2310 -1191 -2306
rect -1171 -2289 -1167 -2285
rect -1181 -2296 -1177 -2292
rect -1157 -2310 -1153 -2306
rect -1139 -2281 -1135 -2277
rect -1129 -2296 -1125 -2292
rect -1139 -2303 -1135 -2299
rect -1115 -2281 -1111 -2277
rect -1111 -2289 -1107 -2285
rect -1097 -2296 -1093 -2292
rect -1087 -2303 -1083 -2299
rect -1073 -2289 -1069 -2285
rect -928 -2289 -924 -2285
rect -924 -2303 -920 -2299
rect -908 -2281 -904 -2277
rect -908 -2310 -904 -2306
rect -894 -2289 -890 -2285
rect -884 -2296 -880 -2292
rect -870 -2281 -866 -2277
rect -866 -2310 -862 -2306
rect -842 -2289 -838 -2285
rect -852 -2296 -848 -2292
rect -828 -2310 -824 -2306
rect -810 -2281 -806 -2277
rect -800 -2296 -796 -2292
rect -810 -2303 -806 -2299
rect -786 -2281 -782 -2277
rect -782 -2289 -778 -2285
rect -768 -2296 -764 -2292
rect -758 -2303 -754 -2299
rect -744 -2289 -740 -2285
rect -570 -2289 -566 -2285
rect -566 -2303 -562 -2299
rect -550 -2281 -546 -2277
rect -550 -2310 -546 -2306
rect -536 -2289 -532 -2285
rect -526 -2296 -522 -2292
rect -512 -2281 -508 -2277
rect -508 -2310 -504 -2306
rect -484 -2289 -480 -2285
rect -494 -2296 -490 -2292
rect -470 -2310 -466 -2306
rect -452 -2281 -448 -2277
rect -442 -2296 -438 -2292
rect -452 -2303 -448 -2299
rect -428 -2281 -424 -2277
rect -424 -2289 -420 -2285
rect -410 -2296 -406 -2292
rect -400 -2303 -396 -2299
rect -386 -2289 -382 -2285
rect -212 -2289 -208 -2285
rect -208 -2303 -204 -2299
rect -192 -2281 -188 -2277
rect -192 -2310 -188 -2306
rect -178 -2289 -174 -2285
rect -168 -2296 -164 -2292
rect -154 -2281 -150 -2277
rect -150 -2310 -146 -2306
rect -126 -2289 -122 -2285
rect -136 -2296 -132 -2292
rect -112 -2310 -108 -2306
rect -94 -2281 -90 -2277
rect -84 -2296 -80 -2292
rect -94 -2303 -90 -2299
rect -70 -2281 -66 -2277
rect -66 -2289 -62 -2285
rect -52 -2296 -48 -2292
rect -42 -2303 -38 -2299
rect -28 -2289 -24 -2285
rect 216 -2289 220 -2285
rect 220 -2303 224 -2299
rect 236 -2281 240 -2277
rect 236 -2310 240 -2306
rect 250 -2289 254 -2285
rect 260 -2296 264 -2292
rect 274 -2281 278 -2277
rect 278 -2310 282 -2306
rect 302 -2289 306 -2285
rect 292 -2296 296 -2292
rect 316 -2310 320 -2306
rect 334 -2281 338 -2277
rect 344 -2296 348 -2292
rect 334 -2303 338 -2299
rect 358 -2281 362 -2277
rect 362 -2289 366 -2285
rect 376 -2296 380 -2292
rect 386 -2303 390 -2299
rect 400 -2289 404 -2285
rect 572 -2289 576 -2285
rect 576 -2303 580 -2299
rect 592 -2281 596 -2277
rect 592 -2310 596 -2306
rect 606 -2289 610 -2285
rect 616 -2296 620 -2292
rect 630 -2281 634 -2277
rect 634 -2310 638 -2306
rect 658 -2289 662 -2285
rect 648 -2296 652 -2292
rect 672 -2310 676 -2306
rect 690 -2281 694 -2277
rect 700 -2296 704 -2292
rect 690 -2303 694 -2299
rect 714 -2281 718 -2277
rect 718 -2289 722 -2285
rect 732 -2296 736 -2292
rect 742 -2303 746 -2299
rect 756 -2289 760 -2285
rect -1257 -2420 -1253 -2416
rect -1253 -2434 -1249 -2430
rect -1237 -2412 -1233 -2408
rect -1237 -2441 -1233 -2437
rect -1223 -2420 -1219 -2416
rect -1213 -2427 -1209 -2423
rect -1199 -2412 -1195 -2408
rect -1195 -2441 -1191 -2437
rect -1171 -2420 -1167 -2416
rect -1181 -2427 -1177 -2423
rect -1157 -2441 -1153 -2437
rect -1139 -2412 -1135 -2408
rect -1129 -2427 -1125 -2423
rect -1139 -2434 -1135 -2430
rect -1115 -2412 -1111 -2408
rect -1111 -2420 -1107 -2416
rect -1097 -2427 -1093 -2423
rect -1087 -2434 -1083 -2430
rect -1073 -2420 -1069 -2416
rect -928 -2420 -924 -2416
rect -924 -2434 -920 -2430
rect -908 -2412 -904 -2408
rect -908 -2441 -904 -2437
rect -894 -2420 -890 -2416
rect -884 -2427 -880 -2423
rect -870 -2412 -866 -2408
rect -866 -2441 -862 -2437
rect -842 -2420 -838 -2416
rect -852 -2427 -848 -2423
rect -828 -2441 -824 -2437
rect -810 -2412 -806 -2408
rect -800 -2427 -796 -2423
rect -810 -2434 -806 -2430
rect -786 -2412 -782 -2408
rect -782 -2420 -778 -2416
rect -768 -2427 -764 -2423
rect -758 -2434 -754 -2430
rect -744 -2420 -740 -2416
rect -570 -2420 -566 -2416
rect -566 -2434 -562 -2430
rect -550 -2412 -546 -2408
rect -550 -2441 -546 -2437
rect -536 -2420 -532 -2416
rect -526 -2427 -522 -2423
rect -512 -2412 -508 -2408
rect -508 -2441 -504 -2437
rect -484 -2420 -480 -2416
rect -494 -2427 -490 -2423
rect -470 -2441 -466 -2437
rect -452 -2412 -448 -2408
rect -442 -2427 -438 -2423
rect -452 -2434 -448 -2430
rect -428 -2412 -424 -2408
rect -424 -2420 -420 -2416
rect -410 -2427 -406 -2423
rect -400 -2434 -396 -2430
rect -386 -2420 -382 -2416
rect -212 -2420 -208 -2416
rect -208 -2434 -204 -2430
rect -192 -2412 -188 -2408
rect -192 -2441 -188 -2437
rect -178 -2420 -174 -2416
rect -168 -2427 -164 -2423
rect -154 -2412 -150 -2408
rect -150 -2441 -146 -2437
rect -126 -2420 -122 -2416
rect -136 -2427 -132 -2423
rect -112 -2441 -108 -2437
rect -94 -2412 -90 -2408
rect -84 -2427 -80 -2423
rect -94 -2434 -90 -2430
rect -70 -2412 -66 -2408
rect -66 -2420 -62 -2416
rect -52 -2427 -48 -2423
rect -42 -2434 -38 -2430
rect -28 -2420 -24 -2416
rect 216 -2420 220 -2416
rect 220 -2434 224 -2430
rect 236 -2412 240 -2408
rect 236 -2441 240 -2437
rect 250 -2420 254 -2416
rect 260 -2427 264 -2423
rect 274 -2412 278 -2408
rect 278 -2441 282 -2437
rect 302 -2420 306 -2416
rect 292 -2427 296 -2423
rect 316 -2441 320 -2437
rect 334 -2412 338 -2408
rect 344 -2427 348 -2423
rect 334 -2434 338 -2430
rect 358 -2412 362 -2408
rect 362 -2420 366 -2416
rect 376 -2427 380 -2423
rect 386 -2434 390 -2430
rect 400 -2420 404 -2416
rect 572 -2420 576 -2416
rect 576 -2434 580 -2430
rect 592 -2412 596 -2408
rect 592 -2441 596 -2437
rect 606 -2420 610 -2416
rect 616 -2427 620 -2423
rect 630 -2412 634 -2408
rect 634 -2441 638 -2437
rect 658 -2420 662 -2416
rect 648 -2427 652 -2423
rect 672 -2441 676 -2437
rect 690 -2412 694 -2408
rect 700 -2427 704 -2423
rect 690 -2434 694 -2430
rect 714 -2412 718 -2408
rect 718 -2420 722 -2416
rect 732 -2427 736 -2423
rect 742 -2434 746 -2430
rect 756 -2420 760 -2416
rect 970 -2420 974 -2416
rect 974 -2434 978 -2430
rect 990 -2412 994 -2408
rect 990 -2441 994 -2437
rect 1004 -2420 1008 -2416
rect 1014 -2427 1018 -2423
rect 1028 -2412 1032 -2408
rect 1032 -2441 1036 -2437
rect 1056 -2420 1060 -2416
rect 1046 -2427 1050 -2423
rect 1070 -2441 1074 -2437
rect 1088 -2412 1092 -2408
rect 1098 -2427 1102 -2423
rect 1088 -2434 1092 -2430
rect 1112 -2412 1116 -2408
rect 1116 -2420 1120 -2416
rect 1130 -2427 1134 -2423
rect 1140 -2434 1144 -2430
rect 1154 -2420 1158 -2416
rect 1328 -2420 1332 -2416
rect 1332 -2434 1336 -2430
rect 1348 -2412 1352 -2408
rect 1348 -2441 1352 -2437
rect 1362 -2420 1366 -2416
rect 1372 -2427 1376 -2423
rect 1386 -2412 1390 -2408
rect 1390 -2441 1394 -2437
rect 1414 -2420 1418 -2416
rect 1404 -2427 1408 -2423
rect 1428 -2441 1432 -2437
rect 1446 -2412 1450 -2408
rect 1456 -2427 1460 -2423
rect 1446 -2434 1450 -2430
rect 1470 -2412 1474 -2408
rect 1474 -2420 1478 -2416
rect 1488 -2427 1492 -2423
rect 1498 -2434 1502 -2430
rect 1512 -2420 1516 -2416
rect -1257 -2551 -1253 -2547
rect -1253 -2565 -1249 -2561
rect -1237 -2543 -1233 -2539
rect -1237 -2572 -1233 -2568
rect -1223 -2551 -1219 -2547
rect -1213 -2558 -1209 -2554
rect -1199 -2543 -1195 -2539
rect -1195 -2572 -1191 -2568
rect -1171 -2551 -1167 -2547
rect -1181 -2558 -1177 -2554
rect -1157 -2572 -1153 -2568
rect -1139 -2543 -1135 -2539
rect -1129 -2558 -1125 -2554
rect -1139 -2565 -1135 -2561
rect -1115 -2543 -1111 -2539
rect -1111 -2551 -1107 -2547
rect -1097 -2558 -1093 -2554
rect -1087 -2565 -1083 -2561
rect -1073 -2551 -1069 -2547
rect -928 -2551 -924 -2547
rect -924 -2565 -920 -2561
rect -908 -2543 -904 -2539
rect -908 -2572 -904 -2568
rect -894 -2551 -890 -2547
rect -884 -2558 -880 -2554
rect -870 -2543 -866 -2539
rect -866 -2572 -862 -2568
rect -842 -2551 -838 -2547
rect -852 -2558 -848 -2554
rect -828 -2572 -824 -2568
rect -810 -2543 -806 -2539
rect -800 -2558 -796 -2554
rect -810 -2565 -806 -2561
rect -786 -2543 -782 -2539
rect -782 -2551 -778 -2547
rect -768 -2558 -764 -2554
rect -758 -2565 -754 -2561
rect -744 -2551 -740 -2547
rect -570 -2551 -566 -2547
rect -566 -2565 -562 -2561
rect -550 -2543 -546 -2539
rect -550 -2572 -546 -2568
rect -536 -2551 -532 -2547
rect -526 -2558 -522 -2554
rect -512 -2543 -508 -2539
rect -508 -2572 -504 -2568
rect -484 -2551 -480 -2547
rect -494 -2558 -490 -2554
rect -470 -2572 -466 -2568
rect -452 -2543 -448 -2539
rect -442 -2558 -438 -2554
rect -452 -2565 -448 -2561
rect -428 -2543 -424 -2539
rect -424 -2551 -420 -2547
rect -410 -2558 -406 -2554
rect -400 -2565 -396 -2561
rect -386 -2551 -382 -2547
rect -212 -2551 -208 -2547
rect -208 -2565 -204 -2561
rect -192 -2543 -188 -2539
rect -192 -2572 -188 -2568
rect -178 -2551 -174 -2547
rect -168 -2558 -164 -2554
rect -154 -2543 -150 -2539
rect -150 -2572 -146 -2568
rect -126 -2551 -122 -2547
rect -136 -2558 -132 -2554
rect -112 -2572 -108 -2568
rect -94 -2543 -90 -2539
rect -84 -2558 -80 -2554
rect -94 -2565 -90 -2561
rect -70 -2543 -66 -2539
rect -66 -2551 -62 -2547
rect -52 -2558 -48 -2554
rect -42 -2565 -38 -2561
rect -28 -2551 -24 -2547
rect 91 -2551 95 -2537
rect 216 -2551 220 -2547
rect 220 -2565 224 -2561
rect 236 -2543 240 -2539
rect 236 -2572 240 -2568
rect 250 -2551 254 -2547
rect 260 -2558 264 -2554
rect 274 -2543 278 -2539
rect 278 -2572 282 -2568
rect 302 -2551 306 -2547
rect 292 -2558 296 -2554
rect 316 -2572 320 -2568
rect 334 -2543 338 -2539
rect 344 -2558 348 -2554
rect 334 -2565 338 -2561
rect 358 -2543 362 -2539
rect 362 -2551 366 -2547
rect 376 -2558 380 -2554
rect 386 -2565 390 -2561
rect 400 -2551 404 -2547
rect 572 -2551 576 -2547
rect 576 -2565 580 -2561
rect 592 -2543 596 -2539
rect 592 -2572 596 -2568
rect 606 -2551 610 -2547
rect 616 -2558 620 -2554
rect 630 -2543 634 -2539
rect 634 -2572 638 -2568
rect 658 -2551 662 -2547
rect 648 -2558 652 -2554
rect 672 -2572 676 -2568
rect 690 -2543 694 -2539
rect 700 -2558 704 -2554
rect 690 -2565 694 -2561
rect 714 -2543 718 -2539
rect 718 -2551 722 -2547
rect 732 -2558 736 -2554
rect 742 -2565 746 -2561
rect 756 -2551 760 -2547
rect 970 -2551 974 -2547
rect 974 -2565 978 -2561
rect 990 -2543 994 -2539
rect 990 -2572 994 -2568
rect 1004 -2551 1008 -2547
rect 1014 -2558 1018 -2554
rect 1028 -2543 1032 -2539
rect 1032 -2572 1036 -2568
rect 1056 -2551 1060 -2547
rect 1046 -2558 1050 -2554
rect 1070 -2572 1074 -2568
rect 1088 -2543 1092 -2539
rect 1098 -2558 1102 -2554
rect 1088 -2565 1092 -2561
rect 1112 -2543 1116 -2539
rect 1116 -2551 1120 -2547
rect 1130 -2558 1134 -2554
rect 1140 -2565 1144 -2561
rect 1154 -2551 1158 -2547
rect 1328 -2551 1332 -2547
rect 1332 -2565 1336 -2561
rect 1348 -2543 1352 -2539
rect 1348 -2572 1352 -2568
rect 1362 -2551 1366 -2547
rect 1372 -2558 1376 -2554
rect 1386 -2543 1390 -2539
rect 1390 -2572 1394 -2568
rect 1414 -2551 1418 -2547
rect 1404 -2558 1408 -2554
rect 1428 -2572 1432 -2568
rect 1446 -2543 1450 -2539
rect 1456 -2558 1460 -2554
rect 1446 -2565 1450 -2561
rect 1470 -2543 1474 -2539
rect 1474 -2551 1478 -2547
rect 1488 -2558 1492 -2554
rect 1498 -2565 1502 -2561
rect 1512 -2551 1516 -2547
rect -1257 -2663 -1253 -2659
rect -1253 -2677 -1249 -2673
rect -1237 -2655 -1233 -2651
rect -1237 -2684 -1233 -2680
rect -1223 -2663 -1219 -2659
rect -1213 -2670 -1209 -2666
rect -1199 -2655 -1195 -2651
rect -1195 -2684 -1191 -2680
rect -1171 -2663 -1167 -2659
rect -1181 -2670 -1177 -2666
rect -1157 -2684 -1153 -2680
rect -1139 -2655 -1135 -2651
rect -1129 -2670 -1125 -2666
rect -1139 -2677 -1135 -2673
rect -1115 -2655 -1111 -2651
rect -1111 -2663 -1107 -2659
rect -1097 -2670 -1093 -2666
rect -1087 -2677 -1083 -2673
rect -1073 -2663 -1069 -2659
rect -928 -2663 -924 -2659
rect -924 -2677 -920 -2673
rect -908 -2655 -904 -2651
rect -908 -2684 -904 -2680
rect -894 -2663 -890 -2659
rect -884 -2670 -880 -2666
rect -870 -2655 -866 -2651
rect -866 -2684 -862 -2680
rect -842 -2663 -838 -2659
rect -852 -2670 -848 -2666
rect -828 -2684 -824 -2680
rect -810 -2655 -806 -2651
rect -800 -2670 -796 -2666
rect -810 -2677 -806 -2673
rect -786 -2655 -782 -2651
rect -782 -2663 -778 -2659
rect -768 -2670 -764 -2666
rect -758 -2677 -754 -2673
rect -744 -2663 -740 -2659
rect -1338 -2752 -1334 -2748
rect -1327 -2760 -1323 -2756
rect -1320 -2782 -1316 -2778
rect -934 -2752 -930 -2748
rect -923 -2760 -919 -2756
rect -916 -2782 -912 -2778
rect -576 -2752 -572 -2748
rect -565 -2760 -561 -2756
rect -558 -2782 -554 -2778
rect -218 -2752 -214 -2748
rect -207 -2760 -203 -2756
rect -200 -2782 -196 -2778
rect 210 -2752 214 -2748
rect 221 -2760 225 -2756
rect 228 -2782 232 -2778
rect 566 -2752 570 -2748
rect 577 -2760 581 -2756
rect 584 -2782 588 -2778
rect 964 -2752 968 -2748
rect 975 -2760 979 -2756
rect 982 -2782 986 -2778
rect 1322 -2752 1326 -2748
rect 1333 -2760 1337 -2756
rect 1340 -2782 1344 -2778
rect -1253 -2895 -1249 -2891
rect -1257 -2902 -1253 -2898
rect -1237 -2882 -1233 -2878
rect -1227 -2902 -1223 -2898
rect -1213 -2895 -1209 -2891
rect -1203 -2888 -1199 -2884
rect -1193 -2895 -1189 -2891
rect -1179 -2902 -1175 -2898
rect -1175 -2916 -1171 -2912
rect -924 -2858 -920 -2854
rect -928 -2879 -924 -2875
rect -924 -2894 -920 -2890
rect -928 -2908 -924 -2904
rect -898 -2879 -894 -2875
rect -902 -2887 -898 -2883
rect -902 -2901 -898 -2897
rect -882 -2865 -878 -2861
rect -872 -2908 -868 -2904
rect -858 -2858 -854 -2854
rect -848 -2872 -844 -2868
rect -838 -2908 -834 -2904
rect -824 -2858 -820 -2854
rect -820 -2916 -816 -2912
rect -804 -2887 -800 -2883
rect -794 -2901 -790 -2897
rect -780 -2858 -776 -2854
rect -780 -2879 -776 -2875
rect -776 -2894 -772 -2890
rect -760 -2901 -756 -2897
rect -746 -2858 -742 -2854
rect -736 -2909 -732 -2905
rect -720 -2916 -716 -2912
rect -706 -2872 -702 -2868
rect -702 -2909 -698 -2905
rect -566 -2858 -562 -2854
rect -570 -2879 -566 -2875
rect -566 -2894 -562 -2890
rect -570 -2908 -566 -2904
rect -540 -2879 -536 -2875
rect -544 -2887 -540 -2883
rect -544 -2901 -540 -2897
rect -524 -2865 -520 -2861
rect -514 -2908 -510 -2904
rect -500 -2858 -496 -2854
rect -490 -2872 -486 -2868
rect -480 -2908 -476 -2904
rect -466 -2858 -462 -2854
rect -462 -2916 -458 -2912
rect -446 -2887 -442 -2883
rect -436 -2901 -432 -2897
rect -422 -2858 -418 -2854
rect -422 -2879 -418 -2875
rect -418 -2894 -414 -2890
rect -402 -2901 -398 -2897
rect -388 -2858 -384 -2854
rect -378 -2909 -374 -2905
rect -362 -2916 -358 -2912
rect -348 -2872 -344 -2868
rect -344 -2909 -340 -2905
rect -208 -2858 -204 -2854
rect -212 -2879 -208 -2875
rect -208 -2894 -204 -2890
rect -212 -2908 -208 -2904
rect -182 -2879 -178 -2875
rect -186 -2887 -182 -2883
rect -186 -2901 -182 -2897
rect -166 -2865 -162 -2861
rect -156 -2908 -152 -2904
rect -142 -2858 -138 -2854
rect -132 -2872 -128 -2868
rect -122 -2908 -118 -2904
rect -108 -2858 -104 -2854
rect -104 -2916 -100 -2912
rect -88 -2887 -84 -2883
rect -78 -2901 -74 -2897
rect -64 -2858 -60 -2854
rect -64 -2879 -60 -2875
rect -60 -2894 -56 -2890
rect -44 -2901 -40 -2897
rect -30 -2858 -26 -2854
rect -20 -2909 -16 -2905
rect -4 -2916 0 -2912
rect 10 -2872 14 -2868
rect 14 -2909 18 -2905
rect 220 -2858 224 -2854
rect 216 -2879 220 -2875
rect 220 -2894 224 -2890
rect 216 -2908 220 -2904
rect 246 -2879 250 -2875
rect 242 -2887 246 -2883
rect 242 -2901 246 -2897
rect 262 -2865 266 -2861
rect 272 -2908 276 -2904
rect 286 -2858 290 -2854
rect 296 -2872 300 -2868
rect 306 -2908 310 -2904
rect 320 -2858 324 -2854
rect 324 -2916 328 -2912
rect 340 -2887 344 -2883
rect 350 -2901 354 -2897
rect 364 -2858 368 -2854
rect 364 -2879 368 -2875
rect 368 -2894 372 -2890
rect 384 -2901 388 -2897
rect 398 -2858 402 -2854
rect 408 -2909 412 -2905
rect 424 -2916 428 -2912
rect 438 -2872 442 -2868
rect 442 -2909 446 -2905
rect 576 -2858 580 -2854
rect 572 -2879 576 -2875
rect 576 -2894 580 -2890
rect 572 -2908 576 -2904
rect 602 -2879 606 -2875
rect 598 -2887 602 -2883
rect 598 -2901 602 -2897
rect 618 -2865 622 -2861
rect 628 -2908 632 -2904
rect 642 -2858 646 -2854
rect 652 -2872 656 -2868
rect 662 -2908 666 -2904
rect 676 -2858 680 -2854
rect 680 -2916 684 -2912
rect 696 -2887 700 -2883
rect 706 -2901 710 -2897
rect 720 -2858 724 -2854
rect 720 -2879 724 -2875
rect 724 -2894 728 -2890
rect 740 -2901 744 -2897
rect 754 -2858 758 -2854
rect 764 -2909 768 -2905
rect 780 -2916 784 -2912
rect 794 -2872 798 -2868
rect 798 -2909 802 -2905
rect 974 -2858 978 -2854
rect 970 -2879 974 -2875
rect 974 -2894 978 -2890
rect 970 -2908 974 -2904
rect 1000 -2879 1004 -2875
rect 996 -2887 1000 -2883
rect 996 -2901 1000 -2897
rect 1016 -2865 1020 -2861
rect 1026 -2908 1030 -2904
rect 1040 -2858 1044 -2854
rect 1050 -2872 1054 -2868
rect 1060 -2908 1064 -2904
rect 1074 -2858 1078 -2854
rect 1078 -2916 1082 -2912
rect 1094 -2887 1098 -2883
rect 1104 -2901 1108 -2897
rect 1118 -2858 1122 -2854
rect 1118 -2879 1122 -2875
rect 1122 -2894 1126 -2890
rect 1138 -2901 1142 -2897
rect 1152 -2858 1156 -2854
rect 1162 -2909 1166 -2905
rect 1178 -2916 1182 -2912
rect 1192 -2872 1196 -2868
rect 1196 -2909 1200 -2905
rect 1332 -2858 1336 -2854
rect 1328 -2879 1332 -2875
rect 1332 -2894 1336 -2890
rect 1328 -2908 1332 -2904
rect 1358 -2879 1362 -2875
rect 1354 -2887 1358 -2883
rect 1354 -2901 1358 -2897
rect 1374 -2865 1378 -2861
rect 1384 -2908 1388 -2904
rect 1398 -2858 1402 -2854
rect 1408 -2872 1412 -2868
rect 1418 -2908 1422 -2904
rect 1432 -2858 1436 -2854
rect 1436 -2916 1440 -2912
rect 1452 -2887 1456 -2883
rect 1462 -2901 1466 -2897
rect 1476 -2858 1480 -2854
rect 1476 -2879 1480 -2875
rect 1480 -2894 1484 -2890
rect 1496 -2901 1500 -2897
rect 1510 -2858 1514 -2854
rect 1520 -2909 1524 -2905
rect 1536 -2916 1540 -2912
rect 1550 -2872 1554 -2868
rect 1554 -2909 1558 -2905
rect -1257 -3014 -1253 -3010
rect -1253 -3028 -1249 -3024
rect -1237 -3006 -1233 -3002
rect -1237 -3035 -1233 -3031
rect -1223 -3014 -1219 -3010
rect -1213 -3021 -1209 -3017
rect -1199 -3006 -1195 -3002
rect -1195 -3035 -1191 -3031
rect -1171 -3014 -1167 -3010
rect -1181 -3021 -1177 -3017
rect -1157 -3035 -1153 -3031
rect -1139 -3006 -1135 -3002
rect -1129 -3021 -1125 -3017
rect -1139 -3028 -1135 -3024
rect -1115 -3006 -1111 -3002
rect -1111 -3014 -1107 -3010
rect -1097 -3021 -1093 -3017
rect -1087 -3028 -1083 -3024
rect -1073 -3014 -1069 -3010
rect -1025 -3011 -1021 -3001
rect -928 -3014 -924 -3010
rect -924 -3028 -920 -3024
rect -908 -3006 -904 -3002
rect -908 -3035 -904 -3031
rect -894 -3014 -890 -3010
rect -884 -3021 -880 -3017
rect -870 -3006 -866 -3002
rect -866 -3035 -862 -3031
rect -842 -3014 -838 -3010
rect -852 -3021 -848 -3017
rect -828 -3035 -824 -3031
rect -810 -3006 -806 -3002
rect -800 -3021 -796 -3017
rect -810 -3028 -806 -3024
rect -786 -3006 -782 -3002
rect -782 -3014 -778 -3010
rect -768 -3021 -764 -3017
rect -758 -3028 -754 -3024
rect -671 -3010 -667 -3000
rect -744 -3014 -740 -3010
rect -570 -3014 -566 -3010
rect -566 -3028 -562 -3024
rect -550 -3006 -546 -3002
rect -550 -3035 -546 -3031
rect -536 -3014 -532 -3010
rect -526 -3021 -522 -3017
rect -512 -3006 -508 -3002
rect -508 -3035 -504 -3031
rect -484 -3014 -480 -3010
rect -494 -3021 -490 -3017
rect -470 -3035 -466 -3031
rect -452 -3006 -448 -3002
rect -442 -3021 -438 -3017
rect -452 -3028 -448 -3024
rect -428 -3006 -424 -3002
rect -424 -3014 -420 -3010
rect -410 -3021 -406 -3017
rect -400 -3028 -396 -3024
rect -386 -3014 -382 -3010
rect -328 -3012 -324 -3002
rect -212 -3014 -208 -3010
rect -208 -3028 -204 -3024
rect -192 -3006 -188 -3002
rect -192 -3035 -188 -3031
rect -178 -3014 -174 -3010
rect -168 -3021 -164 -3017
rect -154 -3006 -150 -3002
rect -150 -3035 -146 -3031
rect -126 -3014 -122 -3010
rect -136 -3021 -132 -3017
rect -112 -3035 -108 -3031
rect -94 -3006 -90 -3002
rect -84 -3021 -80 -3017
rect -94 -3028 -90 -3024
rect -70 -3006 -66 -3002
rect -66 -3014 -62 -3010
rect -52 -3021 -48 -3017
rect -42 -3028 -38 -3024
rect -28 -3014 -24 -3010
rect 216 -3014 220 -3010
rect 220 -3028 224 -3024
rect 236 -3006 240 -3002
rect 236 -3035 240 -3031
rect 250 -3014 254 -3010
rect 260 -3021 264 -3017
rect 274 -3006 278 -3002
rect 278 -3035 282 -3031
rect 302 -3014 306 -3010
rect 292 -3021 296 -3017
rect 316 -3035 320 -3031
rect 334 -3006 338 -3002
rect 344 -3021 348 -3017
rect 334 -3028 338 -3024
rect 358 -3006 362 -3002
rect 362 -3014 366 -3010
rect 376 -3021 380 -3017
rect 386 -3028 390 -3024
rect 473 -3010 477 -3000
rect 400 -3014 404 -3010
rect 842 -3010 846 -3000
rect 1200 -3011 1204 -3001
rect -1257 -3130 -1253 -3126
rect -1253 -3144 -1249 -3140
rect -1237 -3122 -1233 -3118
rect -1237 -3151 -1233 -3147
rect -1223 -3130 -1219 -3126
rect -1213 -3137 -1209 -3133
rect -1199 -3122 -1195 -3118
rect -1195 -3151 -1191 -3147
rect -1171 -3130 -1167 -3126
rect -1181 -3137 -1177 -3133
rect -1157 -3151 -1153 -3147
rect -1139 -3122 -1135 -3118
rect -1129 -3137 -1125 -3133
rect -1139 -3144 -1135 -3140
rect -1115 -3122 -1111 -3118
rect -1111 -3130 -1107 -3126
rect -1097 -3137 -1093 -3133
rect -1087 -3144 -1083 -3140
rect -1025 -3126 -1021 -3116
rect -1073 -3130 -1069 -3126
rect -928 -3130 -924 -3126
rect -924 -3144 -920 -3140
rect -908 -3122 -904 -3118
rect -908 -3151 -904 -3147
rect -894 -3130 -890 -3126
rect -884 -3137 -880 -3133
rect -870 -3122 -866 -3118
rect -866 -3151 -862 -3147
rect -842 -3130 -838 -3126
rect -852 -3137 -848 -3133
rect -828 -3151 -824 -3147
rect -810 -3122 -806 -3118
rect -800 -3137 -796 -3133
rect -810 -3144 -806 -3140
rect -786 -3122 -782 -3118
rect -782 -3130 -778 -3126
rect -768 -3137 -764 -3133
rect -758 -3144 -754 -3140
rect -744 -3130 -740 -3126
rect -570 -3130 -566 -3126
rect -566 -3144 -562 -3140
rect -550 -3122 -546 -3118
rect -550 -3151 -546 -3147
rect -536 -3130 -532 -3126
rect -526 -3137 -522 -3133
rect -512 -3122 -508 -3118
rect -508 -3151 -504 -3147
rect -484 -3130 -480 -3126
rect -494 -3137 -490 -3133
rect -470 -3151 -466 -3147
rect -452 -3122 -448 -3118
rect -442 -3137 -438 -3133
rect -452 -3144 -448 -3140
rect -428 -3122 -424 -3118
rect -424 -3130 -420 -3126
rect -410 -3137 -406 -3133
rect -400 -3144 -396 -3140
rect -386 -3130 -382 -3126
rect -328 -3127 -324 -3117
rect -212 -3130 -208 -3126
rect -208 -3144 -204 -3140
rect -192 -3122 -188 -3118
rect -192 -3151 -188 -3147
rect -178 -3130 -174 -3126
rect -168 -3137 -164 -3133
rect -154 -3122 -150 -3118
rect -150 -3151 -146 -3147
rect -126 -3130 -122 -3126
rect -136 -3137 -132 -3133
rect -112 -3151 -108 -3147
rect -94 -3122 -90 -3118
rect -84 -3137 -80 -3133
rect -94 -3144 -90 -3140
rect -70 -3122 -66 -3118
rect -66 -3130 -62 -3126
rect -52 -3137 -48 -3133
rect -42 -3144 -38 -3140
rect -28 -3130 -24 -3126
rect 216 -3130 220 -3126
rect 220 -3144 224 -3140
rect 236 -3122 240 -3118
rect 236 -3151 240 -3147
rect 250 -3130 254 -3126
rect 260 -3137 264 -3133
rect 274 -3122 278 -3118
rect 278 -3151 282 -3147
rect 302 -3130 306 -3126
rect 292 -3137 296 -3133
rect 316 -3151 320 -3147
rect 334 -3122 338 -3118
rect 344 -3137 348 -3133
rect 334 -3144 338 -3140
rect 358 -3122 362 -3118
rect 362 -3130 366 -3126
rect 376 -3137 380 -3133
rect 386 -3144 390 -3140
rect 473 -3126 477 -3116
rect 400 -3130 404 -3126
rect 572 -3130 576 -3126
rect 576 -3144 580 -3140
rect 592 -3122 596 -3118
rect 592 -3151 596 -3147
rect 606 -3130 610 -3126
rect 616 -3137 620 -3133
rect 630 -3122 634 -3118
rect 634 -3151 638 -3147
rect 658 -3130 662 -3126
rect 648 -3137 652 -3133
rect 672 -3151 676 -3147
rect 690 -3122 694 -3118
rect 700 -3137 704 -3133
rect 690 -3144 694 -3140
rect 714 -3122 718 -3118
rect 718 -3130 722 -3126
rect 732 -3137 736 -3133
rect 742 -3144 746 -3140
rect 756 -3130 760 -3126
rect 970 -3130 974 -3126
rect 974 -3144 978 -3140
rect 990 -3122 994 -3118
rect 990 -3151 994 -3147
rect 1004 -3130 1008 -3126
rect 1014 -3137 1018 -3133
rect 1028 -3122 1032 -3118
rect 1032 -3151 1036 -3147
rect 1056 -3130 1060 -3126
rect 1046 -3137 1050 -3133
rect 1070 -3151 1074 -3147
rect 1088 -3122 1092 -3118
rect 1098 -3137 1102 -3133
rect 1088 -3144 1092 -3140
rect 1112 -3122 1116 -3118
rect 1116 -3130 1120 -3126
rect 1130 -3137 1134 -3133
rect 1140 -3144 1144 -3140
rect 1200 -3126 1204 -3116
rect 1154 -3130 1158 -3126
rect 1328 -3130 1332 -3126
rect 1332 -3144 1336 -3140
rect 1348 -3122 1352 -3118
rect 1348 -3151 1352 -3147
rect 1362 -3130 1366 -3126
rect 1372 -3137 1376 -3133
rect 1386 -3122 1390 -3118
rect 1390 -3151 1394 -3147
rect 1414 -3130 1418 -3126
rect 1404 -3137 1408 -3133
rect 1428 -3151 1432 -3147
rect 1446 -3122 1450 -3118
rect 1456 -3137 1460 -3133
rect 1446 -3144 1450 -3140
rect 1470 -3122 1474 -3118
rect 1474 -3130 1478 -3126
rect 1488 -3137 1492 -3133
rect 1498 -3144 1502 -3140
rect 1512 -3130 1516 -3126
rect -1257 -3251 -1253 -3247
rect -1253 -3265 -1249 -3261
rect -1237 -3243 -1233 -3239
rect -1237 -3272 -1233 -3268
rect -1223 -3251 -1219 -3247
rect -1213 -3258 -1209 -3254
rect -1199 -3243 -1195 -3239
rect -1195 -3272 -1191 -3268
rect -1171 -3251 -1167 -3247
rect -1181 -3258 -1177 -3254
rect -1157 -3272 -1153 -3268
rect -1139 -3243 -1135 -3239
rect -1129 -3258 -1125 -3254
rect -1139 -3265 -1135 -3261
rect -1115 -3243 -1111 -3239
rect -1111 -3251 -1107 -3247
rect -1097 -3258 -1093 -3254
rect -1087 -3265 -1083 -3261
rect -1073 -3251 -1069 -3247
rect -928 -3251 -924 -3247
rect -924 -3265 -920 -3261
rect -908 -3243 -904 -3239
rect -908 -3272 -904 -3268
rect -894 -3251 -890 -3247
rect -884 -3258 -880 -3254
rect -870 -3243 -866 -3239
rect -866 -3272 -862 -3268
rect -842 -3251 -838 -3247
rect -852 -3258 -848 -3254
rect -828 -3272 -824 -3268
rect -810 -3243 -806 -3239
rect -800 -3258 -796 -3254
rect -810 -3265 -806 -3261
rect -786 -3243 -782 -3239
rect -782 -3251 -778 -3247
rect -768 -3258 -764 -3254
rect -758 -3265 -754 -3261
rect -744 -3251 -740 -3247
rect -570 -3251 -566 -3247
rect -566 -3265 -562 -3261
rect -550 -3243 -546 -3239
rect -550 -3272 -546 -3268
rect -536 -3251 -532 -3247
rect -526 -3258 -522 -3254
rect -512 -3243 -508 -3239
rect -508 -3272 -504 -3268
rect -484 -3251 -480 -3247
rect -494 -3258 -490 -3254
rect -470 -3272 -466 -3268
rect -452 -3243 -448 -3239
rect -442 -3258 -438 -3254
rect -452 -3265 -448 -3261
rect -428 -3243 -424 -3239
rect -424 -3251 -420 -3247
rect -410 -3258 -406 -3254
rect -400 -3265 -396 -3261
rect -386 -3251 -382 -3247
rect -212 -3251 -208 -3247
rect -208 -3265 -204 -3261
rect -192 -3243 -188 -3239
rect -192 -3272 -188 -3268
rect -178 -3251 -174 -3247
rect -168 -3258 -164 -3254
rect -154 -3243 -150 -3239
rect -150 -3272 -146 -3268
rect -126 -3251 -122 -3247
rect -136 -3258 -132 -3254
rect -112 -3272 -108 -3268
rect -94 -3243 -90 -3239
rect -84 -3258 -80 -3254
rect -94 -3265 -90 -3261
rect -70 -3243 -66 -3239
rect -66 -3251 -62 -3247
rect -52 -3258 -48 -3254
rect -42 -3265 -38 -3261
rect -28 -3251 -24 -3247
rect 216 -3251 220 -3247
rect 220 -3265 224 -3261
rect 236 -3243 240 -3239
rect 236 -3272 240 -3268
rect 250 -3251 254 -3247
rect 260 -3258 264 -3254
rect 274 -3243 278 -3239
rect 278 -3272 282 -3268
rect 302 -3251 306 -3247
rect 292 -3258 296 -3254
rect 316 -3272 320 -3268
rect 334 -3243 338 -3239
rect 344 -3258 348 -3254
rect 334 -3265 338 -3261
rect 358 -3243 362 -3239
rect 362 -3251 366 -3247
rect 376 -3258 380 -3254
rect 386 -3265 390 -3261
rect 400 -3251 404 -3247
rect 572 -3251 576 -3247
rect 576 -3265 580 -3261
rect 592 -3243 596 -3239
rect 592 -3272 596 -3268
rect 606 -3251 610 -3247
rect 616 -3258 620 -3254
rect 630 -3243 634 -3239
rect 634 -3272 638 -3268
rect 658 -3251 662 -3247
rect 648 -3258 652 -3254
rect 672 -3272 676 -3268
rect 690 -3243 694 -3239
rect 700 -3258 704 -3254
rect 690 -3265 694 -3261
rect 714 -3243 718 -3239
rect 718 -3251 722 -3247
rect 732 -3258 736 -3254
rect 742 -3265 746 -3261
rect 756 -3251 760 -3247
rect 970 -3251 974 -3247
rect 974 -3265 978 -3261
rect 990 -3243 994 -3239
rect 990 -3272 994 -3268
rect 1004 -3251 1008 -3247
rect 1014 -3258 1018 -3254
rect 1028 -3243 1032 -3239
rect 1032 -3272 1036 -3268
rect 1056 -3251 1060 -3247
rect 1046 -3258 1050 -3254
rect 1070 -3272 1074 -3268
rect 1088 -3243 1092 -3239
rect 1098 -3258 1102 -3254
rect 1088 -3265 1092 -3261
rect 1112 -3243 1116 -3239
rect 1116 -3251 1120 -3247
rect 1130 -3258 1134 -3254
rect 1140 -3265 1144 -3261
rect 1154 -3251 1158 -3247
rect 1328 -3251 1332 -3247
rect 1332 -3265 1336 -3261
rect 1348 -3243 1352 -3239
rect 1348 -3272 1352 -3268
rect 1362 -3251 1366 -3247
rect 1372 -3258 1376 -3254
rect 1386 -3243 1390 -3239
rect 1390 -3272 1394 -3268
rect 1414 -3251 1418 -3247
rect 1404 -3258 1408 -3254
rect 1428 -3272 1432 -3268
rect 1446 -3243 1450 -3239
rect 1456 -3258 1460 -3254
rect 1446 -3265 1450 -3261
rect 1470 -3243 1474 -3239
rect 1474 -3251 1478 -3247
rect 1488 -3258 1492 -3254
rect 1498 -3265 1502 -3261
rect 1512 -3251 1516 -3247
rect -1257 -3365 -1253 -3361
rect -1253 -3379 -1249 -3375
rect -1237 -3357 -1233 -3353
rect -1237 -3386 -1233 -3382
rect -1223 -3365 -1219 -3361
rect -1213 -3372 -1209 -3368
rect -1199 -3357 -1195 -3353
rect -1195 -3386 -1191 -3382
rect -1171 -3365 -1167 -3361
rect -1181 -3372 -1177 -3368
rect -1157 -3386 -1153 -3382
rect -1139 -3357 -1135 -3353
rect -1129 -3372 -1125 -3368
rect -1139 -3379 -1135 -3375
rect -1115 -3357 -1111 -3353
rect -1111 -3365 -1107 -3361
rect -1097 -3372 -1093 -3368
rect -1087 -3379 -1083 -3375
rect -1073 -3365 -1069 -3361
rect -928 -3365 -924 -3361
rect -924 -3379 -920 -3375
rect -908 -3357 -904 -3353
rect -908 -3386 -904 -3382
rect -894 -3365 -890 -3361
rect -884 -3372 -880 -3368
rect -870 -3357 -866 -3353
rect -866 -3386 -862 -3382
rect -842 -3365 -838 -3361
rect -852 -3372 -848 -3368
rect -828 -3386 -824 -3382
rect -810 -3357 -806 -3353
rect -800 -3372 -796 -3368
rect -810 -3379 -806 -3375
rect -786 -3357 -782 -3353
rect -782 -3365 -778 -3361
rect -768 -3372 -764 -3368
rect -758 -3379 -754 -3375
rect -744 -3365 -740 -3361
rect -570 -3365 -566 -3361
rect -566 -3379 -562 -3375
rect -550 -3357 -546 -3353
rect -550 -3386 -546 -3382
rect -536 -3365 -532 -3361
rect -526 -3372 -522 -3368
rect -512 -3357 -508 -3353
rect -508 -3386 -504 -3382
rect -484 -3365 -480 -3361
rect -494 -3372 -490 -3368
rect -470 -3386 -466 -3382
rect -452 -3357 -448 -3353
rect -442 -3372 -438 -3368
rect -452 -3379 -448 -3375
rect -428 -3357 -424 -3353
rect -424 -3365 -420 -3361
rect -410 -3372 -406 -3368
rect -400 -3379 -396 -3375
rect -386 -3365 -382 -3361
rect -1338 -3458 -1334 -3454
rect -1327 -3466 -1323 -3462
rect -1320 -3488 -1316 -3484
rect -934 -3458 -930 -3454
rect -923 -3466 -919 -3462
rect -916 -3488 -912 -3484
rect -576 -3458 -572 -3454
rect -565 -3466 -561 -3462
rect -558 -3488 -554 -3484
rect -218 -3458 -214 -3454
rect -207 -3466 -203 -3462
rect -200 -3488 -196 -3484
rect 210 -3458 214 -3454
rect 221 -3466 225 -3462
rect 228 -3488 232 -3484
rect 566 -3458 570 -3454
rect 577 -3466 581 -3462
rect 584 -3488 588 -3484
rect 964 -3458 968 -3454
rect 975 -3466 979 -3462
rect 982 -3488 986 -3484
rect 1322 -3458 1326 -3454
rect 1333 -3466 1337 -3462
rect 1340 -3488 1344 -3484
rect -1253 -3606 -1249 -3602
rect -1257 -3613 -1253 -3609
rect -1237 -3593 -1233 -3589
rect -1227 -3613 -1223 -3609
rect -1213 -3606 -1209 -3602
rect -1203 -3599 -1199 -3595
rect -1193 -3606 -1189 -3602
rect -1179 -3613 -1175 -3609
rect -1175 -3627 -1171 -3623
rect -924 -3569 -920 -3565
rect -928 -3590 -924 -3586
rect -924 -3605 -920 -3601
rect -928 -3619 -924 -3615
rect -898 -3590 -894 -3586
rect -902 -3598 -898 -3594
rect -902 -3612 -898 -3608
rect -882 -3576 -878 -3572
rect -872 -3619 -868 -3615
rect -858 -3569 -854 -3565
rect -848 -3583 -844 -3579
rect -838 -3619 -834 -3615
rect -824 -3569 -820 -3565
rect -820 -3627 -816 -3623
rect -804 -3598 -800 -3594
rect -794 -3612 -790 -3608
rect -780 -3569 -776 -3565
rect -780 -3590 -776 -3586
rect -776 -3605 -772 -3601
rect -760 -3612 -756 -3608
rect -746 -3569 -742 -3565
rect -736 -3620 -732 -3616
rect -720 -3627 -716 -3623
rect -706 -3583 -702 -3579
rect -702 -3620 -698 -3616
rect -566 -3569 -562 -3565
rect -570 -3590 -566 -3586
rect -566 -3605 -562 -3601
rect -570 -3619 -566 -3615
rect -540 -3590 -536 -3586
rect -544 -3598 -540 -3594
rect -544 -3612 -540 -3608
rect -524 -3576 -520 -3572
rect -514 -3619 -510 -3615
rect -500 -3569 -496 -3565
rect -490 -3583 -486 -3579
rect -480 -3619 -476 -3615
rect -466 -3569 -462 -3565
rect -462 -3627 -458 -3623
rect -446 -3598 -442 -3594
rect -436 -3612 -432 -3608
rect -422 -3569 -418 -3565
rect -422 -3590 -418 -3586
rect -418 -3605 -414 -3601
rect -402 -3612 -398 -3608
rect -388 -3569 -384 -3565
rect -378 -3620 -374 -3616
rect -362 -3627 -358 -3623
rect -348 -3583 -344 -3579
rect -344 -3620 -340 -3616
rect -208 -3569 -204 -3565
rect -212 -3590 -208 -3586
rect -208 -3605 -204 -3601
rect -212 -3619 -208 -3615
rect -182 -3590 -178 -3586
rect -186 -3598 -182 -3594
rect -186 -3612 -182 -3608
rect -166 -3576 -162 -3572
rect -156 -3619 -152 -3615
rect -142 -3569 -138 -3565
rect -132 -3583 -128 -3579
rect -122 -3619 -118 -3615
rect -108 -3569 -104 -3565
rect -104 -3627 -100 -3623
rect -88 -3598 -84 -3594
rect -78 -3612 -74 -3608
rect -64 -3569 -60 -3565
rect -64 -3590 -60 -3586
rect -60 -3605 -56 -3601
rect -44 -3612 -40 -3608
rect -30 -3569 -26 -3565
rect -20 -3620 -16 -3616
rect -4 -3627 0 -3623
rect 10 -3583 14 -3579
rect 14 -3620 18 -3616
rect 220 -3569 224 -3565
rect 216 -3590 220 -3586
rect 220 -3605 224 -3601
rect 216 -3619 220 -3615
rect 246 -3590 250 -3586
rect 242 -3598 246 -3594
rect 242 -3612 246 -3608
rect 262 -3576 266 -3572
rect 272 -3619 276 -3615
rect 286 -3569 290 -3565
rect 296 -3583 300 -3579
rect 306 -3619 310 -3615
rect 320 -3569 324 -3565
rect 324 -3627 328 -3623
rect 340 -3598 344 -3594
rect 350 -3612 354 -3608
rect 364 -3569 368 -3565
rect 364 -3590 368 -3586
rect 368 -3605 372 -3601
rect 384 -3612 388 -3608
rect 398 -3569 402 -3565
rect 408 -3620 412 -3616
rect 424 -3627 428 -3623
rect 438 -3583 442 -3579
rect 442 -3620 446 -3616
rect 576 -3569 580 -3565
rect 572 -3590 576 -3586
rect 576 -3605 580 -3601
rect 572 -3619 576 -3615
rect 602 -3590 606 -3586
rect 598 -3598 602 -3594
rect 598 -3612 602 -3608
rect 618 -3576 622 -3572
rect 628 -3619 632 -3615
rect 642 -3569 646 -3565
rect 652 -3583 656 -3579
rect 662 -3619 666 -3615
rect 676 -3569 680 -3565
rect 680 -3627 684 -3623
rect 696 -3598 700 -3594
rect 706 -3612 710 -3608
rect 720 -3569 724 -3565
rect 720 -3590 724 -3586
rect 724 -3605 728 -3601
rect 740 -3612 744 -3608
rect 754 -3569 758 -3565
rect 764 -3620 768 -3616
rect 780 -3627 784 -3623
rect 794 -3583 798 -3579
rect 798 -3620 802 -3616
rect 974 -3569 978 -3565
rect 970 -3590 974 -3586
rect 974 -3605 978 -3601
rect 970 -3619 974 -3615
rect 1000 -3590 1004 -3586
rect 996 -3598 1000 -3594
rect 996 -3612 1000 -3608
rect 1016 -3576 1020 -3572
rect 1026 -3619 1030 -3615
rect 1040 -3569 1044 -3565
rect 1050 -3583 1054 -3579
rect 1060 -3619 1064 -3615
rect 1074 -3569 1078 -3565
rect 1078 -3627 1082 -3623
rect 1094 -3598 1098 -3594
rect 1104 -3612 1108 -3608
rect 1118 -3569 1122 -3565
rect 1118 -3590 1122 -3586
rect 1122 -3605 1126 -3601
rect 1138 -3612 1142 -3608
rect 1152 -3569 1156 -3565
rect 1162 -3620 1166 -3616
rect 1178 -3627 1182 -3623
rect 1192 -3583 1196 -3579
rect 1196 -3620 1200 -3616
rect 1332 -3569 1336 -3565
rect 1328 -3590 1332 -3586
rect 1332 -3605 1336 -3601
rect 1328 -3619 1332 -3615
rect 1358 -3590 1362 -3586
rect 1354 -3598 1358 -3594
rect 1354 -3612 1358 -3608
rect 1374 -3576 1378 -3572
rect 1384 -3619 1388 -3615
rect 1398 -3569 1402 -3565
rect 1408 -3583 1412 -3579
rect 1418 -3619 1422 -3615
rect 1432 -3569 1436 -3565
rect 1436 -3627 1440 -3623
rect 1452 -3598 1456 -3594
rect 1462 -3612 1466 -3608
rect 1476 -3569 1480 -3565
rect 1476 -3590 1480 -3586
rect 1480 -3605 1484 -3601
rect 1496 -3612 1500 -3608
rect 1510 -3569 1514 -3565
rect 1520 -3620 1524 -3616
rect 1536 -3627 1540 -3623
rect 1550 -3583 1554 -3579
rect 1554 -3620 1558 -3616
rect -1257 -3736 -1253 -3732
rect -1253 -3750 -1249 -3746
rect -1237 -3728 -1233 -3724
rect -1237 -3757 -1233 -3753
rect -1223 -3736 -1219 -3732
rect -1213 -3743 -1209 -3739
rect -1199 -3728 -1195 -3724
rect -1195 -3757 -1191 -3753
rect -1171 -3736 -1167 -3732
rect -1181 -3743 -1177 -3739
rect -1157 -3757 -1153 -3753
rect -1139 -3728 -1135 -3724
rect -1129 -3743 -1125 -3739
rect -1139 -3750 -1135 -3746
rect -1115 -3728 -1111 -3724
rect -1111 -3736 -1107 -3732
rect -1097 -3743 -1093 -3739
rect -1087 -3750 -1083 -3746
rect -1073 -3736 -1069 -3732
rect -928 -3736 -924 -3732
rect -924 -3750 -920 -3746
rect -908 -3728 -904 -3724
rect -908 -3757 -904 -3753
rect -894 -3736 -890 -3732
rect -884 -3743 -880 -3739
rect -870 -3728 -866 -3724
rect -866 -3757 -862 -3753
rect -842 -3736 -838 -3732
rect -852 -3743 -848 -3739
rect -828 -3757 -824 -3753
rect -810 -3728 -806 -3724
rect -800 -3743 -796 -3739
rect -810 -3750 -806 -3746
rect -786 -3728 -782 -3724
rect -782 -3736 -778 -3732
rect -768 -3743 -764 -3739
rect -758 -3750 -754 -3746
rect -744 -3736 -740 -3732
rect -570 -3736 -566 -3732
rect -566 -3750 -562 -3746
rect -550 -3728 -546 -3724
rect -550 -3757 -546 -3753
rect -536 -3736 -532 -3732
rect -526 -3743 -522 -3739
rect -512 -3728 -508 -3724
rect -508 -3757 -504 -3753
rect -484 -3736 -480 -3732
rect -494 -3743 -490 -3739
rect -470 -3757 -466 -3753
rect -452 -3728 -448 -3724
rect -442 -3743 -438 -3739
rect -452 -3750 -448 -3746
rect -428 -3728 -424 -3724
rect -424 -3736 -420 -3732
rect -410 -3743 -406 -3739
rect -400 -3750 -396 -3746
rect -386 -3736 -382 -3732
rect -212 -3736 -208 -3732
rect -208 -3750 -204 -3746
rect -192 -3728 -188 -3724
rect -192 -3757 -188 -3753
rect -178 -3736 -174 -3732
rect -168 -3743 -164 -3739
rect -154 -3728 -150 -3724
rect -150 -3757 -146 -3753
rect -126 -3736 -122 -3732
rect -136 -3743 -132 -3739
rect -112 -3757 -108 -3753
rect -94 -3728 -90 -3724
rect -84 -3743 -80 -3739
rect -94 -3750 -90 -3746
rect -70 -3728 -66 -3724
rect -66 -3736 -62 -3732
rect -52 -3743 -48 -3739
rect -42 -3750 -38 -3746
rect -28 -3736 -24 -3732
rect 69 -3852 73 -3836
rect -1257 -3967 -1253 -3963
rect -1253 -3981 -1249 -3977
rect -1237 -3959 -1233 -3955
rect -1237 -3988 -1233 -3984
rect -1223 -3967 -1219 -3963
rect -1213 -3974 -1209 -3970
rect -1199 -3959 -1195 -3955
rect -1195 -3988 -1191 -3984
rect -1171 -3967 -1167 -3963
rect -1181 -3974 -1177 -3970
rect -1157 -3988 -1153 -3984
rect -1139 -3959 -1135 -3955
rect -1129 -3974 -1125 -3970
rect -1139 -3981 -1135 -3977
rect -1115 -3959 -1111 -3955
rect -1111 -3967 -1107 -3963
rect -1097 -3974 -1093 -3970
rect -1087 -3981 -1083 -3977
rect -1073 -3967 -1069 -3963
rect -928 -3967 -924 -3963
rect -924 -3981 -920 -3977
rect -908 -3959 -904 -3955
rect -908 -3988 -904 -3984
rect -894 -3967 -890 -3963
rect -884 -3974 -880 -3970
rect -870 -3959 -866 -3955
rect -866 -3988 -862 -3984
rect -842 -3967 -838 -3963
rect -852 -3974 -848 -3970
rect -828 -3988 -824 -3984
rect -810 -3959 -806 -3955
rect -800 -3974 -796 -3970
rect -810 -3981 -806 -3977
rect -786 -3959 -782 -3955
rect -782 -3967 -778 -3963
rect -768 -3974 -764 -3970
rect -758 -3981 -754 -3977
rect -744 -3967 -740 -3963
rect -570 -3967 -566 -3963
rect -566 -3981 -562 -3977
rect -550 -3959 -546 -3955
rect -550 -3988 -546 -3984
rect -536 -3967 -532 -3963
rect -526 -3974 -522 -3970
rect -512 -3959 -508 -3955
rect -508 -3988 -504 -3984
rect -484 -3967 -480 -3963
rect -494 -3974 -490 -3970
rect -470 -3988 -466 -3984
rect -452 -3959 -448 -3955
rect -442 -3974 -438 -3970
rect -452 -3981 -448 -3977
rect -428 -3959 -424 -3955
rect -424 -3967 -420 -3963
rect -410 -3974 -406 -3970
rect -400 -3981 -396 -3977
rect -386 -3967 -382 -3963
rect -212 -3967 -208 -3963
rect -208 -3981 -204 -3977
rect -192 -3959 -188 -3955
rect -192 -3988 -188 -3984
rect -178 -3967 -174 -3963
rect -168 -3974 -164 -3970
rect -154 -3959 -150 -3955
rect -150 -3988 -146 -3984
rect -126 -3967 -122 -3963
rect -136 -3974 -132 -3970
rect -112 -3988 -108 -3984
rect -94 -3959 -90 -3955
rect -84 -3974 -80 -3970
rect -94 -3981 -90 -3977
rect -70 -3959 -66 -3955
rect -66 -3967 -62 -3963
rect -52 -3974 -48 -3970
rect -42 -3981 -38 -3977
rect -28 -3967 -24 -3963
rect 216 -3967 220 -3963
rect 220 -3981 224 -3977
rect 236 -3959 240 -3955
rect 236 -3988 240 -3984
rect 250 -3967 254 -3963
rect 260 -3974 264 -3970
rect 274 -3959 278 -3955
rect 278 -3988 282 -3984
rect 302 -3967 306 -3963
rect 292 -3974 296 -3970
rect 316 -3988 320 -3984
rect 334 -3959 338 -3955
rect 344 -3974 348 -3970
rect 334 -3981 338 -3977
rect 358 -3959 362 -3955
rect 362 -3967 366 -3963
rect 376 -3974 380 -3970
rect 386 -3981 390 -3977
rect 400 -3967 404 -3963
rect 572 -3967 576 -3963
rect 576 -3981 580 -3977
rect 592 -3959 596 -3955
rect 592 -3988 596 -3984
rect 606 -3967 610 -3963
rect 616 -3974 620 -3970
rect 630 -3959 634 -3955
rect 634 -3988 638 -3984
rect 658 -3967 662 -3963
rect 648 -3974 652 -3970
rect 672 -3988 676 -3984
rect 690 -3959 694 -3955
rect 700 -3974 704 -3970
rect 690 -3981 694 -3977
rect 714 -3959 718 -3955
rect 718 -3967 722 -3963
rect 732 -3974 736 -3970
rect 742 -3981 746 -3977
rect 756 -3967 760 -3963
rect 970 -3967 974 -3963
rect 974 -3981 978 -3977
rect 990 -3959 994 -3955
rect 990 -3988 994 -3984
rect 1004 -3967 1008 -3963
rect 1014 -3974 1018 -3970
rect 1028 -3959 1032 -3955
rect 1032 -3988 1036 -3984
rect 1056 -3967 1060 -3963
rect 1046 -3974 1050 -3970
rect 1070 -3988 1074 -3984
rect 1088 -3959 1092 -3955
rect 1098 -3974 1102 -3970
rect 1088 -3981 1092 -3977
rect 1112 -3959 1116 -3955
rect 1116 -3967 1120 -3963
rect 1130 -3974 1134 -3970
rect 1140 -3981 1144 -3977
rect 1154 -3967 1158 -3963
rect 1328 -3967 1332 -3963
rect 1332 -3981 1336 -3977
rect 1348 -3959 1352 -3955
rect 1348 -3988 1352 -3984
rect 1362 -3967 1366 -3963
rect 1372 -3974 1376 -3970
rect 1386 -3959 1390 -3955
rect 1390 -3988 1394 -3984
rect 1414 -3967 1418 -3963
rect 1404 -3974 1408 -3970
rect 1428 -3988 1432 -3984
rect 1446 -3959 1450 -3955
rect 1456 -3974 1460 -3970
rect 1446 -3981 1450 -3977
rect 1470 -3959 1474 -3955
rect 1474 -3967 1478 -3963
rect 1488 -3974 1492 -3970
rect 1498 -3981 1502 -3977
rect 1512 -3967 1516 -3963
rect -1257 -4092 -1253 -4088
rect -1253 -4106 -1249 -4102
rect -1237 -4084 -1233 -4080
rect -1237 -4113 -1233 -4109
rect -1223 -4092 -1219 -4088
rect -1213 -4099 -1209 -4095
rect -1199 -4084 -1195 -4080
rect -1195 -4113 -1191 -4109
rect -1171 -4092 -1167 -4088
rect -1181 -4099 -1177 -4095
rect -1157 -4113 -1153 -4109
rect -1139 -4084 -1135 -4080
rect -1129 -4099 -1125 -4095
rect -1139 -4106 -1135 -4102
rect -1115 -4084 -1111 -4080
rect -1111 -4092 -1107 -4088
rect -1097 -4099 -1093 -4095
rect -1087 -4106 -1083 -4102
rect -1073 -4092 -1069 -4088
rect -928 -4092 -924 -4088
rect -924 -4106 -920 -4102
rect -908 -4084 -904 -4080
rect -908 -4113 -904 -4109
rect -894 -4092 -890 -4088
rect -884 -4099 -880 -4095
rect -870 -4084 -866 -4080
rect -866 -4113 -862 -4109
rect -842 -4092 -838 -4088
rect -852 -4099 -848 -4095
rect -828 -4113 -824 -4109
rect -810 -4084 -806 -4080
rect -800 -4099 -796 -4095
rect -810 -4106 -806 -4102
rect -786 -4084 -782 -4080
rect -782 -4092 -778 -4088
rect -768 -4099 -764 -4095
rect -758 -4106 -754 -4102
rect -744 -4092 -740 -4088
rect -570 -4092 -566 -4088
rect -566 -4106 -562 -4102
rect -550 -4084 -546 -4080
rect -550 -4113 -546 -4109
rect -536 -4092 -532 -4088
rect -526 -4099 -522 -4095
rect -512 -4084 -508 -4080
rect -508 -4113 -504 -4109
rect -484 -4092 -480 -4088
rect -494 -4099 -490 -4095
rect -470 -4113 -466 -4109
rect -452 -4084 -448 -4080
rect -442 -4099 -438 -4095
rect -452 -4106 -448 -4102
rect -428 -4084 -424 -4080
rect -424 -4092 -420 -4088
rect -410 -4099 -406 -4095
rect -400 -4106 -396 -4102
rect -386 -4092 -382 -4088
rect -212 -4092 -208 -4088
rect -208 -4106 -204 -4102
rect -192 -4084 -188 -4080
rect -192 -4113 -188 -4109
rect -178 -4092 -174 -4088
rect -168 -4099 -164 -4095
rect -154 -4084 -150 -4080
rect -150 -4113 -146 -4109
rect -126 -4092 -122 -4088
rect -136 -4099 -132 -4095
rect -112 -4113 -108 -4109
rect -94 -4084 -90 -4080
rect -84 -4099 -80 -4095
rect -94 -4106 -90 -4102
rect -70 -4084 -66 -4080
rect -66 -4092 -62 -4088
rect -52 -4099 -48 -4095
rect -42 -4106 -38 -4102
rect -28 -4092 -24 -4088
rect 216 -4092 220 -4088
rect 220 -4106 224 -4102
rect 236 -4084 240 -4080
rect 236 -4113 240 -4109
rect 250 -4092 254 -4088
rect 260 -4099 264 -4095
rect 274 -4084 278 -4080
rect 278 -4113 282 -4109
rect 302 -4092 306 -4088
rect 292 -4099 296 -4095
rect 316 -4113 320 -4109
rect 334 -4084 338 -4080
rect 344 -4099 348 -4095
rect 334 -4106 338 -4102
rect 358 -4084 362 -4080
rect 362 -4092 366 -4088
rect 376 -4099 380 -4095
rect 386 -4106 390 -4102
rect 400 -4092 404 -4088
rect 572 -4092 576 -4088
rect 576 -4106 580 -4102
rect 592 -4084 596 -4080
rect 592 -4113 596 -4109
rect 606 -4092 610 -4088
rect 616 -4099 620 -4095
rect 630 -4084 634 -4080
rect 634 -4113 638 -4109
rect 658 -4092 662 -4088
rect 648 -4099 652 -4095
rect 672 -4113 676 -4109
rect 690 -4084 694 -4080
rect 700 -4099 704 -4095
rect 690 -4106 694 -4102
rect 714 -4084 718 -4080
rect 718 -4092 722 -4088
rect 732 -4099 736 -4095
rect 742 -4106 746 -4102
rect 756 -4092 760 -4088
rect 970 -4092 974 -4088
rect 974 -4106 978 -4102
rect 990 -4084 994 -4080
rect 990 -4113 994 -4109
rect 1004 -4092 1008 -4088
rect 1014 -4099 1018 -4095
rect 1028 -4084 1032 -4080
rect 1032 -4113 1036 -4109
rect 1056 -4092 1060 -4088
rect 1046 -4099 1050 -4095
rect 1070 -4113 1074 -4109
rect 1088 -4084 1092 -4080
rect 1098 -4099 1102 -4095
rect 1088 -4106 1092 -4102
rect 1112 -4084 1116 -4080
rect 1116 -4092 1120 -4088
rect 1130 -4099 1134 -4095
rect 1140 -4106 1144 -4102
rect 1154 -4092 1158 -4088
rect 1328 -4092 1332 -4088
rect 1332 -4106 1336 -4102
rect 1348 -4084 1352 -4080
rect 1348 -4113 1352 -4109
rect 1362 -4092 1366 -4088
rect 1372 -4099 1376 -4095
rect 1386 -4084 1390 -4080
rect 1390 -4113 1394 -4109
rect 1414 -4092 1418 -4088
rect 1404 -4099 1408 -4095
rect 1428 -4113 1432 -4109
rect 1446 -4084 1450 -4080
rect 1456 -4099 1460 -4095
rect 1446 -4106 1450 -4102
rect 1470 -4084 1474 -4080
rect 1474 -4092 1478 -4088
rect 1488 -4099 1492 -4095
rect 1498 -4106 1502 -4102
rect 1512 -4092 1516 -4088
rect -1257 -4216 -1253 -4212
rect -1253 -4230 -1249 -4226
rect -1237 -4208 -1233 -4204
rect -1237 -4237 -1233 -4233
rect -1223 -4216 -1219 -4212
rect -1213 -4223 -1209 -4219
rect -1199 -4208 -1195 -4204
rect -1195 -4237 -1191 -4233
rect -1171 -4216 -1167 -4212
rect -1181 -4223 -1177 -4219
rect -1157 -4237 -1153 -4233
rect -1139 -4208 -1135 -4204
rect -1129 -4223 -1125 -4219
rect -1139 -4230 -1135 -4226
rect -1115 -4208 -1111 -4204
rect -1111 -4216 -1107 -4212
rect -1097 -4223 -1093 -4219
rect -1087 -4230 -1083 -4226
rect -1028 -4208 -1024 -4198
rect -1073 -4216 -1069 -4212
rect -928 -4216 -924 -4212
rect -924 -4230 -920 -4226
rect -908 -4208 -904 -4204
rect -908 -4237 -904 -4233
rect -894 -4216 -890 -4212
rect -884 -4223 -880 -4219
rect -870 -4208 -866 -4204
rect -866 -4237 -862 -4233
rect -842 -4216 -838 -4212
rect -852 -4223 -848 -4219
rect -828 -4237 -824 -4233
rect -810 -4208 -806 -4204
rect -800 -4223 -796 -4219
rect -810 -4230 -806 -4226
rect -786 -4208 -782 -4204
rect -782 -4216 -778 -4212
rect -768 -4223 -764 -4219
rect -758 -4230 -754 -4226
rect -744 -4216 -740 -4212
rect -570 -4216 -566 -4212
rect -566 -4230 -562 -4226
rect -550 -4208 -546 -4204
rect -550 -4237 -546 -4233
rect -536 -4216 -532 -4212
rect -526 -4223 -522 -4219
rect -512 -4208 -508 -4204
rect -508 -4237 -504 -4233
rect -484 -4216 -480 -4212
rect -494 -4223 -490 -4219
rect -470 -4237 -466 -4233
rect -452 -4208 -448 -4204
rect -442 -4223 -438 -4219
rect -452 -4230 -448 -4226
rect -428 -4208 -424 -4204
rect -424 -4216 -420 -4212
rect -410 -4223 -406 -4219
rect -400 -4230 -396 -4226
rect -331 -4210 -327 -4200
rect -386 -4216 -382 -4212
rect -212 -4216 -208 -4212
rect -208 -4230 -204 -4226
rect -192 -4208 -188 -4204
rect -192 -4237 -188 -4233
rect -178 -4216 -174 -4212
rect -168 -4223 -164 -4219
rect -154 -4208 -150 -4204
rect -150 -4237 -146 -4233
rect -126 -4216 -122 -4212
rect -136 -4223 -132 -4219
rect -112 -4237 -108 -4233
rect -94 -4208 -90 -4204
rect -84 -4223 -80 -4219
rect -94 -4230 -90 -4226
rect -70 -4208 -66 -4204
rect -66 -4216 -62 -4212
rect -52 -4223 -48 -4219
rect -42 -4230 -38 -4226
rect 457 -4208 461 -4198
rect -28 -4216 -24 -4212
rect 1202 -4208 1206 -4198
rect -1338 -4303 -1334 -4299
rect -1327 -4311 -1323 -4307
rect -1320 -4333 -1316 -4329
rect -1028 -4324 -1024 -4314
rect -934 -4303 -930 -4299
rect -923 -4311 -919 -4307
rect -916 -4333 -912 -4329
rect -672 -4324 -668 -4314
rect -576 -4303 -572 -4299
rect -565 -4311 -561 -4307
rect -558 -4333 -554 -4329
rect -331 -4325 -327 -4315
rect -218 -4303 -214 -4299
rect -207 -4311 -203 -4307
rect -200 -4333 -196 -4329
rect 210 -4303 214 -4299
rect 221 -4311 225 -4307
rect 228 -4333 232 -4329
rect 457 -4324 461 -4314
rect 566 -4303 570 -4299
rect 577 -4311 581 -4307
rect 584 -4333 588 -4329
rect 861 -4324 865 -4314
rect 964 -4303 968 -4299
rect 975 -4311 979 -4307
rect 982 -4333 986 -4329
rect 1202 -4324 1206 -4314
rect 1322 -4303 1326 -4299
rect 1333 -4311 1337 -4307
rect 1340 -4333 1344 -4329
rect -1253 -4446 -1249 -4442
rect -1257 -4453 -1253 -4449
rect -1237 -4433 -1233 -4429
rect -1227 -4453 -1223 -4449
rect -1213 -4446 -1209 -4442
rect -1203 -4439 -1199 -4435
rect -1193 -4446 -1189 -4442
rect -1179 -4453 -1175 -4449
rect -1175 -4467 -1171 -4463
rect -924 -4409 -920 -4405
rect -928 -4430 -924 -4426
rect -924 -4445 -920 -4441
rect -928 -4459 -924 -4455
rect -898 -4430 -894 -4426
rect -902 -4438 -898 -4434
rect -902 -4452 -898 -4448
rect -882 -4416 -878 -4412
rect -872 -4459 -868 -4455
rect -858 -4409 -854 -4405
rect -848 -4423 -844 -4419
rect -838 -4459 -834 -4455
rect -824 -4409 -820 -4405
rect -820 -4467 -816 -4463
rect -804 -4438 -800 -4434
rect -794 -4452 -790 -4448
rect -780 -4409 -776 -4405
rect -780 -4430 -776 -4426
rect -776 -4445 -772 -4441
rect -760 -4452 -756 -4448
rect -746 -4409 -742 -4405
rect -736 -4460 -732 -4456
rect -720 -4467 -716 -4463
rect -706 -4423 -702 -4419
rect -702 -4460 -698 -4456
rect -566 -4409 -562 -4405
rect -570 -4430 -566 -4426
rect -566 -4445 -562 -4441
rect -570 -4459 -566 -4455
rect -540 -4430 -536 -4426
rect -544 -4438 -540 -4434
rect -544 -4452 -540 -4448
rect -524 -4416 -520 -4412
rect -514 -4459 -510 -4455
rect -500 -4409 -496 -4405
rect -490 -4423 -486 -4419
rect -480 -4459 -476 -4455
rect -466 -4409 -462 -4405
rect -462 -4467 -458 -4463
rect -446 -4438 -442 -4434
rect -436 -4452 -432 -4448
rect -422 -4409 -418 -4405
rect -422 -4430 -418 -4426
rect -418 -4445 -414 -4441
rect -402 -4452 -398 -4448
rect -388 -4409 -384 -4405
rect -378 -4460 -374 -4456
rect -362 -4467 -358 -4463
rect -348 -4423 -344 -4419
rect -344 -4460 -340 -4456
rect -208 -4409 -204 -4405
rect -212 -4430 -208 -4426
rect -208 -4445 -204 -4441
rect -212 -4459 -208 -4455
rect -182 -4430 -178 -4426
rect -186 -4438 -182 -4434
rect -186 -4452 -182 -4448
rect -166 -4416 -162 -4412
rect -156 -4459 -152 -4455
rect -142 -4409 -138 -4405
rect -132 -4423 -128 -4419
rect -122 -4459 -118 -4455
rect -108 -4409 -104 -4405
rect -104 -4467 -100 -4463
rect -88 -4438 -84 -4434
rect -78 -4452 -74 -4448
rect -64 -4409 -60 -4405
rect -64 -4430 -60 -4426
rect -60 -4445 -56 -4441
rect -44 -4452 -40 -4448
rect -30 -4409 -26 -4405
rect -20 -4460 -16 -4456
rect -4 -4467 0 -4463
rect 10 -4423 14 -4419
rect 14 -4460 18 -4456
rect 220 -4409 224 -4405
rect 216 -4430 220 -4426
rect 220 -4445 224 -4441
rect 216 -4459 220 -4455
rect 246 -4430 250 -4426
rect 242 -4438 246 -4434
rect 242 -4452 246 -4448
rect 262 -4416 266 -4412
rect 272 -4459 276 -4455
rect 286 -4409 290 -4405
rect 296 -4423 300 -4419
rect 306 -4459 310 -4455
rect 320 -4409 324 -4405
rect 324 -4467 328 -4463
rect 340 -4438 344 -4434
rect 350 -4452 354 -4448
rect 364 -4409 368 -4405
rect 364 -4430 368 -4426
rect 368 -4445 372 -4441
rect 384 -4452 388 -4448
rect 398 -4409 402 -4405
rect 408 -4460 412 -4456
rect 424 -4467 428 -4463
rect 438 -4423 442 -4419
rect 442 -4460 446 -4456
rect 576 -4409 580 -4405
rect 572 -4430 576 -4426
rect 576 -4445 580 -4441
rect 572 -4459 576 -4455
rect 602 -4430 606 -4426
rect 598 -4438 602 -4434
rect 598 -4452 602 -4448
rect 618 -4416 622 -4412
rect 628 -4459 632 -4455
rect 642 -4409 646 -4405
rect 652 -4423 656 -4419
rect 662 -4459 666 -4455
rect 676 -4409 680 -4405
rect 680 -4467 684 -4463
rect 696 -4438 700 -4434
rect 706 -4452 710 -4448
rect 720 -4409 724 -4405
rect 720 -4430 724 -4426
rect 724 -4445 728 -4441
rect 740 -4452 744 -4448
rect 754 -4409 758 -4405
rect 764 -4460 768 -4456
rect 780 -4467 784 -4463
rect 794 -4423 798 -4419
rect 798 -4460 802 -4456
rect 974 -4409 978 -4405
rect 970 -4430 974 -4426
rect 974 -4445 978 -4441
rect 970 -4459 974 -4455
rect 1000 -4430 1004 -4426
rect 996 -4438 1000 -4434
rect 996 -4452 1000 -4448
rect 1016 -4416 1020 -4412
rect 1026 -4459 1030 -4455
rect 1040 -4409 1044 -4405
rect 1050 -4423 1054 -4419
rect 1060 -4459 1064 -4455
rect 1074 -4409 1078 -4405
rect 1078 -4467 1082 -4463
rect 1094 -4438 1098 -4434
rect 1104 -4452 1108 -4448
rect 1118 -4409 1122 -4405
rect 1118 -4430 1122 -4426
rect 1122 -4445 1126 -4441
rect 1138 -4452 1142 -4448
rect 1152 -4409 1156 -4405
rect 1162 -4460 1166 -4456
rect 1178 -4467 1182 -4463
rect 1192 -4423 1196 -4419
rect 1196 -4460 1200 -4456
rect 1332 -4409 1336 -4405
rect 1328 -4430 1332 -4426
rect 1332 -4445 1336 -4441
rect 1328 -4459 1332 -4455
rect 1358 -4430 1362 -4426
rect 1354 -4438 1358 -4434
rect 1354 -4452 1358 -4448
rect 1374 -4416 1378 -4412
rect 1384 -4459 1388 -4455
rect 1398 -4409 1402 -4405
rect 1408 -4423 1412 -4419
rect 1418 -4459 1422 -4455
rect 1432 -4409 1436 -4405
rect 1436 -4467 1440 -4463
rect 1452 -4438 1456 -4434
rect 1462 -4452 1466 -4448
rect 1476 -4409 1480 -4405
rect 1476 -4430 1480 -4426
rect 1480 -4445 1484 -4441
rect 1496 -4452 1500 -4448
rect 1510 -4409 1514 -4405
rect 1520 -4460 1524 -4456
rect 1536 -4467 1540 -4463
rect 1550 -4423 1554 -4419
rect 1554 -4460 1558 -4456
rect -1257 -4569 -1253 -4565
rect -1253 -4583 -1249 -4579
rect -1237 -4561 -1233 -4557
rect -1237 -4590 -1233 -4586
rect -1223 -4569 -1219 -4565
rect -1213 -4576 -1209 -4572
rect -1199 -4561 -1195 -4557
rect -1195 -4590 -1191 -4586
rect -1171 -4569 -1167 -4565
rect -1181 -4576 -1177 -4572
rect -1157 -4590 -1153 -4586
rect -1139 -4561 -1135 -4557
rect -1129 -4576 -1125 -4572
rect -1139 -4583 -1135 -4579
rect -1115 -4561 -1111 -4557
rect -1111 -4569 -1107 -4565
rect -1097 -4576 -1093 -4572
rect -1087 -4583 -1083 -4579
rect -1073 -4569 -1069 -4565
rect -928 -4569 -924 -4565
rect -924 -4583 -920 -4579
rect -908 -4561 -904 -4557
rect -908 -4590 -904 -4586
rect -894 -4569 -890 -4565
rect -884 -4576 -880 -4572
rect -870 -4561 -866 -4557
rect -866 -4590 -862 -4586
rect -842 -4569 -838 -4565
rect -852 -4576 -848 -4572
rect -828 -4590 -824 -4586
rect -810 -4561 -806 -4557
rect -800 -4576 -796 -4572
rect -810 -4583 -806 -4579
rect -786 -4561 -782 -4557
rect -782 -4569 -778 -4565
rect -768 -4576 -764 -4572
rect -758 -4583 -754 -4579
rect -744 -4569 -740 -4565
rect -570 -4569 -566 -4565
rect -566 -4583 -562 -4579
rect -550 -4561 -546 -4557
rect -550 -4590 -546 -4586
rect -536 -4569 -532 -4565
rect -526 -4576 -522 -4572
rect -512 -4561 -508 -4557
rect -508 -4590 -504 -4586
rect -484 -4569 -480 -4565
rect -494 -4576 -490 -4572
rect -470 -4590 -466 -4586
rect -452 -4561 -448 -4557
rect -442 -4576 -438 -4572
rect -452 -4583 -448 -4579
rect -428 -4561 -424 -4557
rect -424 -4569 -420 -4565
rect -410 -4576 -406 -4572
rect -400 -4583 -396 -4579
rect -386 -4569 -382 -4565
rect -1257 -4690 -1253 -4686
rect -1253 -4704 -1249 -4700
rect -1237 -4682 -1233 -4678
rect -1237 -4711 -1233 -4707
rect -1223 -4690 -1219 -4686
rect -1213 -4697 -1209 -4693
rect -1199 -4682 -1195 -4678
rect -1195 -4711 -1191 -4707
rect -1171 -4690 -1167 -4686
rect -1181 -4697 -1177 -4693
rect -1157 -4711 -1153 -4707
rect -1139 -4682 -1135 -4678
rect -1129 -4697 -1125 -4693
rect -1139 -4704 -1135 -4700
rect -1115 -4682 -1111 -4678
rect -1111 -4690 -1107 -4686
rect -1097 -4697 -1093 -4693
rect -1087 -4704 -1083 -4700
rect -1073 -4690 -1069 -4686
rect -928 -4690 -924 -4686
rect -924 -4704 -920 -4700
rect -908 -4682 -904 -4678
rect -908 -4711 -904 -4707
rect -894 -4690 -890 -4686
rect -884 -4697 -880 -4693
rect -870 -4682 -866 -4678
rect -866 -4711 -862 -4707
rect -842 -4690 -838 -4686
rect -852 -4697 -848 -4693
rect -828 -4711 -824 -4707
rect -810 -4682 -806 -4678
rect -800 -4697 -796 -4693
rect -810 -4704 -806 -4700
rect -786 -4682 -782 -4678
rect -782 -4690 -778 -4686
rect -768 -4697 -764 -4693
rect -758 -4704 -754 -4700
rect -744 -4690 -740 -4686
rect -570 -4690 -566 -4686
rect -566 -4704 -562 -4700
rect -550 -4682 -546 -4678
rect -550 -4711 -546 -4707
rect -536 -4690 -532 -4686
rect -526 -4697 -522 -4693
rect -512 -4682 -508 -4678
rect -508 -4711 -504 -4707
rect -484 -4690 -480 -4686
rect -494 -4697 -490 -4693
rect -470 -4711 -466 -4707
rect -452 -4682 -448 -4678
rect -442 -4697 -438 -4693
rect -452 -4704 -448 -4700
rect -428 -4682 -424 -4678
rect -424 -4690 -420 -4686
rect -410 -4697 -406 -4693
rect -400 -4704 -396 -4700
rect -386 -4690 -382 -4686
rect -212 -4690 -208 -4686
rect -208 -4704 -204 -4700
rect -192 -4682 -188 -4678
rect -192 -4711 -188 -4707
rect -178 -4690 -174 -4686
rect -168 -4697 -164 -4693
rect -154 -4682 -150 -4678
rect -150 -4711 -146 -4707
rect -126 -4690 -122 -4686
rect -136 -4697 -132 -4693
rect -112 -4711 -108 -4707
rect -94 -4682 -90 -4678
rect -84 -4697 -80 -4693
rect -94 -4704 -90 -4700
rect -70 -4682 -66 -4678
rect -66 -4690 -62 -4686
rect -52 -4697 -48 -4693
rect -42 -4704 -38 -4700
rect -28 -4690 -24 -4686
rect 216 -4690 220 -4686
rect 220 -4704 224 -4700
rect 236 -4682 240 -4678
rect 236 -4711 240 -4707
rect 250 -4690 254 -4686
rect 260 -4697 264 -4693
rect 274 -4682 278 -4678
rect 278 -4711 282 -4707
rect 302 -4690 306 -4686
rect 292 -4697 296 -4693
rect 316 -4711 320 -4707
rect 334 -4682 338 -4678
rect 344 -4697 348 -4693
rect 334 -4704 338 -4700
rect 358 -4682 362 -4678
rect 362 -4690 366 -4686
rect 376 -4697 380 -4693
rect 386 -4704 390 -4700
rect 400 -4690 404 -4686
rect 572 -4690 576 -4686
rect 576 -4704 580 -4700
rect 592 -4682 596 -4678
rect 592 -4711 596 -4707
rect 606 -4690 610 -4686
rect 616 -4697 620 -4693
rect 630 -4682 634 -4678
rect 634 -4711 638 -4707
rect 658 -4690 662 -4686
rect 648 -4697 652 -4693
rect 672 -4711 676 -4707
rect 690 -4682 694 -4678
rect 700 -4697 704 -4693
rect 690 -4704 694 -4700
rect 714 -4682 718 -4678
rect 718 -4690 722 -4686
rect 732 -4697 736 -4693
rect 742 -4704 746 -4700
rect 756 -4690 760 -4686
rect 970 -4690 974 -4686
rect 974 -4704 978 -4700
rect 990 -4682 994 -4678
rect 990 -4711 994 -4707
rect 1004 -4690 1008 -4686
rect 1014 -4697 1018 -4693
rect 1028 -4682 1032 -4678
rect 1032 -4711 1036 -4707
rect 1056 -4690 1060 -4686
rect 1046 -4697 1050 -4693
rect 1070 -4711 1074 -4707
rect 1088 -4682 1092 -4678
rect 1098 -4697 1102 -4693
rect 1088 -4704 1092 -4700
rect 1112 -4682 1116 -4678
rect 1116 -4690 1120 -4686
rect 1130 -4697 1134 -4693
rect 1140 -4704 1144 -4700
rect 1154 -4690 1158 -4686
rect 1328 -4690 1332 -4686
rect 1332 -4704 1336 -4700
rect 1348 -4682 1352 -4678
rect 1348 -4711 1352 -4707
rect 1362 -4690 1366 -4686
rect 1372 -4697 1376 -4693
rect 1386 -4682 1390 -4678
rect 1390 -4711 1394 -4707
rect 1414 -4690 1418 -4686
rect 1404 -4697 1408 -4693
rect 1428 -4711 1432 -4707
rect 1446 -4682 1450 -4678
rect 1456 -4697 1460 -4693
rect 1446 -4704 1450 -4700
rect 1470 -4682 1474 -4678
rect 1474 -4690 1478 -4686
rect 1488 -4697 1492 -4693
rect 1498 -4704 1502 -4700
rect 1512 -4690 1516 -4686
rect -1257 -4811 -1253 -4807
rect -1253 -4825 -1249 -4821
rect -1237 -4803 -1233 -4799
rect -1237 -4832 -1233 -4828
rect -1223 -4811 -1219 -4807
rect -1213 -4818 -1209 -4814
rect -1199 -4803 -1195 -4799
rect -1195 -4832 -1191 -4828
rect -1171 -4811 -1167 -4807
rect -1181 -4818 -1177 -4814
rect -1157 -4832 -1153 -4828
rect -1139 -4803 -1135 -4799
rect -1129 -4818 -1125 -4814
rect -1139 -4825 -1135 -4821
rect -1115 -4803 -1111 -4799
rect -1111 -4811 -1107 -4807
rect -1097 -4818 -1093 -4814
rect -1087 -4825 -1083 -4821
rect -1073 -4811 -1069 -4807
rect -928 -4811 -924 -4807
rect -924 -4825 -920 -4821
rect -908 -4803 -904 -4799
rect -908 -4832 -904 -4828
rect -894 -4811 -890 -4807
rect -884 -4818 -880 -4814
rect -870 -4803 -866 -4799
rect -866 -4832 -862 -4828
rect -842 -4811 -838 -4807
rect -852 -4818 -848 -4814
rect -828 -4832 -824 -4828
rect -810 -4803 -806 -4799
rect -800 -4818 -796 -4814
rect -810 -4825 -806 -4821
rect -786 -4803 -782 -4799
rect -782 -4811 -778 -4807
rect -768 -4818 -764 -4814
rect -758 -4825 -754 -4821
rect -744 -4811 -740 -4807
rect -570 -4811 -566 -4807
rect -566 -4825 -562 -4821
rect -550 -4803 -546 -4799
rect -550 -4832 -546 -4828
rect -536 -4811 -532 -4807
rect -526 -4818 -522 -4814
rect -512 -4803 -508 -4799
rect -508 -4832 -504 -4828
rect -484 -4811 -480 -4807
rect -494 -4818 -490 -4814
rect -470 -4832 -466 -4828
rect -452 -4803 -448 -4799
rect -442 -4818 -438 -4814
rect -452 -4825 -448 -4821
rect -428 -4803 -424 -4799
rect -424 -4811 -420 -4807
rect -410 -4818 -406 -4814
rect -400 -4825 -396 -4821
rect -386 -4811 -382 -4807
rect -212 -4811 -208 -4807
rect -208 -4825 -204 -4821
rect -192 -4803 -188 -4799
rect -192 -4832 -188 -4828
rect -178 -4811 -174 -4807
rect -168 -4818 -164 -4814
rect -154 -4803 -150 -4799
rect -150 -4832 -146 -4828
rect -126 -4811 -122 -4807
rect -136 -4818 -132 -4814
rect -112 -4832 -108 -4828
rect -94 -4803 -90 -4799
rect -84 -4818 -80 -4814
rect -94 -4825 -90 -4821
rect -70 -4803 -66 -4799
rect -66 -4811 -62 -4807
rect -52 -4818 -48 -4814
rect -42 -4825 -38 -4821
rect -28 -4811 -24 -4807
rect 91 -4812 95 -4796
rect 216 -4811 220 -4807
rect 220 -4825 224 -4821
rect 236 -4803 240 -4799
rect 236 -4832 240 -4828
rect 250 -4811 254 -4807
rect 260 -4818 264 -4814
rect 274 -4803 278 -4799
rect 278 -4832 282 -4828
rect 302 -4811 306 -4807
rect 292 -4818 296 -4814
rect 316 -4832 320 -4828
rect 334 -4803 338 -4799
rect 344 -4818 348 -4814
rect 334 -4825 338 -4821
rect 358 -4803 362 -4799
rect 362 -4811 366 -4807
rect 376 -4818 380 -4814
rect 386 -4825 390 -4821
rect 400 -4811 404 -4807
rect 572 -4811 576 -4807
rect 576 -4825 580 -4821
rect 592 -4803 596 -4799
rect 592 -4832 596 -4828
rect 606 -4811 610 -4807
rect 616 -4818 620 -4814
rect 630 -4803 634 -4799
rect 634 -4832 638 -4828
rect 658 -4811 662 -4807
rect 648 -4818 652 -4814
rect 672 -4832 676 -4828
rect 690 -4803 694 -4799
rect 700 -4818 704 -4814
rect 690 -4825 694 -4821
rect 714 -4803 718 -4799
rect 718 -4811 722 -4807
rect 732 -4818 736 -4814
rect 742 -4825 746 -4821
rect 756 -4811 760 -4807
rect 970 -4811 974 -4807
rect 974 -4825 978 -4821
rect 990 -4803 994 -4799
rect 990 -4832 994 -4828
rect 1004 -4811 1008 -4807
rect 1014 -4818 1018 -4814
rect 1028 -4803 1032 -4799
rect 1032 -4832 1036 -4828
rect 1056 -4811 1060 -4807
rect 1046 -4818 1050 -4814
rect 1070 -4832 1074 -4828
rect 1088 -4803 1092 -4799
rect 1098 -4818 1102 -4814
rect 1088 -4825 1092 -4821
rect 1112 -4803 1116 -4799
rect 1116 -4811 1120 -4807
rect 1130 -4818 1134 -4814
rect 1140 -4825 1144 -4821
rect 1154 -4811 1158 -4807
rect 1328 -4811 1332 -4807
rect 1332 -4825 1336 -4821
rect 1348 -4803 1352 -4799
rect 1348 -4832 1352 -4828
rect 1362 -4811 1366 -4807
rect 1372 -4818 1376 -4814
rect 1386 -4803 1390 -4799
rect 1390 -4832 1394 -4828
rect 1414 -4811 1418 -4807
rect 1404 -4818 1408 -4814
rect 1428 -4832 1432 -4828
rect 1446 -4803 1450 -4799
rect 1456 -4818 1460 -4814
rect 1446 -4825 1450 -4821
rect 1470 -4803 1474 -4799
rect 1474 -4811 1478 -4807
rect 1488 -4818 1492 -4814
rect 1498 -4825 1502 -4821
rect 1512 -4811 1516 -4807
rect -1257 -4929 -1253 -4925
rect -1253 -4943 -1249 -4939
rect -1237 -4921 -1233 -4917
rect -1237 -4950 -1233 -4946
rect -1223 -4929 -1219 -4925
rect -1213 -4936 -1209 -4932
rect -1199 -4921 -1195 -4917
rect -1195 -4950 -1191 -4946
rect -1171 -4929 -1167 -4925
rect -1181 -4936 -1177 -4932
rect -1157 -4950 -1153 -4946
rect -1139 -4921 -1135 -4917
rect -1129 -4936 -1125 -4932
rect -1139 -4943 -1135 -4939
rect -1115 -4921 -1111 -4917
rect -1111 -4929 -1107 -4925
rect -1097 -4936 -1093 -4932
rect -1087 -4943 -1083 -4939
rect -1073 -4929 -1069 -4925
rect -928 -4929 -924 -4925
rect -924 -4943 -920 -4939
rect -908 -4921 -904 -4917
rect -908 -4950 -904 -4946
rect -894 -4929 -890 -4925
rect -884 -4936 -880 -4932
rect -870 -4921 -866 -4917
rect -866 -4950 -862 -4946
rect -842 -4929 -838 -4925
rect -852 -4936 -848 -4932
rect -828 -4950 -824 -4946
rect -810 -4921 -806 -4917
rect -800 -4936 -796 -4932
rect -810 -4943 -806 -4939
rect -786 -4921 -782 -4917
rect -782 -4929 -778 -4925
rect -768 -4936 -764 -4932
rect -758 -4943 -754 -4939
rect -744 -4929 -740 -4925
rect -570 -4929 -566 -4925
rect -566 -4943 -562 -4939
rect -550 -4921 -546 -4917
rect -550 -4950 -546 -4946
rect -536 -4929 -532 -4925
rect -526 -4936 -522 -4932
rect -512 -4921 -508 -4917
rect -508 -4950 -504 -4946
rect -484 -4929 -480 -4925
rect -494 -4936 -490 -4932
rect -470 -4950 -466 -4946
rect -452 -4921 -448 -4917
rect -442 -4936 -438 -4932
rect -452 -4943 -448 -4939
rect -428 -4921 -424 -4917
rect -424 -4929 -420 -4925
rect -410 -4936 -406 -4932
rect -400 -4943 -396 -4939
rect -386 -4929 -382 -4925
rect -212 -4929 -208 -4925
rect -208 -4943 -204 -4939
rect -192 -4921 -188 -4917
rect -192 -4950 -188 -4946
rect -178 -4929 -174 -4925
rect -168 -4936 -164 -4932
rect -154 -4921 -150 -4917
rect -150 -4950 -146 -4946
rect -126 -4929 -122 -4925
rect -136 -4936 -132 -4932
rect -112 -4950 -108 -4946
rect -94 -4921 -90 -4917
rect -84 -4936 -80 -4932
rect -94 -4943 -90 -4939
rect -70 -4921 -66 -4917
rect -66 -4929 -62 -4925
rect -52 -4936 -48 -4932
rect -42 -4943 -38 -4939
rect -28 -4929 -24 -4925
rect 216 -4929 220 -4925
rect 220 -4943 224 -4939
rect 236 -4921 240 -4917
rect 236 -4950 240 -4946
rect 250 -4929 254 -4925
rect 260 -4936 264 -4932
rect 274 -4921 278 -4917
rect 278 -4950 282 -4946
rect 302 -4929 306 -4925
rect 292 -4936 296 -4932
rect 316 -4950 320 -4946
rect 334 -4921 338 -4917
rect 344 -4936 348 -4932
rect 334 -4943 338 -4939
rect 358 -4921 362 -4917
rect 362 -4929 366 -4925
rect 376 -4936 380 -4932
rect 386 -4943 390 -4939
rect 400 -4929 404 -4925
rect -1338 -5022 -1334 -5018
rect -1327 -5030 -1323 -5026
rect -1320 -5052 -1316 -5048
rect -934 -5022 -930 -5018
rect -923 -5030 -919 -5026
rect -916 -5052 -912 -5048
rect -576 -5022 -572 -5018
rect -565 -5030 -561 -5026
rect -558 -5052 -554 -5048
rect -218 -5022 -214 -5018
rect -207 -5030 -203 -5026
rect -200 -5052 -196 -5048
rect 210 -5022 214 -5018
rect 221 -5030 225 -5026
rect 228 -5052 232 -5048
rect 566 -5022 570 -5018
rect 577 -5030 581 -5026
rect 584 -5052 588 -5048
rect 964 -5022 968 -5018
rect 975 -5030 979 -5026
rect 982 -5052 986 -5048
rect 1322 -5022 1326 -5018
rect 1333 -5030 1337 -5026
rect 1340 -5052 1344 -5048
rect -1253 -5165 -1249 -5161
rect -1257 -5172 -1253 -5168
rect -1237 -5152 -1233 -5148
rect -1227 -5172 -1223 -5168
rect -1213 -5165 -1209 -5161
rect -1203 -5158 -1199 -5154
rect -1193 -5165 -1189 -5161
rect -1179 -5172 -1175 -5168
rect -1175 -5186 -1171 -5182
rect -924 -5128 -920 -5124
rect -928 -5149 -924 -5145
rect -924 -5164 -920 -5160
rect -928 -5178 -924 -5174
rect -898 -5149 -894 -5145
rect -902 -5157 -898 -5153
rect -902 -5171 -898 -5167
rect -882 -5135 -878 -5131
rect -872 -5178 -868 -5174
rect -858 -5128 -854 -5124
rect -848 -5142 -844 -5138
rect -838 -5178 -834 -5174
rect -824 -5128 -820 -5124
rect -820 -5186 -816 -5182
rect -804 -5157 -800 -5153
rect -794 -5171 -790 -5167
rect -780 -5128 -776 -5124
rect -780 -5149 -776 -5145
rect -776 -5164 -772 -5160
rect -760 -5171 -756 -5167
rect -746 -5128 -742 -5124
rect -736 -5179 -732 -5175
rect -720 -5186 -716 -5182
rect -706 -5142 -702 -5138
rect -702 -5179 -698 -5175
rect -566 -5128 -562 -5124
rect -570 -5149 -566 -5145
rect -566 -5164 -562 -5160
rect -570 -5178 -566 -5174
rect -540 -5149 -536 -5145
rect -544 -5157 -540 -5153
rect -544 -5171 -540 -5167
rect -524 -5135 -520 -5131
rect -514 -5178 -510 -5174
rect -500 -5128 -496 -5124
rect -490 -5142 -486 -5138
rect -480 -5178 -476 -5174
rect -466 -5128 -462 -5124
rect -462 -5186 -458 -5182
rect -446 -5157 -442 -5153
rect -436 -5171 -432 -5167
rect -422 -5128 -418 -5124
rect -422 -5149 -418 -5145
rect -418 -5164 -414 -5160
rect -402 -5171 -398 -5167
rect -388 -5128 -384 -5124
rect -378 -5179 -374 -5175
rect -362 -5186 -358 -5182
rect -348 -5142 -344 -5138
rect -344 -5179 -340 -5175
rect -208 -5128 -204 -5124
rect -212 -5149 -208 -5145
rect -208 -5164 -204 -5160
rect -212 -5178 -208 -5174
rect -182 -5149 -178 -5145
rect -186 -5157 -182 -5153
rect -186 -5171 -182 -5167
rect -166 -5135 -162 -5131
rect -156 -5178 -152 -5174
rect -142 -5128 -138 -5124
rect -132 -5142 -128 -5138
rect -122 -5178 -118 -5174
rect -108 -5128 -104 -5124
rect -104 -5186 -100 -5182
rect -88 -5157 -84 -5153
rect -78 -5171 -74 -5167
rect -64 -5128 -60 -5124
rect -64 -5149 -60 -5145
rect -60 -5164 -56 -5160
rect -44 -5171 -40 -5167
rect -30 -5128 -26 -5124
rect -20 -5179 -16 -5175
rect -4 -5186 0 -5182
rect 10 -5142 14 -5138
rect 14 -5179 18 -5175
rect 220 -5128 224 -5124
rect 216 -5149 220 -5145
rect 220 -5164 224 -5160
rect 216 -5178 220 -5174
rect 246 -5149 250 -5145
rect 242 -5157 246 -5153
rect 242 -5171 246 -5167
rect 262 -5135 266 -5131
rect 272 -5178 276 -5174
rect 286 -5128 290 -5124
rect 296 -5142 300 -5138
rect 306 -5178 310 -5174
rect 320 -5128 324 -5124
rect 324 -5186 328 -5182
rect 340 -5157 344 -5153
rect 350 -5171 354 -5167
rect 364 -5128 368 -5124
rect 364 -5149 368 -5145
rect 368 -5164 372 -5160
rect 384 -5171 388 -5167
rect 398 -5128 402 -5124
rect 408 -5179 412 -5175
rect 424 -5186 428 -5182
rect 438 -5142 442 -5138
rect 442 -5179 446 -5175
rect 576 -5128 580 -5124
rect 572 -5149 576 -5145
rect 576 -5164 580 -5160
rect 572 -5178 576 -5174
rect 602 -5149 606 -5145
rect 598 -5157 602 -5153
rect 598 -5171 602 -5167
rect 618 -5135 622 -5131
rect 628 -5178 632 -5174
rect 642 -5128 646 -5124
rect 652 -5142 656 -5138
rect 662 -5178 666 -5174
rect 676 -5128 680 -5124
rect 680 -5186 684 -5182
rect 696 -5157 700 -5153
rect 706 -5171 710 -5167
rect 720 -5128 724 -5124
rect 720 -5149 724 -5145
rect 724 -5164 728 -5160
rect 740 -5171 744 -5167
rect 754 -5128 758 -5124
rect 764 -5179 768 -5175
rect 780 -5186 784 -5182
rect 794 -5142 798 -5138
rect 798 -5179 802 -5175
rect 974 -5128 978 -5124
rect 970 -5149 974 -5145
rect 974 -5164 978 -5160
rect 970 -5178 974 -5174
rect 1000 -5149 1004 -5145
rect 996 -5157 1000 -5153
rect 996 -5171 1000 -5167
rect 1016 -5135 1020 -5131
rect 1026 -5178 1030 -5174
rect 1040 -5128 1044 -5124
rect 1050 -5142 1054 -5138
rect 1060 -5178 1064 -5174
rect 1074 -5128 1078 -5124
rect 1078 -5186 1082 -5182
rect 1094 -5157 1098 -5153
rect 1104 -5171 1108 -5167
rect 1118 -5128 1122 -5124
rect 1118 -5149 1122 -5145
rect 1122 -5164 1126 -5160
rect 1138 -5171 1142 -5167
rect 1152 -5128 1156 -5124
rect 1162 -5179 1166 -5175
rect 1178 -5186 1182 -5182
rect 1192 -5142 1196 -5138
rect 1196 -5179 1200 -5175
rect 1332 -5128 1336 -5124
rect 1328 -5149 1332 -5145
rect 1332 -5164 1336 -5160
rect 1328 -5178 1332 -5174
rect 1358 -5149 1362 -5145
rect 1354 -5157 1358 -5153
rect 1354 -5171 1358 -5167
rect 1374 -5135 1378 -5131
rect 1384 -5178 1388 -5174
rect 1398 -5128 1402 -5124
rect 1408 -5142 1412 -5138
rect 1418 -5178 1422 -5174
rect 1432 -5128 1436 -5124
rect 1436 -5186 1440 -5182
rect 1452 -5157 1456 -5153
rect 1462 -5171 1466 -5167
rect 1476 -5128 1480 -5124
rect 1476 -5149 1480 -5145
rect 1480 -5164 1484 -5160
rect 1496 -5171 1500 -5167
rect 1510 -5128 1514 -5124
rect 1520 -5179 1524 -5175
rect 1536 -5186 1540 -5182
rect 1550 -5142 1554 -5138
rect 1554 -5179 1558 -5175
rect -1257 -5284 -1253 -5280
rect -1253 -5298 -1249 -5294
rect -1237 -5276 -1233 -5272
rect -1237 -5305 -1233 -5301
rect -1223 -5284 -1219 -5280
rect -1213 -5291 -1209 -5287
rect -1199 -5276 -1195 -5272
rect -1195 -5305 -1191 -5301
rect -1171 -5284 -1167 -5280
rect -1181 -5291 -1177 -5287
rect -1157 -5305 -1153 -5301
rect -1139 -5276 -1135 -5272
rect -1129 -5291 -1125 -5287
rect -1139 -5298 -1135 -5294
rect -1115 -5276 -1111 -5272
rect -1111 -5284 -1107 -5280
rect -1097 -5291 -1093 -5287
rect -1087 -5298 -1083 -5294
rect -1073 -5284 -1069 -5280
rect -928 -5284 -924 -5280
rect -924 -5298 -920 -5294
rect -908 -5276 -904 -5272
rect -908 -5305 -904 -5301
rect -894 -5284 -890 -5280
rect -884 -5291 -880 -5287
rect -870 -5276 -866 -5272
rect -866 -5305 -862 -5301
rect -842 -5284 -838 -5280
rect -852 -5291 -848 -5287
rect -828 -5305 -824 -5301
rect -810 -5276 -806 -5272
rect -800 -5291 -796 -5287
rect -810 -5298 -806 -5294
rect -786 -5276 -782 -5272
rect -782 -5284 -778 -5280
rect -768 -5291 -764 -5287
rect -758 -5298 -754 -5294
rect -744 -5284 -740 -5280
rect -1257 -5405 -1253 -5401
rect -1253 -5419 -1249 -5415
rect -1237 -5397 -1233 -5393
rect -1237 -5426 -1233 -5422
rect -1223 -5405 -1219 -5401
rect -1213 -5412 -1209 -5408
rect -1199 -5397 -1195 -5393
rect -1195 -5426 -1191 -5422
rect -1171 -5405 -1167 -5401
rect -1181 -5412 -1177 -5408
rect -1157 -5426 -1153 -5422
rect -1139 -5397 -1135 -5393
rect -1129 -5412 -1125 -5408
rect -1139 -5419 -1135 -5415
rect -1115 -5397 -1111 -5393
rect -1111 -5405 -1107 -5401
rect -1097 -5412 -1093 -5408
rect -1087 -5419 -1083 -5415
rect -1025 -5397 -1021 -5387
rect -1073 -5405 -1069 -5401
rect -928 -5405 -924 -5401
rect -924 -5419 -920 -5415
rect -908 -5397 -904 -5393
rect -908 -5426 -904 -5422
rect -894 -5405 -890 -5401
rect -884 -5412 -880 -5408
rect -870 -5397 -866 -5393
rect -866 -5426 -862 -5422
rect -842 -5405 -838 -5401
rect -852 -5412 -848 -5408
rect -828 -5426 -824 -5422
rect -810 -5397 -806 -5393
rect -800 -5412 -796 -5408
rect -810 -5419 -806 -5415
rect -786 -5397 -782 -5393
rect -782 -5405 -778 -5401
rect -768 -5412 -764 -5408
rect -758 -5419 -754 -5415
rect -744 -5405 -740 -5401
rect -672 -5402 -668 -5392
rect -570 -5405 -566 -5401
rect -566 -5419 -562 -5415
rect -550 -5397 -546 -5393
rect -550 -5426 -546 -5422
rect -536 -5405 -532 -5401
rect -526 -5412 -522 -5408
rect -512 -5397 -508 -5393
rect -508 -5426 -504 -5422
rect -484 -5405 -480 -5401
rect -494 -5412 -490 -5408
rect -470 -5426 -466 -5422
rect -452 -5397 -448 -5393
rect -442 -5412 -438 -5408
rect -452 -5419 -448 -5415
rect -428 -5397 -424 -5393
rect -424 -5405 -420 -5401
rect -410 -5412 -406 -5408
rect -400 -5419 -396 -5415
rect -386 -5405 -382 -5401
rect -326 -5403 -322 -5393
rect -212 -5405 -208 -5401
rect -208 -5419 -204 -5415
rect -192 -5397 -188 -5393
rect -192 -5426 -188 -5422
rect -178 -5405 -174 -5401
rect -168 -5412 -164 -5408
rect -154 -5397 -150 -5393
rect -150 -5426 -146 -5422
rect -126 -5405 -122 -5401
rect -136 -5412 -132 -5408
rect -112 -5426 -108 -5422
rect -94 -5397 -90 -5393
rect -84 -5412 -80 -5408
rect -94 -5419 -90 -5415
rect -70 -5397 -66 -5393
rect -66 -5405 -62 -5401
rect -52 -5412 -48 -5408
rect -42 -5419 -38 -5415
rect -28 -5405 -24 -5401
rect 216 -5405 220 -5401
rect 220 -5419 224 -5415
rect 236 -5397 240 -5393
rect 236 -5426 240 -5422
rect 250 -5405 254 -5401
rect 260 -5412 264 -5408
rect 274 -5397 278 -5393
rect 278 -5426 282 -5422
rect 302 -5405 306 -5401
rect 292 -5412 296 -5408
rect 316 -5426 320 -5422
rect 334 -5397 338 -5393
rect 344 -5412 348 -5408
rect 334 -5419 338 -5415
rect 358 -5397 362 -5393
rect 362 -5405 366 -5401
rect 376 -5412 380 -5408
rect 386 -5419 390 -5415
rect 467 -5397 471 -5387
rect 400 -5405 404 -5401
rect 572 -5405 576 -5401
rect 576 -5419 580 -5415
rect 592 -5397 596 -5393
rect 592 -5426 596 -5422
rect 606 -5405 610 -5401
rect 616 -5412 620 -5408
rect 630 -5397 634 -5393
rect 634 -5426 638 -5422
rect 658 -5405 662 -5401
rect 648 -5412 652 -5408
rect 672 -5426 676 -5422
rect 690 -5397 694 -5393
rect 700 -5412 704 -5408
rect 690 -5419 694 -5415
rect 714 -5397 718 -5393
rect 718 -5405 722 -5401
rect 732 -5412 736 -5408
rect 742 -5419 746 -5415
rect 756 -5405 760 -5401
rect 868 -5402 872 -5392
rect 970 -5405 974 -5401
rect 974 -5419 978 -5415
rect 990 -5397 994 -5393
rect 990 -5426 994 -5422
rect 1004 -5405 1008 -5401
rect 1014 -5412 1018 -5408
rect 1028 -5397 1032 -5393
rect 1032 -5426 1036 -5422
rect 1056 -5405 1060 -5401
rect 1046 -5412 1050 -5408
rect 1070 -5426 1074 -5422
rect 1088 -5397 1092 -5393
rect 1098 -5412 1102 -5408
rect 1088 -5419 1092 -5415
rect 1112 -5397 1116 -5393
rect 1116 -5405 1120 -5401
rect 1130 -5412 1134 -5408
rect 1140 -5419 1144 -5415
rect 1154 -5405 1158 -5401
rect 1211 -5406 1215 -5396
rect 1328 -5405 1332 -5401
rect 1332 -5419 1336 -5415
rect 1348 -5397 1352 -5393
rect 1348 -5426 1352 -5422
rect 1362 -5405 1366 -5401
rect 1372 -5412 1376 -5408
rect 1386 -5397 1390 -5393
rect 1390 -5426 1394 -5422
rect 1414 -5405 1418 -5401
rect 1404 -5412 1408 -5408
rect 1428 -5426 1432 -5422
rect 1446 -5397 1450 -5393
rect 1456 -5412 1460 -5408
rect 1446 -5419 1450 -5415
rect 1470 -5397 1474 -5393
rect 1474 -5405 1478 -5401
rect 1488 -5412 1492 -5408
rect 1498 -5419 1502 -5415
rect 1512 -5405 1516 -5401
rect -1257 -5525 -1253 -5521
rect -1253 -5539 -1249 -5535
rect -1237 -5517 -1233 -5513
rect -1237 -5546 -1233 -5542
rect -1223 -5525 -1219 -5521
rect -1213 -5532 -1209 -5528
rect -1199 -5517 -1195 -5513
rect -1195 -5546 -1191 -5542
rect -1171 -5525 -1167 -5521
rect -1181 -5532 -1177 -5528
rect -1157 -5546 -1153 -5542
rect -1139 -5517 -1135 -5513
rect -1129 -5532 -1125 -5528
rect -1139 -5539 -1135 -5535
rect -1115 -5517 -1111 -5513
rect -1111 -5525 -1107 -5521
rect -1097 -5532 -1093 -5528
rect -1087 -5539 -1083 -5535
rect -1073 -5525 -1069 -5521
rect -1025 -5522 -1021 -5512
rect -928 -5525 -924 -5521
rect -924 -5539 -920 -5535
rect -908 -5517 -904 -5513
rect -908 -5546 -904 -5542
rect -894 -5525 -890 -5521
rect -884 -5532 -880 -5528
rect -870 -5517 -866 -5513
rect -866 -5546 -862 -5542
rect -842 -5525 -838 -5521
rect -852 -5532 -848 -5528
rect -828 -5546 -824 -5542
rect -810 -5517 -806 -5513
rect -800 -5532 -796 -5528
rect -810 -5539 -806 -5535
rect -786 -5517 -782 -5513
rect -782 -5525 -778 -5521
rect -768 -5532 -764 -5528
rect -758 -5539 -754 -5535
rect -744 -5525 -740 -5521
rect -570 -5525 -566 -5521
rect -566 -5539 -562 -5535
rect -550 -5517 -546 -5513
rect -550 -5546 -546 -5542
rect -536 -5525 -532 -5521
rect -526 -5532 -522 -5528
rect -512 -5517 -508 -5513
rect -508 -5546 -504 -5542
rect -484 -5525 -480 -5521
rect -494 -5532 -490 -5528
rect -470 -5546 -466 -5542
rect -452 -5517 -448 -5513
rect -442 -5532 -438 -5528
rect -452 -5539 -448 -5535
rect -428 -5517 -424 -5513
rect -424 -5525 -420 -5521
rect -410 -5532 -406 -5528
rect -400 -5539 -396 -5535
rect -326 -5518 -322 -5508
rect -386 -5525 -382 -5521
rect -212 -5525 -208 -5521
rect -208 -5539 -204 -5535
rect -192 -5517 -188 -5513
rect -192 -5546 -188 -5542
rect -178 -5525 -174 -5521
rect -168 -5532 -164 -5528
rect -154 -5517 -150 -5513
rect -150 -5546 -146 -5542
rect -126 -5525 -122 -5521
rect -136 -5532 -132 -5528
rect -112 -5546 -108 -5542
rect -94 -5517 -90 -5513
rect -84 -5532 -80 -5528
rect -94 -5539 -90 -5535
rect -70 -5517 -66 -5513
rect -66 -5525 -62 -5521
rect -52 -5532 -48 -5528
rect -42 -5539 -38 -5535
rect -28 -5525 -24 -5521
rect 216 -5525 220 -5521
rect 220 -5539 224 -5535
rect 236 -5517 240 -5513
rect 236 -5546 240 -5542
rect 250 -5525 254 -5521
rect 260 -5532 264 -5528
rect 274 -5517 278 -5513
rect 278 -5546 282 -5542
rect 302 -5525 306 -5521
rect 292 -5532 296 -5528
rect 316 -5546 320 -5542
rect 334 -5517 338 -5513
rect 344 -5532 348 -5528
rect 334 -5539 338 -5535
rect 358 -5517 362 -5513
rect 362 -5525 366 -5521
rect 376 -5532 380 -5528
rect 386 -5539 390 -5535
rect 400 -5525 404 -5521
rect 467 -5522 471 -5512
rect 572 -5525 576 -5521
rect 576 -5539 580 -5535
rect 592 -5517 596 -5513
rect 592 -5546 596 -5542
rect 606 -5525 610 -5521
rect 616 -5532 620 -5528
rect 630 -5517 634 -5513
rect 634 -5546 638 -5542
rect 658 -5525 662 -5521
rect 648 -5532 652 -5528
rect 672 -5546 676 -5542
rect 690 -5517 694 -5513
rect 700 -5532 704 -5528
rect 690 -5539 694 -5535
rect 714 -5517 718 -5513
rect 718 -5525 722 -5521
rect 732 -5532 736 -5528
rect 742 -5539 746 -5535
rect 756 -5525 760 -5521
rect 970 -5525 974 -5521
rect 974 -5539 978 -5535
rect 990 -5517 994 -5513
rect 990 -5546 994 -5542
rect 1004 -5525 1008 -5521
rect 1014 -5532 1018 -5528
rect 1028 -5517 1032 -5513
rect 1032 -5546 1036 -5542
rect 1056 -5525 1060 -5521
rect 1046 -5532 1050 -5528
rect 1070 -5546 1074 -5542
rect 1088 -5517 1092 -5513
rect 1098 -5532 1102 -5528
rect 1088 -5539 1092 -5535
rect 1112 -5517 1116 -5513
rect 1116 -5525 1120 -5521
rect 1130 -5532 1134 -5528
rect 1140 -5539 1144 -5535
rect 1154 -5525 1158 -5521
rect 1211 -5522 1215 -5512
rect 1328 -5525 1332 -5521
rect 1332 -5539 1336 -5535
rect 1348 -5517 1352 -5513
rect 1348 -5546 1352 -5542
rect 1362 -5525 1366 -5521
rect 1372 -5532 1376 -5528
rect 1386 -5517 1390 -5513
rect 1390 -5546 1394 -5542
rect 1414 -5525 1418 -5521
rect 1404 -5532 1408 -5528
rect 1428 -5546 1432 -5542
rect 1446 -5517 1450 -5513
rect 1456 -5532 1460 -5528
rect 1446 -5539 1450 -5535
rect 1470 -5517 1474 -5513
rect 1474 -5525 1478 -5521
rect 1488 -5532 1492 -5528
rect 1498 -5539 1502 -5535
rect 1512 -5525 1516 -5521
rect -1257 -5642 -1253 -5638
rect -1253 -5656 -1249 -5652
rect -1237 -5634 -1233 -5630
rect -1237 -5663 -1233 -5659
rect -1223 -5642 -1219 -5638
rect -1213 -5649 -1209 -5645
rect -1199 -5634 -1195 -5630
rect -1195 -5663 -1191 -5659
rect -1171 -5642 -1167 -5638
rect -1181 -5649 -1177 -5645
rect -1157 -5663 -1153 -5659
rect -1139 -5634 -1135 -5630
rect -1129 -5649 -1125 -5645
rect -1139 -5656 -1135 -5652
rect -1115 -5634 -1111 -5630
rect -1111 -5642 -1107 -5638
rect -1097 -5649 -1093 -5645
rect -1087 -5656 -1083 -5652
rect -1073 -5642 -1069 -5638
rect -928 -5642 -924 -5638
rect -924 -5656 -920 -5652
rect -908 -5634 -904 -5630
rect -908 -5663 -904 -5659
rect -894 -5642 -890 -5638
rect -884 -5649 -880 -5645
rect -870 -5634 -866 -5630
rect -866 -5663 -862 -5659
rect -842 -5642 -838 -5638
rect -852 -5649 -848 -5645
rect -828 -5663 -824 -5659
rect -810 -5634 -806 -5630
rect -800 -5649 -796 -5645
rect -810 -5656 -806 -5652
rect -786 -5634 -782 -5630
rect -782 -5642 -778 -5638
rect -768 -5649 -764 -5645
rect -758 -5656 -754 -5652
rect -744 -5642 -740 -5638
rect -570 -5642 -566 -5638
rect -566 -5656 -562 -5652
rect -550 -5634 -546 -5630
rect -550 -5663 -546 -5659
rect -536 -5642 -532 -5638
rect -526 -5649 -522 -5645
rect -512 -5634 -508 -5630
rect -508 -5663 -504 -5659
rect -484 -5642 -480 -5638
rect -494 -5649 -490 -5645
rect -470 -5663 -466 -5659
rect -452 -5634 -448 -5630
rect -442 -5649 -438 -5645
rect -452 -5656 -448 -5652
rect -428 -5634 -424 -5630
rect -424 -5642 -420 -5638
rect -410 -5649 -406 -5645
rect -400 -5656 -396 -5652
rect -386 -5642 -382 -5638
rect -212 -5642 -208 -5638
rect -208 -5656 -204 -5652
rect -192 -5634 -188 -5630
rect -192 -5663 -188 -5659
rect -178 -5642 -174 -5638
rect -168 -5649 -164 -5645
rect -154 -5634 -150 -5630
rect -150 -5663 -146 -5659
rect -126 -5642 -122 -5638
rect -136 -5649 -132 -5645
rect -112 -5663 -108 -5659
rect -94 -5634 -90 -5630
rect -84 -5649 -80 -5645
rect -94 -5656 -90 -5652
rect -70 -5634 -66 -5630
rect -66 -5642 -62 -5638
rect -52 -5649 -48 -5645
rect -42 -5656 -38 -5652
rect -28 -5642 -24 -5638
rect 216 -5642 220 -5638
rect 220 -5656 224 -5652
rect 236 -5634 240 -5630
rect 236 -5663 240 -5659
rect 250 -5642 254 -5638
rect 260 -5649 264 -5645
rect 274 -5634 278 -5630
rect 278 -5663 282 -5659
rect 302 -5642 306 -5638
rect 292 -5649 296 -5645
rect 316 -5663 320 -5659
rect 334 -5634 338 -5630
rect 344 -5649 348 -5645
rect 334 -5656 338 -5652
rect 358 -5634 362 -5630
rect 362 -5642 366 -5638
rect 376 -5649 380 -5645
rect 386 -5656 390 -5652
rect 400 -5642 404 -5638
rect 572 -5642 576 -5638
rect 576 -5656 580 -5652
rect 592 -5634 596 -5630
rect 592 -5663 596 -5659
rect 606 -5642 610 -5638
rect 616 -5649 620 -5645
rect 630 -5634 634 -5630
rect 634 -5663 638 -5659
rect 658 -5642 662 -5638
rect 648 -5649 652 -5645
rect 672 -5663 676 -5659
rect 690 -5634 694 -5630
rect 700 -5649 704 -5645
rect 690 -5656 694 -5652
rect 714 -5634 718 -5630
rect 718 -5642 722 -5638
rect 732 -5649 736 -5645
rect 742 -5656 746 -5652
rect 756 -5642 760 -5638
rect -1338 -5735 -1334 -5731
rect -1327 -5743 -1323 -5739
rect -1320 -5765 -1316 -5761
rect -934 -5735 -930 -5731
rect -923 -5743 -919 -5739
rect -916 -5765 -912 -5761
rect -576 -5735 -572 -5731
rect -565 -5743 -561 -5739
rect -558 -5765 -554 -5761
rect -218 -5735 -214 -5731
rect -207 -5743 -203 -5739
rect -200 -5765 -196 -5761
rect 210 -5735 214 -5731
rect 221 -5743 225 -5739
rect 228 -5765 232 -5761
rect 566 -5735 570 -5731
rect 577 -5743 581 -5739
rect 584 -5765 588 -5761
rect 964 -5735 968 -5731
rect 975 -5743 979 -5739
rect 982 -5765 986 -5761
rect 1322 -5735 1326 -5731
rect 1333 -5743 1337 -5739
rect 1340 -5765 1344 -5761
rect -1253 -5878 -1249 -5874
rect -1257 -5885 -1253 -5881
rect -1237 -5865 -1233 -5861
rect -1227 -5885 -1223 -5881
rect -1213 -5878 -1209 -5874
rect -1203 -5871 -1199 -5867
rect -1193 -5878 -1189 -5874
rect -1179 -5885 -1175 -5881
rect -1175 -5899 -1171 -5895
rect -924 -5841 -920 -5837
rect -928 -5862 -924 -5858
rect -924 -5877 -920 -5873
rect -928 -5891 -924 -5887
rect -898 -5862 -894 -5858
rect -902 -5870 -898 -5866
rect -902 -5884 -898 -5880
rect -882 -5848 -878 -5844
rect -872 -5891 -868 -5887
rect -858 -5841 -854 -5837
rect -848 -5855 -844 -5851
rect -838 -5891 -834 -5887
rect -824 -5841 -820 -5837
rect -820 -5899 -816 -5895
rect -804 -5870 -800 -5866
rect -794 -5884 -790 -5880
rect -780 -5841 -776 -5837
rect -780 -5862 -776 -5858
rect -776 -5877 -772 -5873
rect -760 -5884 -756 -5880
rect -746 -5841 -742 -5837
rect -736 -5892 -732 -5888
rect -720 -5899 -716 -5895
rect -706 -5855 -702 -5851
rect -702 -5892 -698 -5888
rect -566 -5841 -562 -5837
rect -570 -5862 -566 -5858
rect -566 -5877 -562 -5873
rect -570 -5891 -566 -5887
rect -540 -5862 -536 -5858
rect -544 -5870 -540 -5866
rect -544 -5884 -540 -5880
rect -524 -5848 -520 -5844
rect -514 -5891 -510 -5887
rect -500 -5841 -496 -5837
rect -490 -5855 -486 -5851
rect -480 -5891 -476 -5887
rect -466 -5841 -462 -5837
rect -462 -5899 -458 -5895
rect -446 -5870 -442 -5866
rect -436 -5884 -432 -5880
rect -422 -5841 -418 -5837
rect -422 -5862 -418 -5858
rect -418 -5877 -414 -5873
rect -402 -5884 -398 -5880
rect -388 -5841 -384 -5837
rect -378 -5892 -374 -5888
rect -362 -5899 -358 -5895
rect -348 -5855 -344 -5851
rect -344 -5892 -340 -5888
rect -208 -5841 -204 -5837
rect -212 -5862 -208 -5858
rect -208 -5877 -204 -5873
rect -212 -5891 -208 -5887
rect -182 -5862 -178 -5858
rect -186 -5870 -182 -5866
rect -186 -5884 -182 -5880
rect -166 -5848 -162 -5844
rect -156 -5891 -152 -5887
rect -142 -5841 -138 -5837
rect -132 -5855 -128 -5851
rect -122 -5891 -118 -5887
rect -108 -5841 -104 -5837
rect -104 -5899 -100 -5895
rect -88 -5870 -84 -5866
rect -78 -5884 -74 -5880
rect -64 -5841 -60 -5837
rect -64 -5862 -60 -5858
rect -60 -5877 -56 -5873
rect -44 -5884 -40 -5880
rect -30 -5841 -26 -5837
rect -20 -5892 -16 -5888
rect -4 -5899 0 -5895
rect 10 -5855 14 -5851
rect 14 -5892 18 -5888
rect 220 -5841 224 -5837
rect 216 -5862 220 -5858
rect 220 -5877 224 -5873
rect 216 -5891 220 -5887
rect 246 -5862 250 -5858
rect 242 -5870 246 -5866
rect 242 -5884 246 -5880
rect 262 -5848 266 -5844
rect 272 -5891 276 -5887
rect 286 -5841 290 -5837
rect 296 -5855 300 -5851
rect 306 -5891 310 -5887
rect 320 -5841 324 -5837
rect 324 -5899 328 -5895
rect 340 -5870 344 -5866
rect 350 -5884 354 -5880
rect 364 -5841 368 -5837
rect 364 -5862 368 -5858
rect 368 -5877 372 -5873
rect 384 -5884 388 -5880
rect 398 -5841 402 -5837
rect 408 -5892 412 -5888
rect 424 -5899 428 -5895
rect 438 -5855 442 -5851
rect 442 -5892 446 -5888
rect 576 -5841 580 -5837
rect 572 -5862 576 -5858
rect 576 -5877 580 -5873
rect 572 -5891 576 -5887
rect 602 -5862 606 -5858
rect 598 -5870 602 -5866
rect 598 -5884 602 -5880
rect 618 -5848 622 -5844
rect 628 -5891 632 -5887
rect 642 -5841 646 -5837
rect 652 -5855 656 -5851
rect 662 -5891 666 -5887
rect 676 -5841 680 -5837
rect 680 -5899 684 -5895
rect 696 -5870 700 -5866
rect 706 -5884 710 -5880
rect 720 -5841 724 -5837
rect 720 -5862 724 -5858
rect 724 -5877 728 -5873
rect 740 -5884 744 -5880
rect 754 -5841 758 -5837
rect 764 -5892 768 -5888
rect 780 -5899 784 -5895
rect 794 -5855 798 -5851
rect 798 -5892 802 -5888
rect 974 -5841 978 -5837
rect 970 -5862 974 -5858
rect 974 -5877 978 -5873
rect 970 -5891 974 -5887
rect 1000 -5862 1004 -5858
rect 996 -5870 1000 -5866
rect 996 -5884 1000 -5880
rect 1016 -5848 1020 -5844
rect 1026 -5891 1030 -5887
rect 1040 -5841 1044 -5837
rect 1050 -5855 1054 -5851
rect 1060 -5891 1064 -5887
rect 1074 -5841 1078 -5837
rect 1078 -5899 1082 -5895
rect 1094 -5870 1098 -5866
rect 1104 -5884 1108 -5880
rect 1118 -5841 1122 -5837
rect 1118 -5862 1122 -5858
rect 1122 -5877 1126 -5873
rect 1138 -5884 1142 -5880
rect 1152 -5841 1156 -5837
rect 1162 -5892 1166 -5888
rect 1178 -5899 1182 -5895
rect 1192 -5855 1196 -5851
rect 1196 -5892 1200 -5888
rect 1332 -5841 1336 -5837
rect 1328 -5862 1332 -5858
rect 1332 -5877 1336 -5873
rect 1328 -5891 1332 -5887
rect 1358 -5862 1362 -5858
rect 1354 -5870 1358 -5866
rect 1354 -5884 1358 -5880
rect 1374 -5848 1378 -5844
rect 1384 -5891 1388 -5887
rect 1398 -5841 1402 -5837
rect 1408 -5855 1412 -5851
rect 1418 -5891 1422 -5887
rect 1432 -5841 1436 -5837
rect 1436 -5899 1440 -5895
rect 1452 -5870 1456 -5866
rect 1462 -5884 1466 -5880
rect 1476 -5841 1480 -5837
rect 1476 -5862 1480 -5858
rect 1480 -5877 1484 -5873
rect 1496 -5884 1500 -5880
rect 1510 -5841 1514 -5837
rect 1520 -5892 1524 -5888
rect 1536 -5899 1540 -5895
rect 1550 -5855 1554 -5851
rect 1554 -5892 1558 -5888
rect -1257 -6001 -1253 -5997
rect -1253 -6015 -1249 -6011
rect -1237 -5993 -1233 -5989
rect -1237 -6022 -1233 -6018
rect -1223 -6001 -1219 -5997
rect -1213 -6008 -1209 -6004
rect -1199 -5993 -1195 -5989
rect -1195 -6022 -1191 -6018
rect -1171 -6001 -1167 -5997
rect -1181 -6008 -1177 -6004
rect -1157 -6022 -1153 -6018
rect -1139 -5993 -1135 -5989
rect -1129 -6008 -1125 -6004
rect -1139 -6015 -1135 -6011
rect -1115 -5993 -1111 -5989
rect -1111 -6001 -1107 -5997
rect -1097 -6008 -1093 -6004
rect -1087 -6015 -1083 -6011
rect -1073 -6001 -1069 -5997
rect -928 -6001 -924 -5997
rect -924 -6015 -920 -6011
rect -908 -5993 -904 -5989
rect -908 -6022 -904 -6018
rect -894 -6001 -890 -5997
rect -884 -6008 -880 -6004
rect -870 -5993 -866 -5989
rect -866 -6022 -862 -6018
rect -842 -6001 -838 -5997
rect -852 -6008 -848 -6004
rect -828 -6022 -824 -6018
rect -810 -5993 -806 -5989
rect -800 -6008 -796 -6004
rect -810 -6015 -806 -6011
rect -786 -5993 -782 -5989
rect -782 -6001 -778 -5997
rect -768 -6008 -764 -6004
rect -758 -6015 -754 -6011
rect -744 -6001 -740 -5997
rect -570 -6001 -566 -5997
rect -566 -6015 -562 -6011
rect -550 -5993 -546 -5989
rect -550 -6022 -546 -6018
rect -536 -6001 -532 -5997
rect -526 -6008 -522 -6004
rect -512 -5993 -508 -5989
rect -508 -6022 -504 -6018
rect -484 -6001 -480 -5997
rect -494 -6008 -490 -6004
rect -470 -6022 -466 -6018
rect -452 -5993 -448 -5989
rect -442 -6008 -438 -6004
rect -452 -6015 -448 -6011
rect -428 -5993 -424 -5989
rect -424 -6001 -420 -5997
rect -410 -6008 -406 -6004
rect -400 -6015 -396 -6011
rect -386 -6001 -382 -5997
rect -212 -6001 -208 -5997
rect -208 -6015 -204 -6011
rect -192 -5993 -188 -5989
rect -192 -6022 -188 -6018
rect -178 -6001 -174 -5997
rect -168 -6008 -164 -6004
rect -154 -5993 -150 -5989
rect -150 -6022 -146 -6018
rect -126 -6001 -122 -5997
rect -136 -6008 -132 -6004
rect -112 -6022 -108 -6018
rect -94 -5993 -90 -5989
rect -84 -6008 -80 -6004
rect -94 -6015 -90 -6011
rect -70 -5993 -66 -5989
rect -66 -6001 -62 -5997
rect -52 -6008 -48 -6004
rect -42 -6015 -38 -6011
rect -28 -6001 -24 -5997
rect 216 -6001 220 -5997
rect 220 -6015 224 -6011
rect 236 -5993 240 -5989
rect 236 -6022 240 -6018
rect 250 -6001 254 -5997
rect 260 -6008 264 -6004
rect 274 -5993 278 -5989
rect 278 -6022 282 -6018
rect 302 -6001 306 -5997
rect 292 -6008 296 -6004
rect 316 -6022 320 -6018
rect 334 -5993 338 -5989
rect 344 -6008 348 -6004
rect 334 -6015 338 -6011
rect 358 -5993 362 -5989
rect 362 -6001 366 -5997
rect 376 -6008 380 -6004
rect 386 -6015 390 -6011
rect 400 -6001 404 -5997
rect 572 -6001 576 -5997
rect 576 -6015 580 -6011
rect 592 -5993 596 -5989
rect 592 -6022 596 -6018
rect 606 -6001 610 -5997
rect 616 -6008 620 -6004
rect 630 -5993 634 -5989
rect 634 -6022 638 -6018
rect 658 -6001 662 -5997
rect 648 -6008 652 -6004
rect 672 -6022 676 -6018
rect 690 -5993 694 -5989
rect 700 -6008 704 -6004
rect 690 -6015 694 -6011
rect 714 -5993 718 -5989
rect 718 -6001 722 -5997
rect 732 -6008 736 -6004
rect 742 -6015 746 -6011
rect 756 -6001 760 -5997
rect 970 -6001 974 -5997
rect 974 -6015 978 -6011
rect 990 -5993 994 -5989
rect 990 -6022 994 -6018
rect 1004 -6001 1008 -5997
rect 1014 -6008 1018 -6004
rect 1028 -5993 1032 -5989
rect 1032 -6022 1036 -6018
rect 1056 -6001 1060 -5997
rect 1046 -6008 1050 -6004
rect 1070 -6022 1074 -6018
rect 1088 -5993 1092 -5989
rect 1098 -6008 1102 -6004
rect 1088 -6015 1092 -6011
rect 1112 -5993 1116 -5989
rect 1116 -6001 1120 -5997
rect 1130 -6008 1134 -6004
rect 1140 -6015 1144 -6011
rect 1154 -6001 1158 -5997
rect 1328 -6001 1332 -5997
rect 1332 -6015 1336 -6011
rect 1348 -5993 1352 -5989
rect 1348 -6022 1352 -6018
rect 1362 -6001 1366 -5997
rect 1372 -6008 1376 -6004
rect 1386 -5993 1390 -5989
rect 1390 -6022 1394 -6018
rect 1414 -6001 1418 -5997
rect 1404 -6008 1408 -6004
rect 1428 -6022 1432 -6018
rect 1446 -5993 1450 -5989
rect 1456 -6008 1460 -6004
rect 1446 -6015 1450 -6011
rect 1470 -5993 1474 -5989
rect 1474 -6001 1478 -5997
rect 1488 -6008 1492 -6004
rect 1498 -6015 1502 -6011
rect 1512 -6001 1516 -5997
rect 1328 -6119 1332 -6115
rect 1332 -6133 1336 -6129
rect 1348 -6111 1352 -6107
rect 1348 -6140 1352 -6136
rect 1362 -6119 1366 -6115
rect 1372 -6126 1376 -6122
rect 1386 -6111 1390 -6107
rect 1390 -6140 1394 -6136
rect 1414 -6119 1418 -6115
rect 1404 -6126 1408 -6122
rect 1428 -6140 1432 -6136
rect 1446 -6111 1450 -6107
rect 1456 -6126 1460 -6122
rect 1446 -6133 1450 -6129
rect 1470 -6111 1474 -6107
rect 1474 -6119 1478 -6115
rect 1488 -6126 1492 -6122
rect 1498 -6133 1502 -6129
rect 1512 -6119 1516 -6115
<< ndcontact >>
rect -1337 -1118 -1333 -1114
rect -1320 -1118 -1316 -1114
rect -1311 -1118 -1307 -1114
rect -936 -1118 -932 -1114
rect -919 -1118 -915 -1114
rect -910 -1118 -906 -1114
rect -577 -1118 -573 -1114
rect -560 -1118 -556 -1114
rect -551 -1118 -547 -1114
rect -219 -1118 -215 -1114
rect -202 -1118 -198 -1114
rect -193 -1118 -189 -1114
rect 209 -1118 213 -1114
rect 226 -1118 230 -1114
rect 235 -1118 239 -1114
rect 565 -1118 569 -1114
rect 582 -1118 586 -1114
rect 591 -1118 595 -1114
rect 963 -1118 967 -1114
rect 980 -1118 984 -1114
rect 989 -1118 993 -1114
rect 1321 -1118 1325 -1114
rect 1338 -1118 1342 -1114
rect 1347 -1118 1351 -1114
rect -1260 -1232 -1256 -1228
rect -1251 -1232 -1247 -1228
rect -1242 -1232 -1238 -1228
rect -1234 -1232 -1230 -1228
rect -1218 -1232 -1214 -1228
rect -1210 -1232 -1206 -1228
rect -1193 -1232 -1189 -1228
rect -1176 -1232 -1172 -1228
rect -1168 -1232 -1164 -1228
rect -1151 -1232 -1147 -1228
rect -1134 -1232 -1130 -1228
rect -1126 -1232 -1122 -1228
rect -1109 -1232 -1105 -1228
rect -1092 -1232 -1088 -1228
rect -1084 -1232 -1080 -1228
rect -1068 -1232 -1064 -1228
rect -935 -1232 -931 -1228
rect -926 -1232 -922 -1228
rect -917 -1232 -913 -1228
rect -909 -1232 -905 -1228
rect -893 -1232 -889 -1228
rect -885 -1232 -881 -1228
rect -868 -1232 -864 -1228
rect -851 -1232 -847 -1228
rect -843 -1232 -839 -1228
rect -826 -1232 -822 -1228
rect -809 -1232 -805 -1228
rect -801 -1232 -797 -1228
rect -784 -1232 -780 -1228
rect -767 -1232 -763 -1228
rect -759 -1232 -755 -1228
rect -743 -1232 -739 -1228
rect -577 -1232 -573 -1228
rect -568 -1232 -564 -1228
rect -559 -1232 -555 -1228
rect -551 -1232 -547 -1228
rect -535 -1232 -531 -1228
rect -527 -1232 -523 -1228
rect -510 -1232 -506 -1228
rect -493 -1232 -489 -1228
rect -485 -1232 -481 -1228
rect -468 -1232 -464 -1228
rect -451 -1232 -447 -1228
rect -443 -1232 -439 -1228
rect -426 -1232 -422 -1228
rect -409 -1232 -405 -1228
rect -401 -1232 -397 -1228
rect -385 -1232 -381 -1228
rect -219 -1232 -215 -1228
rect -210 -1232 -206 -1228
rect -201 -1232 -197 -1228
rect -193 -1232 -189 -1228
rect -177 -1232 -173 -1228
rect -169 -1232 -165 -1228
rect -152 -1232 -148 -1228
rect -135 -1232 -131 -1228
rect -127 -1232 -123 -1228
rect -110 -1232 -106 -1228
rect -93 -1232 -89 -1228
rect -85 -1232 -81 -1228
rect -68 -1232 -64 -1228
rect -51 -1232 -47 -1228
rect -43 -1232 -39 -1228
rect -27 -1232 -23 -1228
rect 209 -1232 213 -1228
rect 218 -1232 222 -1228
rect 227 -1232 231 -1228
rect 235 -1232 239 -1228
rect 251 -1232 255 -1228
rect 259 -1232 263 -1228
rect 276 -1232 280 -1228
rect 293 -1232 297 -1228
rect 301 -1232 305 -1228
rect 318 -1232 322 -1228
rect 335 -1232 339 -1228
rect 343 -1232 347 -1228
rect 360 -1232 364 -1228
rect 377 -1232 381 -1228
rect 385 -1232 389 -1228
rect 401 -1232 405 -1228
rect 565 -1232 569 -1228
rect 574 -1232 578 -1228
rect 583 -1232 587 -1228
rect 591 -1232 595 -1228
rect 607 -1232 611 -1228
rect 615 -1232 619 -1228
rect 632 -1232 636 -1228
rect 649 -1232 653 -1228
rect 657 -1232 661 -1228
rect 674 -1232 678 -1228
rect 691 -1232 695 -1228
rect 699 -1232 703 -1228
rect 716 -1232 720 -1228
rect 733 -1232 737 -1228
rect 741 -1232 745 -1228
rect 757 -1232 761 -1228
rect 963 -1232 967 -1228
rect 972 -1232 976 -1228
rect 981 -1232 985 -1228
rect 989 -1232 993 -1228
rect 1005 -1232 1009 -1228
rect 1013 -1232 1017 -1228
rect 1030 -1232 1034 -1228
rect 1047 -1232 1051 -1228
rect 1055 -1232 1059 -1228
rect 1072 -1232 1076 -1228
rect 1089 -1232 1093 -1228
rect 1097 -1232 1101 -1228
rect 1114 -1232 1118 -1228
rect 1131 -1232 1135 -1228
rect 1139 -1232 1143 -1228
rect 1155 -1232 1159 -1228
rect -1339 -1348 -1335 -1344
rect -1322 -1348 -1318 -1344
rect -1313 -1348 -1309 -1344
rect -935 -1348 -931 -1344
rect -918 -1348 -914 -1344
rect -909 -1348 -905 -1344
rect -577 -1348 -573 -1344
rect -560 -1348 -556 -1344
rect -551 -1348 -547 -1344
rect -219 -1348 -215 -1344
rect -202 -1348 -198 -1344
rect -193 -1348 -189 -1344
rect 209 -1348 213 -1344
rect 226 -1348 230 -1344
rect 235 -1348 239 -1344
rect 565 -1348 569 -1344
rect 582 -1348 586 -1344
rect 591 -1348 595 -1344
rect 963 -1348 967 -1344
rect 980 -1348 984 -1344
rect 989 -1348 993 -1344
rect 1321 -1348 1325 -1344
rect 1338 -1348 1342 -1344
rect 1347 -1348 1351 -1344
rect -1260 -1462 -1256 -1458
rect -1251 -1462 -1247 -1458
rect -1242 -1462 -1238 -1458
rect -1234 -1462 -1230 -1458
rect -1225 -1462 -1221 -1458
rect -1207 -1462 -1203 -1458
rect -1198 -1462 -1194 -1458
rect -1190 -1462 -1186 -1458
rect -1173 -1462 -1169 -1458
rect -1164 -1462 -1160 -1458
rect -935 -1462 -931 -1458
rect -926 -1462 -922 -1458
rect -917 -1462 -913 -1458
rect -909 -1462 -905 -1458
rect -900 -1462 -896 -1458
rect -891 -1462 -887 -1458
rect -883 -1462 -879 -1458
rect -875 -1462 -871 -1458
rect -857 -1462 -853 -1458
rect -847 -1462 -843 -1458
rect -839 -1462 -835 -1458
rect -822 -1462 -818 -1458
rect -813 -1462 -809 -1458
rect -805 -1462 -801 -1458
rect -796 -1462 -792 -1458
rect -778 -1462 -774 -1458
rect -769 -1462 -765 -1458
rect -761 -1462 -757 -1458
rect -745 -1462 -741 -1458
rect -737 -1462 -733 -1458
rect -725 -1462 -721 -1458
rect -713 -1462 -709 -1458
rect -704 -1462 -700 -1458
rect -695 -1462 -691 -1458
rect -577 -1462 -573 -1458
rect -568 -1462 -564 -1458
rect -559 -1462 -555 -1458
rect -551 -1462 -547 -1458
rect -542 -1462 -538 -1458
rect -533 -1462 -529 -1458
rect -525 -1462 -521 -1458
rect -517 -1462 -513 -1458
rect -499 -1462 -495 -1458
rect -489 -1462 -485 -1458
rect -481 -1462 -477 -1458
rect -464 -1462 -460 -1458
rect -455 -1462 -451 -1458
rect -447 -1462 -443 -1458
rect -438 -1462 -434 -1458
rect -420 -1462 -416 -1458
rect -411 -1462 -407 -1458
rect -403 -1462 -399 -1458
rect -387 -1462 -383 -1458
rect -379 -1462 -375 -1458
rect -367 -1462 -363 -1458
rect -355 -1462 -351 -1458
rect -346 -1462 -342 -1458
rect -337 -1462 -333 -1458
rect -219 -1462 -215 -1458
rect -210 -1462 -206 -1458
rect -201 -1462 -197 -1458
rect -193 -1462 -189 -1458
rect -184 -1462 -180 -1458
rect -175 -1462 -171 -1458
rect -167 -1462 -163 -1458
rect -159 -1462 -155 -1458
rect -141 -1462 -137 -1458
rect -131 -1462 -127 -1458
rect -123 -1462 -119 -1458
rect -106 -1462 -102 -1458
rect -97 -1462 -93 -1458
rect -89 -1462 -85 -1458
rect -80 -1462 -76 -1458
rect -62 -1462 -58 -1458
rect -53 -1462 -49 -1458
rect -45 -1462 -41 -1458
rect -29 -1462 -25 -1458
rect -21 -1462 -17 -1458
rect -9 -1462 -5 -1458
rect 3 -1462 7 -1458
rect 12 -1462 16 -1458
rect 21 -1462 25 -1458
rect 209 -1462 213 -1458
rect 218 -1462 222 -1458
rect 227 -1462 231 -1458
rect 235 -1462 239 -1458
rect 244 -1462 248 -1458
rect 253 -1462 257 -1458
rect 261 -1462 265 -1458
rect 269 -1462 273 -1458
rect 287 -1462 291 -1458
rect 297 -1462 301 -1458
rect 305 -1462 309 -1458
rect 322 -1462 326 -1458
rect 331 -1462 335 -1458
rect 339 -1462 343 -1458
rect 348 -1462 352 -1458
rect 366 -1462 370 -1458
rect 375 -1462 379 -1458
rect 383 -1462 387 -1458
rect 399 -1462 403 -1458
rect 407 -1462 411 -1458
rect 419 -1462 423 -1458
rect 431 -1462 435 -1458
rect 440 -1462 444 -1458
rect 449 -1462 453 -1458
rect 565 -1462 569 -1458
rect 574 -1462 578 -1458
rect 583 -1462 587 -1458
rect 591 -1462 595 -1458
rect 600 -1462 604 -1458
rect 609 -1462 613 -1458
rect 617 -1462 621 -1458
rect 625 -1462 629 -1458
rect 643 -1462 647 -1458
rect 653 -1462 657 -1458
rect 661 -1462 665 -1458
rect 678 -1462 682 -1458
rect 687 -1462 691 -1458
rect 695 -1462 699 -1458
rect 704 -1462 708 -1458
rect 722 -1462 726 -1458
rect 731 -1462 735 -1458
rect 739 -1462 743 -1458
rect 755 -1462 759 -1458
rect 763 -1462 767 -1458
rect 775 -1462 779 -1458
rect 787 -1462 791 -1458
rect 796 -1462 800 -1458
rect 805 -1462 809 -1458
rect 963 -1462 967 -1458
rect 972 -1462 976 -1458
rect 981 -1462 985 -1458
rect 989 -1462 993 -1458
rect 998 -1462 1002 -1458
rect 1007 -1462 1011 -1458
rect 1015 -1462 1019 -1458
rect 1023 -1462 1027 -1458
rect 1041 -1462 1045 -1458
rect 1051 -1462 1055 -1458
rect 1059 -1462 1063 -1458
rect 1076 -1462 1080 -1458
rect 1085 -1462 1089 -1458
rect 1093 -1462 1097 -1458
rect 1102 -1462 1106 -1458
rect 1120 -1462 1124 -1458
rect 1129 -1462 1133 -1458
rect 1137 -1462 1141 -1458
rect 1153 -1462 1157 -1458
rect 1161 -1462 1165 -1458
rect 1173 -1462 1177 -1458
rect 1185 -1462 1189 -1458
rect 1194 -1462 1198 -1458
rect 1203 -1462 1207 -1458
rect 1321 -1462 1325 -1458
rect 1330 -1462 1334 -1458
rect 1339 -1462 1343 -1458
rect 1347 -1462 1351 -1458
rect 1356 -1462 1360 -1458
rect 1374 -1462 1378 -1458
rect 1383 -1462 1387 -1458
rect 1391 -1462 1395 -1458
rect 1408 -1462 1412 -1458
rect 1417 -1462 1421 -1458
rect -1260 -1585 -1256 -1581
rect -1251 -1585 -1247 -1581
rect -1242 -1585 -1238 -1581
rect -1234 -1585 -1230 -1581
rect -1218 -1585 -1214 -1581
rect -1210 -1585 -1206 -1581
rect -1193 -1585 -1189 -1581
rect -1176 -1585 -1172 -1581
rect -1168 -1585 -1164 -1581
rect -1151 -1585 -1147 -1581
rect -1134 -1585 -1130 -1581
rect -1126 -1585 -1122 -1581
rect -1109 -1585 -1105 -1581
rect -1092 -1585 -1088 -1581
rect -1084 -1585 -1080 -1581
rect -1068 -1585 -1064 -1581
rect -935 -1585 -931 -1581
rect -926 -1585 -922 -1581
rect -917 -1585 -913 -1581
rect -909 -1585 -905 -1581
rect -893 -1585 -889 -1581
rect -885 -1585 -881 -1581
rect -868 -1585 -864 -1581
rect -851 -1585 -847 -1581
rect -843 -1585 -839 -1581
rect -826 -1585 -822 -1581
rect -809 -1585 -805 -1581
rect -801 -1585 -797 -1581
rect -784 -1585 -780 -1581
rect -767 -1585 -763 -1581
rect -759 -1585 -755 -1581
rect -743 -1585 -739 -1581
rect -577 -1585 -573 -1581
rect -568 -1585 -564 -1581
rect -559 -1585 -555 -1581
rect -551 -1585 -547 -1581
rect -535 -1585 -531 -1581
rect -527 -1585 -523 -1581
rect -510 -1585 -506 -1581
rect -493 -1585 -489 -1581
rect -485 -1585 -481 -1581
rect -468 -1585 -464 -1581
rect -451 -1585 -447 -1581
rect -443 -1585 -439 -1581
rect -426 -1585 -422 -1581
rect -409 -1585 -405 -1581
rect -401 -1585 -397 -1581
rect -385 -1585 -381 -1581
rect -219 -1585 -215 -1581
rect -210 -1585 -206 -1581
rect -201 -1585 -197 -1581
rect -193 -1585 -189 -1581
rect -177 -1585 -173 -1581
rect -169 -1585 -165 -1581
rect -152 -1585 -148 -1581
rect -135 -1585 -131 -1581
rect -127 -1585 -123 -1581
rect -110 -1585 -106 -1581
rect -93 -1585 -89 -1581
rect -85 -1585 -81 -1581
rect -68 -1585 -64 -1581
rect -51 -1585 -47 -1581
rect -43 -1585 -39 -1581
rect -27 -1585 -23 -1581
rect 209 -1585 213 -1581
rect 218 -1585 222 -1581
rect 227 -1585 231 -1581
rect 235 -1585 239 -1581
rect 251 -1585 255 -1581
rect 259 -1585 263 -1581
rect 276 -1585 280 -1581
rect 293 -1585 297 -1581
rect 301 -1585 305 -1581
rect 318 -1585 322 -1581
rect 335 -1585 339 -1581
rect 343 -1585 347 -1581
rect 360 -1585 364 -1581
rect 377 -1585 381 -1581
rect 385 -1585 389 -1581
rect 401 -1585 405 -1581
rect 565 -1585 569 -1581
rect 574 -1585 578 -1581
rect 583 -1585 587 -1581
rect 591 -1585 595 -1581
rect 607 -1585 611 -1581
rect 615 -1585 619 -1581
rect 632 -1585 636 -1581
rect 649 -1585 653 -1581
rect 657 -1585 661 -1581
rect 674 -1585 678 -1581
rect 691 -1585 695 -1581
rect 699 -1585 703 -1581
rect 716 -1585 720 -1581
rect 733 -1585 737 -1581
rect 741 -1585 745 -1581
rect 757 -1585 761 -1581
rect 963 -1585 967 -1581
rect 972 -1585 976 -1581
rect 981 -1585 985 -1581
rect 989 -1585 993 -1581
rect 1005 -1585 1009 -1581
rect 1013 -1585 1017 -1581
rect 1030 -1585 1034 -1581
rect 1047 -1585 1051 -1581
rect 1055 -1585 1059 -1581
rect 1072 -1585 1076 -1581
rect 1089 -1585 1093 -1581
rect 1097 -1585 1101 -1581
rect 1114 -1585 1118 -1581
rect 1131 -1585 1135 -1581
rect 1139 -1585 1143 -1581
rect 1155 -1585 1159 -1581
rect -1260 -1706 -1256 -1702
rect -1251 -1706 -1247 -1702
rect -1242 -1706 -1238 -1702
rect -1234 -1706 -1230 -1702
rect -1218 -1706 -1214 -1702
rect -1210 -1706 -1206 -1702
rect -1193 -1706 -1189 -1702
rect -1176 -1706 -1172 -1702
rect -1168 -1706 -1164 -1702
rect -1151 -1706 -1147 -1702
rect -1134 -1706 -1130 -1702
rect -1126 -1706 -1122 -1702
rect -1109 -1706 -1105 -1702
rect -1092 -1706 -1088 -1702
rect -1084 -1706 -1080 -1702
rect -1068 -1706 -1064 -1702
rect -935 -1706 -931 -1702
rect -926 -1706 -922 -1702
rect -917 -1706 -913 -1702
rect -909 -1706 -905 -1702
rect -893 -1706 -889 -1702
rect -885 -1706 -881 -1702
rect -868 -1706 -864 -1702
rect -851 -1706 -847 -1702
rect -843 -1706 -839 -1702
rect -826 -1706 -822 -1702
rect -809 -1706 -805 -1702
rect -801 -1706 -797 -1702
rect -784 -1706 -780 -1702
rect -767 -1706 -763 -1702
rect -759 -1706 -755 -1702
rect -743 -1706 -739 -1702
rect -577 -1706 -573 -1702
rect -568 -1706 -564 -1702
rect -559 -1706 -555 -1702
rect -551 -1706 -547 -1702
rect -535 -1706 -531 -1702
rect -527 -1706 -523 -1702
rect -510 -1706 -506 -1702
rect -493 -1706 -489 -1702
rect -485 -1706 -481 -1702
rect -468 -1706 -464 -1702
rect -451 -1706 -447 -1702
rect -443 -1706 -439 -1702
rect -426 -1706 -422 -1702
rect -409 -1706 -405 -1702
rect -401 -1706 -397 -1702
rect -385 -1706 -381 -1702
rect -219 -1706 -215 -1702
rect -210 -1706 -206 -1702
rect -201 -1706 -197 -1702
rect -193 -1706 -189 -1702
rect -177 -1706 -173 -1702
rect -169 -1706 -165 -1702
rect -152 -1706 -148 -1702
rect -135 -1706 -131 -1702
rect -127 -1706 -123 -1702
rect -110 -1706 -106 -1702
rect -93 -1706 -89 -1702
rect -85 -1706 -81 -1702
rect -68 -1706 -64 -1702
rect -51 -1706 -47 -1702
rect -43 -1706 -39 -1702
rect -27 -1706 -23 -1702
rect 209 -1706 213 -1702
rect 218 -1706 222 -1702
rect 227 -1706 231 -1702
rect 235 -1706 239 -1702
rect 251 -1706 255 -1702
rect 259 -1706 263 -1702
rect 276 -1706 280 -1702
rect 293 -1706 297 -1702
rect 301 -1706 305 -1702
rect 318 -1706 322 -1702
rect 335 -1706 339 -1702
rect 343 -1706 347 -1702
rect 360 -1706 364 -1702
rect 377 -1706 381 -1702
rect 385 -1706 389 -1702
rect 401 -1706 405 -1702
rect 565 -1706 569 -1702
rect 574 -1706 578 -1702
rect 583 -1706 587 -1702
rect 591 -1706 595 -1702
rect 607 -1706 611 -1702
rect 615 -1706 619 -1702
rect 632 -1706 636 -1702
rect 649 -1706 653 -1702
rect 657 -1706 661 -1702
rect 674 -1706 678 -1702
rect 691 -1706 695 -1702
rect 699 -1706 703 -1702
rect 716 -1706 720 -1702
rect 733 -1706 737 -1702
rect 741 -1706 745 -1702
rect 757 -1706 761 -1702
rect 963 -1706 967 -1702
rect 972 -1706 976 -1702
rect 981 -1706 985 -1702
rect 989 -1706 993 -1702
rect 1005 -1706 1009 -1702
rect 1013 -1706 1017 -1702
rect 1030 -1706 1034 -1702
rect 1047 -1706 1051 -1702
rect 1055 -1706 1059 -1702
rect 1072 -1706 1076 -1702
rect 1089 -1706 1093 -1702
rect 1097 -1706 1101 -1702
rect 1114 -1706 1118 -1702
rect 1131 -1706 1135 -1702
rect 1139 -1706 1143 -1702
rect 1155 -1706 1159 -1702
rect 1321 -1706 1325 -1702
rect 1330 -1706 1334 -1702
rect 1339 -1706 1343 -1702
rect 1347 -1706 1351 -1702
rect 1363 -1706 1367 -1702
rect 1371 -1706 1375 -1702
rect 1388 -1706 1392 -1702
rect 1405 -1706 1409 -1702
rect 1413 -1706 1417 -1702
rect 1430 -1706 1434 -1702
rect 1447 -1706 1451 -1702
rect 1455 -1706 1459 -1702
rect 1472 -1706 1476 -1702
rect 1489 -1706 1493 -1702
rect 1497 -1706 1501 -1702
rect 1513 -1706 1517 -1702
rect -1260 -1827 -1256 -1823
rect -1251 -1827 -1247 -1823
rect -1242 -1827 -1238 -1823
rect -1234 -1827 -1230 -1823
rect -1218 -1827 -1214 -1823
rect -1210 -1827 -1206 -1823
rect -1193 -1827 -1189 -1823
rect -1176 -1827 -1172 -1823
rect -1168 -1827 -1164 -1823
rect -1151 -1827 -1147 -1823
rect -1134 -1827 -1130 -1823
rect -1126 -1827 -1122 -1823
rect -1109 -1827 -1105 -1823
rect -1092 -1827 -1088 -1823
rect -1084 -1827 -1080 -1823
rect -1068 -1827 -1064 -1823
rect -1029 -1827 -1025 -1823
rect -1021 -1827 -1017 -1823
rect -935 -1827 -931 -1823
rect -926 -1827 -922 -1823
rect -917 -1827 -913 -1823
rect -909 -1827 -905 -1823
rect -893 -1827 -889 -1823
rect -885 -1827 -881 -1823
rect -868 -1827 -864 -1823
rect -851 -1827 -847 -1823
rect -843 -1827 -839 -1823
rect -826 -1827 -822 -1823
rect -809 -1827 -805 -1823
rect -801 -1827 -797 -1823
rect -784 -1827 -780 -1823
rect -767 -1827 -763 -1823
rect -759 -1827 -755 -1823
rect -743 -1827 -739 -1823
rect -577 -1827 -573 -1823
rect -568 -1827 -564 -1823
rect -559 -1827 -555 -1823
rect -551 -1827 -547 -1823
rect -535 -1827 -531 -1823
rect -527 -1827 -523 -1823
rect -510 -1827 -506 -1823
rect -493 -1827 -489 -1823
rect -485 -1827 -481 -1823
rect -468 -1827 -464 -1823
rect -451 -1827 -447 -1823
rect -443 -1827 -439 -1823
rect -426 -1827 -422 -1823
rect -409 -1827 -405 -1823
rect -401 -1827 -397 -1823
rect -385 -1827 -381 -1823
rect -332 -1827 -328 -1823
rect -324 -1827 -320 -1823
rect -219 -1827 -215 -1823
rect -210 -1827 -206 -1823
rect -201 -1827 -197 -1823
rect -193 -1827 -189 -1823
rect -177 -1827 -173 -1823
rect -169 -1827 -165 -1823
rect -152 -1827 -148 -1823
rect -135 -1827 -131 -1823
rect -127 -1827 -123 -1823
rect -110 -1827 -106 -1823
rect -93 -1827 -89 -1823
rect -85 -1827 -81 -1823
rect -68 -1827 -64 -1823
rect -51 -1827 -47 -1823
rect -43 -1827 -39 -1823
rect -27 -1827 -23 -1823
rect 209 -1827 213 -1823
rect 218 -1827 222 -1823
rect 227 -1827 231 -1823
rect 235 -1827 239 -1823
rect 251 -1827 255 -1823
rect 259 -1827 263 -1823
rect 276 -1827 280 -1823
rect 293 -1827 297 -1823
rect 301 -1827 305 -1823
rect 318 -1827 322 -1823
rect 335 -1827 339 -1823
rect 343 -1827 347 -1823
rect 360 -1827 364 -1823
rect 377 -1827 381 -1823
rect 385 -1827 389 -1823
rect 401 -1827 405 -1823
rect 464 -1827 468 -1823
rect 472 -1827 476 -1823
rect 565 -1827 569 -1823
rect 574 -1827 578 -1823
rect 583 -1827 587 -1823
rect 591 -1827 595 -1823
rect 607 -1827 611 -1823
rect 615 -1827 619 -1823
rect 632 -1827 636 -1823
rect 649 -1827 653 -1823
rect 657 -1827 661 -1823
rect 674 -1827 678 -1823
rect 691 -1827 695 -1823
rect 699 -1827 703 -1823
rect 716 -1827 720 -1823
rect 733 -1827 737 -1823
rect 741 -1827 745 -1823
rect 757 -1827 761 -1823
rect 963 -1827 967 -1823
rect 972 -1827 976 -1823
rect 981 -1827 985 -1823
rect 989 -1827 993 -1823
rect 1005 -1827 1009 -1823
rect 1013 -1827 1017 -1823
rect 1030 -1827 1034 -1823
rect 1047 -1827 1051 -1823
rect 1055 -1827 1059 -1823
rect 1072 -1827 1076 -1823
rect 1089 -1827 1093 -1823
rect 1097 -1827 1101 -1823
rect 1114 -1827 1118 -1823
rect 1131 -1827 1135 -1823
rect 1139 -1827 1143 -1823
rect 1155 -1827 1159 -1823
rect 1203 -1827 1207 -1823
rect 1211 -1827 1215 -1823
rect 1321 -1827 1325 -1823
rect 1330 -1827 1334 -1823
rect 1339 -1827 1343 -1823
rect 1347 -1827 1351 -1823
rect 1363 -1827 1367 -1823
rect 1371 -1827 1375 -1823
rect 1388 -1827 1392 -1823
rect 1405 -1827 1409 -1823
rect 1413 -1827 1417 -1823
rect 1430 -1827 1434 -1823
rect 1447 -1827 1451 -1823
rect 1455 -1827 1459 -1823
rect 1472 -1827 1476 -1823
rect 1489 -1827 1493 -1823
rect 1497 -1827 1501 -1823
rect 1513 -1827 1517 -1823
rect -1260 -1942 -1256 -1938
rect -1251 -1942 -1247 -1938
rect -1242 -1942 -1238 -1938
rect -1234 -1942 -1230 -1938
rect -1218 -1942 -1214 -1938
rect -1210 -1942 -1206 -1938
rect -1193 -1942 -1189 -1938
rect -1176 -1942 -1172 -1938
rect -1168 -1942 -1164 -1938
rect -1151 -1942 -1147 -1938
rect -1134 -1942 -1130 -1938
rect -1126 -1942 -1122 -1938
rect -1109 -1942 -1105 -1938
rect -1092 -1942 -1088 -1938
rect -1084 -1942 -1080 -1938
rect -1068 -1942 -1064 -1938
rect -1029 -1942 -1025 -1938
rect -1021 -1942 -1017 -1938
rect -673 -1942 -669 -1934
rect -665 -1942 -661 -1934
rect -332 -1942 -328 -1938
rect -324 -1942 -320 -1938
rect 464 -1942 468 -1938
rect 472 -1942 476 -1938
rect 841 -1942 845 -1934
rect 849 -1942 853 -1934
rect 1203 -1942 1207 -1938
rect 1211 -1942 1215 -1938
rect -1339 -2054 -1335 -2050
rect -1322 -2054 -1318 -2050
rect -1313 -2054 -1309 -2050
rect -935 -2054 -931 -2050
rect -918 -2054 -914 -2050
rect -909 -2054 -905 -2050
rect -577 -2054 -573 -2050
rect -560 -2054 -556 -2050
rect -551 -2054 -547 -2050
rect -219 -2054 -215 -2050
rect -202 -2054 -198 -2050
rect -193 -2054 -189 -2050
rect 209 -2054 213 -2050
rect 226 -2054 230 -2050
rect 235 -2054 239 -2050
rect 565 -2054 569 -2050
rect 582 -2054 586 -2050
rect 591 -2054 595 -2050
rect 963 -2054 967 -2050
rect 980 -2054 984 -2050
rect 989 -2054 993 -2050
rect 1321 -2054 1325 -2050
rect 1338 -2054 1342 -2050
rect 1347 -2054 1351 -2050
rect -1260 -2173 -1256 -2169
rect -1251 -2173 -1247 -2169
rect -1242 -2173 -1238 -2169
rect -1234 -2173 -1230 -2169
rect -1225 -2173 -1221 -2169
rect -1207 -2173 -1203 -2169
rect -1198 -2173 -1194 -2169
rect -1190 -2173 -1186 -2169
rect -1173 -2173 -1169 -2169
rect -1164 -2173 -1160 -2169
rect -935 -2173 -931 -2169
rect -926 -2173 -922 -2169
rect -917 -2173 -913 -2169
rect -909 -2173 -905 -2169
rect -900 -2173 -896 -2169
rect -891 -2173 -887 -2169
rect -883 -2173 -879 -2169
rect -875 -2173 -871 -2169
rect -857 -2173 -853 -2169
rect -847 -2173 -843 -2169
rect -839 -2173 -835 -2169
rect -822 -2173 -818 -2169
rect -813 -2173 -809 -2169
rect -805 -2173 -801 -2169
rect -796 -2173 -792 -2169
rect -778 -2173 -774 -2169
rect -769 -2173 -765 -2169
rect -761 -2173 -757 -2169
rect -745 -2173 -741 -2169
rect -737 -2173 -733 -2169
rect -725 -2173 -721 -2169
rect -713 -2173 -709 -2169
rect -704 -2173 -700 -2169
rect -695 -2173 -691 -2169
rect -577 -2173 -573 -2169
rect -568 -2173 -564 -2169
rect -559 -2173 -555 -2169
rect -551 -2173 -547 -2169
rect -542 -2173 -538 -2169
rect -533 -2173 -529 -2169
rect -525 -2173 -521 -2169
rect -517 -2173 -513 -2169
rect -499 -2173 -495 -2169
rect -489 -2173 -485 -2169
rect -481 -2173 -477 -2169
rect -464 -2173 -460 -2169
rect -455 -2173 -451 -2169
rect -447 -2173 -443 -2169
rect -438 -2173 -434 -2169
rect -420 -2173 -416 -2169
rect -411 -2173 -407 -2169
rect -403 -2173 -399 -2169
rect -387 -2173 -383 -2169
rect -379 -2173 -375 -2169
rect -367 -2173 -363 -2169
rect -355 -2173 -351 -2169
rect -346 -2173 -342 -2169
rect -337 -2173 -333 -2169
rect -219 -2173 -215 -2169
rect -210 -2173 -206 -2169
rect -201 -2173 -197 -2169
rect -193 -2173 -189 -2169
rect -184 -2173 -180 -2169
rect -175 -2173 -171 -2169
rect -167 -2173 -163 -2169
rect -159 -2173 -155 -2169
rect -141 -2173 -137 -2169
rect -131 -2173 -127 -2169
rect -123 -2173 -119 -2169
rect -106 -2173 -102 -2169
rect -97 -2173 -93 -2169
rect -89 -2173 -85 -2169
rect -80 -2173 -76 -2169
rect -62 -2173 -58 -2169
rect -53 -2173 -49 -2169
rect -45 -2173 -41 -2169
rect -29 -2173 -25 -2169
rect -21 -2173 -17 -2169
rect -9 -2173 -5 -2169
rect 3 -2173 7 -2169
rect 12 -2173 16 -2169
rect 21 -2173 25 -2169
rect 209 -2173 213 -2169
rect 218 -2173 222 -2169
rect 227 -2173 231 -2169
rect 235 -2173 239 -2169
rect 244 -2173 248 -2169
rect 253 -2173 257 -2169
rect 261 -2173 265 -2169
rect 269 -2173 273 -2169
rect 287 -2173 291 -2169
rect 297 -2173 301 -2169
rect 305 -2173 309 -2169
rect 322 -2173 326 -2169
rect 331 -2173 335 -2169
rect 339 -2173 343 -2169
rect 348 -2173 352 -2169
rect 366 -2173 370 -2169
rect 375 -2173 379 -2169
rect 383 -2173 387 -2169
rect 399 -2173 403 -2169
rect 407 -2173 411 -2169
rect 419 -2173 423 -2169
rect 431 -2173 435 -2169
rect 440 -2173 444 -2169
rect 449 -2173 453 -2169
rect 565 -2173 569 -2169
rect 574 -2173 578 -2169
rect 583 -2173 587 -2169
rect 591 -2173 595 -2169
rect 600 -2173 604 -2169
rect 609 -2173 613 -2169
rect 617 -2173 621 -2169
rect 625 -2173 629 -2169
rect 643 -2173 647 -2169
rect 653 -2173 657 -2169
rect 661 -2173 665 -2169
rect 678 -2173 682 -2169
rect 687 -2173 691 -2169
rect 695 -2173 699 -2169
rect 704 -2173 708 -2169
rect 722 -2173 726 -2169
rect 731 -2173 735 -2169
rect 739 -2173 743 -2169
rect 755 -2173 759 -2169
rect 763 -2173 767 -2169
rect 775 -2173 779 -2169
rect 787 -2173 791 -2169
rect 796 -2173 800 -2169
rect 805 -2173 809 -2169
rect 963 -2173 967 -2169
rect 972 -2173 976 -2169
rect 981 -2173 985 -2169
rect 989 -2173 993 -2169
rect 998 -2173 1002 -2169
rect 1007 -2173 1011 -2169
rect 1015 -2173 1019 -2169
rect 1023 -2173 1027 -2169
rect 1041 -2173 1045 -2169
rect 1051 -2173 1055 -2169
rect 1059 -2173 1063 -2169
rect 1076 -2173 1080 -2169
rect 1085 -2173 1089 -2169
rect 1093 -2173 1097 -2169
rect 1102 -2173 1106 -2169
rect 1120 -2173 1124 -2169
rect 1129 -2173 1133 -2169
rect 1137 -2173 1141 -2169
rect 1153 -2173 1157 -2169
rect 1161 -2173 1165 -2169
rect 1173 -2173 1177 -2169
rect 1185 -2173 1189 -2169
rect 1194 -2173 1198 -2169
rect 1203 -2173 1207 -2169
rect 1321 -2173 1325 -2169
rect 1330 -2173 1334 -2169
rect 1339 -2173 1343 -2169
rect 1347 -2173 1351 -2169
rect 1356 -2173 1360 -2169
rect 1365 -2173 1369 -2169
rect 1373 -2173 1377 -2169
rect 1381 -2173 1385 -2169
rect 1399 -2173 1403 -2169
rect 1409 -2173 1413 -2169
rect 1417 -2173 1421 -2169
rect 1434 -2173 1438 -2169
rect 1443 -2173 1447 -2169
rect 1451 -2173 1455 -2169
rect 1460 -2173 1464 -2169
rect 1478 -2173 1482 -2169
rect 1487 -2173 1491 -2169
rect 1495 -2173 1499 -2169
rect 1511 -2173 1515 -2169
rect 1519 -2173 1523 -2169
rect 1531 -2173 1535 -2169
rect 1543 -2173 1547 -2169
rect 1552 -2173 1556 -2169
rect 1561 -2173 1565 -2169
rect -1264 -2317 -1260 -2313
rect -1255 -2317 -1251 -2313
rect -1246 -2317 -1242 -2313
rect -1238 -2317 -1234 -2313
rect -1222 -2317 -1218 -2313
rect -1214 -2317 -1210 -2313
rect -1197 -2317 -1193 -2313
rect -1180 -2317 -1176 -2313
rect -1172 -2317 -1168 -2313
rect -1155 -2317 -1151 -2313
rect -1138 -2317 -1134 -2313
rect -1130 -2317 -1126 -2313
rect -1113 -2317 -1109 -2313
rect -1096 -2317 -1092 -2313
rect -1088 -2317 -1084 -2313
rect -1072 -2317 -1068 -2313
rect -935 -2317 -931 -2313
rect -926 -2317 -922 -2313
rect -917 -2317 -913 -2313
rect -909 -2317 -905 -2313
rect -893 -2317 -889 -2313
rect -885 -2317 -881 -2313
rect -868 -2317 -864 -2313
rect -851 -2317 -847 -2313
rect -843 -2317 -839 -2313
rect -826 -2317 -822 -2313
rect -809 -2317 -805 -2313
rect -801 -2317 -797 -2313
rect -784 -2317 -780 -2313
rect -767 -2317 -763 -2313
rect -759 -2317 -755 -2313
rect -743 -2317 -739 -2313
rect -577 -2317 -573 -2313
rect -568 -2317 -564 -2313
rect -559 -2317 -555 -2313
rect -551 -2317 -547 -2313
rect -535 -2317 -531 -2313
rect -527 -2317 -523 -2313
rect -510 -2317 -506 -2313
rect -493 -2317 -489 -2313
rect -485 -2317 -481 -2313
rect -468 -2317 -464 -2313
rect -451 -2317 -447 -2313
rect -443 -2317 -439 -2313
rect -426 -2317 -422 -2313
rect -409 -2317 -405 -2313
rect -401 -2317 -397 -2313
rect -385 -2317 -381 -2313
rect -219 -2317 -215 -2313
rect -210 -2317 -206 -2313
rect -201 -2317 -197 -2313
rect -193 -2317 -189 -2313
rect -177 -2317 -173 -2313
rect -169 -2317 -165 -2313
rect -152 -2317 -148 -2313
rect -135 -2317 -131 -2313
rect -127 -2317 -123 -2313
rect -110 -2317 -106 -2313
rect -93 -2317 -89 -2313
rect -85 -2317 -81 -2313
rect -68 -2317 -64 -2313
rect -51 -2317 -47 -2313
rect -43 -2317 -39 -2313
rect -27 -2317 -23 -2313
rect 209 -2317 213 -2313
rect 218 -2317 222 -2313
rect 227 -2317 231 -2313
rect 235 -2317 239 -2313
rect 251 -2317 255 -2313
rect 259 -2317 263 -2313
rect 276 -2317 280 -2313
rect 293 -2317 297 -2313
rect 301 -2317 305 -2313
rect 318 -2317 322 -2313
rect 335 -2317 339 -2313
rect 343 -2317 347 -2313
rect 360 -2317 364 -2313
rect 377 -2317 381 -2313
rect 385 -2317 389 -2313
rect 401 -2317 405 -2313
rect 565 -2317 569 -2313
rect 574 -2317 578 -2313
rect 583 -2317 587 -2313
rect 591 -2317 595 -2313
rect 607 -2317 611 -2313
rect 615 -2317 619 -2313
rect 632 -2317 636 -2313
rect 649 -2317 653 -2313
rect 657 -2317 661 -2313
rect 674 -2317 678 -2313
rect 691 -2317 695 -2313
rect 699 -2317 703 -2313
rect 716 -2317 720 -2313
rect 733 -2317 737 -2313
rect 741 -2317 745 -2313
rect 757 -2317 761 -2313
rect -1264 -2448 -1260 -2444
rect -1255 -2448 -1251 -2444
rect -1246 -2448 -1242 -2444
rect -1238 -2448 -1234 -2444
rect -1222 -2448 -1218 -2444
rect -1214 -2448 -1210 -2444
rect -1197 -2448 -1193 -2444
rect -1180 -2448 -1176 -2444
rect -1172 -2448 -1168 -2444
rect -1155 -2448 -1151 -2444
rect -1138 -2448 -1134 -2444
rect -1130 -2448 -1126 -2444
rect -1113 -2448 -1109 -2444
rect -1096 -2448 -1092 -2444
rect -1088 -2448 -1084 -2444
rect -1072 -2448 -1068 -2444
rect -935 -2448 -931 -2444
rect -926 -2448 -922 -2444
rect -917 -2448 -913 -2444
rect -909 -2448 -905 -2444
rect -893 -2448 -889 -2444
rect -885 -2448 -881 -2444
rect -868 -2448 -864 -2444
rect -851 -2448 -847 -2444
rect -843 -2448 -839 -2444
rect -826 -2448 -822 -2444
rect -809 -2448 -805 -2444
rect -801 -2448 -797 -2444
rect -784 -2448 -780 -2444
rect -767 -2448 -763 -2444
rect -759 -2448 -755 -2444
rect -743 -2448 -739 -2444
rect -577 -2448 -573 -2444
rect -568 -2448 -564 -2444
rect -559 -2448 -555 -2444
rect -551 -2448 -547 -2444
rect -535 -2448 -531 -2444
rect -527 -2448 -523 -2444
rect -510 -2448 -506 -2444
rect -493 -2448 -489 -2444
rect -485 -2448 -481 -2444
rect -468 -2448 -464 -2444
rect -451 -2448 -447 -2444
rect -443 -2448 -439 -2444
rect -426 -2448 -422 -2444
rect -409 -2448 -405 -2444
rect -401 -2448 -397 -2444
rect -385 -2448 -381 -2444
rect -219 -2448 -215 -2444
rect -210 -2448 -206 -2444
rect -201 -2448 -197 -2444
rect -193 -2448 -189 -2444
rect -177 -2448 -173 -2444
rect -169 -2448 -165 -2444
rect -152 -2448 -148 -2444
rect -135 -2448 -131 -2444
rect -127 -2448 -123 -2444
rect -110 -2448 -106 -2444
rect -93 -2448 -89 -2444
rect -85 -2448 -81 -2444
rect -68 -2448 -64 -2444
rect -51 -2448 -47 -2444
rect -43 -2448 -39 -2444
rect -27 -2448 -23 -2444
rect 209 -2448 213 -2444
rect 218 -2448 222 -2444
rect 227 -2448 231 -2444
rect 235 -2448 239 -2444
rect 251 -2448 255 -2444
rect 259 -2448 263 -2444
rect 276 -2448 280 -2444
rect 293 -2448 297 -2444
rect 301 -2448 305 -2444
rect 318 -2448 322 -2444
rect 335 -2448 339 -2444
rect 343 -2448 347 -2444
rect 360 -2448 364 -2444
rect 377 -2448 381 -2444
rect 385 -2448 389 -2444
rect 401 -2448 405 -2444
rect 565 -2448 569 -2444
rect 574 -2448 578 -2444
rect 583 -2448 587 -2444
rect 591 -2448 595 -2444
rect 607 -2448 611 -2444
rect 615 -2448 619 -2444
rect 632 -2448 636 -2444
rect 649 -2448 653 -2444
rect 657 -2448 661 -2444
rect 674 -2448 678 -2444
rect 691 -2448 695 -2444
rect 699 -2448 703 -2444
rect 716 -2448 720 -2444
rect 733 -2448 737 -2444
rect 741 -2448 745 -2444
rect 757 -2448 761 -2444
rect 963 -2448 967 -2444
rect 972 -2448 976 -2444
rect 981 -2448 985 -2444
rect 989 -2448 993 -2444
rect 1005 -2448 1009 -2444
rect 1013 -2448 1017 -2444
rect 1030 -2448 1034 -2444
rect 1047 -2448 1051 -2444
rect 1055 -2448 1059 -2444
rect 1072 -2448 1076 -2444
rect 1089 -2448 1093 -2444
rect 1097 -2448 1101 -2444
rect 1114 -2448 1118 -2444
rect 1131 -2448 1135 -2444
rect 1139 -2448 1143 -2444
rect 1155 -2448 1159 -2444
rect 1321 -2448 1325 -2444
rect 1330 -2448 1334 -2444
rect 1339 -2448 1343 -2444
rect 1347 -2448 1351 -2444
rect 1363 -2448 1367 -2444
rect 1371 -2448 1375 -2444
rect 1388 -2448 1392 -2444
rect 1405 -2448 1409 -2444
rect 1413 -2448 1417 -2444
rect 1430 -2448 1434 -2444
rect 1447 -2448 1451 -2444
rect 1455 -2448 1459 -2444
rect 1472 -2448 1476 -2444
rect 1489 -2448 1493 -2444
rect 1497 -2448 1501 -2444
rect 1513 -2448 1517 -2444
rect -1264 -2579 -1260 -2575
rect -1255 -2579 -1251 -2575
rect -1246 -2579 -1242 -2575
rect -1238 -2579 -1234 -2575
rect -1222 -2579 -1218 -2575
rect -1214 -2579 -1210 -2575
rect -1197 -2579 -1193 -2575
rect -1180 -2579 -1176 -2575
rect -1172 -2579 -1168 -2575
rect -1155 -2579 -1151 -2575
rect -1138 -2579 -1134 -2575
rect -1130 -2579 -1126 -2575
rect -1113 -2579 -1109 -2575
rect -1096 -2579 -1092 -2575
rect -1088 -2579 -1084 -2575
rect -1072 -2579 -1068 -2575
rect -935 -2579 -931 -2575
rect -926 -2579 -922 -2575
rect -917 -2579 -913 -2575
rect -909 -2579 -905 -2575
rect -893 -2579 -889 -2575
rect -885 -2579 -881 -2575
rect -868 -2579 -864 -2575
rect -851 -2579 -847 -2575
rect -843 -2579 -839 -2575
rect -826 -2579 -822 -2575
rect -809 -2579 -805 -2575
rect -801 -2579 -797 -2575
rect -784 -2579 -780 -2575
rect -767 -2579 -763 -2575
rect -759 -2579 -755 -2575
rect -743 -2579 -739 -2575
rect -577 -2579 -573 -2575
rect -568 -2579 -564 -2575
rect -559 -2579 -555 -2575
rect -551 -2579 -547 -2575
rect -535 -2579 -531 -2575
rect -527 -2579 -523 -2575
rect -510 -2579 -506 -2575
rect -493 -2579 -489 -2575
rect -485 -2579 -481 -2575
rect -468 -2579 -464 -2575
rect -451 -2579 -447 -2575
rect -443 -2579 -439 -2575
rect -426 -2579 -422 -2575
rect -409 -2579 -405 -2575
rect -401 -2579 -397 -2575
rect -385 -2579 -381 -2575
rect -219 -2579 -215 -2575
rect -210 -2579 -206 -2575
rect -201 -2579 -197 -2575
rect -193 -2579 -189 -2575
rect -177 -2579 -173 -2575
rect -169 -2579 -165 -2575
rect -152 -2579 -148 -2575
rect -135 -2579 -131 -2575
rect -127 -2579 -123 -2575
rect -110 -2579 -106 -2575
rect -93 -2579 -89 -2575
rect -85 -2579 -81 -2575
rect -68 -2579 -64 -2575
rect -51 -2579 -47 -2575
rect -43 -2579 -39 -2575
rect -27 -2579 -23 -2575
rect 90 -2579 94 -2563
rect 98 -2579 102 -2563
rect 209 -2579 213 -2575
rect 218 -2579 222 -2575
rect 227 -2579 231 -2575
rect 235 -2579 239 -2575
rect 251 -2579 255 -2575
rect 259 -2579 263 -2575
rect 276 -2579 280 -2575
rect 293 -2579 297 -2575
rect 301 -2579 305 -2575
rect 318 -2579 322 -2575
rect 335 -2579 339 -2575
rect 343 -2579 347 -2575
rect 360 -2579 364 -2575
rect 377 -2579 381 -2575
rect 385 -2579 389 -2575
rect 401 -2579 405 -2575
rect 565 -2579 569 -2575
rect 574 -2579 578 -2575
rect 583 -2579 587 -2575
rect 591 -2579 595 -2575
rect 607 -2579 611 -2575
rect 615 -2579 619 -2575
rect 632 -2579 636 -2575
rect 649 -2579 653 -2575
rect 657 -2579 661 -2575
rect 674 -2579 678 -2575
rect 691 -2579 695 -2575
rect 699 -2579 703 -2575
rect 716 -2579 720 -2575
rect 733 -2579 737 -2575
rect 741 -2579 745 -2575
rect 757 -2579 761 -2575
rect 963 -2579 967 -2575
rect 972 -2579 976 -2575
rect 981 -2579 985 -2575
rect 989 -2579 993 -2575
rect 1005 -2579 1009 -2575
rect 1013 -2579 1017 -2575
rect 1030 -2579 1034 -2575
rect 1047 -2579 1051 -2575
rect 1055 -2579 1059 -2575
rect 1072 -2579 1076 -2575
rect 1089 -2579 1093 -2575
rect 1097 -2579 1101 -2575
rect 1114 -2579 1118 -2575
rect 1131 -2579 1135 -2575
rect 1139 -2579 1143 -2575
rect 1155 -2579 1159 -2575
rect 1321 -2579 1325 -2575
rect 1330 -2579 1334 -2575
rect 1339 -2579 1343 -2575
rect 1347 -2579 1351 -2575
rect 1363 -2579 1367 -2575
rect 1371 -2579 1375 -2575
rect 1388 -2579 1392 -2575
rect 1405 -2579 1409 -2575
rect 1413 -2579 1417 -2575
rect 1430 -2579 1434 -2575
rect 1447 -2579 1451 -2575
rect 1455 -2579 1459 -2575
rect 1472 -2579 1476 -2575
rect 1489 -2579 1493 -2575
rect 1497 -2579 1501 -2575
rect 1513 -2579 1517 -2575
rect -1264 -2691 -1260 -2687
rect -1255 -2691 -1251 -2687
rect -1246 -2691 -1242 -2687
rect -1238 -2691 -1234 -2687
rect -1222 -2691 -1218 -2687
rect -1214 -2691 -1210 -2687
rect -1197 -2691 -1193 -2687
rect -1180 -2691 -1176 -2687
rect -1172 -2691 -1168 -2687
rect -1155 -2691 -1151 -2687
rect -1138 -2691 -1134 -2687
rect -1130 -2691 -1126 -2687
rect -1113 -2691 -1109 -2687
rect -1096 -2691 -1092 -2687
rect -1088 -2691 -1084 -2687
rect -1072 -2691 -1068 -2687
rect -935 -2691 -931 -2687
rect -926 -2691 -922 -2687
rect -917 -2691 -913 -2687
rect -909 -2691 -905 -2687
rect -893 -2691 -889 -2687
rect -885 -2691 -881 -2687
rect -868 -2691 -864 -2687
rect -851 -2691 -847 -2687
rect -843 -2691 -839 -2687
rect -826 -2691 -822 -2687
rect -809 -2691 -805 -2687
rect -801 -2691 -797 -2687
rect -784 -2691 -780 -2687
rect -767 -2691 -763 -2687
rect -759 -2691 -755 -2687
rect -743 -2691 -739 -2687
rect -1339 -2804 -1335 -2800
rect -1322 -2804 -1318 -2800
rect -1313 -2804 -1309 -2800
rect -935 -2804 -931 -2800
rect -918 -2804 -914 -2800
rect -909 -2804 -905 -2800
rect -577 -2804 -573 -2800
rect -560 -2804 -556 -2800
rect -551 -2804 -547 -2800
rect -219 -2804 -215 -2800
rect -202 -2804 -198 -2800
rect -193 -2804 -189 -2800
rect 209 -2804 213 -2800
rect 226 -2804 230 -2800
rect 235 -2804 239 -2800
rect 565 -2804 569 -2800
rect 582 -2804 586 -2800
rect 591 -2804 595 -2800
rect 963 -2804 967 -2800
rect 980 -2804 984 -2800
rect 989 -2804 993 -2800
rect 1321 -2804 1325 -2800
rect 1338 -2804 1342 -2800
rect 1347 -2804 1351 -2800
rect -1264 -2923 -1260 -2919
rect -1255 -2923 -1251 -2919
rect -1246 -2923 -1242 -2919
rect -1238 -2923 -1234 -2919
rect -1229 -2923 -1225 -2919
rect -1211 -2923 -1207 -2919
rect -1202 -2923 -1198 -2919
rect -1194 -2923 -1190 -2919
rect -1177 -2923 -1173 -2919
rect -1168 -2923 -1164 -2919
rect -935 -2923 -931 -2919
rect -926 -2923 -922 -2919
rect -917 -2923 -913 -2919
rect -909 -2923 -905 -2919
rect -900 -2923 -896 -2919
rect -891 -2923 -887 -2919
rect -883 -2923 -879 -2919
rect -875 -2923 -871 -2919
rect -857 -2923 -853 -2919
rect -847 -2923 -843 -2919
rect -839 -2923 -835 -2919
rect -822 -2923 -818 -2919
rect -813 -2923 -809 -2919
rect -805 -2923 -801 -2919
rect -796 -2923 -792 -2919
rect -778 -2923 -774 -2919
rect -769 -2923 -765 -2919
rect -761 -2923 -757 -2919
rect -745 -2923 -741 -2919
rect -737 -2923 -733 -2919
rect -725 -2923 -721 -2919
rect -713 -2923 -709 -2919
rect -704 -2923 -700 -2919
rect -695 -2923 -691 -2919
rect -577 -2923 -573 -2919
rect -568 -2923 -564 -2919
rect -559 -2923 -555 -2919
rect -551 -2923 -547 -2919
rect -542 -2923 -538 -2919
rect -533 -2923 -529 -2919
rect -525 -2923 -521 -2919
rect -517 -2923 -513 -2919
rect -499 -2923 -495 -2919
rect -489 -2923 -485 -2919
rect -481 -2923 -477 -2919
rect -464 -2923 -460 -2919
rect -455 -2923 -451 -2919
rect -447 -2923 -443 -2919
rect -438 -2923 -434 -2919
rect -420 -2923 -416 -2919
rect -411 -2923 -407 -2919
rect -403 -2923 -399 -2919
rect -387 -2923 -383 -2919
rect -379 -2923 -375 -2919
rect -367 -2923 -363 -2919
rect -355 -2923 -351 -2919
rect -346 -2923 -342 -2919
rect -337 -2923 -333 -2919
rect -219 -2923 -215 -2919
rect -210 -2923 -206 -2919
rect -201 -2923 -197 -2919
rect -193 -2923 -189 -2919
rect -184 -2923 -180 -2919
rect -175 -2923 -171 -2919
rect -167 -2923 -163 -2919
rect -159 -2923 -155 -2919
rect -141 -2923 -137 -2919
rect -131 -2923 -127 -2919
rect -123 -2923 -119 -2919
rect -106 -2923 -102 -2919
rect -97 -2923 -93 -2919
rect -89 -2923 -85 -2919
rect -80 -2923 -76 -2919
rect -62 -2923 -58 -2919
rect -53 -2923 -49 -2919
rect -45 -2923 -41 -2919
rect -29 -2923 -25 -2919
rect -21 -2923 -17 -2919
rect -9 -2923 -5 -2919
rect 3 -2923 7 -2919
rect 12 -2923 16 -2919
rect 21 -2923 25 -2919
rect 209 -2923 213 -2919
rect 218 -2923 222 -2919
rect 227 -2923 231 -2919
rect 235 -2923 239 -2919
rect 244 -2923 248 -2919
rect 253 -2923 257 -2919
rect 261 -2923 265 -2919
rect 269 -2923 273 -2919
rect 287 -2923 291 -2919
rect 297 -2923 301 -2919
rect 305 -2923 309 -2919
rect 322 -2923 326 -2919
rect 331 -2923 335 -2919
rect 339 -2923 343 -2919
rect 348 -2923 352 -2919
rect 366 -2923 370 -2919
rect 375 -2923 379 -2919
rect 383 -2923 387 -2919
rect 399 -2923 403 -2919
rect 407 -2923 411 -2919
rect 419 -2923 423 -2919
rect 431 -2923 435 -2919
rect 440 -2923 444 -2919
rect 449 -2923 453 -2919
rect 565 -2923 569 -2919
rect 574 -2923 578 -2919
rect 583 -2923 587 -2919
rect 591 -2923 595 -2919
rect 600 -2923 604 -2919
rect 609 -2923 613 -2919
rect 617 -2923 621 -2919
rect 625 -2923 629 -2919
rect 643 -2923 647 -2919
rect 653 -2923 657 -2919
rect 661 -2923 665 -2919
rect 678 -2923 682 -2919
rect 687 -2923 691 -2919
rect 695 -2923 699 -2919
rect 704 -2923 708 -2919
rect 722 -2923 726 -2919
rect 731 -2923 735 -2919
rect 739 -2923 743 -2919
rect 755 -2923 759 -2919
rect 763 -2923 767 -2919
rect 775 -2923 779 -2919
rect 787 -2923 791 -2919
rect 796 -2923 800 -2919
rect 805 -2923 809 -2919
rect 963 -2923 967 -2919
rect 972 -2923 976 -2919
rect 981 -2923 985 -2919
rect 989 -2923 993 -2919
rect 998 -2923 1002 -2919
rect 1007 -2923 1011 -2919
rect 1015 -2923 1019 -2919
rect 1023 -2923 1027 -2919
rect 1041 -2923 1045 -2919
rect 1051 -2923 1055 -2919
rect 1059 -2923 1063 -2919
rect 1076 -2923 1080 -2919
rect 1085 -2923 1089 -2919
rect 1093 -2923 1097 -2919
rect 1102 -2923 1106 -2919
rect 1120 -2923 1124 -2919
rect 1129 -2923 1133 -2919
rect 1137 -2923 1141 -2919
rect 1153 -2923 1157 -2919
rect 1161 -2923 1165 -2919
rect 1173 -2923 1177 -2919
rect 1185 -2923 1189 -2919
rect 1194 -2923 1198 -2919
rect 1203 -2923 1207 -2919
rect 1321 -2923 1325 -2919
rect 1330 -2923 1334 -2919
rect 1339 -2923 1343 -2919
rect 1347 -2923 1351 -2919
rect 1356 -2923 1360 -2919
rect 1365 -2923 1369 -2919
rect 1373 -2923 1377 -2919
rect 1381 -2923 1385 -2919
rect 1399 -2923 1403 -2919
rect 1409 -2923 1413 -2919
rect 1417 -2923 1421 -2919
rect 1434 -2923 1438 -2919
rect 1443 -2923 1447 -2919
rect 1451 -2923 1455 -2919
rect 1460 -2923 1464 -2919
rect 1478 -2923 1482 -2919
rect 1487 -2923 1491 -2919
rect 1495 -2923 1499 -2919
rect 1511 -2923 1515 -2919
rect 1519 -2923 1523 -2919
rect 1531 -2923 1535 -2919
rect 1543 -2923 1547 -2919
rect 1552 -2923 1556 -2919
rect 1561 -2923 1565 -2919
rect -1264 -3042 -1260 -3038
rect -1255 -3042 -1251 -3038
rect -1246 -3042 -1242 -3038
rect -1238 -3042 -1234 -3038
rect -1222 -3042 -1218 -3038
rect -1214 -3042 -1210 -3038
rect -1197 -3042 -1193 -3038
rect -1180 -3042 -1176 -3038
rect -1172 -3042 -1168 -3038
rect -1155 -3042 -1151 -3038
rect -1138 -3042 -1134 -3038
rect -1130 -3042 -1126 -3038
rect -1113 -3042 -1109 -3038
rect -1096 -3042 -1092 -3038
rect -1088 -3042 -1084 -3038
rect -1072 -3042 -1068 -3038
rect -1026 -3042 -1022 -3038
rect -1018 -3042 -1014 -3038
rect -935 -3042 -931 -3038
rect -926 -3042 -922 -3038
rect -917 -3042 -913 -3038
rect -909 -3042 -905 -3038
rect -893 -3042 -889 -3038
rect -885 -3042 -881 -3038
rect -868 -3042 -864 -3038
rect -851 -3042 -847 -3038
rect -843 -3042 -839 -3038
rect -826 -3042 -822 -3038
rect -809 -3042 -805 -3038
rect -801 -3042 -797 -3038
rect -784 -3042 -780 -3038
rect -767 -3042 -763 -3038
rect -759 -3042 -755 -3038
rect -743 -3042 -739 -3038
rect -672 -3042 -668 -3034
rect -664 -3042 -660 -3034
rect -577 -3042 -573 -3038
rect -568 -3042 -564 -3038
rect -559 -3042 -555 -3038
rect -551 -3042 -547 -3038
rect -535 -3042 -531 -3038
rect -527 -3042 -523 -3038
rect -510 -3042 -506 -3038
rect -493 -3042 -489 -3038
rect -485 -3042 -481 -3038
rect -468 -3042 -464 -3038
rect -451 -3042 -447 -3038
rect -443 -3042 -439 -3038
rect -426 -3042 -422 -3038
rect -409 -3042 -405 -3038
rect -401 -3042 -397 -3038
rect -385 -3042 -381 -3038
rect -329 -3042 -325 -3038
rect -321 -3042 -317 -3038
rect -219 -3042 -215 -3038
rect -210 -3042 -206 -3038
rect -201 -3042 -197 -3038
rect -193 -3042 -189 -3038
rect -177 -3042 -173 -3038
rect -169 -3042 -165 -3038
rect -152 -3042 -148 -3038
rect -135 -3042 -131 -3038
rect -127 -3042 -123 -3038
rect -110 -3042 -106 -3038
rect -93 -3042 -89 -3038
rect -85 -3042 -81 -3038
rect -68 -3042 -64 -3038
rect -51 -3042 -47 -3038
rect -43 -3042 -39 -3038
rect -27 -3042 -23 -3038
rect 209 -3042 213 -3038
rect 218 -3042 222 -3038
rect 227 -3042 231 -3038
rect 235 -3042 239 -3038
rect 251 -3042 255 -3038
rect 259 -3042 263 -3038
rect 276 -3042 280 -3038
rect 293 -3042 297 -3038
rect 301 -3042 305 -3038
rect 318 -3042 322 -3038
rect 335 -3042 339 -3038
rect 343 -3042 347 -3038
rect 360 -3042 364 -3038
rect 377 -3042 381 -3038
rect 385 -3042 389 -3038
rect 401 -3042 405 -3038
rect 472 -3042 476 -3038
rect 480 -3042 484 -3038
rect 841 -3042 845 -3034
rect 849 -3042 853 -3034
rect 1199 -3042 1203 -3038
rect 1207 -3042 1211 -3038
rect -1264 -3158 -1260 -3154
rect -1255 -3158 -1251 -3154
rect -1246 -3158 -1242 -3154
rect -1238 -3158 -1234 -3154
rect -1222 -3158 -1218 -3154
rect -1214 -3158 -1210 -3154
rect -1197 -3158 -1193 -3154
rect -1180 -3158 -1176 -3154
rect -1172 -3158 -1168 -3154
rect -1155 -3158 -1151 -3154
rect -1138 -3158 -1134 -3154
rect -1130 -3158 -1126 -3154
rect -1113 -3158 -1109 -3154
rect -1096 -3158 -1092 -3154
rect -1088 -3158 -1084 -3154
rect -1072 -3158 -1068 -3154
rect -1026 -3158 -1022 -3154
rect -1018 -3158 -1014 -3154
rect -935 -3158 -931 -3154
rect -926 -3158 -922 -3154
rect -917 -3158 -913 -3154
rect -909 -3158 -905 -3154
rect -893 -3158 -889 -3154
rect -885 -3158 -881 -3154
rect -868 -3158 -864 -3154
rect -851 -3158 -847 -3154
rect -843 -3158 -839 -3154
rect -826 -3158 -822 -3154
rect -809 -3158 -805 -3154
rect -801 -3158 -797 -3154
rect -784 -3158 -780 -3154
rect -767 -3158 -763 -3154
rect -759 -3158 -755 -3154
rect -743 -3158 -739 -3154
rect -577 -3158 -573 -3154
rect -568 -3158 -564 -3154
rect -559 -3158 -555 -3154
rect -551 -3158 -547 -3154
rect -535 -3158 -531 -3154
rect -527 -3158 -523 -3154
rect -510 -3158 -506 -3154
rect -493 -3158 -489 -3154
rect -485 -3158 -481 -3154
rect -468 -3158 -464 -3154
rect -451 -3158 -447 -3154
rect -443 -3158 -439 -3154
rect -426 -3158 -422 -3154
rect -409 -3158 -405 -3154
rect -401 -3158 -397 -3154
rect -385 -3158 -381 -3154
rect -329 -3158 -325 -3154
rect -321 -3158 -317 -3154
rect -219 -3158 -215 -3154
rect -210 -3158 -206 -3154
rect -201 -3158 -197 -3154
rect -193 -3158 -189 -3154
rect -177 -3158 -173 -3154
rect -169 -3158 -165 -3154
rect -152 -3158 -148 -3154
rect -135 -3158 -131 -3154
rect -127 -3158 -123 -3154
rect -110 -3158 -106 -3154
rect -93 -3158 -89 -3154
rect -85 -3158 -81 -3154
rect -68 -3158 -64 -3154
rect -51 -3158 -47 -3154
rect -43 -3158 -39 -3154
rect -27 -3158 -23 -3154
rect 209 -3158 213 -3154
rect 218 -3158 222 -3154
rect 227 -3158 231 -3154
rect 235 -3158 239 -3154
rect 251 -3158 255 -3154
rect 259 -3158 263 -3154
rect 276 -3158 280 -3154
rect 293 -3158 297 -3154
rect 301 -3158 305 -3154
rect 318 -3158 322 -3154
rect 335 -3158 339 -3154
rect 343 -3158 347 -3154
rect 360 -3158 364 -3154
rect 377 -3158 381 -3154
rect 385 -3158 389 -3154
rect 401 -3158 405 -3154
rect 472 -3158 476 -3154
rect 480 -3158 484 -3154
rect 565 -3158 569 -3154
rect 574 -3158 578 -3154
rect 583 -3158 587 -3154
rect 591 -3158 595 -3154
rect 607 -3158 611 -3154
rect 615 -3158 619 -3154
rect 632 -3158 636 -3154
rect 649 -3158 653 -3154
rect 657 -3158 661 -3154
rect 674 -3158 678 -3154
rect 691 -3158 695 -3154
rect 699 -3158 703 -3154
rect 716 -3158 720 -3154
rect 733 -3158 737 -3154
rect 741 -3158 745 -3154
rect 757 -3158 761 -3154
rect 963 -3158 967 -3154
rect 972 -3158 976 -3154
rect 981 -3158 985 -3154
rect 989 -3158 993 -3154
rect 1005 -3158 1009 -3154
rect 1013 -3158 1017 -3154
rect 1030 -3158 1034 -3154
rect 1047 -3158 1051 -3154
rect 1055 -3158 1059 -3154
rect 1072 -3158 1076 -3154
rect 1089 -3158 1093 -3154
rect 1097 -3158 1101 -3154
rect 1114 -3158 1118 -3154
rect 1131 -3158 1135 -3154
rect 1139 -3158 1143 -3154
rect 1155 -3158 1159 -3154
rect 1199 -3158 1203 -3154
rect 1207 -3158 1211 -3154
rect 1321 -3158 1325 -3154
rect 1330 -3158 1334 -3154
rect 1339 -3158 1343 -3154
rect 1347 -3158 1351 -3154
rect 1363 -3158 1367 -3154
rect 1371 -3158 1375 -3154
rect 1388 -3158 1392 -3154
rect 1405 -3158 1409 -3154
rect 1413 -3158 1417 -3154
rect 1430 -3158 1434 -3154
rect 1447 -3158 1451 -3154
rect 1455 -3158 1459 -3154
rect 1472 -3158 1476 -3154
rect 1489 -3158 1493 -3154
rect 1497 -3158 1501 -3154
rect 1513 -3158 1517 -3154
rect -1264 -3279 -1260 -3275
rect -1255 -3279 -1251 -3275
rect -1246 -3279 -1242 -3275
rect -1238 -3279 -1234 -3275
rect -1222 -3279 -1218 -3275
rect -1214 -3279 -1210 -3275
rect -1197 -3279 -1193 -3275
rect -1180 -3279 -1176 -3275
rect -1172 -3279 -1168 -3275
rect -1155 -3279 -1151 -3275
rect -1138 -3279 -1134 -3275
rect -1130 -3279 -1126 -3275
rect -1113 -3279 -1109 -3275
rect -1096 -3279 -1092 -3275
rect -1088 -3279 -1084 -3275
rect -1072 -3279 -1068 -3275
rect -935 -3279 -931 -3275
rect -926 -3279 -922 -3275
rect -917 -3279 -913 -3275
rect -909 -3279 -905 -3275
rect -893 -3279 -889 -3275
rect -885 -3279 -881 -3275
rect -868 -3279 -864 -3275
rect -851 -3279 -847 -3275
rect -843 -3279 -839 -3275
rect -826 -3279 -822 -3275
rect -809 -3279 -805 -3275
rect -801 -3279 -797 -3275
rect -784 -3279 -780 -3275
rect -767 -3279 -763 -3275
rect -759 -3279 -755 -3275
rect -743 -3279 -739 -3275
rect -577 -3279 -573 -3275
rect -568 -3279 -564 -3275
rect -559 -3279 -555 -3275
rect -551 -3279 -547 -3275
rect -535 -3279 -531 -3275
rect -527 -3279 -523 -3275
rect -510 -3279 -506 -3275
rect -493 -3279 -489 -3275
rect -485 -3279 -481 -3275
rect -468 -3279 -464 -3275
rect -451 -3279 -447 -3275
rect -443 -3279 -439 -3275
rect -426 -3279 -422 -3275
rect -409 -3279 -405 -3275
rect -401 -3279 -397 -3275
rect -385 -3279 -381 -3275
rect -219 -3279 -215 -3275
rect -210 -3279 -206 -3275
rect -201 -3279 -197 -3275
rect -193 -3279 -189 -3275
rect -177 -3279 -173 -3275
rect -169 -3279 -165 -3275
rect -152 -3279 -148 -3275
rect -135 -3279 -131 -3275
rect -127 -3279 -123 -3275
rect -110 -3279 -106 -3275
rect -93 -3279 -89 -3275
rect -85 -3279 -81 -3275
rect -68 -3279 -64 -3275
rect -51 -3279 -47 -3275
rect -43 -3279 -39 -3275
rect -27 -3279 -23 -3275
rect 209 -3279 213 -3275
rect 218 -3279 222 -3275
rect 227 -3279 231 -3275
rect 235 -3279 239 -3275
rect 251 -3279 255 -3275
rect 259 -3279 263 -3275
rect 276 -3279 280 -3275
rect 293 -3279 297 -3275
rect 301 -3279 305 -3275
rect 318 -3279 322 -3275
rect 335 -3279 339 -3275
rect 343 -3279 347 -3275
rect 360 -3279 364 -3275
rect 377 -3279 381 -3275
rect 385 -3279 389 -3275
rect 401 -3279 405 -3275
rect 565 -3279 569 -3275
rect 574 -3279 578 -3275
rect 583 -3279 587 -3275
rect 591 -3279 595 -3275
rect 607 -3279 611 -3275
rect 615 -3279 619 -3275
rect 632 -3279 636 -3275
rect 649 -3279 653 -3275
rect 657 -3279 661 -3275
rect 674 -3279 678 -3275
rect 691 -3279 695 -3275
rect 699 -3279 703 -3275
rect 716 -3279 720 -3275
rect 733 -3279 737 -3275
rect 741 -3279 745 -3275
rect 757 -3279 761 -3275
rect 963 -3279 967 -3275
rect 972 -3279 976 -3275
rect 981 -3279 985 -3275
rect 989 -3279 993 -3275
rect 1005 -3279 1009 -3275
rect 1013 -3279 1017 -3275
rect 1030 -3279 1034 -3275
rect 1047 -3279 1051 -3275
rect 1055 -3279 1059 -3275
rect 1072 -3279 1076 -3275
rect 1089 -3279 1093 -3275
rect 1097 -3279 1101 -3275
rect 1114 -3279 1118 -3275
rect 1131 -3279 1135 -3275
rect 1139 -3279 1143 -3275
rect 1155 -3279 1159 -3275
rect 1321 -3279 1325 -3275
rect 1330 -3279 1334 -3275
rect 1339 -3279 1343 -3275
rect 1347 -3279 1351 -3275
rect 1363 -3279 1367 -3275
rect 1371 -3279 1375 -3275
rect 1388 -3279 1392 -3275
rect 1405 -3279 1409 -3275
rect 1413 -3279 1417 -3275
rect 1430 -3279 1434 -3275
rect 1447 -3279 1451 -3275
rect 1455 -3279 1459 -3275
rect 1472 -3279 1476 -3275
rect 1489 -3279 1493 -3275
rect 1497 -3279 1501 -3275
rect 1513 -3279 1517 -3275
rect -1264 -3393 -1260 -3389
rect -1255 -3393 -1251 -3389
rect -1246 -3393 -1242 -3389
rect -1238 -3393 -1234 -3389
rect -1222 -3393 -1218 -3389
rect -1214 -3393 -1210 -3389
rect -1197 -3393 -1193 -3389
rect -1180 -3393 -1176 -3389
rect -1172 -3393 -1168 -3389
rect -1155 -3393 -1151 -3389
rect -1138 -3393 -1134 -3389
rect -1130 -3393 -1126 -3389
rect -1113 -3393 -1109 -3389
rect -1096 -3393 -1092 -3389
rect -1088 -3393 -1084 -3389
rect -1072 -3393 -1068 -3389
rect -935 -3393 -931 -3389
rect -926 -3393 -922 -3389
rect -917 -3393 -913 -3389
rect -909 -3393 -905 -3389
rect -893 -3393 -889 -3389
rect -885 -3393 -881 -3389
rect -868 -3393 -864 -3389
rect -851 -3393 -847 -3389
rect -843 -3393 -839 -3389
rect -826 -3393 -822 -3389
rect -809 -3393 -805 -3389
rect -801 -3393 -797 -3389
rect -784 -3393 -780 -3389
rect -767 -3393 -763 -3389
rect -759 -3393 -755 -3389
rect -743 -3393 -739 -3389
rect -577 -3393 -573 -3389
rect -568 -3393 -564 -3389
rect -559 -3393 -555 -3389
rect -551 -3393 -547 -3389
rect -535 -3393 -531 -3389
rect -527 -3393 -523 -3389
rect -510 -3393 -506 -3389
rect -493 -3393 -489 -3389
rect -485 -3393 -481 -3389
rect -468 -3393 -464 -3389
rect -451 -3393 -447 -3389
rect -443 -3393 -439 -3389
rect -426 -3393 -422 -3389
rect -409 -3393 -405 -3389
rect -401 -3393 -397 -3389
rect -385 -3393 -381 -3389
rect -1339 -3510 -1335 -3506
rect -1322 -3510 -1318 -3506
rect -1313 -3510 -1309 -3506
rect -935 -3510 -931 -3506
rect -918 -3510 -914 -3506
rect -909 -3510 -905 -3506
rect -577 -3510 -573 -3506
rect -560 -3510 -556 -3506
rect -551 -3510 -547 -3506
rect -219 -3510 -215 -3506
rect -202 -3510 -198 -3506
rect -193 -3510 -189 -3506
rect 209 -3510 213 -3506
rect 226 -3510 230 -3506
rect 235 -3510 239 -3506
rect 565 -3510 569 -3506
rect 582 -3510 586 -3506
rect 591 -3510 595 -3506
rect 963 -3510 967 -3506
rect 980 -3510 984 -3506
rect 989 -3510 993 -3506
rect 1321 -3510 1325 -3506
rect 1338 -3510 1342 -3506
rect 1347 -3510 1351 -3506
rect -1264 -3634 -1260 -3630
rect -1255 -3634 -1251 -3630
rect -1246 -3634 -1242 -3630
rect -1238 -3634 -1234 -3630
rect -1229 -3634 -1225 -3630
rect -1211 -3634 -1207 -3630
rect -1202 -3634 -1198 -3630
rect -1194 -3634 -1190 -3630
rect -1177 -3634 -1173 -3630
rect -1168 -3634 -1164 -3630
rect -935 -3634 -931 -3630
rect -926 -3634 -922 -3630
rect -917 -3634 -913 -3630
rect -909 -3634 -905 -3630
rect -900 -3634 -896 -3630
rect -891 -3634 -887 -3630
rect -883 -3634 -879 -3630
rect -875 -3634 -871 -3630
rect -857 -3634 -853 -3630
rect -847 -3634 -843 -3630
rect -839 -3634 -835 -3630
rect -822 -3634 -818 -3630
rect -813 -3634 -809 -3630
rect -805 -3634 -801 -3630
rect -796 -3634 -792 -3630
rect -778 -3634 -774 -3630
rect -769 -3634 -765 -3630
rect -761 -3634 -757 -3630
rect -745 -3634 -741 -3630
rect -737 -3634 -733 -3630
rect -725 -3634 -721 -3630
rect -713 -3634 -709 -3630
rect -704 -3634 -700 -3630
rect -695 -3634 -691 -3630
rect -577 -3634 -573 -3630
rect -568 -3634 -564 -3630
rect -559 -3634 -555 -3630
rect -551 -3634 -547 -3630
rect -542 -3634 -538 -3630
rect -533 -3634 -529 -3630
rect -525 -3634 -521 -3630
rect -517 -3634 -513 -3630
rect -499 -3634 -495 -3630
rect -489 -3634 -485 -3630
rect -481 -3634 -477 -3630
rect -464 -3634 -460 -3630
rect -455 -3634 -451 -3630
rect -447 -3634 -443 -3630
rect -438 -3634 -434 -3630
rect -420 -3634 -416 -3630
rect -411 -3634 -407 -3630
rect -403 -3634 -399 -3630
rect -387 -3634 -383 -3630
rect -379 -3634 -375 -3630
rect -367 -3634 -363 -3630
rect -355 -3634 -351 -3630
rect -346 -3634 -342 -3630
rect -337 -3634 -333 -3630
rect -219 -3634 -215 -3630
rect -210 -3634 -206 -3630
rect -201 -3634 -197 -3630
rect -193 -3634 -189 -3630
rect -184 -3634 -180 -3630
rect -175 -3634 -171 -3630
rect -167 -3634 -163 -3630
rect -159 -3634 -155 -3630
rect -141 -3634 -137 -3630
rect -131 -3634 -127 -3630
rect -123 -3634 -119 -3630
rect -106 -3634 -102 -3630
rect -97 -3634 -93 -3630
rect -89 -3634 -85 -3630
rect -80 -3634 -76 -3630
rect -62 -3634 -58 -3630
rect -53 -3634 -49 -3630
rect -45 -3634 -41 -3630
rect -29 -3634 -25 -3630
rect -21 -3634 -17 -3630
rect -9 -3634 -5 -3630
rect 3 -3634 7 -3630
rect 12 -3634 16 -3630
rect 21 -3634 25 -3630
rect 209 -3634 213 -3630
rect 218 -3634 222 -3630
rect 227 -3634 231 -3630
rect 235 -3634 239 -3630
rect 244 -3634 248 -3630
rect 253 -3634 257 -3630
rect 261 -3634 265 -3630
rect 269 -3634 273 -3630
rect 287 -3634 291 -3630
rect 297 -3634 301 -3630
rect 305 -3634 309 -3630
rect 322 -3634 326 -3630
rect 331 -3634 335 -3630
rect 339 -3634 343 -3630
rect 348 -3634 352 -3630
rect 366 -3634 370 -3630
rect 375 -3634 379 -3630
rect 383 -3634 387 -3630
rect 399 -3634 403 -3630
rect 407 -3634 411 -3630
rect 419 -3634 423 -3630
rect 431 -3634 435 -3630
rect 440 -3634 444 -3630
rect 449 -3634 453 -3630
rect 565 -3634 569 -3630
rect 574 -3634 578 -3630
rect 583 -3634 587 -3630
rect 591 -3634 595 -3630
rect 600 -3634 604 -3630
rect 609 -3634 613 -3630
rect 617 -3634 621 -3630
rect 625 -3634 629 -3630
rect 643 -3634 647 -3630
rect 653 -3634 657 -3630
rect 661 -3634 665 -3630
rect 678 -3634 682 -3630
rect 687 -3634 691 -3630
rect 695 -3634 699 -3630
rect 704 -3634 708 -3630
rect 722 -3634 726 -3630
rect 731 -3634 735 -3630
rect 739 -3634 743 -3630
rect 755 -3634 759 -3630
rect 763 -3634 767 -3630
rect 775 -3634 779 -3630
rect 787 -3634 791 -3630
rect 796 -3634 800 -3630
rect 805 -3634 809 -3630
rect 963 -3634 967 -3630
rect 972 -3634 976 -3630
rect 981 -3634 985 -3630
rect 989 -3634 993 -3630
rect 998 -3634 1002 -3630
rect 1007 -3634 1011 -3630
rect 1015 -3634 1019 -3630
rect 1023 -3634 1027 -3630
rect 1041 -3634 1045 -3630
rect 1051 -3634 1055 -3630
rect 1059 -3634 1063 -3630
rect 1076 -3634 1080 -3630
rect 1085 -3634 1089 -3630
rect 1093 -3634 1097 -3630
rect 1102 -3634 1106 -3630
rect 1120 -3634 1124 -3630
rect 1129 -3634 1133 -3630
rect 1137 -3634 1141 -3630
rect 1153 -3634 1157 -3630
rect 1161 -3634 1165 -3630
rect 1173 -3634 1177 -3630
rect 1185 -3634 1189 -3630
rect 1194 -3634 1198 -3630
rect 1203 -3634 1207 -3630
rect 1321 -3634 1325 -3630
rect 1330 -3634 1334 -3630
rect 1339 -3634 1343 -3630
rect 1347 -3634 1351 -3630
rect 1356 -3634 1360 -3630
rect 1365 -3634 1369 -3630
rect 1373 -3634 1377 -3630
rect 1381 -3634 1385 -3630
rect 1399 -3634 1403 -3630
rect 1409 -3634 1413 -3630
rect 1417 -3634 1421 -3630
rect 1434 -3634 1438 -3630
rect 1443 -3634 1447 -3630
rect 1451 -3634 1455 -3630
rect 1460 -3634 1464 -3630
rect 1478 -3634 1482 -3630
rect 1487 -3634 1491 -3630
rect 1495 -3634 1499 -3630
rect 1511 -3634 1515 -3630
rect 1519 -3634 1523 -3630
rect 1531 -3634 1535 -3630
rect 1543 -3634 1547 -3630
rect 1552 -3634 1556 -3630
rect 1561 -3634 1565 -3630
rect -1264 -3764 -1260 -3760
rect -1255 -3764 -1251 -3760
rect -1246 -3764 -1242 -3760
rect -1238 -3764 -1234 -3760
rect -1222 -3764 -1218 -3760
rect -1214 -3764 -1210 -3760
rect -1197 -3764 -1193 -3760
rect -1180 -3764 -1176 -3760
rect -1172 -3764 -1168 -3760
rect -1155 -3764 -1151 -3760
rect -1138 -3764 -1134 -3760
rect -1130 -3764 -1126 -3760
rect -1113 -3764 -1109 -3760
rect -1096 -3764 -1092 -3760
rect -1088 -3764 -1084 -3760
rect -1072 -3764 -1068 -3760
rect -935 -3764 -931 -3760
rect -926 -3764 -922 -3760
rect -917 -3764 -913 -3760
rect -909 -3764 -905 -3760
rect -893 -3764 -889 -3760
rect -885 -3764 -881 -3760
rect -868 -3764 -864 -3760
rect -851 -3764 -847 -3760
rect -843 -3764 -839 -3760
rect -826 -3764 -822 -3760
rect -809 -3764 -805 -3760
rect -801 -3764 -797 -3760
rect -784 -3764 -780 -3760
rect -767 -3764 -763 -3760
rect -759 -3764 -755 -3760
rect -743 -3764 -739 -3760
rect -577 -3764 -573 -3760
rect -568 -3764 -564 -3760
rect -559 -3764 -555 -3760
rect -551 -3764 -547 -3760
rect -535 -3764 -531 -3760
rect -527 -3764 -523 -3760
rect -510 -3764 -506 -3760
rect -493 -3764 -489 -3760
rect -485 -3764 -481 -3760
rect -468 -3764 -464 -3760
rect -451 -3764 -447 -3760
rect -443 -3764 -439 -3760
rect -426 -3764 -422 -3760
rect -409 -3764 -405 -3760
rect -401 -3764 -397 -3760
rect -385 -3764 -381 -3760
rect -219 -3764 -215 -3760
rect -210 -3764 -206 -3760
rect -201 -3764 -197 -3760
rect -193 -3764 -189 -3760
rect -177 -3764 -173 -3760
rect -169 -3764 -165 -3760
rect -152 -3764 -148 -3760
rect -135 -3764 -131 -3760
rect -127 -3764 -123 -3760
rect -110 -3764 -106 -3760
rect -93 -3764 -89 -3760
rect -85 -3764 -81 -3760
rect -68 -3764 -64 -3760
rect -51 -3764 -47 -3760
rect -43 -3764 -39 -3760
rect -27 -3764 -23 -3760
rect 68 -3879 72 -3863
rect 76 -3879 80 -3863
rect -1264 -3995 -1260 -3991
rect -1255 -3995 -1251 -3991
rect -1246 -3995 -1242 -3991
rect -1238 -3995 -1234 -3991
rect -1222 -3995 -1218 -3991
rect -1214 -3995 -1210 -3991
rect -1197 -3995 -1193 -3991
rect -1180 -3995 -1176 -3991
rect -1172 -3995 -1168 -3991
rect -1155 -3995 -1151 -3991
rect -1138 -3995 -1134 -3991
rect -1130 -3995 -1126 -3991
rect -1113 -3995 -1109 -3991
rect -1096 -3995 -1092 -3991
rect -1088 -3995 -1084 -3991
rect -1072 -3995 -1068 -3991
rect -935 -3995 -931 -3991
rect -926 -3995 -922 -3991
rect -917 -3995 -913 -3991
rect -909 -3995 -905 -3991
rect -893 -3995 -889 -3991
rect -885 -3995 -881 -3991
rect -868 -3995 -864 -3991
rect -851 -3995 -847 -3991
rect -843 -3995 -839 -3991
rect -826 -3995 -822 -3991
rect -809 -3995 -805 -3991
rect -801 -3995 -797 -3991
rect -784 -3995 -780 -3991
rect -767 -3995 -763 -3991
rect -759 -3995 -755 -3991
rect -743 -3995 -739 -3991
rect -577 -3995 -573 -3991
rect -568 -3995 -564 -3991
rect -559 -3995 -555 -3991
rect -551 -3995 -547 -3991
rect -535 -3995 -531 -3991
rect -527 -3995 -523 -3991
rect -510 -3995 -506 -3991
rect -493 -3995 -489 -3991
rect -485 -3995 -481 -3991
rect -468 -3995 -464 -3991
rect -451 -3995 -447 -3991
rect -443 -3995 -439 -3991
rect -426 -3995 -422 -3991
rect -409 -3995 -405 -3991
rect -401 -3995 -397 -3991
rect -385 -3995 -381 -3991
rect -219 -3995 -215 -3991
rect -210 -3995 -206 -3991
rect -201 -3995 -197 -3991
rect -193 -3995 -189 -3991
rect -177 -3995 -173 -3991
rect -169 -3995 -165 -3991
rect -152 -3995 -148 -3991
rect -135 -3995 -131 -3991
rect -127 -3995 -123 -3991
rect -110 -3995 -106 -3991
rect -93 -3995 -89 -3991
rect -85 -3995 -81 -3991
rect -68 -3995 -64 -3991
rect -51 -3995 -47 -3991
rect -43 -3995 -39 -3991
rect -27 -3995 -23 -3991
rect 209 -3995 213 -3991
rect 218 -3995 222 -3991
rect 227 -3995 231 -3991
rect 235 -3995 239 -3991
rect 251 -3995 255 -3991
rect 259 -3995 263 -3991
rect 276 -3995 280 -3991
rect 293 -3995 297 -3991
rect 301 -3995 305 -3991
rect 318 -3995 322 -3991
rect 335 -3995 339 -3991
rect 343 -3995 347 -3991
rect 360 -3995 364 -3991
rect 377 -3995 381 -3991
rect 385 -3995 389 -3991
rect 401 -3995 405 -3991
rect 565 -3995 569 -3991
rect 574 -3995 578 -3991
rect 583 -3995 587 -3991
rect 591 -3995 595 -3991
rect 607 -3995 611 -3991
rect 615 -3995 619 -3991
rect 632 -3995 636 -3991
rect 649 -3995 653 -3991
rect 657 -3995 661 -3991
rect 674 -3995 678 -3991
rect 691 -3995 695 -3991
rect 699 -3995 703 -3991
rect 716 -3995 720 -3991
rect 733 -3995 737 -3991
rect 741 -3995 745 -3991
rect 757 -3995 761 -3991
rect 963 -3995 967 -3991
rect 972 -3995 976 -3991
rect 981 -3995 985 -3991
rect 989 -3995 993 -3991
rect 1005 -3995 1009 -3991
rect 1013 -3995 1017 -3991
rect 1030 -3995 1034 -3991
rect 1047 -3995 1051 -3991
rect 1055 -3995 1059 -3991
rect 1072 -3995 1076 -3991
rect 1089 -3995 1093 -3991
rect 1097 -3995 1101 -3991
rect 1114 -3995 1118 -3991
rect 1131 -3995 1135 -3991
rect 1139 -3995 1143 -3991
rect 1155 -3995 1159 -3991
rect 1321 -3995 1325 -3991
rect 1330 -3995 1334 -3991
rect 1339 -3995 1343 -3991
rect 1347 -3995 1351 -3991
rect 1363 -3995 1367 -3991
rect 1371 -3995 1375 -3991
rect 1388 -3995 1392 -3991
rect 1405 -3995 1409 -3991
rect 1413 -3995 1417 -3991
rect 1430 -3995 1434 -3991
rect 1447 -3995 1451 -3991
rect 1455 -3995 1459 -3991
rect 1472 -3995 1476 -3991
rect 1489 -3995 1493 -3991
rect 1497 -3995 1501 -3991
rect 1513 -3995 1517 -3991
rect -1264 -4120 -1260 -4116
rect -1255 -4120 -1251 -4116
rect -1246 -4120 -1242 -4116
rect -1238 -4120 -1234 -4116
rect -1222 -4120 -1218 -4116
rect -1214 -4120 -1210 -4116
rect -1197 -4120 -1193 -4116
rect -1180 -4120 -1176 -4116
rect -1172 -4120 -1168 -4116
rect -1155 -4120 -1151 -4116
rect -1138 -4120 -1134 -4116
rect -1130 -4120 -1126 -4116
rect -1113 -4120 -1109 -4116
rect -1096 -4120 -1092 -4116
rect -1088 -4120 -1084 -4116
rect -1072 -4120 -1068 -4116
rect -935 -4120 -931 -4116
rect -926 -4120 -922 -4116
rect -917 -4120 -913 -4116
rect -909 -4120 -905 -4116
rect -893 -4120 -889 -4116
rect -885 -4120 -881 -4116
rect -868 -4120 -864 -4116
rect -851 -4120 -847 -4116
rect -843 -4120 -839 -4116
rect -826 -4120 -822 -4116
rect -809 -4120 -805 -4116
rect -801 -4120 -797 -4116
rect -784 -4120 -780 -4116
rect -767 -4120 -763 -4116
rect -759 -4120 -755 -4116
rect -743 -4120 -739 -4116
rect -577 -4120 -573 -4116
rect -568 -4120 -564 -4116
rect -559 -4120 -555 -4116
rect -551 -4120 -547 -4116
rect -535 -4120 -531 -4116
rect -527 -4120 -523 -4116
rect -510 -4120 -506 -4116
rect -493 -4120 -489 -4116
rect -485 -4120 -481 -4116
rect -468 -4120 -464 -4116
rect -451 -4120 -447 -4116
rect -443 -4120 -439 -4116
rect -426 -4120 -422 -4116
rect -409 -4120 -405 -4116
rect -401 -4120 -397 -4116
rect -385 -4120 -381 -4116
rect -219 -4120 -215 -4116
rect -210 -4120 -206 -4116
rect -201 -4120 -197 -4116
rect -193 -4120 -189 -4116
rect -177 -4120 -173 -4116
rect -169 -4120 -165 -4116
rect -152 -4120 -148 -4116
rect -135 -4120 -131 -4116
rect -127 -4120 -123 -4116
rect -110 -4120 -106 -4116
rect -93 -4120 -89 -4116
rect -85 -4120 -81 -4116
rect -68 -4120 -64 -4116
rect -51 -4120 -47 -4116
rect -43 -4120 -39 -4116
rect -27 -4120 -23 -4116
rect 209 -4120 213 -4116
rect 218 -4120 222 -4116
rect 227 -4120 231 -4116
rect 235 -4120 239 -4116
rect 251 -4120 255 -4116
rect 259 -4120 263 -4116
rect 276 -4120 280 -4116
rect 293 -4120 297 -4116
rect 301 -4120 305 -4116
rect 318 -4120 322 -4116
rect 335 -4120 339 -4116
rect 343 -4120 347 -4116
rect 360 -4120 364 -4116
rect 377 -4120 381 -4116
rect 385 -4120 389 -4116
rect 401 -4120 405 -4116
rect 565 -4120 569 -4116
rect 574 -4120 578 -4116
rect 583 -4120 587 -4116
rect 591 -4120 595 -4116
rect 607 -4120 611 -4116
rect 615 -4120 619 -4116
rect 632 -4120 636 -4116
rect 649 -4120 653 -4116
rect 657 -4120 661 -4116
rect 674 -4120 678 -4116
rect 691 -4120 695 -4116
rect 699 -4120 703 -4116
rect 716 -4120 720 -4116
rect 733 -4120 737 -4116
rect 741 -4120 745 -4116
rect 757 -4120 761 -4116
rect 963 -4120 967 -4116
rect 972 -4120 976 -4116
rect 981 -4120 985 -4116
rect 989 -4120 993 -4116
rect 1005 -4120 1009 -4116
rect 1013 -4120 1017 -4116
rect 1030 -4120 1034 -4116
rect 1047 -4120 1051 -4116
rect 1055 -4120 1059 -4116
rect 1072 -4120 1076 -4116
rect 1089 -4120 1093 -4116
rect 1097 -4120 1101 -4116
rect 1114 -4120 1118 -4116
rect 1131 -4120 1135 -4116
rect 1139 -4120 1143 -4116
rect 1155 -4120 1159 -4116
rect 1321 -4120 1325 -4116
rect 1330 -4120 1334 -4116
rect 1339 -4120 1343 -4116
rect 1347 -4120 1351 -4116
rect 1363 -4120 1367 -4116
rect 1371 -4120 1375 -4116
rect 1388 -4120 1392 -4116
rect 1405 -4120 1409 -4116
rect 1413 -4120 1417 -4116
rect 1430 -4120 1434 -4116
rect 1447 -4120 1451 -4116
rect 1455 -4120 1459 -4116
rect 1472 -4120 1476 -4116
rect 1489 -4120 1493 -4116
rect 1497 -4120 1501 -4116
rect 1513 -4120 1517 -4116
rect -1264 -4244 -1260 -4240
rect -1255 -4244 -1251 -4240
rect -1246 -4244 -1242 -4240
rect -1238 -4244 -1234 -4240
rect -1222 -4244 -1218 -4240
rect -1214 -4244 -1210 -4240
rect -1197 -4244 -1193 -4240
rect -1180 -4244 -1176 -4240
rect -1172 -4244 -1168 -4240
rect -1155 -4244 -1151 -4240
rect -1138 -4244 -1134 -4240
rect -1130 -4244 -1126 -4240
rect -1113 -4244 -1109 -4240
rect -1096 -4244 -1092 -4240
rect -1088 -4244 -1084 -4240
rect -1072 -4244 -1068 -4240
rect -1029 -4244 -1025 -4240
rect -1021 -4244 -1017 -4240
rect -935 -4244 -931 -4240
rect -926 -4244 -922 -4240
rect -917 -4244 -913 -4240
rect -909 -4244 -905 -4240
rect -893 -4244 -889 -4240
rect -885 -4244 -881 -4240
rect -868 -4244 -864 -4240
rect -851 -4244 -847 -4240
rect -843 -4244 -839 -4240
rect -826 -4244 -822 -4240
rect -809 -4244 -805 -4240
rect -801 -4244 -797 -4240
rect -784 -4244 -780 -4240
rect -767 -4244 -763 -4240
rect -759 -4244 -755 -4240
rect -743 -4244 -739 -4240
rect -577 -4244 -573 -4240
rect -568 -4244 -564 -4240
rect -559 -4244 -555 -4240
rect -551 -4244 -547 -4240
rect -535 -4244 -531 -4240
rect -527 -4244 -523 -4240
rect -510 -4244 -506 -4240
rect -493 -4244 -489 -4240
rect -485 -4244 -481 -4240
rect -468 -4244 -464 -4240
rect -451 -4244 -447 -4240
rect -443 -4244 -439 -4240
rect -426 -4244 -422 -4240
rect -409 -4244 -405 -4240
rect -401 -4244 -397 -4240
rect -385 -4244 -381 -4240
rect -332 -4244 -328 -4240
rect -324 -4244 -320 -4240
rect -219 -4244 -215 -4240
rect -210 -4244 -206 -4240
rect -201 -4244 -197 -4240
rect -193 -4244 -189 -4240
rect -177 -4244 -173 -4240
rect -169 -4244 -165 -4240
rect -152 -4244 -148 -4240
rect -135 -4244 -131 -4240
rect -127 -4244 -123 -4240
rect -110 -4244 -106 -4240
rect -93 -4244 -89 -4240
rect -85 -4244 -81 -4240
rect -68 -4244 -64 -4240
rect -51 -4244 -47 -4240
rect -43 -4244 -39 -4240
rect -27 -4244 -23 -4240
rect 456 -4244 460 -4240
rect 464 -4244 468 -4240
rect 1201 -4244 1205 -4240
rect 1209 -4244 1213 -4240
rect -1339 -4355 -1335 -4351
rect -1322 -4355 -1318 -4351
rect -1313 -4355 -1309 -4351
rect -1029 -4355 -1025 -4351
rect -1021 -4355 -1017 -4351
rect -935 -4355 -931 -4351
rect -918 -4355 -914 -4351
rect -909 -4355 -905 -4351
rect -673 -4355 -669 -4347
rect -665 -4355 -661 -4347
rect -577 -4355 -573 -4351
rect -560 -4355 -556 -4351
rect -551 -4355 -547 -4351
rect -332 -4355 -328 -4351
rect -324 -4355 -320 -4351
rect -219 -4355 -215 -4351
rect -202 -4355 -198 -4351
rect -193 -4355 -189 -4351
rect 209 -4355 213 -4351
rect 226 -4355 230 -4351
rect 235 -4355 239 -4351
rect 456 -4355 460 -4351
rect 464 -4355 468 -4351
rect 565 -4355 569 -4351
rect 582 -4355 586 -4351
rect 591 -4355 595 -4351
rect 860 -4355 864 -4347
rect 868 -4355 872 -4347
rect 963 -4355 967 -4351
rect 980 -4355 984 -4351
rect 989 -4355 993 -4351
rect 1201 -4355 1205 -4351
rect 1209 -4355 1213 -4351
rect 1321 -4355 1325 -4351
rect 1338 -4355 1342 -4351
rect 1347 -4355 1351 -4351
rect -1264 -4474 -1260 -4470
rect -1255 -4474 -1251 -4470
rect -1246 -4474 -1242 -4470
rect -1238 -4474 -1234 -4470
rect -1229 -4474 -1225 -4470
rect -1211 -4474 -1207 -4470
rect -1202 -4474 -1198 -4470
rect -1194 -4474 -1190 -4470
rect -1177 -4474 -1173 -4470
rect -1168 -4474 -1164 -4470
rect -935 -4474 -931 -4470
rect -926 -4474 -922 -4470
rect -917 -4474 -913 -4470
rect -909 -4474 -905 -4470
rect -900 -4474 -896 -4470
rect -891 -4474 -887 -4470
rect -883 -4474 -879 -4470
rect -875 -4474 -871 -4470
rect -857 -4474 -853 -4470
rect -847 -4474 -843 -4470
rect -839 -4474 -835 -4470
rect -822 -4474 -818 -4470
rect -813 -4474 -809 -4470
rect -805 -4474 -801 -4470
rect -796 -4474 -792 -4470
rect -778 -4474 -774 -4470
rect -769 -4474 -765 -4470
rect -761 -4474 -757 -4470
rect -745 -4474 -741 -4470
rect -737 -4474 -733 -4470
rect -725 -4474 -721 -4470
rect -713 -4474 -709 -4470
rect -704 -4474 -700 -4470
rect -695 -4474 -691 -4470
rect -577 -4474 -573 -4470
rect -568 -4474 -564 -4470
rect -559 -4474 -555 -4470
rect -551 -4474 -547 -4470
rect -542 -4474 -538 -4470
rect -533 -4474 -529 -4470
rect -525 -4474 -521 -4470
rect -517 -4474 -513 -4470
rect -499 -4474 -495 -4470
rect -489 -4474 -485 -4470
rect -481 -4474 -477 -4470
rect -464 -4474 -460 -4470
rect -455 -4474 -451 -4470
rect -447 -4474 -443 -4470
rect -438 -4474 -434 -4470
rect -420 -4474 -416 -4470
rect -411 -4474 -407 -4470
rect -403 -4474 -399 -4470
rect -387 -4474 -383 -4470
rect -379 -4474 -375 -4470
rect -367 -4474 -363 -4470
rect -355 -4474 -351 -4470
rect -346 -4474 -342 -4470
rect -337 -4474 -333 -4470
rect -219 -4474 -215 -4470
rect -210 -4474 -206 -4470
rect -201 -4474 -197 -4470
rect -193 -4474 -189 -4470
rect -184 -4474 -180 -4470
rect -175 -4474 -171 -4470
rect -167 -4474 -163 -4470
rect -159 -4474 -155 -4470
rect -141 -4474 -137 -4470
rect -131 -4474 -127 -4470
rect -123 -4474 -119 -4470
rect -106 -4474 -102 -4470
rect -97 -4474 -93 -4470
rect -89 -4474 -85 -4470
rect -80 -4474 -76 -4470
rect -62 -4474 -58 -4470
rect -53 -4474 -49 -4470
rect -45 -4474 -41 -4470
rect -29 -4474 -25 -4470
rect -21 -4474 -17 -4470
rect -9 -4474 -5 -4470
rect 3 -4474 7 -4470
rect 12 -4474 16 -4470
rect 21 -4474 25 -4470
rect 209 -4474 213 -4470
rect 218 -4474 222 -4470
rect 227 -4474 231 -4470
rect 235 -4474 239 -4470
rect 244 -4474 248 -4470
rect 253 -4474 257 -4470
rect 261 -4474 265 -4470
rect 269 -4474 273 -4470
rect 287 -4474 291 -4470
rect 297 -4474 301 -4470
rect 305 -4474 309 -4470
rect 322 -4474 326 -4470
rect 331 -4474 335 -4470
rect 339 -4474 343 -4470
rect 348 -4474 352 -4470
rect 366 -4474 370 -4470
rect 375 -4474 379 -4470
rect 383 -4474 387 -4470
rect 399 -4474 403 -4470
rect 407 -4474 411 -4470
rect 419 -4474 423 -4470
rect 431 -4474 435 -4470
rect 440 -4474 444 -4470
rect 449 -4474 453 -4470
rect 565 -4474 569 -4470
rect 574 -4474 578 -4470
rect 583 -4474 587 -4470
rect 591 -4474 595 -4470
rect 600 -4474 604 -4470
rect 609 -4474 613 -4470
rect 617 -4474 621 -4470
rect 625 -4474 629 -4470
rect 643 -4474 647 -4470
rect 653 -4474 657 -4470
rect 661 -4474 665 -4470
rect 678 -4474 682 -4470
rect 687 -4474 691 -4470
rect 695 -4474 699 -4470
rect 704 -4474 708 -4470
rect 722 -4474 726 -4470
rect 731 -4474 735 -4470
rect 739 -4474 743 -4470
rect 755 -4474 759 -4470
rect 763 -4474 767 -4470
rect 775 -4474 779 -4470
rect 787 -4474 791 -4470
rect 796 -4474 800 -4470
rect 805 -4474 809 -4470
rect 963 -4474 967 -4470
rect 972 -4474 976 -4470
rect 981 -4474 985 -4470
rect 989 -4474 993 -4470
rect 998 -4474 1002 -4470
rect 1007 -4474 1011 -4470
rect 1015 -4474 1019 -4470
rect 1023 -4474 1027 -4470
rect 1041 -4474 1045 -4470
rect 1051 -4474 1055 -4470
rect 1059 -4474 1063 -4470
rect 1076 -4474 1080 -4470
rect 1085 -4474 1089 -4470
rect 1093 -4474 1097 -4470
rect 1102 -4474 1106 -4470
rect 1120 -4474 1124 -4470
rect 1129 -4474 1133 -4470
rect 1137 -4474 1141 -4470
rect 1153 -4474 1157 -4470
rect 1161 -4474 1165 -4470
rect 1173 -4474 1177 -4470
rect 1185 -4474 1189 -4470
rect 1194 -4474 1198 -4470
rect 1203 -4474 1207 -4470
rect 1321 -4474 1325 -4470
rect 1330 -4474 1334 -4470
rect 1339 -4474 1343 -4470
rect 1347 -4474 1351 -4470
rect 1356 -4474 1360 -4470
rect 1365 -4474 1369 -4470
rect 1373 -4474 1377 -4470
rect 1381 -4474 1385 -4470
rect 1399 -4474 1403 -4470
rect 1409 -4474 1413 -4470
rect 1417 -4474 1421 -4470
rect 1434 -4474 1438 -4470
rect 1443 -4474 1447 -4470
rect 1451 -4474 1455 -4470
rect 1460 -4474 1464 -4470
rect 1478 -4474 1482 -4470
rect 1487 -4474 1491 -4470
rect 1495 -4474 1499 -4470
rect 1511 -4474 1515 -4470
rect 1519 -4474 1523 -4470
rect 1531 -4474 1535 -4470
rect 1543 -4474 1547 -4470
rect 1552 -4474 1556 -4470
rect 1561 -4474 1565 -4470
rect -1264 -4597 -1260 -4593
rect -1255 -4597 -1251 -4593
rect -1246 -4597 -1242 -4593
rect -1238 -4597 -1234 -4593
rect -1222 -4597 -1218 -4593
rect -1214 -4597 -1210 -4593
rect -1197 -4597 -1193 -4593
rect -1180 -4597 -1176 -4593
rect -1172 -4597 -1168 -4593
rect -1155 -4597 -1151 -4593
rect -1138 -4597 -1134 -4593
rect -1130 -4597 -1126 -4593
rect -1113 -4597 -1109 -4593
rect -1096 -4597 -1092 -4593
rect -1088 -4597 -1084 -4593
rect -1072 -4597 -1068 -4593
rect -935 -4597 -931 -4593
rect -926 -4597 -922 -4593
rect -917 -4597 -913 -4593
rect -909 -4597 -905 -4593
rect -893 -4597 -889 -4593
rect -885 -4597 -881 -4593
rect -868 -4597 -864 -4593
rect -851 -4597 -847 -4593
rect -843 -4597 -839 -4593
rect -826 -4597 -822 -4593
rect -809 -4597 -805 -4593
rect -801 -4597 -797 -4593
rect -784 -4597 -780 -4593
rect -767 -4597 -763 -4593
rect -759 -4597 -755 -4593
rect -743 -4597 -739 -4593
rect -577 -4597 -573 -4593
rect -568 -4597 -564 -4593
rect -559 -4597 -555 -4593
rect -551 -4597 -547 -4593
rect -535 -4597 -531 -4593
rect -527 -4597 -523 -4593
rect -510 -4597 -506 -4593
rect -493 -4597 -489 -4593
rect -485 -4597 -481 -4593
rect -468 -4597 -464 -4593
rect -451 -4597 -447 -4593
rect -443 -4597 -439 -4593
rect -426 -4597 -422 -4593
rect -409 -4597 -405 -4593
rect -401 -4597 -397 -4593
rect -385 -4597 -381 -4593
rect -1264 -4718 -1260 -4714
rect -1255 -4718 -1251 -4714
rect -1246 -4718 -1242 -4714
rect -1238 -4718 -1234 -4714
rect -1222 -4718 -1218 -4714
rect -1214 -4718 -1210 -4714
rect -1197 -4718 -1193 -4714
rect -1180 -4718 -1176 -4714
rect -1172 -4718 -1168 -4714
rect -1155 -4718 -1151 -4714
rect -1138 -4718 -1134 -4714
rect -1130 -4718 -1126 -4714
rect -1113 -4718 -1109 -4714
rect -1096 -4718 -1092 -4714
rect -1088 -4718 -1084 -4714
rect -1072 -4718 -1068 -4714
rect -935 -4718 -931 -4714
rect -926 -4718 -922 -4714
rect -917 -4718 -913 -4714
rect -909 -4718 -905 -4714
rect -893 -4718 -889 -4714
rect -885 -4718 -881 -4714
rect -868 -4718 -864 -4714
rect -851 -4718 -847 -4714
rect -843 -4718 -839 -4714
rect -826 -4718 -822 -4714
rect -809 -4718 -805 -4714
rect -801 -4718 -797 -4714
rect -784 -4718 -780 -4714
rect -767 -4718 -763 -4714
rect -759 -4718 -755 -4714
rect -743 -4718 -739 -4714
rect -577 -4718 -573 -4714
rect -568 -4718 -564 -4714
rect -559 -4718 -555 -4714
rect -551 -4718 -547 -4714
rect -535 -4718 -531 -4714
rect -527 -4718 -523 -4714
rect -510 -4718 -506 -4714
rect -493 -4718 -489 -4714
rect -485 -4718 -481 -4714
rect -468 -4718 -464 -4714
rect -451 -4718 -447 -4714
rect -443 -4718 -439 -4714
rect -426 -4718 -422 -4714
rect -409 -4718 -405 -4714
rect -401 -4718 -397 -4714
rect -385 -4718 -381 -4714
rect -219 -4718 -215 -4714
rect -210 -4718 -206 -4714
rect -201 -4718 -197 -4714
rect -193 -4718 -189 -4714
rect -177 -4718 -173 -4714
rect -169 -4718 -165 -4714
rect -152 -4718 -148 -4714
rect -135 -4718 -131 -4714
rect -127 -4718 -123 -4714
rect -110 -4718 -106 -4714
rect -93 -4718 -89 -4714
rect -85 -4718 -81 -4714
rect -68 -4718 -64 -4714
rect -51 -4718 -47 -4714
rect -43 -4718 -39 -4714
rect -27 -4718 -23 -4714
rect 209 -4718 213 -4714
rect 218 -4718 222 -4714
rect 227 -4718 231 -4714
rect 235 -4718 239 -4714
rect 251 -4718 255 -4714
rect 259 -4718 263 -4714
rect 276 -4718 280 -4714
rect 293 -4718 297 -4714
rect 301 -4718 305 -4714
rect 318 -4718 322 -4714
rect 335 -4718 339 -4714
rect 343 -4718 347 -4714
rect 360 -4718 364 -4714
rect 377 -4718 381 -4714
rect 385 -4718 389 -4714
rect 401 -4718 405 -4714
rect 565 -4718 569 -4714
rect 574 -4718 578 -4714
rect 583 -4718 587 -4714
rect 591 -4718 595 -4714
rect 607 -4718 611 -4714
rect 615 -4718 619 -4714
rect 632 -4718 636 -4714
rect 649 -4718 653 -4714
rect 657 -4718 661 -4714
rect 674 -4718 678 -4714
rect 691 -4718 695 -4714
rect 699 -4718 703 -4714
rect 716 -4718 720 -4714
rect 733 -4718 737 -4714
rect 741 -4718 745 -4714
rect 757 -4718 761 -4714
rect 963 -4718 967 -4714
rect 972 -4718 976 -4714
rect 981 -4718 985 -4714
rect 989 -4718 993 -4714
rect 1005 -4718 1009 -4714
rect 1013 -4718 1017 -4714
rect 1030 -4718 1034 -4714
rect 1047 -4718 1051 -4714
rect 1055 -4718 1059 -4714
rect 1072 -4718 1076 -4714
rect 1089 -4718 1093 -4714
rect 1097 -4718 1101 -4714
rect 1114 -4718 1118 -4714
rect 1131 -4718 1135 -4714
rect 1139 -4718 1143 -4714
rect 1155 -4718 1159 -4714
rect 1321 -4718 1325 -4714
rect 1330 -4718 1334 -4714
rect 1339 -4718 1343 -4714
rect 1347 -4718 1351 -4714
rect 1363 -4718 1367 -4714
rect 1371 -4718 1375 -4714
rect 1388 -4718 1392 -4714
rect 1405 -4718 1409 -4714
rect 1413 -4718 1417 -4714
rect 1430 -4718 1434 -4714
rect 1447 -4718 1451 -4714
rect 1455 -4718 1459 -4714
rect 1472 -4718 1476 -4714
rect 1489 -4718 1493 -4714
rect 1497 -4718 1501 -4714
rect 1513 -4718 1517 -4714
rect -1264 -4839 -1260 -4835
rect -1255 -4839 -1251 -4835
rect -1246 -4839 -1242 -4835
rect -1238 -4839 -1234 -4835
rect -1222 -4839 -1218 -4835
rect -1214 -4839 -1210 -4835
rect -1197 -4839 -1193 -4835
rect -1180 -4839 -1176 -4835
rect -1172 -4839 -1168 -4835
rect -1155 -4839 -1151 -4835
rect -1138 -4839 -1134 -4835
rect -1130 -4839 -1126 -4835
rect -1113 -4839 -1109 -4835
rect -1096 -4839 -1092 -4835
rect -1088 -4839 -1084 -4835
rect -1072 -4839 -1068 -4835
rect -935 -4839 -931 -4835
rect -926 -4839 -922 -4835
rect -917 -4839 -913 -4835
rect -909 -4839 -905 -4835
rect -893 -4839 -889 -4835
rect -885 -4839 -881 -4835
rect -868 -4839 -864 -4835
rect -851 -4839 -847 -4835
rect -843 -4839 -839 -4835
rect -826 -4839 -822 -4835
rect -809 -4839 -805 -4835
rect -801 -4839 -797 -4835
rect -784 -4839 -780 -4835
rect -767 -4839 -763 -4835
rect -759 -4839 -755 -4835
rect -743 -4839 -739 -4835
rect -577 -4839 -573 -4835
rect -568 -4839 -564 -4835
rect -559 -4839 -555 -4835
rect -551 -4839 -547 -4835
rect -535 -4839 -531 -4835
rect -527 -4839 -523 -4835
rect -510 -4839 -506 -4835
rect -493 -4839 -489 -4835
rect -485 -4839 -481 -4835
rect -468 -4839 -464 -4835
rect -451 -4839 -447 -4835
rect -443 -4839 -439 -4835
rect -426 -4839 -422 -4835
rect -409 -4839 -405 -4835
rect -401 -4839 -397 -4835
rect -385 -4839 -381 -4835
rect -219 -4839 -215 -4835
rect -210 -4839 -206 -4835
rect -201 -4839 -197 -4835
rect -193 -4839 -189 -4835
rect -177 -4839 -173 -4835
rect -169 -4839 -165 -4835
rect -152 -4839 -148 -4835
rect -135 -4839 -131 -4835
rect -127 -4839 -123 -4835
rect -110 -4839 -106 -4835
rect -93 -4839 -89 -4835
rect -85 -4839 -81 -4835
rect -68 -4839 -64 -4835
rect -51 -4839 -47 -4835
rect -43 -4839 -39 -4835
rect -27 -4839 -23 -4835
rect 90 -4839 94 -4823
rect 98 -4839 102 -4823
rect 209 -4839 213 -4835
rect 218 -4839 222 -4835
rect 227 -4839 231 -4835
rect 235 -4839 239 -4835
rect 251 -4839 255 -4835
rect 259 -4839 263 -4835
rect 276 -4839 280 -4835
rect 293 -4839 297 -4835
rect 301 -4839 305 -4835
rect 318 -4839 322 -4835
rect 335 -4839 339 -4835
rect 343 -4839 347 -4835
rect 360 -4839 364 -4835
rect 377 -4839 381 -4835
rect 385 -4839 389 -4835
rect 401 -4839 405 -4835
rect 565 -4839 569 -4835
rect 574 -4839 578 -4835
rect 583 -4839 587 -4835
rect 591 -4839 595 -4835
rect 607 -4839 611 -4835
rect 615 -4839 619 -4835
rect 632 -4839 636 -4835
rect 649 -4839 653 -4835
rect 657 -4839 661 -4835
rect 674 -4839 678 -4835
rect 691 -4839 695 -4835
rect 699 -4839 703 -4835
rect 716 -4839 720 -4835
rect 733 -4839 737 -4835
rect 741 -4839 745 -4835
rect 757 -4839 761 -4835
rect 963 -4839 967 -4835
rect 972 -4839 976 -4835
rect 981 -4839 985 -4835
rect 989 -4839 993 -4835
rect 1005 -4839 1009 -4835
rect 1013 -4839 1017 -4835
rect 1030 -4839 1034 -4835
rect 1047 -4839 1051 -4835
rect 1055 -4839 1059 -4835
rect 1072 -4839 1076 -4835
rect 1089 -4839 1093 -4835
rect 1097 -4839 1101 -4835
rect 1114 -4839 1118 -4835
rect 1131 -4839 1135 -4835
rect 1139 -4839 1143 -4835
rect 1155 -4839 1159 -4835
rect 1321 -4839 1325 -4835
rect 1330 -4839 1334 -4835
rect 1339 -4839 1343 -4835
rect 1347 -4839 1351 -4835
rect 1363 -4839 1367 -4835
rect 1371 -4839 1375 -4835
rect 1388 -4839 1392 -4835
rect 1405 -4839 1409 -4835
rect 1413 -4839 1417 -4835
rect 1430 -4839 1434 -4835
rect 1447 -4839 1451 -4835
rect 1455 -4839 1459 -4835
rect 1472 -4839 1476 -4835
rect 1489 -4839 1493 -4835
rect 1497 -4839 1501 -4835
rect 1513 -4839 1517 -4835
rect -1264 -4957 -1260 -4953
rect -1255 -4957 -1251 -4953
rect -1246 -4957 -1242 -4953
rect -1238 -4957 -1234 -4953
rect -1222 -4957 -1218 -4953
rect -1214 -4957 -1210 -4953
rect -1197 -4957 -1193 -4953
rect -1180 -4957 -1176 -4953
rect -1172 -4957 -1168 -4953
rect -1155 -4957 -1151 -4953
rect -1138 -4957 -1134 -4953
rect -1130 -4957 -1126 -4953
rect -1113 -4957 -1109 -4953
rect -1096 -4957 -1092 -4953
rect -1088 -4957 -1084 -4953
rect -1072 -4957 -1068 -4953
rect -935 -4957 -931 -4953
rect -926 -4957 -922 -4953
rect -917 -4957 -913 -4953
rect -909 -4957 -905 -4953
rect -893 -4957 -889 -4953
rect -885 -4957 -881 -4953
rect -868 -4957 -864 -4953
rect -851 -4957 -847 -4953
rect -843 -4957 -839 -4953
rect -826 -4957 -822 -4953
rect -809 -4957 -805 -4953
rect -801 -4957 -797 -4953
rect -784 -4957 -780 -4953
rect -767 -4957 -763 -4953
rect -759 -4957 -755 -4953
rect -743 -4957 -739 -4953
rect -577 -4957 -573 -4953
rect -568 -4957 -564 -4953
rect -559 -4957 -555 -4953
rect -551 -4957 -547 -4953
rect -535 -4957 -531 -4953
rect -527 -4957 -523 -4953
rect -510 -4957 -506 -4953
rect -493 -4957 -489 -4953
rect -485 -4957 -481 -4953
rect -468 -4957 -464 -4953
rect -451 -4957 -447 -4953
rect -443 -4957 -439 -4953
rect -426 -4957 -422 -4953
rect -409 -4957 -405 -4953
rect -401 -4957 -397 -4953
rect -385 -4957 -381 -4953
rect -219 -4957 -215 -4953
rect -210 -4957 -206 -4953
rect -201 -4957 -197 -4953
rect -193 -4957 -189 -4953
rect -177 -4957 -173 -4953
rect -169 -4957 -165 -4953
rect -152 -4957 -148 -4953
rect -135 -4957 -131 -4953
rect -127 -4957 -123 -4953
rect -110 -4957 -106 -4953
rect -93 -4957 -89 -4953
rect -85 -4957 -81 -4953
rect -68 -4957 -64 -4953
rect -51 -4957 -47 -4953
rect -43 -4957 -39 -4953
rect -27 -4957 -23 -4953
rect 209 -4957 213 -4953
rect 218 -4957 222 -4953
rect 227 -4957 231 -4953
rect 235 -4957 239 -4953
rect 251 -4957 255 -4953
rect 259 -4957 263 -4953
rect 276 -4957 280 -4953
rect 293 -4957 297 -4953
rect 301 -4957 305 -4953
rect 318 -4957 322 -4953
rect 335 -4957 339 -4953
rect 343 -4957 347 -4953
rect 360 -4957 364 -4953
rect 377 -4957 381 -4953
rect 385 -4957 389 -4953
rect 401 -4957 405 -4953
rect -1339 -5074 -1335 -5070
rect -1322 -5074 -1318 -5070
rect -1313 -5074 -1309 -5070
rect -935 -5074 -931 -5070
rect -918 -5074 -914 -5070
rect -909 -5074 -905 -5070
rect -577 -5074 -573 -5070
rect -560 -5074 -556 -5070
rect -551 -5074 -547 -5070
rect -219 -5074 -215 -5070
rect -202 -5074 -198 -5070
rect -193 -5074 -189 -5070
rect 209 -5074 213 -5070
rect 226 -5074 230 -5070
rect 235 -5074 239 -5070
rect 565 -5074 569 -5070
rect 582 -5074 586 -5070
rect 591 -5074 595 -5070
rect 963 -5074 967 -5070
rect 980 -5074 984 -5070
rect 989 -5074 993 -5070
rect 1321 -5074 1325 -5070
rect 1338 -5074 1342 -5070
rect 1347 -5074 1351 -5070
rect -1264 -5193 -1260 -5189
rect -1255 -5193 -1251 -5189
rect -1246 -5193 -1242 -5189
rect -1238 -5193 -1234 -5189
rect -1229 -5193 -1225 -5189
rect -1211 -5193 -1207 -5189
rect -1202 -5193 -1198 -5189
rect -1194 -5193 -1190 -5189
rect -1177 -5193 -1173 -5189
rect -1168 -5193 -1164 -5189
rect -935 -5193 -931 -5189
rect -926 -5193 -922 -5189
rect -917 -5193 -913 -5189
rect -909 -5193 -905 -5189
rect -900 -5193 -896 -5189
rect -891 -5193 -887 -5189
rect -883 -5193 -879 -5189
rect -875 -5193 -871 -5189
rect -857 -5193 -853 -5189
rect -847 -5193 -843 -5189
rect -839 -5193 -835 -5189
rect -822 -5193 -818 -5189
rect -813 -5193 -809 -5189
rect -805 -5193 -801 -5189
rect -796 -5193 -792 -5189
rect -778 -5193 -774 -5189
rect -769 -5193 -765 -5189
rect -761 -5193 -757 -5189
rect -745 -5193 -741 -5189
rect -737 -5193 -733 -5189
rect -725 -5193 -721 -5189
rect -713 -5193 -709 -5189
rect -704 -5193 -700 -5189
rect -695 -5193 -691 -5189
rect -577 -5193 -573 -5189
rect -568 -5193 -564 -5189
rect -559 -5193 -555 -5189
rect -551 -5193 -547 -5189
rect -542 -5193 -538 -5189
rect -533 -5193 -529 -5189
rect -525 -5193 -521 -5189
rect -517 -5193 -513 -5189
rect -499 -5193 -495 -5189
rect -489 -5193 -485 -5189
rect -481 -5193 -477 -5189
rect -464 -5193 -460 -5189
rect -455 -5193 -451 -5189
rect -447 -5193 -443 -5189
rect -438 -5193 -434 -5189
rect -420 -5193 -416 -5189
rect -411 -5193 -407 -5189
rect -403 -5193 -399 -5189
rect -387 -5193 -383 -5189
rect -379 -5193 -375 -5189
rect -367 -5193 -363 -5189
rect -355 -5193 -351 -5189
rect -346 -5193 -342 -5189
rect -337 -5193 -333 -5189
rect -219 -5193 -215 -5189
rect -210 -5193 -206 -5189
rect -201 -5193 -197 -5189
rect -193 -5193 -189 -5189
rect -184 -5193 -180 -5189
rect -175 -5193 -171 -5189
rect -167 -5193 -163 -5189
rect -159 -5193 -155 -5189
rect -141 -5193 -137 -5189
rect -131 -5193 -127 -5189
rect -123 -5193 -119 -5189
rect -106 -5193 -102 -5189
rect -97 -5193 -93 -5189
rect -89 -5193 -85 -5189
rect -80 -5193 -76 -5189
rect -62 -5193 -58 -5189
rect -53 -5193 -49 -5189
rect -45 -5193 -41 -5189
rect -29 -5193 -25 -5189
rect -21 -5193 -17 -5189
rect -9 -5193 -5 -5189
rect 3 -5193 7 -5189
rect 12 -5193 16 -5189
rect 21 -5193 25 -5189
rect 209 -5193 213 -5189
rect 218 -5193 222 -5189
rect 227 -5193 231 -5189
rect 235 -5193 239 -5189
rect 244 -5193 248 -5189
rect 253 -5193 257 -5189
rect 261 -5193 265 -5189
rect 269 -5193 273 -5189
rect 287 -5193 291 -5189
rect 297 -5193 301 -5189
rect 305 -5193 309 -5189
rect 322 -5193 326 -5189
rect 331 -5193 335 -5189
rect 339 -5193 343 -5189
rect 348 -5193 352 -5189
rect 366 -5193 370 -5189
rect 375 -5193 379 -5189
rect 383 -5193 387 -5189
rect 399 -5193 403 -5189
rect 407 -5193 411 -5189
rect 419 -5193 423 -5189
rect 431 -5193 435 -5189
rect 440 -5193 444 -5189
rect 449 -5193 453 -5189
rect 565 -5193 569 -5189
rect 574 -5193 578 -5189
rect 583 -5193 587 -5189
rect 591 -5193 595 -5189
rect 600 -5193 604 -5189
rect 609 -5193 613 -5189
rect 617 -5193 621 -5189
rect 625 -5193 629 -5189
rect 643 -5193 647 -5189
rect 653 -5193 657 -5189
rect 661 -5193 665 -5189
rect 678 -5193 682 -5189
rect 687 -5193 691 -5189
rect 695 -5193 699 -5189
rect 704 -5193 708 -5189
rect 722 -5193 726 -5189
rect 731 -5193 735 -5189
rect 739 -5193 743 -5189
rect 755 -5193 759 -5189
rect 763 -5193 767 -5189
rect 775 -5193 779 -5189
rect 787 -5193 791 -5189
rect 796 -5193 800 -5189
rect 805 -5193 809 -5189
rect 963 -5193 967 -5189
rect 972 -5193 976 -5189
rect 981 -5193 985 -5189
rect 989 -5193 993 -5189
rect 998 -5193 1002 -5189
rect 1007 -5193 1011 -5189
rect 1015 -5193 1019 -5189
rect 1023 -5193 1027 -5189
rect 1041 -5193 1045 -5189
rect 1051 -5193 1055 -5189
rect 1059 -5193 1063 -5189
rect 1076 -5193 1080 -5189
rect 1085 -5193 1089 -5189
rect 1093 -5193 1097 -5189
rect 1102 -5193 1106 -5189
rect 1120 -5193 1124 -5189
rect 1129 -5193 1133 -5189
rect 1137 -5193 1141 -5189
rect 1153 -5193 1157 -5189
rect 1161 -5193 1165 -5189
rect 1173 -5193 1177 -5189
rect 1185 -5193 1189 -5189
rect 1194 -5193 1198 -5189
rect 1203 -5193 1207 -5189
rect 1321 -5193 1325 -5189
rect 1330 -5193 1334 -5189
rect 1339 -5193 1343 -5189
rect 1347 -5193 1351 -5189
rect 1356 -5193 1360 -5189
rect 1365 -5193 1369 -5189
rect 1373 -5193 1377 -5189
rect 1381 -5193 1385 -5189
rect 1399 -5193 1403 -5189
rect 1409 -5193 1413 -5189
rect 1417 -5193 1421 -5189
rect 1434 -5193 1438 -5189
rect 1443 -5193 1447 -5189
rect 1451 -5193 1455 -5189
rect 1460 -5193 1464 -5189
rect 1478 -5193 1482 -5189
rect 1487 -5193 1491 -5189
rect 1495 -5193 1499 -5189
rect 1511 -5193 1515 -5189
rect 1519 -5193 1523 -5189
rect 1531 -5193 1535 -5189
rect 1543 -5193 1547 -5189
rect 1552 -5193 1556 -5189
rect 1561 -5193 1565 -5189
rect -1264 -5312 -1260 -5308
rect -1255 -5312 -1251 -5308
rect -1246 -5312 -1242 -5308
rect -1238 -5312 -1234 -5308
rect -1222 -5312 -1218 -5308
rect -1214 -5312 -1210 -5308
rect -1197 -5312 -1193 -5308
rect -1180 -5312 -1176 -5308
rect -1172 -5312 -1168 -5308
rect -1155 -5312 -1151 -5308
rect -1138 -5312 -1134 -5308
rect -1130 -5312 -1126 -5308
rect -1113 -5312 -1109 -5308
rect -1096 -5312 -1092 -5308
rect -1088 -5312 -1084 -5308
rect -1072 -5312 -1068 -5308
rect -935 -5312 -931 -5308
rect -926 -5312 -922 -5308
rect -917 -5312 -913 -5308
rect -909 -5312 -905 -5308
rect -893 -5312 -889 -5308
rect -885 -5312 -881 -5308
rect -868 -5312 -864 -5308
rect -851 -5312 -847 -5308
rect -843 -5312 -839 -5308
rect -826 -5312 -822 -5308
rect -809 -5312 -805 -5308
rect -801 -5312 -797 -5308
rect -784 -5312 -780 -5308
rect -767 -5312 -763 -5308
rect -759 -5312 -755 -5308
rect -743 -5312 -739 -5308
rect -1264 -5433 -1260 -5429
rect -1255 -5433 -1251 -5429
rect -1246 -5433 -1242 -5429
rect -1238 -5433 -1234 -5429
rect -1222 -5433 -1218 -5429
rect -1214 -5433 -1210 -5429
rect -1197 -5433 -1193 -5429
rect -1180 -5433 -1176 -5429
rect -1172 -5433 -1168 -5429
rect -1155 -5433 -1151 -5429
rect -1138 -5433 -1134 -5429
rect -1130 -5433 -1126 -5429
rect -1113 -5433 -1109 -5429
rect -1096 -5433 -1092 -5429
rect -1088 -5433 -1084 -5429
rect -1072 -5433 -1068 -5429
rect -1026 -5433 -1022 -5429
rect -1018 -5433 -1014 -5429
rect -935 -5433 -931 -5429
rect -926 -5433 -922 -5429
rect -917 -5433 -913 -5429
rect -909 -5433 -905 -5429
rect -893 -5433 -889 -5429
rect -885 -5433 -881 -5429
rect -868 -5433 -864 -5429
rect -851 -5433 -847 -5429
rect -843 -5433 -839 -5429
rect -826 -5433 -822 -5429
rect -809 -5433 -805 -5429
rect -801 -5433 -797 -5429
rect -784 -5433 -780 -5429
rect -767 -5433 -763 -5429
rect -759 -5433 -755 -5429
rect -743 -5433 -739 -5429
rect -673 -5433 -669 -5425
rect -665 -5433 -661 -5425
rect -577 -5433 -573 -5429
rect -568 -5433 -564 -5429
rect -559 -5433 -555 -5429
rect -551 -5433 -547 -5429
rect -535 -5433 -531 -5429
rect -527 -5433 -523 -5429
rect -510 -5433 -506 -5429
rect -493 -5433 -489 -5429
rect -485 -5433 -481 -5429
rect -468 -5433 -464 -5429
rect -451 -5433 -447 -5429
rect -443 -5433 -439 -5429
rect -426 -5433 -422 -5429
rect -409 -5433 -405 -5429
rect -401 -5433 -397 -5429
rect -385 -5433 -381 -5429
rect -327 -5433 -323 -5429
rect -319 -5433 -315 -5429
rect -219 -5433 -215 -5429
rect -210 -5433 -206 -5429
rect -201 -5433 -197 -5429
rect -193 -5433 -189 -5429
rect -177 -5433 -173 -5429
rect -169 -5433 -165 -5429
rect -152 -5433 -148 -5429
rect -135 -5433 -131 -5429
rect -127 -5433 -123 -5429
rect -110 -5433 -106 -5429
rect -93 -5433 -89 -5429
rect -85 -5433 -81 -5429
rect -68 -5433 -64 -5429
rect -51 -5433 -47 -5429
rect -43 -5433 -39 -5429
rect -27 -5433 -23 -5429
rect 209 -5433 213 -5429
rect 218 -5433 222 -5429
rect 227 -5433 231 -5429
rect 235 -5433 239 -5429
rect 251 -5433 255 -5429
rect 259 -5433 263 -5429
rect 276 -5433 280 -5429
rect 293 -5433 297 -5429
rect 301 -5433 305 -5429
rect 318 -5433 322 -5429
rect 335 -5433 339 -5429
rect 343 -5433 347 -5429
rect 360 -5433 364 -5429
rect 377 -5433 381 -5429
rect 385 -5433 389 -5429
rect 401 -5433 405 -5429
rect 466 -5433 470 -5429
rect 474 -5433 478 -5429
rect 565 -5433 569 -5429
rect 574 -5433 578 -5429
rect 583 -5433 587 -5429
rect 591 -5433 595 -5429
rect 607 -5433 611 -5429
rect 615 -5433 619 -5429
rect 632 -5433 636 -5429
rect 649 -5433 653 -5429
rect 657 -5433 661 -5429
rect 674 -5433 678 -5429
rect 691 -5433 695 -5429
rect 699 -5433 703 -5429
rect 716 -5433 720 -5429
rect 733 -5433 737 -5429
rect 741 -5433 745 -5429
rect 757 -5433 761 -5429
rect 867 -5433 871 -5425
rect 875 -5433 879 -5425
rect 963 -5433 967 -5429
rect 972 -5433 976 -5429
rect 981 -5433 985 -5429
rect 989 -5433 993 -5429
rect 1005 -5433 1009 -5429
rect 1013 -5433 1017 -5429
rect 1030 -5433 1034 -5429
rect 1047 -5433 1051 -5429
rect 1055 -5433 1059 -5429
rect 1072 -5433 1076 -5429
rect 1089 -5433 1093 -5429
rect 1097 -5433 1101 -5429
rect 1114 -5433 1118 -5429
rect 1131 -5433 1135 -5429
rect 1139 -5433 1143 -5429
rect 1155 -5433 1159 -5429
rect 1210 -5433 1214 -5429
rect 1218 -5433 1222 -5429
rect 1321 -5433 1325 -5429
rect 1330 -5433 1334 -5429
rect 1339 -5433 1343 -5429
rect 1347 -5433 1351 -5429
rect 1363 -5433 1367 -5429
rect 1371 -5433 1375 -5429
rect 1388 -5433 1392 -5429
rect 1405 -5433 1409 -5429
rect 1413 -5433 1417 -5429
rect 1430 -5433 1434 -5429
rect 1447 -5433 1451 -5429
rect 1455 -5433 1459 -5429
rect 1472 -5433 1476 -5429
rect 1489 -5433 1493 -5429
rect 1497 -5433 1501 -5429
rect 1513 -5433 1517 -5429
rect -1264 -5553 -1260 -5549
rect -1255 -5553 -1251 -5549
rect -1246 -5553 -1242 -5549
rect -1238 -5553 -1234 -5549
rect -1222 -5553 -1218 -5549
rect -1214 -5553 -1210 -5549
rect -1197 -5553 -1193 -5549
rect -1180 -5553 -1176 -5549
rect -1172 -5553 -1168 -5549
rect -1155 -5553 -1151 -5549
rect -1138 -5553 -1134 -5549
rect -1130 -5553 -1126 -5549
rect -1113 -5553 -1109 -5549
rect -1096 -5553 -1092 -5549
rect -1088 -5553 -1084 -5549
rect -1072 -5553 -1068 -5549
rect -1026 -5553 -1022 -5549
rect -1018 -5553 -1014 -5549
rect -935 -5553 -931 -5549
rect -926 -5553 -922 -5549
rect -917 -5553 -913 -5549
rect -909 -5553 -905 -5549
rect -893 -5553 -889 -5549
rect -885 -5553 -881 -5549
rect -868 -5553 -864 -5549
rect -851 -5553 -847 -5549
rect -843 -5553 -839 -5549
rect -826 -5553 -822 -5549
rect -809 -5553 -805 -5549
rect -801 -5553 -797 -5549
rect -784 -5553 -780 -5549
rect -767 -5553 -763 -5549
rect -759 -5553 -755 -5549
rect -743 -5553 -739 -5549
rect -577 -5553 -573 -5549
rect -568 -5553 -564 -5549
rect -559 -5553 -555 -5549
rect -551 -5553 -547 -5549
rect -535 -5553 -531 -5549
rect -527 -5553 -523 -5549
rect -510 -5553 -506 -5549
rect -493 -5553 -489 -5549
rect -485 -5553 -481 -5549
rect -468 -5553 -464 -5549
rect -451 -5553 -447 -5549
rect -443 -5553 -439 -5549
rect -426 -5553 -422 -5549
rect -409 -5553 -405 -5549
rect -401 -5553 -397 -5549
rect -385 -5553 -381 -5549
rect -327 -5553 -323 -5549
rect -319 -5553 -315 -5549
rect -219 -5553 -215 -5549
rect -210 -5553 -206 -5549
rect -201 -5553 -197 -5549
rect -193 -5553 -189 -5549
rect -177 -5553 -173 -5549
rect -169 -5553 -165 -5549
rect -152 -5553 -148 -5549
rect -135 -5553 -131 -5549
rect -127 -5553 -123 -5549
rect -110 -5553 -106 -5549
rect -93 -5553 -89 -5549
rect -85 -5553 -81 -5549
rect -68 -5553 -64 -5549
rect -51 -5553 -47 -5549
rect -43 -5553 -39 -5549
rect -27 -5553 -23 -5549
rect 209 -5553 213 -5549
rect 218 -5553 222 -5549
rect 227 -5553 231 -5549
rect 235 -5553 239 -5549
rect 251 -5553 255 -5549
rect 259 -5553 263 -5549
rect 276 -5553 280 -5549
rect 293 -5553 297 -5549
rect 301 -5553 305 -5549
rect 318 -5553 322 -5549
rect 335 -5553 339 -5549
rect 343 -5553 347 -5549
rect 360 -5553 364 -5549
rect 377 -5553 381 -5549
rect 385 -5553 389 -5549
rect 401 -5553 405 -5549
rect 466 -5553 470 -5549
rect 474 -5553 478 -5549
rect 565 -5553 569 -5549
rect 574 -5553 578 -5549
rect 583 -5553 587 -5549
rect 591 -5553 595 -5549
rect 607 -5553 611 -5549
rect 615 -5553 619 -5549
rect 632 -5553 636 -5549
rect 649 -5553 653 -5549
rect 657 -5553 661 -5549
rect 674 -5553 678 -5549
rect 691 -5553 695 -5549
rect 699 -5553 703 -5549
rect 716 -5553 720 -5549
rect 733 -5553 737 -5549
rect 741 -5553 745 -5549
rect 757 -5553 761 -5549
rect 963 -5553 967 -5549
rect 972 -5553 976 -5549
rect 981 -5553 985 -5549
rect 989 -5553 993 -5549
rect 1005 -5553 1009 -5549
rect 1013 -5553 1017 -5549
rect 1030 -5553 1034 -5549
rect 1047 -5553 1051 -5549
rect 1055 -5553 1059 -5549
rect 1072 -5553 1076 -5549
rect 1089 -5553 1093 -5549
rect 1097 -5553 1101 -5549
rect 1114 -5553 1118 -5549
rect 1131 -5553 1135 -5549
rect 1139 -5553 1143 -5549
rect 1155 -5553 1159 -5549
rect 1210 -5553 1214 -5549
rect 1218 -5553 1222 -5549
rect 1321 -5553 1325 -5549
rect 1330 -5553 1334 -5549
rect 1339 -5553 1343 -5549
rect 1347 -5553 1351 -5549
rect 1363 -5553 1367 -5549
rect 1371 -5553 1375 -5549
rect 1388 -5553 1392 -5549
rect 1405 -5553 1409 -5549
rect 1413 -5553 1417 -5549
rect 1430 -5553 1434 -5549
rect 1447 -5553 1451 -5549
rect 1455 -5553 1459 -5549
rect 1472 -5553 1476 -5549
rect 1489 -5553 1493 -5549
rect 1497 -5553 1501 -5549
rect 1513 -5553 1517 -5549
rect -1264 -5670 -1260 -5666
rect -1255 -5670 -1251 -5666
rect -1246 -5670 -1242 -5666
rect -1238 -5670 -1234 -5666
rect -1222 -5670 -1218 -5666
rect -1214 -5670 -1210 -5666
rect -1197 -5670 -1193 -5666
rect -1180 -5670 -1176 -5666
rect -1172 -5670 -1168 -5666
rect -1155 -5670 -1151 -5666
rect -1138 -5670 -1134 -5666
rect -1130 -5670 -1126 -5666
rect -1113 -5670 -1109 -5666
rect -1096 -5670 -1092 -5666
rect -1088 -5670 -1084 -5666
rect -1072 -5670 -1068 -5666
rect -935 -5670 -931 -5666
rect -926 -5670 -922 -5666
rect -917 -5670 -913 -5666
rect -909 -5670 -905 -5666
rect -893 -5670 -889 -5666
rect -885 -5670 -881 -5666
rect -868 -5670 -864 -5666
rect -851 -5670 -847 -5666
rect -843 -5670 -839 -5666
rect -826 -5670 -822 -5666
rect -809 -5670 -805 -5666
rect -801 -5670 -797 -5666
rect -784 -5670 -780 -5666
rect -767 -5670 -763 -5666
rect -759 -5670 -755 -5666
rect -743 -5670 -739 -5666
rect -577 -5670 -573 -5666
rect -568 -5670 -564 -5666
rect -559 -5670 -555 -5666
rect -551 -5670 -547 -5666
rect -535 -5670 -531 -5666
rect -527 -5670 -523 -5666
rect -510 -5670 -506 -5666
rect -493 -5670 -489 -5666
rect -485 -5670 -481 -5666
rect -468 -5670 -464 -5666
rect -451 -5670 -447 -5666
rect -443 -5670 -439 -5666
rect -426 -5670 -422 -5666
rect -409 -5670 -405 -5666
rect -401 -5670 -397 -5666
rect -385 -5670 -381 -5666
rect -219 -5670 -215 -5666
rect -210 -5670 -206 -5666
rect -201 -5670 -197 -5666
rect -193 -5670 -189 -5666
rect -177 -5670 -173 -5666
rect -169 -5670 -165 -5666
rect -152 -5670 -148 -5666
rect -135 -5670 -131 -5666
rect -127 -5670 -123 -5666
rect -110 -5670 -106 -5666
rect -93 -5670 -89 -5666
rect -85 -5670 -81 -5666
rect -68 -5670 -64 -5666
rect -51 -5670 -47 -5666
rect -43 -5670 -39 -5666
rect -27 -5670 -23 -5666
rect 209 -5670 213 -5666
rect 218 -5670 222 -5666
rect 227 -5670 231 -5666
rect 235 -5670 239 -5666
rect 251 -5670 255 -5666
rect 259 -5670 263 -5666
rect 276 -5670 280 -5666
rect 293 -5670 297 -5666
rect 301 -5670 305 -5666
rect 318 -5670 322 -5666
rect 335 -5670 339 -5666
rect 343 -5670 347 -5666
rect 360 -5670 364 -5666
rect 377 -5670 381 -5666
rect 385 -5670 389 -5666
rect 401 -5670 405 -5666
rect 565 -5670 569 -5666
rect 574 -5670 578 -5666
rect 583 -5670 587 -5666
rect 591 -5670 595 -5666
rect 607 -5670 611 -5666
rect 615 -5670 619 -5666
rect 632 -5670 636 -5666
rect 649 -5670 653 -5666
rect 657 -5670 661 -5666
rect 674 -5670 678 -5666
rect 691 -5670 695 -5666
rect 699 -5670 703 -5666
rect 716 -5670 720 -5666
rect 733 -5670 737 -5666
rect 741 -5670 745 -5666
rect 757 -5670 761 -5666
rect -1339 -5787 -1335 -5783
rect -1322 -5787 -1318 -5783
rect -1313 -5787 -1309 -5783
rect -935 -5787 -931 -5783
rect -918 -5787 -914 -5783
rect -909 -5787 -905 -5783
rect -577 -5787 -573 -5783
rect -560 -5787 -556 -5783
rect -551 -5787 -547 -5783
rect -219 -5787 -215 -5783
rect -202 -5787 -198 -5783
rect -193 -5787 -189 -5783
rect 209 -5787 213 -5783
rect 226 -5787 230 -5783
rect 235 -5787 239 -5783
rect 565 -5787 569 -5783
rect 582 -5787 586 -5783
rect 591 -5787 595 -5783
rect 963 -5787 967 -5783
rect 980 -5787 984 -5783
rect 989 -5787 993 -5783
rect 1321 -5787 1325 -5783
rect 1338 -5787 1342 -5783
rect 1347 -5787 1351 -5783
rect -1264 -5906 -1260 -5902
rect -1255 -5906 -1251 -5902
rect -1246 -5906 -1242 -5902
rect -1238 -5906 -1234 -5902
rect -1229 -5906 -1225 -5902
rect -1211 -5906 -1207 -5902
rect -1202 -5906 -1198 -5902
rect -1194 -5906 -1190 -5902
rect -1177 -5906 -1173 -5902
rect -1168 -5906 -1164 -5902
rect -935 -5906 -931 -5902
rect -926 -5906 -922 -5902
rect -917 -5906 -913 -5902
rect -909 -5906 -905 -5902
rect -900 -5906 -896 -5902
rect -891 -5906 -887 -5902
rect -883 -5906 -879 -5902
rect -875 -5906 -871 -5902
rect -857 -5906 -853 -5902
rect -847 -5906 -843 -5902
rect -839 -5906 -835 -5902
rect -822 -5906 -818 -5902
rect -813 -5906 -809 -5902
rect -805 -5906 -801 -5902
rect -796 -5906 -792 -5902
rect -778 -5906 -774 -5902
rect -769 -5906 -765 -5902
rect -761 -5906 -757 -5902
rect -745 -5906 -741 -5902
rect -737 -5906 -733 -5902
rect -725 -5906 -721 -5902
rect -713 -5906 -709 -5902
rect -704 -5906 -700 -5902
rect -695 -5906 -691 -5902
rect -577 -5906 -573 -5902
rect -568 -5906 -564 -5902
rect -559 -5906 -555 -5902
rect -551 -5906 -547 -5902
rect -542 -5906 -538 -5902
rect -533 -5906 -529 -5902
rect -525 -5906 -521 -5902
rect -517 -5906 -513 -5902
rect -499 -5906 -495 -5902
rect -489 -5906 -485 -5902
rect -481 -5906 -477 -5902
rect -464 -5906 -460 -5902
rect -455 -5906 -451 -5902
rect -447 -5906 -443 -5902
rect -438 -5906 -434 -5902
rect -420 -5906 -416 -5902
rect -411 -5906 -407 -5902
rect -403 -5906 -399 -5902
rect -387 -5906 -383 -5902
rect -379 -5906 -375 -5902
rect -367 -5906 -363 -5902
rect -355 -5906 -351 -5902
rect -346 -5906 -342 -5902
rect -337 -5906 -333 -5902
rect -219 -5906 -215 -5902
rect -210 -5906 -206 -5902
rect -201 -5906 -197 -5902
rect -193 -5906 -189 -5902
rect -184 -5906 -180 -5902
rect -175 -5906 -171 -5902
rect -167 -5906 -163 -5902
rect -159 -5906 -155 -5902
rect -141 -5906 -137 -5902
rect -131 -5906 -127 -5902
rect -123 -5906 -119 -5902
rect -106 -5906 -102 -5902
rect -97 -5906 -93 -5902
rect -89 -5906 -85 -5902
rect -80 -5906 -76 -5902
rect -62 -5906 -58 -5902
rect -53 -5906 -49 -5902
rect -45 -5906 -41 -5902
rect -29 -5906 -25 -5902
rect -21 -5906 -17 -5902
rect -9 -5906 -5 -5902
rect 3 -5906 7 -5902
rect 12 -5906 16 -5902
rect 21 -5906 25 -5902
rect 209 -5906 213 -5902
rect 218 -5906 222 -5902
rect 227 -5906 231 -5902
rect 235 -5906 239 -5902
rect 244 -5906 248 -5902
rect 253 -5906 257 -5902
rect 261 -5906 265 -5902
rect 269 -5906 273 -5902
rect 287 -5906 291 -5902
rect 297 -5906 301 -5902
rect 305 -5906 309 -5902
rect 322 -5906 326 -5902
rect 331 -5906 335 -5902
rect 339 -5906 343 -5902
rect 348 -5906 352 -5902
rect 366 -5906 370 -5902
rect 375 -5906 379 -5902
rect 383 -5906 387 -5902
rect 399 -5906 403 -5902
rect 407 -5906 411 -5902
rect 419 -5906 423 -5902
rect 431 -5906 435 -5902
rect 440 -5906 444 -5902
rect 449 -5906 453 -5902
rect 565 -5906 569 -5902
rect 574 -5906 578 -5902
rect 583 -5906 587 -5902
rect 591 -5906 595 -5902
rect 600 -5906 604 -5902
rect 609 -5906 613 -5902
rect 617 -5906 621 -5902
rect 625 -5906 629 -5902
rect 643 -5906 647 -5902
rect 653 -5906 657 -5902
rect 661 -5906 665 -5902
rect 678 -5906 682 -5902
rect 687 -5906 691 -5902
rect 695 -5906 699 -5902
rect 704 -5906 708 -5902
rect 722 -5906 726 -5902
rect 731 -5906 735 -5902
rect 739 -5906 743 -5902
rect 755 -5906 759 -5902
rect 763 -5906 767 -5902
rect 775 -5906 779 -5902
rect 787 -5906 791 -5902
rect 796 -5906 800 -5902
rect 805 -5906 809 -5902
rect 963 -5906 967 -5902
rect 972 -5906 976 -5902
rect 981 -5906 985 -5902
rect 989 -5906 993 -5902
rect 998 -5906 1002 -5902
rect 1007 -5906 1011 -5902
rect 1015 -5906 1019 -5902
rect 1023 -5906 1027 -5902
rect 1041 -5906 1045 -5902
rect 1051 -5906 1055 -5902
rect 1059 -5906 1063 -5902
rect 1076 -5906 1080 -5902
rect 1085 -5906 1089 -5902
rect 1093 -5906 1097 -5902
rect 1102 -5906 1106 -5902
rect 1120 -5906 1124 -5902
rect 1129 -5906 1133 -5902
rect 1137 -5906 1141 -5902
rect 1153 -5906 1157 -5902
rect 1161 -5906 1165 -5902
rect 1173 -5906 1177 -5902
rect 1185 -5906 1189 -5902
rect 1194 -5906 1198 -5902
rect 1203 -5906 1207 -5902
rect 1321 -5906 1325 -5902
rect 1330 -5906 1334 -5902
rect 1339 -5906 1343 -5902
rect 1347 -5906 1351 -5902
rect 1356 -5906 1360 -5902
rect 1365 -5906 1369 -5902
rect 1373 -5906 1377 -5902
rect 1381 -5906 1385 -5902
rect 1399 -5906 1403 -5902
rect 1409 -5906 1413 -5902
rect 1417 -5906 1421 -5902
rect 1434 -5906 1438 -5902
rect 1443 -5906 1447 -5902
rect 1451 -5906 1455 -5902
rect 1460 -5906 1464 -5902
rect 1478 -5906 1482 -5902
rect 1487 -5906 1491 -5902
rect 1495 -5906 1499 -5902
rect 1511 -5906 1515 -5902
rect 1519 -5906 1523 -5902
rect 1531 -5906 1535 -5902
rect 1543 -5906 1547 -5902
rect 1552 -5906 1556 -5902
rect 1561 -5906 1565 -5902
rect -1264 -6029 -1260 -6025
rect -1255 -6029 -1251 -6025
rect -1246 -6029 -1242 -6025
rect -1238 -6029 -1234 -6025
rect -1222 -6029 -1218 -6025
rect -1214 -6029 -1210 -6025
rect -1197 -6029 -1193 -6025
rect -1180 -6029 -1176 -6025
rect -1172 -6029 -1168 -6025
rect -1155 -6029 -1151 -6025
rect -1138 -6029 -1134 -6025
rect -1130 -6029 -1126 -6025
rect -1113 -6029 -1109 -6025
rect -1096 -6029 -1092 -6025
rect -1088 -6029 -1084 -6025
rect -1072 -6029 -1068 -6025
rect -935 -6029 -931 -6025
rect -926 -6029 -922 -6025
rect -917 -6029 -913 -6025
rect -909 -6029 -905 -6025
rect -893 -6029 -889 -6025
rect -885 -6029 -881 -6025
rect -868 -6029 -864 -6025
rect -851 -6029 -847 -6025
rect -843 -6029 -839 -6025
rect -826 -6029 -822 -6025
rect -809 -6029 -805 -6025
rect -801 -6029 -797 -6025
rect -784 -6029 -780 -6025
rect -767 -6029 -763 -6025
rect -759 -6029 -755 -6025
rect -743 -6029 -739 -6025
rect -577 -6029 -573 -6025
rect -568 -6029 -564 -6025
rect -559 -6029 -555 -6025
rect -551 -6029 -547 -6025
rect -535 -6029 -531 -6025
rect -527 -6029 -523 -6025
rect -510 -6029 -506 -6025
rect -493 -6029 -489 -6025
rect -485 -6029 -481 -6025
rect -468 -6029 -464 -6025
rect -451 -6029 -447 -6025
rect -443 -6029 -439 -6025
rect -426 -6029 -422 -6025
rect -409 -6029 -405 -6025
rect -401 -6029 -397 -6025
rect -385 -6029 -381 -6025
rect -219 -6029 -215 -6025
rect -210 -6029 -206 -6025
rect -201 -6029 -197 -6025
rect -193 -6029 -189 -6025
rect -177 -6029 -173 -6025
rect -169 -6029 -165 -6025
rect -152 -6029 -148 -6025
rect -135 -6029 -131 -6025
rect -127 -6029 -123 -6025
rect -110 -6029 -106 -6025
rect -93 -6029 -89 -6025
rect -85 -6029 -81 -6025
rect -68 -6029 -64 -6025
rect -51 -6029 -47 -6025
rect -43 -6029 -39 -6025
rect -27 -6029 -23 -6025
rect 209 -6029 213 -6025
rect 218 -6029 222 -6025
rect 227 -6029 231 -6025
rect 235 -6029 239 -6025
rect 251 -6029 255 -6025
rect 259 -6029 263 -6025
rect 276 -6029 280 -6025
rect 293 -6029 297 -6025
rect 301 -6029 305 -6025
rect 318 -6029 322 -6025
rect 335 -6029 339 -6025
rect 343 -6029 347 -6025
rect 360 -6029 364 -6025
rect 377 -6029 381 -6025
rect 385 -6029 389 -6025
rect 401 -6029 405 -6025
rect 565 -6029 569 -6025
rect 574 -6029 578 -6025
rect 583 -6029 587 -6025
rect 591 -6029 595 -6025
rect 607 -6029 611 -6025
rect 615 -6029 619 -6025
rect 632 -6029 636 -6025
rect 649 -6029 653 -6025
rect 657 -6029 661 -6025
rect 674 -6029 678 -6025
rect 691 -6029 695 -6025
rect 699 -6029 703 -6025
rect 716 -6029 720 -6025
rect 733 -6029 737 -6025
rect 741 -6029 745 -6025
rect 757 -6029 761 -6025
rect 963 -6029 967 -6025
rect 972 -6029 976 -6025
rect 981 -6029 985 -6025
rect 989 -6029 993 -6025
rect 1005 -6029 1009 -6025
rect 1013 -6029 1017 -6025
rect 1030 -6029 1034 -6025
rect 1047 -6029 1051 -6025
rect 1055 -6029 1059 -6025
rect 1072 -6029 1076 -6025
rect 1089 -6029 1093 -6025
rect 1097 -6029 1101 -6025
rect 1114 -6029 1118 -6025
rect 1131 -6029 1135 -6025
rect 1139 -6029 1143 -6025
rect 1155 -6029 1159 -6025
rect 1321 -6029 1325 -6025
rect 1330 -6029 1334 -6025
rect 1339 -6029 1343 -6025
rect 1347 -6029 1351 -6025
rect 1363 -6029 1367 -6025
rect 1371 -6029 1375 -6025
rect 1388 -6029 1392 -6025
rect 1405 -6029 1409 -6025
rect 1413 -6029 1417 -6025
rect 1430 -6029 1434 -6025
rect 1447 -6029 1451 -6025
rect 1455 -6029 1459 -6025
rect 1472 -6029 1476 -6025
rect 1489 -6029 1493 -6025
rect 1497 -6029 1501 -6025
rect 1513 -6029 1517 -6025
rect 1321 -6147 1325 -6143
rect 1330 -6147 1334 -6143
rect 1339 -6147 1343 -6143
rect 1347 -6147 1351 -6143
rect 1363 -6147 1367 -6143
rect 1371 -6147 1375 -6143
rect 1388 -6147 1392 -6143
rect 1405 -6147 1409 -6143
rect 1413 -6147 1417 -6143
rect 1430 -6147 1434 -6143
rect 1447 -6147 1451 -6143
rect 1455 -6147 1459 -6143
rect 1472 -6147 1476 -6143
rect 1489 -6147 1493 -6143
rect 1497 -6147 1501 -6143
rect 1513 -6147 1517 -6143
<< pdcontact >>
rect -1337 -1046 -1333 -1038
rect -1329 -1046 -1325 -1038
rect -1320 -1046 -1316 -1038
rect -1311 -1046 -1307 -1038
rect -936 -1046 -932 -1038
rect -928 -1046 -924 -1038
rect -919 -1046 -915 -1038
rect -910 -1046 -906 -1038
rect -577 -1046 -573 -1038
rect -569 -1046 -565 -1038
rect -560 -1046 -556 -1038
rect -551 -1046 -547 -1038
rect -219 -1046 -215 -1038
rect -211 -1046 -207 -1038
rect -202 -1046 -198 -1038
rect -193 -1046 -189 -1038
rect 209 -1046 213 -1038
rect 217 -1046 221 -1038
rect 226 -1046 230 -1038
rect 235 -1046 239 -1038
rect 565 -1046 569 -1038
rect 573 -1046 577 -1038
rect 582 -1046 586 -1038
rect 591 -1046 595 -1038
rect 963 -1046 967 -1038
rect 971 -1046 975 -1038
rect 980 -1046 984 -1038
rect 989 -1046 993 -1038
rect 1321 -1046 1325 -1038
rect 1329 -1046 1333 -1038
rect 1338 -1046 1342 -1038
rect 1347 -1046 1351 -1038
rect -1260 -1160 -1256 -1152
rect -1251 -1160 -1247 -1152
rect -1242 -1160 -1238 -1152
rect -1234 -1160 -1230 -1152
rect -1226 -1160 -1222 -1152
rect -1214 -1160 -1210 -1152
rect -1202 -1160 -1198 -1152
rect -1193 -1160 -1189 -1152
rect -1184 -1160 -1180 -1152
rect -1172 -1160 -1168 -1152
rect -1160 -1160 -1156 -1152
rect -1151 -1160 -1147 -1152
rect -1142 -1160 -1138 -1152
rect -1130 -1160 -1126 -1152
rect -1118 -1160 -1114 -1152
rect -1109 -1160 -1105 -1152
rect -1100 -1160 -1096 -1152
rect -1088 -1160 -1084 -1152
rect -1076 -1160 -1072 -1152
rect -1068 -1160 -1064 -1152
rect -935 -1160 -931 -1152
rect -926 -1160 -922 -1152
rect -917 -1160 -913 -1152
rect -909 -1160 -905 -1152
rect -901 -1160 -897 -1152
rect -889 -1160 -885 -1152
rect -877 -1160 -873 -1152
rect -868 -1160 -864 -1152
rect -859 -1160 -855 -1152
rect -847 -1160 -843 -1152
rect -835 -1160 -831 -1152
rect -826 -1160 -822 -1152
rect -817 -1160 -813 -1152
rect -805 -1160 -801 -1152
rect -793 -1160 -789 -1152
rect -784 -1160 -780 -1152
rect -775 -1160 -771 -1152
rect -763 -1160 -759 -1152
rect -751 -1160 -747 -1152
rect -743 -1160 -739 -1152
rect -577 -1160 -573 -1152
rect -568 -1160 -564 -1152
rect -559 -1160 -555 -1152
rect -551 -1160 -547 -1152
rect -543 -1160 -539 -1152
rect -531 -1160 -527 -1152
rect -519 -1160 -515 -1152
rect -510 -1160 -506 -1152
rect -501 -1160 -497 -1152
rect -489 -1160 -485 -1152
rect -477 -1160 -473 -1152
rect -468 -1160 -464 -1152
rect -459 -1160 -455 -1152
rect -447 -1160 -443 -1152
rect -435 -1160 -431 -1152
rect -426 -1160 -422 -1152
rect -417 -1160 -413 -1152
rect -405 -1160 -401 -1152
rect -393 -1160 -389 -1152
rect -385 -1160 -381 -1152
rect -219 -1160 -215 -1152
rect -210 -1160 -206 -1152
rect -201 -1160 -197 -1152
rect -193 -1160 -189 -1152
rect -185 -1160 -181 -1152
rect -173 -1160 -169 -1152
rect -161 -1160 -157 -1152
rect -152 -1160 -148 -1152
rect -143 -1160 -139 -1152
rect -131 -1160 -127 -1152
rect -119 -1160 -115 -1152
rect -110 -1160 -106 -1152
rect -101 -1160 -97 -1152
rect -89 -1160 -85 -1152
rect -77 -1160 -73 -1152
rect -68 -1160 -64 -1152
rect -59 -1160 -55 -1152
rect -47 -1160 -43 -1152
rect -35 -1160 -31 -1152
rect -27 -1160 -23 -1152
rect 209 -1160 213 -1152
rect 218 -1160 222 -1152
rect 227 -1160 231 -1152
rect 235 -1160 239 -1152
rect 243 -1160 247 -1152
rect 255 -1160 259 -1152
rect 267 -1160 271 -1152
rect 276 -1160 280 -1152
rect 285 -1160 289 -1152
rect 297 -1160 301 -1152
rect 309 -1160 313 -1152
rect 318 -1160 322 -1152
rect 327 -1160 331 -1152
rect 339 -1160 343 -1152
rect 351 -1160 355 -1152
rect 360 -1160 364 -1152
rect 369 -1160 373 -1152
rect 381 -1160 385 -1152
rect 393 -1160 397 -1152
rect 401 -1160 405 -1152
rect 565 -1160 569 -1152
rect 574 -1160 578 -1152
rect 583 -1160 587 -1152
rect 591 -1160 595 -1152
rect 599 -1160 603 -1152
rect 611 -1160 615 -1152
rect 623 -1160 627 -1152
rect 632 -1160 636 -1152
rect 641 -1160 645 -1152
rect 653 -1160 657 -1152
rect 665 -1160 669 -1152
rect 674 -1160 678 -1152
rect 683 -1160 687 -1152
rect 695 -1160 699 -1152
rect 707 -1160 711 -1152
rect 716 -1160 720 -1152
rect 725 -1160 729 -1152
rect 737 -1160 741 -1152
rect 749 -1160 753 -1152
rect 757 -1160 761 -1152
rect 963 -1160 967 -1152
rect 972 -1160 976 -1152
rect 981 -1160 985 -1152
rect 989 -1160 993 -1152
rect 997 -1160 1001 -1152
rect 1009 -1160 1013 -1152
rect 1021 -1160 1025 -1152
rect 1030 -1160 1034 -1152
rect 1039 -1160 1043 -1152
rect 1051 -1160 1055 -1152
rect 1063 -1160 1067 -1152
rect 1072 -1160 1076 -1152
rect 1081 -1160 1085 -1152
rect 1093 -1160 1097 -1152
rect 1105 -1160 1109 -1152
rect 1114 -1160 1118 -1152
rect 1123 -1160 1127 -1152
rect 1135 -1160 1139 -1152
rect 1147 -1160 1151 -1152
rect 1155 -1160 1159 -1152
rect -1339 -1276 -1335 -1268
rect -1331 -1276 -1327 -1268
rect -1322 -1276 -1318 -1268
rect -1313 -1276 -1309 -1268
rect -935 -1276 -931 -1268
rect -927 -1276 -923 -1268
rect -918 -1276 -914 -1268
rect -909 -1276 -905 -1268
rect -577 -1276 -573 -1268
rect -569 -1276 -565 -1268
rect -560 -1276 -556 -1268
rect -551 -1276 -547 -1268
rect -219 -1276 -215 -1268
rect -211 -1276 -207 -1268
rect -202 -1276 -198 -1268
rect -193 -1276 -189 -1268
rect 209 -1276 213 -1268
rect 217 -1276 221 -1268
rect 226 -1276 230 -1268
rect 235 -1276 239 -1268
rect 565 -1276 569 -1268
rect 573 -1276 577 -1268
rect 582 -1276 586 -1268
rect 591 -1276 595 -1268
rect 963 -1276 967 -1268
rect 971 -1276 975 -1268
rect 980 -1276 984 -1268
rect 989 -1276 993 -1268
rect 1321 -1276 1325 -1268
rect 1329 -1276 1333 -1268
rect 1338 -1276 1342 -1268
rect 1347 -1276 1351 -1268
rect -1260 -1390 -1256 -1382
rect -1251 -1390 -1247 -1382
rect -1242 -1390 -1238 -1382
rect -1234 -1390 -1230 -1382
rect -1216 -1390 -1212 -1382
rect -1194 -1390 -1190 -1382
rect -1182 -1390 -1178 -1382
rect -1173 -1390 -1169 -1382
rect -1164 -1390 -1160 -1382
rect -935 -1390 -931 -1382
rect -926 -1390 -922 -1382
rect -917 -1390 -913 -1382
rect -909 -1390 -905 -1382
rect -900 -1390 -896 -1382
rect -891 -1390 -887 -1382
rect -883 -1390 -879 -1382
rect -865 -1390 -861 -1382
rect -843 -1390 -839 -1382
rect -831 -1390 -827 -1382
rect -822 -1390 -818 -1382
rect -813 -1390 -809 -1382
rect -805 -1390 -801 -1382
rect -787 -1390 -783 -1382
rect -765 -1390 -761 -1382
rect -753 -1390 -749 -1382
rect -741 -1390 -737 -1382
rect -729 -1390 -725 -1382
rect -721 -1390 -717 -1382
rect -704 -1390 -700 -1382
rect -695 -1390 -691 -1382
rect -577 -1390 -573 -1382
rect -568 -1390 -564 -1382
rect -559 -1390 -555 -1382
rect -551 -1390 -547 -1382
rect -542 -1390 -538 -1382
rect -533 -1390 -529 -1382
rect -525 -1390 -521 -1382
rect -507 -1390 -503 -1382
rect -485 -1390 -481 -1382
rect -473 -1390 -469 -1382
rect -464 -1390 -460 -1382
rect -455 -1390 -451 -1382
rect -447 -1390 -443 -1382
rect -429 -1390 -425 -1382
rect -407 -1390 -403 -1382
rect -395 -1390 -391 -1382
rect -383 -1390 -379 -1382
rect -371 -1390 -367 -1382
rect -363 -1390 -359 -1382
rect -346 -1390 -342 -1382
rect -337 -1390 -333 -1382
rect -219 -1390 -215 -1382
rect -210 -1390 -206 -1382
rect -201 -1390 -197 -1382
rect -193 -1390 -189 -1382
rect -184 -1390 -180 -1382
rect -175 -1390 -171 -1382
rect -167 -1390 -163 -1382
rect -149 -1390 -145 -1382
rect -127 -1390 -123 -1382
rect -115 -1390 -111 -1382
rect -106 -1390 -102 -1382
rect -97 -1390 -93 -1382
rect -89 -1390 -85 -1382
rect -71 -1390 -67 -1382
rect -49 -1390 -45 -1382
rect -37 -1390 -33 -1382
rect -25 -1390 -21 -1382
rect -13 -1390 -9 -1382
rect -5 -1390 -1 -1382
rect 12 -1390 16 -1382
rect 21 -1390 25 -1382
rect 209 -1390 213 -1382
rect 218 -1390 222 -1382
rect 227 -1390 231 -1382
rect 235 -1390 239 -1382
rect 244 -1390 248 -1382
rect 253 -1390 257 -1382
rect 261 -1390 265 -1382
rect 279 -1390 283 -1382
rect 301 -1390 305 -1382
rect 313 -1390 317 -1382
rect 322 -1390 326 -1382
rect 331 -1390 335 -1382
rect 339 -1390 343 -1382
rect 357 -1390 361 -1382
rect 379 -1390 383 -1382
rect 391 -1390 395 -1382
rect 403 -1390 407 -1382
rect 415 -1390 419 -1382
rect 423 -1390 427 -1382
rect 440 -1390 444 -1382
rect 449 -1390 453 -1382
rect 565 -1390 569 -1382
rect 574 -1390 578 -1382
rect 583 -1390 587 -1382
rect 591 -1390 595 -1382
rect 600 -1390 604 -1382
rect 609 -1390 613 -1382
rect 617 -1390 621 -1382
rect 635 -1390 639 -1382
rect 657 -1390 661 -1382
rect 669 -1390 673 -1382
rect 678 -1390 682 -1382
rect 687 -1390 691 -1382
rect 695 -1390 699 -1382
rect 713 -1390 717 -1382
rect 735 -1390 739 -1382
rect 747 -1390 751 -1382
rect 759 -1390 763 -1382
rect 771 -1390 775 -1382
rect 779 -1390 783 -1382
rect 796 -1390 800 -1382
rect 805 -1390 809 -1382
rect 963 -1390 967 -1382
rect 972 -1390 976 -1382
rect 981 -1390 985 -1382
rect 989 -1390 993 -1382
rect 998 -1390 1002 -1382
rect 1007 -1390 1011 -1382
rect 1015 -1390 1019 -1382
rect 1033 -1390 1037 -1382
rect 1055 -1390 1059 -1382
rect 1067 -1390 1071 -1382
rect 1076 -1390 1080 -1382
rect 1085 -1390 1089 -1382
rect 1093 -1390 1097 -1382
rect 1111 -1390 1115 -1382
rect 1133 -1390 1137 -1382
rect 1145 -1390 1149 -1382
rect 1157 -1390 1161 -1382
rect 1169 -1390 1173 -1382
rect 1177 -1390 1181 -1382
rect 1194 -1390 1198 -1382
rect 1203 -1390 1207 -1382
rect 1321 -1390 1325 -1382
rect 1330 -1390 1334 -1382
rect 1339 -1390 1343 -1382
rect 1347 -1390 1351 -1382
rect 1365 -1390 1369 -1382
rect 1387 -1390 1391 -1382
rect 1399 -1390 1403 -1382
rect 1408 -1390 1412 -1382
rect 1417 -1390 1421 -1382
rect -1260 -1513 -1256 -1505
rect -1251 -1513 -1247 -1505
rect -1242 -1513 -1238 -1505
rect -1234 -1513 -1230 -1505
rect -1226 -1513 -1222 -1505
rect -1214 -1513 -1210 -1505
rect -1202 -1513 -1198 -1505
rect -1193 -1513 -1189 -1505
rect -1184 -1513 -1180 -1505
rect -1172 -1513 -1168 -1505
rect -1160 -1513 -1156 -1505
rect -1151 -1513 -1147 -1505
rect -1142 -1513 -1138 -1505
rect -1130 -1513 -1126 -1505
rect -1118 -1513 -1114 -1505
rect -1109 -1513 -1105 -1505
rect -1100 -1513 -1096 -1505
rect -1088 -1513 -1084 -1505
rect -1076 -1513 -1072 -1505
rect -1068 -1513 -1064 -1505
rect -935 -1513 -931 -1505
rect -926 -1513 -922 -1505
rect -917 -1513 -913 -1505
rect -909 -1513 -905 -1505
rect -901 -1513 -897 -1505
rect -889 -1513 -885 -1505
rect -877 -1513 -873 -1505
rect -868 -1513 -864 -1505
rect -859 -1513 -855 -1505
rect -847 -1513 -843 -1505
rect -835 -1513 -831 -1505
rect -826 -1513 -822 -1505
rect -817 -1513 -813 -1505
rect -805 -1513 -801 -1505
rect -793 -1513 -789 -1505
rect -784 -1513 -780 -1505
rect -775 -1513 -771 -1505
rect -763 -1513 -759 -1505
rect -751 -1513 -747 -1505
rect -743 -1513 -739 -1505
rect -577 -1513 -573 -1505
rect -568 -1513 -564 -1505
rect -559 -1513 -555 -1505
rect -551 -1513 -547 -1505
rect -543 -1513 -539 -1505
rect -531 -1513 -527 -1505
rect -519 -1513 -515 -1505
rect -510 -1513 -506 -1505
rect -501 -1513 -497 -1505
rect -489 -1513 -485 -1505
rect -477 -1513 -473 -1505
rect -468 -1513 -464 -1505
rect -459 -1513 -455 -1505
rect -447 -1513 -443 -1505
rect -435 -1513 -431 -1505
rect -426 -1513 -422 -1505
rect -417 -1513 -413 -1505
rect -405 -1513 -401 -1505
rect -393 -1513 -389 -1505
rect -385 -1513 -381 -1505
rect -219 -1513 -215 -1505
rect -210 -1513 -206 -1505
rect -201 -1513 -197 -1505
rect -193 -1513 -189 -1505
rect -185 -1513 -181 -1505
rect -173 -1513 -169 -1505
rect -161 -1513 -157 -1505
rect -152 -1513 -148 -1505
rect -143 -1513 -139 -1505
rect -131 -1513 -127 -1505
rect -119 -1513 -115 -1505
rect -110 -1513 -106 -1505
rect -101 -1513 -97 -1505
rect -89 -1513 -85 -1505
rect -77 -1513 -73 -1505
rect -68 -1513 -64 -1505
rect -59 -1513 -55 -1505
rect -47 -1513 -43 -1505
rect -35 -1513 -31 -1505
rect -27 -1513 -23 -1505
rect 209 -1513 213 -1505
rect 218 -1513 222 -1505
rect 227 -1513 231 -1505
rect 235 -1513 239 -1505
rect 243 -1513 247 -1505
rect 255 -1513 259 -1505
rect 267 -1513 271 -1505
rect 276 -1513 280 -1505
rect 285 -1513 289 -1505
rect 297 -1513 301 -1505
rect 309 -1513 313 -1505
rect 318 -1513 322 -1505
rect 327 -1513 331 -1505
rect 339 -1513 343 -1505
rect 351 -1513 355 -1505
rect 360 -1513 364 -1505
rect 369 -1513 373 -1505
rect 381 -1513 385 -1505
rect 393 -1513 397 -1505
rect 401 -1513 405 -1505
rect 565 -1513 569 -1505
rect 574 -1513 578 -1505
rect 583 -1513 587 -1505
rect 591 -1513 595 -1505
rect 599 -1513 603 -1505
rect 611 -1513 615 -1505
rect 623 -1513 627 -1505
rect 632 -1513 636 -1505
rect 641 -1513 645 -1505
rect 653 -1513 657 -1505
rect 665 -1513 669 -1505
rect 674 -1513 678 -1505
rect 683 -1513 687 -1505
rect 695 -1513 699 -1505
rect 707 -1513 711 -1505
rect 716 -1513 720 -1505
rect 725 -1513 729 -1505
rect 737 -1513 741 -1505
rect 749 -1513 753 -1505
rect 757 -1513 761 -1505
rect 963 -1513 967 -1505
rect 972 -1513 976 -1505
rect 981 -1513 985 -1505
rect 989 -1513 993 -1505
rect 997 -1513 1001 -1505
rect 1009 -1513 1013 -1505
rect 1021 -1513 1025 -1505
rect 1030 -1513 1034 -1505
rect 1039 -1513 1043 -1505
rect 1051 -1513 1055 -1505
rect 1063 -1513 1067 -1505
rect 1072 -1513 1076 -1505
rect 1081 -1513 1085 -1505
rect 1093 -1513 1097 -1505
rect 1105 -1513 1109 -1505
rect 1114 -1513 1118 -1505
rect 1123 -1513 1127 -1505
rect 1135 -1513 1139 -1505
rect 1147 -1513 1151 -1505
rect 1155 -1513 1159 -1505
rect -1260 -1634 -1256 -1626
rect -1251 -1634 -1247 -1626
rect -1242 -1634 -1238 -1626
rect -1234 -1634 -1230 -1626
rect -1226 -1634 -1222 -1626
rect -1214 -1634 -1210 -1626
rect -1202 -1634 -1198 -1626
rect -1193 -1634 -1189 -1626
rect -1184 -1634 -1180 -1626
rect -1172 -1634 -1168 -1626
rect -1160 -1634 -1156 -1626
rect -1151 -1634 -1147 -1626
rect -1142 -1634 -1138 -1626
rect -1130 -1634 -1126 -1626
rect -1118 -1634 -1114 -1626
rect -1109 -1634 -1105 -1626
rect -1100 -1634 -1096 -1626
rect -1088 -1634 -1084 -1626
rect -1076 -1634 -1072 -1626
rect -1068 -1634 -1064 -1626
rect -935 -1634 -931 -1626
rect -926 -1634 -922 -1626
rect -917 -1634 -913 -1626
rect -909 -1634 -905 -1626
rect -901 -1634 -897 -1626
rect -889 -1634 -885 -1626
rect -877 -1634 -873 -1626
rect -868 -1634 -864 -1626
rect -859 -1634 -855 -1626
rect -847 -1634 -843 -1626
rect -835 -1634 -831 -1626
rect -826 -1634 -822 -1626
rect -817 -1634 -813 -1626
rect -805 -1634 -801 -1626
rect -793 -1634 -789 -1626
rect -784 -1634 -780 -1626
rect -775 -1634 -771 -1626
rect -763 -1634 -759 -1626
rect -751 -1634 -747 -1626
rect -743 -1634 -739 -1626
rect -577 -1634 -573 -1626
rect -568 -1634 -564 -1626
rect -559 -1634 -555 -1626
rect -551 -1634 -547 -1626
rect -543 -1634 -539 -1626
rect -531 -1634 -527 -1626
rect -519 -1634 -515 -1626
rect -510 -1634 -506 -1626
rect -501 -1634 -497 -1626
rect -489 -1634 -485 -1626
rect -477 -1634 -473 -1626
rect -468 -1634 -464 -1626
rect -459 -1634 -455 -1626
rect -447 -1634 -443 -1626
rect -435 -1634 -431 -1626
rect -426 -1634 -422 -1626
rect -417 -1634 -413 -1626
rect -405 -1634 -401 -1626
rect -393 -1634 -389 -1626
rect -385 -1634 -381 -1626
rect -219 -1634 -215 -1626
rect -210 -1634 -206 -1626
rect -201 -1634 -197 -1626
rect -193 -1634 -189 -1626
rect -185 -1634 -181 -1626
rect -173 -1634 -169 -1626
rect -161 -1634 -157 -1626
rect -152 -1634 -148 -1626
rect -143 -1634 -139 -1626
rect -131 -1634 -127 -1626
rect -119 -1634 -115 -1626
rect -110 -1634 -106 -1626
rect -101 -1634 -97 -1626
rect -89 -1634 -85 -1626
rect -77 -1634 -73 -1626
rect -68 -1634 -64 -1626
rect -59 -1634 -55 -1626
rect -47 -1634 -43 -1626
rect -35 -1634 -31 -1626
rect -27 -1634 -23 -1626
rect 209 -1634 213 -1626
rect 218 -1634 222 -1626
rect 227 -1634 231 -1626
rect 235 -1634 239 -1626
rect 243 -1634 247 -1626
rect 255 -1634 259 -1626
rect 267 -1634 271 -1626
rect 276 -1634 280 -1626
rect 285 -1634 289 -1626
rect 297 -1634 301 -1626
rect 309 -1634 313 -1626
rect 318 -1634 322 -1626
rect 327 -1634 331 -1626
rect 339 -1634 343 -1626
rect 351 -1634 355 -1626
rect 360 -1634 364 -1626
rect 369 -1634 373 -1626
rect 381 -1634 385 -1626
rect 393 -1634 397 -1626
rect 401 -1634 405 -1626
rect 565 -1634 569 -1626
rect 574 -1634 578 -1626
rect 583 -1634 587 -1626
rect 591 -1634 595 -1626
rect 599 -1634 603 -1626
rect 611 -1634 615 -1626
rect 623 -1634 627 -1626
rect 632 -1634 636 -1626
rect 641 -1634 645 -1626
rect 653 -1634 657 -1626
rect 665 -1634 669 -1626
rect 674 -1634 678 -1626
rect 683 -1634 687 -1626
rect 695 -1634 699 -1626
rect 707 -1634 711 -1626
rect 716 -1634 720 -1626
rect 725 -1634 729 -1626
rect 737 -1634 741 -1626
rect 749 -1634 753 -1626
rect 757 -1634 761 -1626
rect 963 -1634 967 -1626
rect 972 -1634 976 -1626
rect 981 -1634 985 -1626
rect 989 -1634 993 -1626
rect 997 -1634 1001 -1626
rect 1009 -1634 1013 -1626
rect 1021 -1634 1025 -1626
rect 1030 -1634 1034 -1626
rect 1039 -1634 1043 -1626
rect 1051 -1634 1055 -1626
rect 1063 -1634 1067 -1626
rect 1072 -1634 1076 -1626
rect 1081 -1634 1085 -1626
rect 1093 -1634 1097 -1626
rect 1105 -1634 1109 -1626
rect 1114 -1634 1118 -1626
rect 1123 -1634 1127 -1626
rect 1135 -1634 1139 -1626
rect 1147 -1634 1151 -1626
rect 1155 -1634 1159 -1626
rect 1321 -1634 1325 -1626
rect 1330 -1634 1334 -1626
rect 1339 -1634 1343 -1626
rect 1347 -1634 1351 -1626
rect 1355 -1634 1359 -1626
rect 1367 -1634 1371 -1626
rect 1379 -1634 1383 -1626
rect 1388 -1634 1392 -1626
rect 1397 -1634 1401 -1626
rect 1409 -1634 1413 -1626
rect 1421 -1634 1425 -1626
rect 1430 -1634 1434 -1626
rect 1439 -1634 1443 -1626
rect 1451 -1634 1455 -1626
rect 1463 -1634 1467 -1626
rect 1472 -1634 1476 -1626
rect 1481 -1634 1485 -1626
rect 1493 -1634 1497 -1626
rect 1505 -1634 1509 -1626
rect 1513 -1634 1517 -1626
rect -1260 -1755 -1256 -1747
rect -1251 -1755 -1247 -1747
rect -1242 -1755 -1238 -1747
rect -1234 -1755 -1230 -1747
rect -1226 -1755 -1222 -1747
rect -1214 -1755 -1210 -1747
rect -1202 -1755 -1198 -1747
rect -1193 -1755 -1189 -1747
rect -1184 -1755 -1180 -1747
rect -1172 -1755 -1168 -1747
rect -1160 -1755 -1156 -1747
rect -1151 -1755 -1147 -1747
rect -1142 -1755 -1138 -1747
rect -1130 -1755 -1126 -1747
rect -1118 -1755 -1114 -1747
rect -1109 -1755 -1105 -1747
rect -1100 -1755 -1096 -1747
rect -1088 -1755 -1084 -1747
rect -1076 -1755 -1072 -1747
rect -1068 -1755 -1064 -1747
rect -1029 -1755 -1025 -1747
rect -1021 -1755 -1017 -1747
rect -935 -1755 -931 -1747
rect -926 -1755 -922 -1747
rect -917 -1755 -913 -1747
rect -909 -1755 -905 -1747
rect -901 -1755 -897 -1747
rect -889 -1755 -885 -1747
rect -877 -1755 -873 -1747
rect -868 -1755 -864 -1747
rect -859 -1755 -855 -1747
rect -847 -1755 -843 -1747
rect -835 -1755 -831 -1747
rect -826 -1755 -822 -1747
rect -817 -1755 -813 -1747
rect -805 -1755 -801 -1747
rect -793 -1755 -789 -1747
rect -784 -1755 -780 -1747
rect -775 -1755 -771 -1747
rect -763 -1755 -759 -1747
rect -751 -1755 -747 -1747
rect -743 -1755 -739 -1747
rect -577 -1755 -573 -1747
rect -568 -1755 -564 -1747
rect -559 -1755 -555 -1747
rect -551 -1755 -547 -1747
rect -543 -1755 -539 -1747
rect -531 -1755 -527 -1747
rect -519 -1755 -515 -1747
rect -510 -1755 -506 -1747
rect -501 -1755 -497 -1747
rect -489 -1755 -485 -1747
rect -477 -1755 -473 -1747
rect -468 -1755 -464 -1747
rect -459 -1755 -455 -1747
rect -447 -1755 -443 -1747
rect -435 -1755 -431 -1747
rect -426 -1755 -422 -1747
rect -417 -1755 -413 -1747
rect -405 -1755 -401 -1747
rect -393 -1755 -389 -1747
rect -385 -1755 -381 -1747
rect -332 -1755 -328 -1747
rect -324 -1755 -320 -1747
rect -219 -1755 -215 -1747
rect -210 -1755 -206 -1747
rect -201 -1755 -197 -1747
rect -193 -1755 -189 -1747
rect -185 -1755 -181 -1747
rect -173 -1755 -169 -1747
rect -161 -1755 -157 -1747
rect -152 -1755 -148 -1747
rect -143 -1755 -139 -1747
rect -131 -1755 -127 -1747
rect -119 -1755 -115 -1747
rect -110 -1755 -106 -1747
rect -101 -1755 -97 -1747
rect -89 -1755 -85 -1747
rect -77 -1755 -73 -1747
rect -68 -1755 -64 -1747
rect -59 -1755 -55 -1747
rect -47 -1755 -43 -1747
rect -35 -1755 -31 -1747
rect -27 -1755 -23 -1747
rect 209 -1755 213 -1747
rect 218 -1755 222 -1747
rect 227 -1755 231 -1747
rect 235 -1755 239 -1747
rect 243 -1755 247 -1747
rect 255 -1755 259 -1747
rect 267 -1755 271 -1747
rect 276 -1755 280 -1747
rect 285 -1755 289 -1747
rect 297 -1755 301 -1747
rect 309 -1755 313 -1747
rect 318 -1755 322 -1747
rect 327 -1755 331 -1747
rect 339 -1755 343 -1747
rect 351 -1755 355 -1747
rect 360 -1755 364 -1747
rect 369 -1755 373 -1747
rect 381 -1755 385 -1747
rect 393 -1755 397 -1747
rect 401 -1755 405 -1747
rect 464 -1755 468 -1747
rect 472 -1755 476 -1747
rect 565 -1755 569 -1747
rect 574 -1755 578 -1747
rect 583 -1755 587 -1747
rect 591 -1755 595 -1747
rect 599 -1755 603 -1747
rect 611 -1755 615 -1747
rect 623 -1755 627 -1747
rect 632 -1755 636 -1747
rect 641 -1755 645 -1747
rect 653 -1755 657 -1747
rect 665 -1755 669 -1747
rect 674 -1755 678 -1747
rect 683 -1755 687 -1747
rect 695 -1755 699 -1747
rect 707 -1755 711 -1747
rect 716 -1755 720 -1747
rect 725 -1755 729 -1747
rect 737 -1755 741 -1747
rect 749 -1755 753 -1747
rect 757 -1755 761 -1747
rect 963 -1755 967 -1747
rect 972 -1755 976 -1747
rect 981 -1755 985 -1747
rect 989 -1755 993 -1747
rect 997 -1755 1001 -1747
rect 1009 -1755 1013 -1747
rect 1021 -1755 1025 -1747
rect 1030 -1755 1034 -1747
rect 1039 -1755 1043 -1747
rect 1051 -1755 1055 -1747
rect 1063 -1755 1067 -1747
rect 1072 -1755 1076 -1747
rect 1081 -1755 1085 -1747
rect 1093 -1755 1097 -1747
rect 1105 -1755 1109 -1747
rect 1114 -1755 1118 -1747
rect 1123 -1755 1127 -1747
rect 1135 -1755 1139 -1747
rect 1147 -1755 1151 -1747
rect 1155 -1755 1159 -1747
rect 1203 -1755 1207 -1747
rect 1211 -1755 1215 -1747
rect 1321 -1755 1325 -1747
rect 1330 -1755 1334 -1747
rect 1339 -1755 1343 -1747
rect 1347 -1755 1351 -1747
rect 1355 -1755 1359 -1747
rect 1367 -1755 1371 -1747
rect 1379 -1755 1383 -1747
rect 1388 -1755 1392 -1747
rect 1397 -1755 1401 -1747
rect 1409 -1755 1413 -1747
rect 1421 -1755 1425 -1747
rect 1430 -1755 1434 -1747
rect 1439 -1755 1443 -1747
rect 1451 -1755 1455 -1747
rect 1463 -1755 1467 -1747
rect 1472 -1755 1476 -1747
rect 1481 -1755 1485 -1747
rect 1493 -1755 1497 -1747
rect 1505 -1755 1509 -1747
rect 1513 -1755 1517 -1747
rect -1260 -1870 -1256 -1862
rect -1251 -1870 -1247 -1862
rect -1242 -1870 -1238 -1862
rect -1234 -1870 -1230 -1862
rect -1226 -1870 -1222 -1862
rect -1214 -1870 -1210 -1862
rect -1202 -1870 -1198 -1862
rect -1193 -1870 -1189 -1862
rect -1184 -1870 -1180 -1862
rect -1172 -1870 -1168 -1862
rect -1160 -1870 -1156 -1862
rect -1151 -1870 -1147 -1862
rect -1142 -1870 -1138 -1862
rect -1130 -1870 -1126 -1862
rect -1118 -1870 -1114 -1862
rect -1109 -1870 -1105 -1862
rect -1100 -1870 -1096 -1862
rect -1088 -1870 -1084 -1862
rect -1076 -1870 -1072 -1862
rect -1068 -1870 -1064 -1862
rect -1029 -1870 -1025 -1862
rect -1021 -1870 -1017 -1862
rect -673 -1878 -669 -1862
rect -665 -1878 -661 -1862
rect -332 -1870 -328 -1862
rect -324 -1870 -320 -1862
rect 464 -1870 468 -1862
rect 472 -1870 476 -1862
rect 841 -1878 845 -1862
rect 849 -1878 853 -1862
rect 1203 -1870 1207 -1862
rect 1211 -1870 1215 -1862
rect -1339 -1982 -1335 -1974
rect -1331 -1982 -1327 -1974
rect -1322 -1982 -1318 -1974
rect -1313 -1982 -1309 -1974
rect -935 -1982 -931 -1974
rect -927 -1982 -923 -1974
rect -918 -1982 -914 -1974
rect -909 -1982 -905 -1974
rect -577 -1982 -573 -1974
rect -569 -1982 -565 -1974
rect -560 -1982 -556 -1974
rect -551 -1982 -547 -1974
rect -219 -1982 -215 -1974
rect -211 -1982 -207 -1974
rect -202 -1982 -198 -1974
rect -193 -1982 -189 -1974
rect 209 -1982 213 -1974
rect 217 -1982 221 -1974
rect 226 -1982 230 -1974
rect 235 -1982 239 -1974
rect 565 -1982 569 -1974
rect 573 -1982 577 -1974
rect 582 -1982 586 -1974
rect 591 -1982 595 -1974
rect 963 -1982 967 -1974
rect 971 -1982 975 -1974
rect 980 -1982 984 -1974
rect 989 -1982 993 -1974
rect 1321 -1982 1325 -1974
rect 1329 -1982 1333 -1974
rect 1338 -1982 1342 -1974
rect 1347 -1982 1351 -1974
rect -1260 -2101 -1256 -2093
rect -1251 -2101 -1247 -2093
rect -1242 -2101 -1238 -2093
rect -1234 -2101 -1230 -2093
rect -1216 -2101 -1212 -2093
rect -1194 -2101 -1190 -2093
rect -1182 -2101 -1178 -2093
rect -1173 -2101 -1169 -2093
rect -1164 -2101 -1160 -2093
rect -935 -2101 -931 -2093
rect -926 -2101 -922 -2093
rect -917 -2101 -913 -2093
rect -909 -2101 -905 -2093
rect -900 -2101 -896 -2093
rect -891 -2101 -887 -2093
rect -883 -2101 -879 -2093
rect -865 -2101 -861 -2093
rect -843 -2101 -839 -2093
rect -831 -2101 -827 -2093
rect -822 -2101 -818 -2093
rect -813 -2101 -809 -2093
rect -805 -2101 -801 -2093
rect -787 -2101 -783 -2093
rect -765 -2101 -761 -2093
rect -753 -2101 -749 -2093
rect -741 -2101 -737 -2093
rect -729 -2101 -725 -2093
rect -721 -2101 -717 -2093
rect -704 -2101 -700 -2093
rect -695 -2101 -691 -2093
rect -577 -2101 -573 -2093
rect -568 -2101 -564 -2093
rect -559 -2101 -555 -2093
rect -551 -2101 -547 -2093
rect -542 -2101 -538 -2093
rect -533 -2101 -529 -2093
rect -525 -2101 -521 -2093
rect -507 -2101 -503 -2093
rect -485 -2101 -481 -2093
rect -473 -2101 -469 -2093
rect -464 -2101 -460 -2093
rect -455 -2101 -451 -2093
rect -447 -2101 -443 -2093
rect -429 -2101 -425 -2093
rect -407 -2101 -403 -2093
rect -395 -2101 -391 -2093
rect -383 -2101 -379 -2093
rect -371 -2101 -367 -2093
rect -363 -2101 -359 -2093
rect -346 -2101 -342 -2093
rect -337 -2101 -333 -2093
rect -219 -2101 -215 -2093
rect -210 -2101 -206 -2093
rect -201 -2101 -197 -2093
rect -193 -2101 -189 -2093
rect -184 -2101 -180 -2093
rect -175 -2101 -171 -2093
rect -167 -2101 -163 -2093
rect -149 -2101 -145 -2093
rect -127 -2101 -123 -2093
rect -115 -2101 -111 -2093
rect -106 -2101 -102 -2093
rect -97 -2101 -93 -2093
rect -89 -2101 -85 -2093
rect -71 -2101 -67 -2093
rect -49 -2101 -45 -2093
rect -37 -2101 -33 -2093
rect -25 -2101 -21 -2093
rect -13 -2101 -9 -2093
rect -5 -2101 -1 -2093
rect 12 -2101 16 -2093
rect 21 -2101 25 -2093
rect 209 -2101 213 -2093
rect 218 -2101 222 -2093
rect 227 -2101 231 -2093
rect 235 -2101 239 -2093
rect 244 -2101 248 -2093
rect 253 -2101 257 -2093
rect 261 -2101 265 -2093
rect 279 -2101 283 -2093
rect 301 -2101 305 -2093
rect 313 -2101 317 -2093
rect 322 -2101 326 -2093
rect 331 -2101 335 -2093
rect 339 -2101 343 -2093
rect 357 -2101 361 -2093
rect 379 -2101 383 -2093
rect 391 -2101 395 -2093
rect 403 -2101 407 -2093
rect 415 -2101 419 -2093
rect 423 -2101 427 -2093
rect 440 -2101 444 -2093
rect 449 -2101 453 -2093
rect 565 -2101 569 -2093
rect 574 -2101 578 -2093
rect 583 -2101 587 -2093
rect 591 -2101 595 -2093
rect 600 -2101 604 -2093
rect 609 -2101 613 -2093
rect 617 -2101 621 -2093
rect 635 -2101 639 -2093
rect 657 -2101 661 -2093
rect 669 -2101 673 -2093
rect 678 -2101 682 -2093
rect 687 -2101 691 -2093
rect 695 -2101 699 -2093
rect 713 -2101 717 -2093
rect 735 -2101 739 -2093
rect 747 -2101 751 -2093
rect 759 -2101 763 -2093
rect 771 -2101 775 -2093
rect 779 -2101 783 -2093
rect 796 -2101 800 -2093
rect 805 -2101 809 -2093
rect 963 -2101 967 -2093
rect 972 -2101 976 -2093
rect 981 -2101 985 -2093
rect 989 -2101 993 -2093
rect 998 -2101 1002 -2093
rect 1007 -2101 1011 -2093
rect 1015 -2101 1019 -2093
rect 1033 -2101 1037 -2093
rect 1055 -2101 1059 -2093
rect 1067 -2101 1071 -2093
rect 1076 -2101 1080 -2093
rect 1085 -2101 1089 -2093
rect 1093 -2101 1097 -2093
rect 1111 -2101 1115 -2093
rect 1133 -2101 1137 -2093
rect 1145 -2101 1149 -2093
rect 1157 -2101 1161 -2093
rect 1169 -2101 1173 -2093
rect 1177 -2101 1181 -2093
rect 1194 -2101 1198 -2093
rect 1203 -2101 1207 -2093
rect 1321 -2101 1325 -2093
rect 1330 -2101 1334 -2093
rect 1339 -2101 1343 -2093
rect 1347 -2101 1351 -2093
rect 1356 -2101 1360 -2093
rect 1365 -2101 1369 -2093
rect 1373 -2101 1377 -2093
rect 1391 -2101 1395 -2093
rect 1413 -2101 1417 -2093
rect 1425 -2101 1429 -2093
rect 1434 -2101 1438 -2093
rect 1443 -2101 1447 -2093
rect 1451 -2101 1455 -2093
rect 1469 -2101 1473 -2093
rect 1491 -2101 1495 -2093
rect 1503 -2101 1507 -2093
rect 1515 -2101 1519 -2093
rect 1527 -2101 1531 -2093
rect 1535 -2101 1539 -2093
rect 1552 -2101 1556 -2093
rect 1561 -2101 1565 -2093
rect -1264 -2245 -1260 -2237
rect -1255 -2245 -1251 -2237
rect -1246 -2245 -1242 -2237
rect -1238 -2245 -1234 -2237
rect -1230 -2245 -1226 -2237
rect -1218 -2245 -1214 -2237
rect -1206 -2245 -1202 -2237
rect -1197 -2245 -1193 -2237
rect -1188 -2245 -1184 -2237
rect -1176 -2245 -1172 -2237
rect -1164 -2245 -1160 -2237
rect -1155 -2245 -1151 -2237
rect -1146 -2245 -1142 -2237
rect -1134 -2245 -1130 -2237
rect -1122 -2245 -1118 -2237
rect -1113 -2245 -1109 -2237
rect -1104 -2245 -1100 -2237
rect -1092 -2245 -1088 -2237
rect -1080 -2245 -1076 -2237
rect -1072 -2245 -1068 -2237
rect -935 -2245 -931 -2237
rect -926 -2245 -922 -2237
rect -917 -2245 -913 -2237
rect -909 -2245 -905 -2237
rect -901 -2245 -897 -2237
rect -889 -2245 -885 -2237
rect -877 -2245 -873 -2237
rect -868 -2245 -864 -2237
rect -859 -2245 -855 -2237
rect -847 -2245 -843 -2237
rect -835 -2245 -831 -2237
rect -826 -2245 -822 -2237
rect -817 -2245 -813 -2237
rect -805 -2245 -801 -2237
rect -793 -2245 -789 -2237
rect -784 -2245 -780 -2237
rect -775 -2245 -771 -2237
rect -763 -2245 -759 -2237
rect -751 -2245 -747 -2237
rect -743 -2245 -739 -2237
rect -577 -2245 -573 -2237
rect -568 -2245 -564 -2237
rect -559 -2245 -555 -2237
rect -551 -2245 -547 -2237
rect -543 -2245 -539 -2237
rect -531 -2245 -527 -2237
rect -519 -2245 -515 -2237
rect -510 -2245 -506 -2237
rect -501 -2245 -497 -2237
rect -489 -2245 -485 -2237
rect -477 -2245 -473 -2237
rect -468 -2245 -464 -2237
rect -459 -2245 -455 -2237
rect -447 -2245 -443 -2237
rect -435 -2245 -431 -2237
rect -426 -2245 -422 -2237
rect -417 -2245 -413 -2237
rect -405 -2245 -401 -2237
rect -393 -2245 -389 -2237
rect -385 -2245 -381 -2237
rect -219 -2245 -215 -2237
rect -210 -2245 -206 -2237
rect -201 -2245 -197 -2237
rect -193 -2245 -189 -2237
rect -185 -2245 -181 -2237
rect -173 -2245 -169 -2237
rect -161 -2245 -157 -2237
rect -152 -2245 -148 -2237
rect -143 -2245 -139 -2237
rect -131 -2245 -127 -2237
rect -119 -2245 -115 -2237
rect -110 -2245 -106 -2237
rect -101 -2245 -97 -2237
rect -89 -2245 -85 -2237
rect -77 -2245 -73 -2237
rect -68 -2245 -64 -2237
rect -59 -2245 -55 -2237
rect -47 -2245 -43 -2237
rect -35 -2245 -31 -2237
rect -27 -2245 -23 -2237
rect 209 -2245 213 -2237
rect 218 -2245 222 -2237
rect 227 -2245 231 -2237
rect 235 -2245 239 -2237
rect 243 -2245 247 -2237
rect 255 -2245 259 -2237
rect 267 -2245 271 -2237
rect 276 -2245 280 -2237
rect 285 -2245 289 -2237
rect 297 -2245 301 -2237
rect 309 -2245 313 -2237
rect 318 -2245 322 -2237
rect 327 -2245 331 -2237
rect 339 -2245 343 -2237
rect 351 -2245 355 -2237
rect 360 -2245 364 -2237
rect 369 -2245 373 -2237
rect 381 -2245 385 -2237
rect 393 -2245 397 -2237
rect 401 -2245 405 -2237
rect 565 -2245 569 -2237
rect 574 -2245 578 -2237
rect 583 -2245 587 -2237
rect 591 -2245 595 -2237
rect 599 -2245 603 -2237
rect 611 -2245 615 -2237
rect 623 -2245 627 -2237
rect 632 -2245 636 -2237
rect 641 -2245 645 -2237
rect 653 -2245 657 -2237
rect 665 -2245 669 -2237
rect 674 -2245 678 -2237
rect 683 -2245 687 -2237
rect 695 -2245 699 -2237
rect 707 -2245 711 -2237
rect 716 -2245 720 -2237
rect 725 -2245 729 -2237
rect 737 -2245 741 -2237
rect 749 -2245 753 -2237
rect 757 -2245 761 -2237
rect -1264 -2376 -1260 -2368
rect -1255 -2376 -1251 -2368
rect -1246 -2376 -1242 -2368
rect -1238 -2376 -1234 -2368
rect -1230 -2376 -1226 -2368
rect -1218 -2376 -1214 -2368
rect -1206 -2376 -1202 -2368
rect -1197 -2376 -1193 -2368
rect -1188 -2376 -1184 -2368
rect -1176 -2376 -1172 -2368
rect -1164 -2376 -1160 -2368
rect -1155 -2376 -1151 -2368
rect -1146 -2376 -1142 -2368
rect -1134 -2376 -1130 -2368
rect -1122 -2376 -1118 -2368
rect -1113 -2376 -1109 -2368
rect -1104 -2376 -1100 -2368
rect -1092 -2376 -1088 -2368
rect -1080 -2376 -1076 -2368
rect -1072 -2376 -1068 -2368
rect -935 -2376 -931 -2368
rect -926 -2376 -922 -2368
rect -917 -2376 -913 -2368
rect -909 -2376 -905 -2368
rect -901 -2376 -897 -2368
rect -889 -2376 -885 -2368
rect -877 -2376 -873 -2368
rect -868 -2376 -864 -2368
rect -859 -2376 -855 -2368
rect -847 -2376 -843 -2368
rect -835 -2376 -831 -2368
rect -826 -2376 -822 -2368
rect -817 -2376 -813 -2368
rect -805 -2376 -801 -2368
rect -793 -2376 -789 -2368
rect -784 -2376 -780 -2368
rect -775 -2376 -771 -2368
rect -763 -2376 -759 -2368
rect -751 -2376 -747 -2368
rect -743 -2376 -739 -2368
rect -577 -2376 -573 -2368
rect -568 -2376 -564 -2368
rect -559 -2376 -555 -2368
rect -551 -2376 -547 -2368
rect -543 -2376 -539 -2368
rect -531 -2376 -527 -2368
rect -519 -2376 -515 -2368
rect -510 -2376 -506 -2368
rect -501 -2376 -497 -2368
rect -489 -2376 -485 -2368
rect -477 -2376 -473 -2368
rect -468 -2376 -464 -2368
rect -459 -2376 -455 -2368
rect -447 -2376 -443 -2368
rect -435 -2376 -431 -2368
rect -426 -2376 -422 -2368
rect -417 -2376 -413 -2368
rect -405 -2376 -401 -2368
rect -393 -2376 -389 -2368
rect -385 -2376 -381 -2368
rect -219 -2376 -215 -2368
rect -210 -2376 -206 -2368
rect -201 -2376 -197 -2368
rect -193 -2376 -189 -2368
rect -185 -2376 -181 -2368
rect -173 -2376 -169 -2368
rect -161 -2376 -157 -2368
rect -152 -2376 -148 -2368
rect -143 -2376 -139 -2368
rect -131 -2376 -127 -2368
rect -119 -2376 -115 -2368
rect -110 -2376 -106 -2368
rect -101 -2376 -97 -2368
rect -89 -2376 -85 -2368
rect -77 -2376 -73 -2368
rect -68 -2376 -64 -2368
rect -59 -2376 -55 -2368
rect -47 -2376 -43 -2368
rect -35 -2376 -31 -2368
rect -27 -2376 -23 -2368
rect 209 -2376 213 -2368
rect 218 -2376 222 -2368
rect 227 -2376 231 -2368
rect 235 -2376 239 -2368
rect 243 -2376 247 -2368
rect 255 -2376 259 -2368
rect 267 -2376 271 -2368
rect 276 -2376 280 -2368
rect 285 -2376 289 -2368
rect 297 -2376 301 -2368
rect 309 -2376 313 -2368
rect 318 -2376 322 -2368
rect 327 -2376 331 -2368
rect 339 -2376 343 -2368
rect 351 -2376 355 -2368
rect 360 -2376 364 -2368
rect 369 -2376 373 -2368
rect 381 -2376 385 -2368
rect 393 -2376 397 -2368
rect 401 -2376 405 -2368
rect 565 -2376 569 -2368
rect 574 -2376 578 -2368
rect 583 -2376 587 -2368
rect 591 -2376 595 -2368
rect 599 -2376 603 -2368
rect 611 -2376 615 -2368
rect 623 -2376 627 -2368
rect 632 -2376 636 -2368
rect 641 -2376 645 -2368
rect 653 -2376 657 -2368
rect 665 -2376 669 -2368
rect 674 -2376 678 -2368
rect 683 -2376 687 -2368
rect 695 -2376 699 -2368
rect 707 -2376 711 -2368
rect 716 -2376 720 -2368
rect 725 -2376 729 -2368
rect 737 -2376 741 -2368
rect 749 -2376 753 -2368
rect 757 -2376 761 -2368
rect 963 -2376 967 -2368
rect 972 -2376 976 -2368
rect 981 -2376 985 -2368
rect 989 -2376 993 -2368
rect 997 -2376 1001 -2368
rect 1009 -2376 1013 -2368
rect 1021 -2376 1025 -2368
rect 1030 -2376 1034 -2368
rect 1039 -2376 1043 -2368
rect 1051 -2376 1055 -2368
rect 1063 -2376 1067 -2368
rect 1072 -2376 1076 -2368
rect 1081 -2376 1085 -2368
rect 1093 -2376 1097 -2368
rect 1105 -2376 1109 -2368
rect 1114 -2376 1118 -2368
rect 1123 -2376 1127 -2368
rect 1135 -2376 1139 -2368
rect 1147 -2376 1151 -2368
rect 1155 -2376 1159 -2368
rect 1321 -2376 1325 -2368
rect 1330 -2376 1334 -2368
rect 1339 -2376 1343 -2368
rect 1347 -2376 1351 -2368
rect 1355 -2376 1359 -2368
rect 1367 -2376 1371 -2368
rect 1379 -2376 1383 -2368
rect 1388 -2376 1392 -2368
rect 1397 -2376 1401 -2368
rect 1409 -2376 1413 -2368
rect 1421 -2376 1425 -2368
rect 1430 -2376 1434 -2368
rect 1439 -2376 1443 -2368
rect 1451 -2376 1455 -2368
rect 1463 -2376 1467 -2368
rect 1472 -2376 1476 -2368
rect 1481 -2376 1485 -2368
rect 1493 -2376 1497 -2368
rect 1505 -2376 1509 -2368
rect 1513 -2376 1517 -2368
rect -1264 -2507 -1260 -2499
rect -1255 -2507 -1251 -2499
rect -1246 -2507 -1242 -2499
rect -1238 -2507 -1234 -2499
rect -1230 -2507 -1226 -2499
rect -1218 -2507 -1214 -2499
rect -1206 -2507 -1202 -2499
rect -1197 -2507 -1193 -2499
rect -1188 -2507 -1184 -2499
rect -1176 -2507 -1172 -2499
rect -1164 -2507 -1160 -2499
rect -1155 -2507 -1151 -2499
rect -1146 -2507 -1142 -2499
rect -1134 -2507 -1130 -2499
rect -1122 -2507 -1118 -2499
rect -1113 -2507 -1109 -2499
rect -1104 -2507 -1100 -2499
rect -1092 -2507 -1088 -2499
rect -1080 -2507 -1076 -2499
rect -1072 -2507 -1068 -2499
rect -935 -2507 -931 -2499
rect -926 -2507 -922 -2499
rect -917 -2507 -913 -2499
rect -909 -2507 -905 -2499
rect -901 -2507 -897 -2499
rect -889 -2507 -885 -2499
rect -877 -2507 -873 -2499
rect -868 -2507 -864 -2499
rect -859 -2507 -855 -2499
rect -847 -2507 -843 -2499
rect -835 -2507 -831 -2499
rect -826 -2507 -822 -2499
rect -817 -2507 -813 -2499
rect -805 -2507 -801 -2499
rect -793 -2507 -789 -2499
rect -784 -2507 -780 -2499
rect -775 -2507 -771 -2499
rect -763 -2507 -759 -2499
rect -751 -2507 -747 -2499
rect -743 -2507 -739 -2499
rect -577 -2507 -573 -2499
rect -568 -2507 -564 -2499
rect -559 -2507 -555 -2499
rect -551 -2507 -547 -2499
rect -543 -2507 -539 -2499
rect -531 -2507 -527 -2499
rect -519 -2507 -515 -2499
rect -510 -2507 -506 -2499
rect -501 -2507 -497 -2499
rect -489 -2507 -485 -2499
rect -477 -2507 -473 -2499
rect -468 -2507 -464 -2499
rect -459 -2507 -455 -2499
rect -447 -2507 -443 -2499
rect -435 -2507 -431 -2499
rect -426 -2507 -422 -2499
rect -417 -2507 -413 -2499
rect -405 -2507 -401 -2499
rect -393 -2507 -389 -2499
rect -385 -2507 -381 -2499
rect -219 -2507 -215 -2499
rect -210 -2507 -206 -2499
rect -201 -2507 -197 -2499
rect -193 -2507 -189 -2499
rect -185 -2507 -181 -2499
rect -173 -2507 -169 -2499
rect -161 -2507 -157 -2499
rect -152 -2507 -148 -2499
rect -143 -2507 -139 -2499
rect -131 -2507 -127 -2499
rect -119 -2507 -115 -2499
rect -110 -2507 -106 -2499
rect -101 -2507 -97 -2499
rect -89 -2507 -85 -2499
rect -77 -2507 -73 -2499
rect -68 -2507 -64 -2499
rect -59 -2507 -55 -2499
rect -47 -2507 -43 -2499
rect -35 -2507 -31 -2499
rect -27 -2507 -23 -2499
rect 90 -2531 94 -2499
rect 98 -2531 102 -2499
rect 209 -2507 213 -2499
rect 218 -2507 222 -2499
rect 227 -2507 231 -2499
rect 235 -2507 239 -2499
rect 243 -2507 247 -2499
rect 255 -2507 259 -2499
rect 267 -2507 271 -2499
rect 276 -2507 280 -2499
rect 285 -2507 289 -2499
rect 297 -2507 301 -2499
rect 309 -2507 313 -2499
rect 318 -2507 322 -2499
rect 327 -2507 331 -2499
rect 339 -2507 343 -2499
rect 351 -2507 355 -2499
rect 360 -2507 364 -2499
rect 369 -2507 373 -2499
rect 381 -2507 385 -2499
rect 393 -2507 397 -2499
rect 401 -2507 405 -2499
rect 565 -2507 569 -2499
rect 574 -2507 578 -2499
rect 583 -2507 587 -2499
rect 591 -2507 595 -2499
rect 599 -2507 603 -2499
rect 611 -2507 615 -2499
rect 623 -2507 627 -2499
rect 632 -2507 636 -2499
rect 641 -2507 645 -2499
rect 653 -2507 657 -2499
rect 665 -2507 669 -2499
rect 674 -2507 678 -2499
rect 683 -2507 687 -2499
rect 695 -2507 699 -2499
rect 707 -2507 711 -2499
rect 716 -2507 720 -2499
rect 725 -2507 729 -2499
rect 737 -2507 741 -2499
rect 749 -2507 753 -2499
rect 757 -2507 761 -2499
rect 963 -2507 967 -2499
rect 972 -2507 976 -2499
rect 981 -2507 985 -2499
rect 989 -2507 993 -2499
rect 997 -2507 1001 -2499
rect 1009 -2507 1013 -2499
rect 1021 -2507 1025 -2499
rect 1030 -2507 1034 -2499
rect 1039 -2507 1043 -2499
rect 1051 -2507 1055 -2499
rect 1063 -2507 1067 -2499
rect 1072 -2507 1076 -2499
rect 1081 -2507 1085 -2499
rect 1093 -2507 1097 -2499
rect 1105 -2507 1109 -2499
rect 1114 -2507 1118 -2499
rect 1123 -2507 1127 -2499
rect 1135 -2507 1139 -2499
rect 1147 -2507 1151 -2499
rect 1155 -2507 1159 -2499
rect 1321 -2507 1325 -2499
rect 1330 -2507 1334 -2499
rect 1339 -2507 1343 -2499
rect 1347 -2507 1351 -2499
rect 1355 -2507 1359 -2499
rect 1367 -2507 1371 -2499
rect 1379 -2507 1383 -2499
rect 1388 -2507 1392 -2499
rect 1397 -2507 1401 -2499
rect 1409 -2507 1413 -2499
rect 1421 -2507 1425 -2499
rect 1430 -2507 1434 -2499
rect 1439 -2507 1443 -2499
rect 1451 -2507 1455 -2499
rect 1463 -2507 1467 -2499
rect 1472 -2507 1476 -2499
rect 1481 -2507 1485 -2499
rect 1493 -2507 1497 -2499
rect 1505 -2507 1509 -2499
rect 1513 -2507 1517 -2499
rect -1264 -2619 -1260 -2611
rect -1255 -2619 -1251 -2611
rect -1246 -2619 -1242 -2611
rect -1238 -2619 -1234 -2611
rect -1230 -2619 -1226 -2611
rect -1218 -2619 -1214 -2611
rect -1206 -2619 -1202 -2611
rect -1197 -2619 -1193 -2611
rect -1188 -2619 -1184 -2611
rect -1176 -2619 -1172 -2611
rect -1164 -2619 -1160 -2611
rect -1155 -2619 -1151 -2611
rect -1146 -2619 -1142 -2611
rect -1134 -2619 -1130 -2611
rect -1122 -2619 -1118 -2611
rect -1113 -2619 -1109 -2611
rect -1104 -2619 -1100 -2611
rect -1092 -2619 -1088 -2611
rect -1080 -2619 -1076 -2611
rect -1072 -2619 -1068 -2611
rect -935 -2619 -931 -2611
rect -926 -2619 -922 -2611
rect -917 -2619 -913 -2611
rect -909 -2619 -905 -2611
rect -901 -2619 -897 -2611
rect -889 -2619 -885 -2611
rect -877 -2619 -873 -2611
rect -868 -2619 -864 -2611
rect -859 -2619 -855 -2611
rect -847 -2619 -843 -2611
rect -835 -2619 -831 -2611
rect -826 -2619 -822 -2611
rect -817 -2619 -813 -2611
rect -805 -2619 -801 -2611
rect -793 -2619 -789 -2611
rect -784 -2619 -780 -2611
rect -775 -2619 -771 -2611
rect -763 -2619 -759 -2611
rect -751 -2619 -747 -2611
rect -743 -2619 -739 -2611
rect -1339 -2732 -1335 -2724
rect -1331 -2732 -1327 -2724
rect -1322 -2732 -1318 -2724
rect -1313 -2732 -1309 -2724
rect -935 -2732 -931 -2724
rect -927 -2732 -923 -2724
rect -918 -2732 -914 -2724
rect -909 -2732 -905 -2724
rect -577 -2732 -573 -2724
rect -569 -2732 -565 -2724
rect -560 -2732 -556 -2724
rect -551 -2732 -547 -2724
rect -219 -2732 -215 -2724
rect -211 -2732 -207 -2724
rect -202 -2732 -198 -2724
rect -193 -2732 -189 -2724
rect 209 -2732 213 -2724
rect 217 -2732 221 -2724
rect 226 -2732 230 -2724
rect 235 -2732 239 -2724
rect 565 -2732 569 -2724
rect 573 -2732 577 -2724
rect 582 -2732 586 -2724
rect 591 -2732 595 -2724
rect 963 -2732 967 -2724
rect 971 -2732 975 -2724
rect 980 -2732 984 -2724
rect 989 -2732 993 -2724
rect 1321 -2732 1325 -2724
rect 1329 -2732 1333 -2724
rect 1338 -2732 1342 -2724
rect 1347 -2732 1351 -2724
rect -1264 -2851 -1260 -2843
rect -1255 -2851 -1251 -2843
rect -1246 -2851 -1242 -2843
rect -1238 -2851 -1234 -2843
rect -1220 -2851 -1216 -2843
rect -1198 -2851 -1194 -2843
rect -1186 -2851 -1182 -2843
rect -1177 -2851 -1173 -2843
rect -1168 -2851 -1164 -2843
rect -935 -2851 -931 -2843
rect -926 -2851 -922 -2843
rect -917 -2851 -913 -2843
rect -909 -2851 -905 -2843
rect -900 -2851 -896 -2843
rect -891 -2851 -887 -2843
rect -883 -2851 -879 -2843
rect -865 -2851 -861 -2843
rect -843 -2851 -839 -2843
rect -831 -2851 -827 -2843
rect -822 -2851 -818 -2843
rect -813 -2851 -809 -2843
rect -805 -2851 -801 -2843
rect -787 -2851 -783 -2843
rect -765 -2851 -761 -2843
rect -753 -2851 -749 -2843
rect -741 -2851 -737 -2843
rect -729 -2851 -725 -2843
rect -721 -2851 -717 -2843
rect -704 -2851 -700 -2843
rect -695 -2851 -691 -2843
rect -577 -2851 -573 -2843
rect -568 -2851 -564 -2843
rect -559 -2851 -555 -2843
rect -551 -2851 -547 -2843
rect -542 -2851 -538 -2843
rect -533 -2851 -529 -2843
rect -525 -2851 -521 -2843
rect -507 -2851 -503 -2843
rect -485 -2851 -481 -2843
rect -473 -2851 -469 -2843
rect -464 -2851 -460 -2843
rect -455 -2851 -451 -2843
rect -447 -2851 -443 -2843
rect -429 -2851 -425 -2843
rect -407 -2851 -403 -2843
rect -395 -2851 -391 -2843
rect -383 -2851 -379 -2843
rect -371 -2851 -367 -2843
rect -363 -2851 -359 -2843
rect -346 -2851 -342 -2843
rect -337 -2851 -333 -2843
rect -219 -2851 -215 -2843
rect -210 -2851 -206 -2843
rect -201 -2851 -197 -2843
rect -193 -2851 -189 -2843
rect -184 -2851 -180 -2843
rect -175 -2851 -171 -2843
rect -167 -2851 -163 -2843
rect -149 -2851 -145 -2843
rect -127 -2851 -123 -2843
rect -115 -2851 -111 -2843
rect -106 -2851 -102 -2843
rect -97 -2851 -93 -2843
rect -89 -2851 -85 -2843
rect -71 -2851 -67 -2843
rect -49 -2851 -45 -2843
rect -37 -2851 -33 -2843
rect -25 -2851 -21 -2843
rect -13 -2851 -9 -2843
rect -5 -2851 -1 -2843
rect 12 -2851 16 -2843
rect 21 -2851 25 -2843
rect 209 -2851 213 -2843
rect 218 -2851 222 -2843
rect 227 -2851 231 -2843
rect 235 -2851 239 -2843
rect 244 -2851 248 -2843
rect 253 -2851 257 -2843
rect 261 -2851 265 -2843
rect 279 -2851 283 -2843
rect 301 -2851 305 -2843
rect 313 -2851 317 -2843
rect 322 -2851 326 -2843
rect 331 -2851 335 -2843
rect 339 -2851 343 -2843
rect 357 -2851 361 -2843
rect 379 -2851 383 -2843
rect 391 -2851 395 -2843
rect 403 -2851 407 -2843
rect 415 -2851 419 -2843
rect 423 -2851 427 -2843
rect 440 -2851 444 -2843
rect 449 -2851 453 -2843
rect 565 -2851 569 -2843
rect 574 -2851 578 -2843
rect 583 -2851 587 -2843
rect 591 -2851 595 -2843
rect 600 -2851 604 -2843
rect 609 -2851 613 -2843
rect 617 -2851 621 -2843
rect 635 -2851 639 -2843
rect 657 -2851 661 -2843
rect 669 -2851 673 -2843
rect 678 -2851 682 -2843
rect 687 -2851 691 -2843
rect 695 -2851 699 -2843
rect 713 -2851 717 -2843
rect 735 -2851 739 -2843
rect 747 -2851 751 -2843
rect 759 -2851 763 -2843
rect 771 -2851 775 -2843
rect 779 -2851 783 -2843
rect 796 -2851 800 -2843
rect 805 -2851 809 -2843
rect 963 -2851 967 -2843
rect 972 -2851 976 -2843
rect 981 -2851 985 -2843
rect 989 -2851 993 -2843
rect 998 -2851 1002 -2843
rect 1007 -2851 1011 -2843
rect 1015 -2851 1019 -2843
rect 1033 -2851 1037 -2843
rect 1055 -2851 1059 -2843
rect 1067 -2851 1071 -2843
rect 1076 -2851 1080 -2843
rect 1085 -2851 1089 -2843
rect 1093 -2851 1097 -2843
rect 1111 -2851 1115 -2843
rect 1133 -2851 1137 -2843
rect 1145 -2851 1149 -2843
rect 1157 -2851 1161 -2843
rect 1169 -2851 1173 -2843
rect 1177 -2851 1181 -2843
rect 1194 -2851 1198 -2843
rect 1203 -2851 1207 -2843
rect 1321 -2851 1325 -2843
rect 1330 -2851 1334 -2843
rect 1339 -2851 1343 -2843
rect 1347 -2851 1351 -2843
rect 1356 -2851 1360 -2843
rect 1365 -2851 1369 -2843
rect 1373 -2851 1377 -2843
rect 1391 -2851 1395 -2843
rect 1413 -2851 1417 -2843
rect 1425 -2851 1429 -2843
rect 1434 -2851 1438 -2843
rect 1443 -2851 1447 -2843
rect 1451 -2851 1455 -2843
rect 1469 -2851 1473 -2843
rect 1491 -2851 1495 -2843
rect 1503 -2851 1507 -2843
rect 1515 -2851 1519 -2843
rect 1527 -2851 1531 -2843
rect 1535 -2851 1539 -2843
rect 1552 -2851 1556 -2843
rect 1561 -2851 1565 -2843
rect -1264 -2970 -1260 -2962
rect -1255 -2970 -1251 -2962
rect -1246 -2970 -1242 -2962
rect -1238 -2970 -1234 -2962
rect -1230 -2970 -1226 -2962
rect -1218 -2970 -1214 -2962
rect -1206 -2970 -1202 -2962
rect -1197 -2970 -1193 -2962
rect -1188 -2970 -1184 -2962
rect -1176 -2970 -1172 -2962
rect -1164 -2970 -1160 -2962
rect -1155 -2970 -1151 -2962
rect -1146 -2970 -1142 -2962
rect -1134 -2970 -1130 -2962
rect -1122 -2970 -1118 -2962
rect -1113 -2970 -1109 -2962
rect -1104 -2970 -1100 -2962
rect -1092 -2970 -1088 -2962
rect -1080 -2970 -1076 -2962
rect -1072 -2970 -1068 -2962
rect -1026 -2970 -1022 -2962
rect -1018 -2970 -1014 -2962
rect -935 -2970 -931 -2962
rect -926 -2970 -922 -2962
rect -917 -2970 -913 -2962
rect -909 -2970 -905 -2962
rect -901 -2970 -897 -2962
rect -889 -2970 -885 -2962
rect -877 -2970 -873 -2962
rect -868 -2970 -864 -2962
rect -859 -2970 -855 -2962
rect -847 -2970 -843 -2962
rect -835 -2970 -831 -2962
rect -826 -2970 -822 -2962
rect -817 -2970 -813 -2962
rect -805 -2970 -801 -2962
rect -793 -2970 -789 -2962
rect -784 -2970 -780 -2962
rect -775 -2970 -771 -2962
rect -763 -2970 -759 -2962
rect -751 -2970 -747 -2962
rect -743 -2970 -739 -2962
rect -672 -2978 -668 -2962
rect -664 -2978 -660 -2962
rect -577 -2970 -573 -2962
rect -568 -2970 -564 -2962
rect -559 -2970 -555 -2962
rect -551 -2970 -547 -2962
rect -543 -2970 -539 -2962
rect -531 -2970 -527 -2962
rect -519 -2970 -515 -2962
rect -510 -2970 -506 -2962
rect -501 -2970 -497 -2962
rect -489 -2970 -485 -2962
rect -477 -2970 -473 -2962
rect -468 -2970 -464 -2962
rect -459 -2970 -455 -2962
rect -447 -2970 -443 -2962
rect -435 -2970 -431 -2962
rect -426 -2970 -422 -2962
rect -417 -2970 -413 -2962
rect -405 -2970 -401 -2962
rect -393 -2970 -389 -2962
rect -385 -2970 -381 -2962
rect -329 -2970 -325 -2962
rect -321 -2970 -317 -2962
rect -219 -2970 -215 -2962
rect -210 -2970 -206 -2962
rect -201 -2970 -197 -2962
rect -193 -2970 -189 -2962
rect -185 -2970 -181 -2962
rect -173 -2970 -169 -2962
rect -161 -2970 -157 -2962
rect -152 -2970 -148 -2962
rect -143 -2970 -139 -2962
rect -131 -2970 -127 -2962
rect -119 -2970 -115 -2962
rect -110 -2970 -106 -2962
rect -101 -2970 -97 -2962
rect -89 -2970 -85 -2962
rect -77 -2970 -73 -2962
rect -68 -2970 -64 -2962
rect -59 -2970 -55 -2962
rect -47 -2970 -43 -2962
rect -35 -2970 -31 -2962
rect -27 -2970 -23 -2962
rect 209 -2970 213 -2962
rect 218 -2970 222 -2962
rect 227 -2970 231 -2962
rect 235 -2970 239 -2962
rect 243 -2970 247 -2962
rect 255 -2970 259 -2962
rect 267 -2970 271 -2962
rect 276 -2970 280 -2962
rect 285 -2970 289 -2962
rect 297 -2970 301 -2962
rect 309 -2970 313 -2962
rect 318 -2970 322 -2962
rect 327 -2970 331 -2962
rect 339 -2970 343 -2962
rect 351 -2970 355 -2962
rect 360 -2970 364 -2962
rect 369 -2970 373 -2962
rect 381 -2970 385 -2962
rect 393 -2970 397 -2962
rect 401 -2970 405 -2962
rect 472 -2970 476 -2962
rect 480 -2970 484 -2962
rect 841 -2978 845 -2962
rect 849 -2978 853 -2962
rect 1199 -2970 1203 -2962
rect 1207 -2970 1211 -2962
rect -1264 -3086 -1260 -3078
rect -1255 -3086 -1251 -3078
rect -1246 -3086 -1242 -3078
rect -1238 -3086 -1234 -3078
rect -1230 -3086 -1226 -3078
rect -1218 -3086 -1214 -3078
rect -1206 -3086 -1202 -3078
rect -1197 -3086 -1193 -3078
rect -1188 -3086 -1184 -3078
rect -1176 -3086 -1172 -3078
rect -1164 -3086 -1160 -3078
rect -1155 -3086 -1151 -3078
rect -1146 -3086 -1142 -3078
rect -1134 -3086 -1130 -3078
rect -1122 -3086 -1118 -3078
rect -1113 -3086 -1109 -3078
rect -1104 -3086 -1100 -3078
rect -1092 -3086 -1088 -3078
rect -1080 -3086 -1076 -3078
rect -1072 -3086 -1068 -3078
rect -1026 -3086 -1022 -3078
rect -1018 -3086 -1014 -3078
rect -935 -3086 -931 -3078
rect -926 -3086 -922 -3078
rect -917 -3086 -913 -3078
rect -909 -3086 -905 -3078
rect -901 -3086 -897 -3078
rect -889 -3086 -885 -3078
rect -877 -3086 -873 -3078
rect -868 -3086 -864 -3078
rect -859 -3086 -855 -3078
rect -847 -3086 -843 -3078
rect -835 -3086 -831 -3078
rect -826 -3086 -822 -3078
rect -817 -3086 -813 -3078
rect -805 -3086 -801 -3078
rect -793 -3086 -789 -3078
rect -784 -3086 -780 -3078
rect -775 -3086 -771 -3078
rect -763 -3086 -759 -3078
rect -751 -3086 -747 -3078
rect -743 -3086 -739 -3078
rect -577 -3086 -573 -3078
rect -568 -3086 -564 -3078
rect -559 -3086 -555 -3078
rect -551 -3086 -547 -3078
rect -543 -3086 -539 -3078
rect -531 -3086 -527 -3078
rect -519 -3086 -515 -3078
rect -510 -3086 -506 -3078
rect -501 -3086 -497 -3078
rect -489 -3086 -485 -3078
rect -477 -3086 -473 -3078
rect -468 -3086 -464 -3078
rect -459 -3086 -455 -3078
rect -447 -3086 -443 -3078
rect -435 -3086 -431 -3078
rect -426 -3086 -422 -3078
rect -417 -3086 -413 -3078
rect -405 -3086 -401 -3078
rect -393 -3086 -389 -3078
rect -385 -3086 -381 -3078
rect -329 -3086 -325 -3078
rect -321 -3086 -317 -3078
rect -219 -3086 -215 -3078
rect -210 -3086 -206 -3078
rect -201 -3086 -197 -3078
rect -193 -3086 -189 -3078
rect -185 -3086 -181 -3078
rect -173 -3086 -169 -3078
rect -161 -3086 -157 -3078
rect -152 -3086 -148 -3078
rect -143 -3086 -139 -3078
rect -131 -3086 -127 -3078
rect -119 -3086 -115 -3078
rect -110 -3086 -106 -3078
rect -101 -3086 -97 -3078
rect -89 -3086 -85 -3078
rect -77 -3086 -73 -3078
rect -68 -3086 -64 -3078
rect -59 -3086 -55 -3078
rect -47 -3086 -43 -3078
rect -35 -3086 -31 -3078
rect -27 -3086 -23 -3078
rect 209 -3086 213 -3078
rect 218 -3086 222 -3078
rect 227 -3086 231 -3078
rect 235 -3086 239 -3078
rect 243 -3086 247 -3078
rect 255 -3086 259 -3078
rect 267 -3086 271 -3078
rect 276 -3086 280 -3078
rect 285 -3086 289 -3078
rect 297 -3086 301 -3078
rect 309 -3086 313 -3078
rect 318 -3086 322 -3078
rect 327 -3086 331 -3078
rect 339 -3086 343 -3078
rect 351 -3086 355 -3078
rect 360 -3086 364 -3078
rect 369 -3086 373 -3078
rect 381 -3086 385 -3078
rect 393 -3086 397 -3078
rect 401 -3086 405 -3078
rect 472 -3086 476 -3078
rect 480 -3086 484 -3078
rect 565 -3086 569 -3078
rect 574 -3086 578 -3078
rect 583 -3086 587 -3078
rect 591 -3086 595 -3078
rect 599 -3086 603 -3078
rect 611 -3086 615 -3078
rect 623 -3086 627 -3078
rect 632 -3086 636 -3078
rect 641 -3086 645 -3078
rect 653 -3086 657 -3078
rect 665 -3086 669 -3078
rect 674 -3086 678 -3078
rect 683 -3086 687 -3078
rect 695 -3086 699 -3078
rect 707 -3086 711 -3078
rect 716 -3086 720 -3078
rect 725 -3086 729 -3078
rect 737 -3086 741 -3078
rect 749 -3086 753 -3078
rect 757 -3086 761 -3078
rect 963 -3086 967 -3078
rect 972 -3086 976 -3078
rect 981 -3086 985 -3078
rect 989 -3086 993 -3078
rect 997 -3086 1001 -3078
rect 1009 -3086 1013 -3078
rect 1021 -3086 1025 -3078
rect 1030 -3086 1034 -3078
rect 1039 -3086 1043 -3078
rect 1051 -3086 1055 -3078
rect 1063 -3086 1067 -3078
rect 1072 -3086 1076 -3078
rect 1081 -3086 1085 -3078
rect 1093 -3086 1097 -3078
rect 1105 -3086 1109 -3078
rect 1114 -3086 1118 -3078
rect 1123 -3086 1127 -3078
rect 1135 -3086 1139 -3078
rect 1147 -3086 1151 -3078
rect 1155 -3086 1159 -3078
rect 1199 -3086 1203 -3078
rect 1207 -3086 1211 -3078
rect 1321 -3086 1325 -3078
rect 1330 -3086 1334 -3078
rect 1339 -3086 1343 -3078
rect 1347 -3086 1351 -3078
rect 1355 -3086 1359 -3078
rect 1367 -3086 1371 -3078
rect 1379 -3086 1383 -3078
rect 1388 -3086 1392 -3078
rect 1397 -3086 1401 -3078
rect 1409 -3086 1413 -3078
rect 1421 -3086 1425 -3078
rect 1430 -3086 1434 -3078
rect 1439 -3086 1443 -3078
rect 1451 -3086 1455 -3078
rect 1463 -3086 1467 -3078
rect 1472 -3086 1476 -3078
rect 1481 -3086 1485 -3078
rect 1493 -3086 1497 -3078
rect 1505 -3086 1509 -3078
rect 1513 -3086 1517 -3078
rect -1264 -3207 -1260 -3199
rect -1255 -3207 -1251 -3199
rect -1246 -3207 -1242 -3199
rect -1238 -3207 -1234 -3199
rect -1230 -3207 -1226 -3199
rect -1218 -3207 -1214 -3199
rect -1206 -3207 -1202 -3199
rect -1197 -3207 -1193 -3199
rect -1188 -3207 -1184 -3199
rect -1176 -3207 -1172 -3199
rect -1164 -3207 -1160 -3199
rect -1155 -3207 -1151 -3199
rect -1146 -3207 -1142 -3199
rect -1134 -3207 -1130 -3199
rect -1122 -3207 -1118 -3199
rect -1113 -3207 -1109 -3199
rect -1104 -3207 -1100 -3199
rect -1092 -3207 -1088 -3199
rect -1080 -3207 -1076 -3199
rect -1072 -3207 -1068 -3199
rect -935 -3207 -931 -3199
rect -926 -3207 -922 -3199
rect -917 -3207 -913 -3199
rect -909 -3207 -905 -3199
rect -901 -3207 -897 -3199
rect -889 -3207 -885 -3199
rect -877 -3207 -873 -3199
rect -868 -3207 -864 -3199
rect -859 -3207 -855 -3199
rect -847 -3207 -843 -3199
rect -835 -3207 -831 -3199
rect -826 -3207 -822 -3199
rect -817 -3207 -813 -3199
rect -805 -3207 -801 -3199
rect -793 -3207 -789 -3199
rect -784 -3207 -780 -3199
rect -775 -3207 -771 -3199
rect -763 -3207 -759 -3199
rect -751 -3207 -747 -3199
rect -743 -3207 -739 -3199
rect -577 -3207 -573 -3199
rect -568 -3207 -564 -3199
rect -559 -3207 -555 -3199
rect -551 -3207 -547 -3199
rect -543 -3207 -539 -3199
rect -531 -3207 -527 -3199
rect -519 -3207 -515 -3199
rect -510 -3207 -506 -3199
rect -501 -3207 -497 -3199
rect -489 -3207 -485 -3199
rect -477 -3207 -473 -3199
rect -468 -3207 -464 -3199
rect -459 -3207 -455 -3199
rect -447 -3207 -443 -3199
rect -435 -3207 -431 -3199
rect -426 -3207 -422 -3199
rect -417 -3207 -413 -3199
rect -405 -3207 -401 -3199
rect -393 -3207 -389 -3199
rect -385 -3207 -381 -3199
rect -219 -3207 -215 -3199
rect -210 -3207 -206 -3199
rect -201 -3207 -197 -3199
rect -193 -3207 -189 -3199
rect -185 -3207 -181 -3199
rect -173 -3207 -169 -3199
rect -161 -3207 -157 -3199
rect -152 -3207 -148 -3199
rect -143 -3207 -139 -3199
rect -131 -3207 -127 -3199
rect -119 -3207 -115 -3199
rect -110 -3207 -106 -3199
rect -101 -3207 -97 -3199
rect -89 -3207 -85 -3199
rect -77 -3207 -73 -3199
rect -68 -3207 -64 -3199
rect -59 -3207 -55 -3199
rect -47 -3207 -43 -3199
rect -35 -3207 -31 -3199
rect -27 -3207 -23 -3199
rect 209 -3207 213 -3199
rect 218 -3207 222 -3199
rect 227 -3207 231 -3199
rect 235 -3207 239 -3199
rect 243 -3207 247 -3199
rect 255 -3207 259 -3199
rect 267 -3207 271 -3199
rect 276 -3207 280 -3199
rect 285 -3207 289 -3199
rect 297 -3207 301 -3199
rect 309 -3207 313 -3199
rect 318 -3207 322 -3199
rect 327 -3207 331 -3199
rect 339 -3207 343 -3199
rect 351 -3207 355 -3199
rect 360 -3207 364 -3199
rect 369 -3207 373 -3199
rect 381 -3207 385 -3199
rect 393 -3207 397 -3199
rect 401 -3207 405 -3199
rect 565 -3207 569 -3199
rect 574 -3207 578 -3199
rect 583 -3207 587 -3199
rect 591 -3207 595 -3199
rect 599 -3207 603 -3199
rect 611 -3207 615 -3199
rect 623 -3207 627 -3199
rect 632 -3207 636 -3199
rect 641 -3207 645 -3199
rect 653 -3207 657 -3199
rect 665 -3207 669 -3199
rect 674 -3207 678 -3199
rect 683 -3207 687 -3199
rect 695 -3207 699 -3199
rect 707 -3207 711 -3199
rect 716 -3207 720 -3199
rect 725 -3207 729 -3199
rect 737 -3207 741 -3199
rect 749 -3207 753 -3199
rect 757 -3207 761 -3199
rect 963 -3207 967 -3199
rect 972 -3207 976 -3199
rect 981 -3207 985 -3199
rect 989 -3207 993 -3199
rect 997 -3207 1001 -3199
rect 1009 -3207 1013 -3199
rect 1021 -3207 1025 -3199
rect 1030 -3207 1034 -3199
rect 1039 -3207 1043 -3199
rect 1051 -3207 1055 -3199
rect 1063 -3207 1067 -3199
rect 1072 -3207 1076 -3199
rect 1081 -3207 1085 -3199
rect 1093 -3207 1097 -3199
rect 1105 -3207 1109 -3199
rect 1114 -3207 1118 -3199
rect 1123 -3207 1127 -3199
rect 1135 -3207 1139 -3199
rect 1147 -3207 1151 -3199
rect 1155 -3207 1159 -3199
rect 1321 -3207 1325 -3199
rect 1330 -3207 1334 -3199
rect 1339 -3207 1343 -3199
rect 1347 -3207 1351 -3199
rect 1355 -3207 1359 -3199
rect 1367 -3207 1371 -3199
rect 1379 -3207 1383 -3199
rect 1388 -3207 1392 -3199
rect 1397 -3207 1401 -3199
rect 1409 -3207 1413 -3199
rect 1421 -3207 1425 -3199
rect 1430 -3207 1434 -3199
rect 1439 -3207 1443 -3199
rect 1451 -3207 1455 -3199
rect 1463 -3207 1467 -3199
rect 1472 -3207 1476 -3199
rect 1481 -3207 1485 -3199
rect 1493 -3207 1497 -3199
rect 1505 -3207 1509 -3199
rect 1513 -3207 1517 -3199
rect -1264 -3321 -1260 -3313
rect -1255 -3321 -1251 -3313
rect -1246 -3321 -1242 -3313
rect -1238 -3321 -1234 -3313
rect -1230 -3321 -1226 -3313
rect -1218 -3321 -1214 -3313
rect -1206 -3321 -1202 -3313
rect -1197 -3321 -1193 -3313
rect -1188 -3321 -1184 -3313
rect -1176 -3321 -1172 -3313
rect -1164 -3321 -1160 -3313
rect -1155 -3321 -1151 -3313
rect -1146 -3321 -1142 -3313
rect -1134 -3321 -1130 -3313
rect -1122 -3321 -1118 -3313
rect -1113 -3321 -1109 -3313
rect -1104 -3321 -1100 -3313
rect -1092 -3321 -1088 -3313
rect -1080 -3321 -1076 -3313
rect -1072 -3321 -1068 -3313
rect -935 -3321 -931 -3313
rect -926 -3321 -922 -3313
rect -917 -3321 -913 -3313
rect -909 -3321 -905 -3313
rect -901 -3321 -897 -3313
rect -889 -3321 -885 -3313
rect -877 -3321 -873 -3313
rect -868 -3321 -864 -3313
rect -859 -3321 -855 -3313
rect -847 -3321 -843 -3313
rect -835 -3321 -831 -3313
rect -826 -3321 -822 -3313
rect -817 -3321 -813 -3313
rect -805 -3321 -801 -3313
rect -793 -3321 -789 -3313
rect -784 -3321 -780 -3313
rect -775 -3321 -771 -3313
rect -763 -3321 -759 -3313
rect -751 -3321 -747 -3313
rect -743 -3321 -739 -3313
rect -577 -3321 -573 -3313
rect -568 -3321 -564 -3313
rect -559 -3321 -555 -3313
rect -551 -3321 -547 -3313
rect -543 -3321 -539 -3313
rect -531 -3321 -527 -3313
rect -519 -3321 -515 -3313
rect -510 -3321 -506 -3313
rect -501 -3321 -497 -3313
rect -489 -3321 -485 -3313
rect -477 -3321 -473 -3313
rect -468 -3321 -464 -3313
rect -459 -3321 -455 -3313
rect -447 -3321 -443 -3313
rect -435 -3321 -431 -3313
rect -426 -3321 -422 -3313
rect -417 -3321 -413 -3313
rect -405 -3321 -401 -3313
rect -393 -3321 -389 -3313
rect -385 -3321 -381 -3313
rect -1339 -3438 -1335 -3430
rect -1331 -3438 -1327 -3430
rect -1322 -3438 -1318 -3430
rect -1313 -3438 -1309 -3430
rect -935 -3438 -931 -3430
rect -927 -3438 -923 -3430
rect -918 -3438 -914 -3430
rect -909 -3438 -905 -3430
rect -577 -3438 -573 -3430
rect -569 -3438 -565 -3430
rect -560 -3438 -556 -3430
rect -551 -3438 -547 -3430
rect -219 -3438 -215 -3430
rect -211 -3438 -207 -3430
rect -202 -3438 -198 -3430
rect -193 -3438 -189 -3430
rect 209 -3438 213 -3430
rect 217 -3438 221 -3430
rect 226 -3438 230 -3430
rect 235 -3438 239 -3430
rect 565 -3438 569 -3430
rect 573 -3438 577 -3430
rect 582 -3438 586 -3430
rect 591 -3438 595 -3430
rect 963 -3438 967 -3430
rect 971 -3438 975 -3430
rect 980 -3438 984 -3430
rect 989 -3438 993 -3430
rect 1321 -3438 1325 -3430
rect 1329 -3438 1333 -3430
rect 1338 -3438 1342 -3430
rect 1347 -3438 1351 -3430
rect -1264 -3562 -1260 -3554
rect -1255 -3562 -1251 -3554
rect -1246 -3562 -1242 -3554
rect -1238 -3562 -1234 -3554
rect -1220 -3562 -1216 -3554
rect -1198 -3562 -1194 -3554
rect -1186 -3562 -1182 -3554
rect -1177 -3562 -1173 -3554
rect -1168 -3562 -1164 -3554
rect -935 -3562 -931 -3554
rect -926 -3562 -922 -3554
rect -917 -3562 -913 -3554
rect -909 -3562 -905 -3554
rect -900 -3562 -896 -3554
rect -891 -3562 -887 -3554
rect -883 -3562 -879 -3554
rect -865 -3562 -861 -3554
rect -843 -3562 -839 -3554
rect -831 -3562 -827 -3554
rect -822 -3562 -818 -3554
rect -813 -3562 -809 -3554
rect -805 -3562 -801 -3554
rect -787 -3562 -783 -3554
rect -765 -3562 -761 -3554
rect -753 -3562 -749 -3554
rect -741 -3562 -737 -3554
rect -729 -3562 -725 -3554
rect -721 -3562 -717 -3554
rect -704 -3562 -700 -3554
rect -695 -3562 -691 -3554
rect -577 -3562 -573 -3554
rect -568 -3562 -564 -3554
rect -559 -3562 -555 -3554
rect -551 -3562 -547 -3554
rect -542 -3562 -538 -3554
rect -533 -3562 -529 -3554
rect -525 -3562 -521 -3554
rect -507 -3562 -503 -3554
rect -485 -3562 -481 -3554
rect -473 -3562 -469 -3554
rect -464 -3562 -460 -3554
rect -455 -3562 -451 -3554
rect -447 -3562 -443 -3554
rect -429 -3562 -425 -3554
rect -407 -3562 -403 -3554
rect -395 -3562 -391 -3554
rect -383 -3562 -379 -3554
rect -371 -3562 -367 -3554
rect -363 -3562 -359 -3554
rect -346 -3562 -342 -3554
rect -337 -3562 -333 -3554
rect -219 -3562 -215 -3554
rect -210 -3562 -206 -3554
rect -201 -3562 -197 -3554
rect -193 -3562 -189 -3554
rect -184 -3562 -180 -3554
rect -175 -3562 -171 -3554
rect -167 -3562 -163 -3554
rect -149 -3562 -145 -3554
rect -127 -3562 -123 -3554
rect -115 -3562 -111 -3554
rect -106 -3562 -102 -3554
rect -97 -3562 -93 -3554
rect -89 -3562 -85 -3554
rect -71 -3562 -67 -3554
rect -49 -3562 -45 -3554
rect -37 -3562 -33 -3554
rect -25 -3562 -21 -3554
rect -13 -3562 -9 -3554
rect -5 -3562 -1 -3554
rect 12 -3562 16 -3554
rect 21 -3562 25 -3554
rect 209 -3562 213 -3554
rect 218 -3562 222 -3554
rect 227 -3562 231 -3554
rect 235 -3562 239 -3554
rect 244 -3562 248 -3554
rect 253 -3562 257 -3554
rect 261 -3562 265 -3554
rect 279 -3562 283 -3554
rect 301 -3562 305 -3554
rect 313 -3562 317 -3554
rect 322 -3562 326 -3554
rect 331 -3562 335 -3554
rect 339 -3562 343 -3554
rect 357 -3562 361 -3554
rect 379 -3562 383 -3554
rect 391 -3562 395 -3554
rect 403 -3562 407 -3554
rect 415 -3562 419 -3554
rect 423 -3562 427 -3554
rect 440 -3562 444 -3554
rect 449 -3562 453 -3554
rect 565 -3562 569 -3554
rect 574 -3562 578 -3554
rect 583 -3562 587 -3554
rect 591 -3562 595 -3554
rect 600 -3562 604 -3554
rect 609 -3562 613 -3554
rect 617 -3562 621 -3554
rect 635 -3562 639 -3554
rect 657 -3562 661 -3554
rect 669 -3562 673 -3554
rect 678 -3562 682 -3554
rect 687 -3562 691 -3554
rect 695 -3562 699 -3554
rect 713 -3562 717 -3554
rect 735 -3562 739 -3554
rect 747 -3562 751 -3554
rect 759 -3562 763 -3554
rect 771 -3562 775 -3554
rect 779 -3562 783 -3554
rect 796 -3562 800 -3554
rect 805 -3562 809 -3554
rect 963 -3562 967 -3554
rect 972 -3562 976 -3554
rect 981 -3562 985 -3554
rect 989 -3562 993 -3554
rect 998 -3562 1002 -3554
rect 1007 -3562 1011 -3554
rect 1015 -3562 1019 -3554
rect 1033 -3562 1037 -3554
rect 1055 -3562 1059 -3554
rect 1067 -3562 1071 -3554
rect 1076 -3562 1080 -3554
rect 1085 -3562 1089 -3554
rect 1093 -3562 1097 -3554
rect 1111 -3562 1115 -3554
rect 1133 -3562 1137 -3554
rect 1145 -3562 1149 -3554
rect 1157 -3562 1161 -3554
rect 1169 -3562 1173 -3554
rect 1177 -3562 1181 -3554
rect 1194 -3562 1198 -3554
rect 1203 -3562 1207 -3554
rect 1321 -3562 1325 -3554
rect 1330 -3562 1334 -3554
rect 1339 -3562 1343 -3554
rect 1347 -3562 1351 -3554
rect 1356 -3562 1360 -3554
rect 1365 -3562 1369 -3554
rect 1373 -3562 1377 -3554
rect 1391 -3562 1395 -3554
rect 1413 -3562 1417 -3554
rect 1425 -3562 1429 -3554
rect 1434 -3562 1438 -3554
rect 1443 -3562 1447 -3554
rect 1451 -3562 1455 -3554
rect 1469 -3562 1473 -3554
rect 1491 -3562 1495 -3554
rect 1503 -3562 1507 -3554
rect 1515 -3562 1519 -3554
rect 1527 -3562 1531 -3554
rect 1535 -3562 1539 -3554
rect 1552 -3562 1556 -3554
rect 1561 -3562 1565 -3554
rect -1264 -3692 -1260 -3684
rect -1255 -3692 -1251 -3684
rect -1246 -3692 -1242 -3684
rect -1238 -3692 -1234 -3684
rect -1230 -3692 -1226 -3684
rect -1218 -3692 -1214 -3684
rect -1206 -3692 -1202 -3684
rect -1197 -3692 -1193 -3684
rect -1188 -3692 -1184 -3684
rect -1176 -3692 -1172 -3684
rect -1164 -3692 -1160 -3684
rect -1155 -3692 -1151 -3684
rect -1146 -3692 -1142 -3684
rect -1134 -3692 -1130 -3684
rect -1122 -3692 -1118 -3684
rect -1113 -3692 -1109 -3684
rect -1104 -3692 -1100 -3684
rect -1092 -3692 -1088 -3684
rect -1080 -3692 -1076 -3684
rect -1072 -3692 -1068 -3684
rect -935 -3692 -931 -3684
rect -926 -3692 -922 -3684
rect -917 -3692 -913 -3684
rect -909 -3692 -905 -3684
rect -901 -3692 -897 -3684
rect -889 -3692 -885 -3684
rect -877 -3692 -873 -3684
rect -868 -3692 -864 -3684
rect -859 -3692 -855 -3684
rect -847 -3692 -843 -3684
rect -835 -3692 -831 -3684
rect -826 -3692 -822 -3684
rect -817 -3692 -813 -3684
rect -805 -3692 -801 -3684
rect -793 -3692 -789 -3684
rect -784 -3692 -780 -3684
rect -775 -3692 -771 -3684
rect -763 -3692 -759 -3684
rect -751 -3692 -747 -3684
rect -743 -3692 -739 -3684
rect -577 -3692 -573 -3684
rect -568 -3692 -564 -3684
rect -559 -3692 -555 -3684
rect -551 -3692 -547 -3684
rect -543 -3692 -539 -3684
rect -531 -3692 -527 -3684
rect -519 -3692 -515 -3684
rect -510 -3692 -506 -3684
rect -501 -3692 -497 -3684
rect -489 -3692 -485 -3684
rect -477 -3692 -473 -3684
rect -468 -3692 -464 -3684
rect -459 -3692 -455 -3684
rect -447 -3692 -443 -3684
rect -435 -3692 -431 -3684
rect -426 -3692 -422 -3684
rect -417 -3692 -413 -3684
rect -405 -3692 -401 -3684
rect -393 -3692 -389 -3684
rect -385 -3692 -381 -3684
rect -219 -3692 -215 -3684
rect -210 -3692 -206 -3684
rect -201 -3692 -197 -3684
rect -193 -3692 -189 -3684
rect -185 -3692 -181 -3684
rect -173 -3692 -169 -3684
rect -161 -3692 -157 -3684
rect -152 -3692 -148 -3684
rect -143 -3692 -139 -3684
rect -131 -3692 -127 -3684
rect -119 -3692 -115 -3684
rect -110 -3692 -106 -3684
rect -101 -3692 -97 -3684
rect -89 -3692 -85 -3684
rect -77 -3692 -73 -3684
rect -68 -3692 -64 -3684
rect -59 -3692 -55 -3684
rect -47 -3692 -43 -3684
rect -35 -3692 -31 -3684
rect -27 -3692 -23 -3684
rect 68 -3831 72 -3799
rect 76 -3831 80 -3799
rect -1264 -3923 -1260 -3915
rect -1255 -3923 -1251 -3915
rect -1246 -3923 -1242 -3915
rect -1238 -3923 -1234 -3915
rect -1230 -3923 -1226 -3915
rect -1218 -3923 -1214 -3915
rect -1206 -3923 -1202 -3915
rect -1197 -3923 -1193 -3915
rect -1188 -3923 -1184 -3915
rect -1176 -3923 -1172 -3915
rect -1164 -3923 -1160 -3915
rect -1155 -3923 -1151 -3915
rect -1146 -3923 -1142 -3915
rect -1134 -3923 -1130 -3915
rect -1122 -3923 -1118 -3915
rect -1113 -3923 -1109 -3915
rect -1104 -3923 -1100 -3915
rect -1092 -3923 -1088 -3915
rect -1080 -3923 -1076 -3915
rect -1072 -3923 -1068 -3915
rect -935 -3923 -931 -3915
rect -926 -3923 -922 -3915
rect -917 -3923 -913 -3915
rect -909 -3923 -905 -3915
rect -901 -3923 -897 -3915
rect -889 -3923 -885 -3915
rect -877 -3923 -873 -3915
rect -868 -3923 -864 -3915
rect -859 -3923 -855 -3915
rect -847 -3923 -843 -3915
rect -835 -3923 -831 -3915
rect -826 -3923 -822 -3915
rect -817 -3923 -813 -3915
rect -805 -3923 -801 -3915
rect -793 -3923 -789 -3915
rect -784 -3923 -780 -3915
rect -775 -3923 -771 -3915
rect -763 -3923 -759 -3915
rect -751 -3923 -747 -3915
rect -743 -3923 -739 -3915
rect -577 -3923 -573 -3915
rect -568 -3923 -564 -3915
rect -559 -3923 -555 -3915
rect -551 -3923 -547 -3915
rect -543 -3923 -539 -3915
rect -531 -3923 -527 -3915
rect -519 -3923 -515 -3915
rect -510 -3923 -506 -3915
rect -501 -3923 -497 -3915
rect -489 -3923 -485 -3915
rect -477 -3923 -473 -3915
rect -468 -3923 -464 -3915
rect -459 -3923 -455 -3915
rect -447 -3923 -443 -3915
rect -435 -3923 -431 -3915
rect -426 -3923 -422 -3915
rect -417 -3923 -413 -3915
rect -405 -3923 -401 -3915
rect -393 -3923 -389 -3915
rect -385 -3923 -381 -3915
rect -219 -3923 -215 -3915
rect -210 -3923 -206 -3915
rect -201 -3923 -197 -3915
rect -193 -3923 -189 -3915
rect -185 -3923 -181 -3915
rect -173 -3923 -169 -3915
rect -161 -3923 -157 -3915
rect -152 -3923 -148 -3915
rect -143 -3923 -139 -3915
rect -131 -3923 -127 -3915
rect -119 -3923 -115 -3915
rect -110 -3923 -106 -3915
rect -101 -3923 -97 -3915
rect -89 -3923 -85 -3915
rect -77 -3923 -73 -3915
rect -68 -3923 -64 -3915
rect -59 -3923 -55 -3915
rect -47 -3923 -43 -3915
rect -35 -3923 -31 -3915
rect -27 -3923 -23 -3915
rect 209 -3923 213 -3915
rect 218 -3923 222 -3915
rect 227 -3923 231 -3915
rect 235 -3923 239 -3915
rect 243 -3923 247 -3915
rect 255 -3923 259 -3915
rect 267 -3923 271 -3915
rect 276 -3923 280 -3915
rect 285 -3923 289 -3915
rect 297 -3923 301 -3915
rect 309 -3923 313 -3915
rect 318 -3923 322 -3915
rect 327 -3923 331 -3915
rect 339 -3923 343 -3915
rect 351 -3923 355 -3915
rect 360 -3923 364 -3915
rect 369 -3923 373 -3915
rect 381 -3923 385 -3915
rect 393 -3923 397 -3915
rect 401 -3923 405 -3915
rect 565 -3923 569 -3915
rect 574 -3923 578 -3915
rect 583 -3923 587 -3915
rect 591 -3923 595 -3915
rect 599 -3923 603 -3915
rect 611 -3923 615 -3915
rect 623 -3923 627 -3915
rect 632 -3923 636 -3915
rect 641 -3923 645 -3915
rect 653 -3923 657 -3915
rect 665 -3923 669 -3915
rect 674 -3923 678 -3915
rect 683 -3923 687 -3915
rect 695 -3923 699 -3915
rect 707 -3923 711 -3915
rect 716 -3923 720 -3915
rect 725 -3923 729 -3915
rect 737 -3923 741 -3915
rect 749 -3923 753 -3915
rect 757 -3923 761 -3915
rect 963 -3923 967 -3915
rect 972 -3923 976 -3915
rect 981 -3923 985 -3915
rect 989 -3923 993 -3915
rect 997 -3923 1001 -3915
rect 1009 -3923 1013 -3915
rect 1021 -3923 1025 -3915
rect 1030 -3923 1034 -3915
rect 1039 -3923 1043 -3915
rect 1051 -3923 1055 -3915
rect 1063 -3923 1067 -3915
rect 1072 -3923 1076 -3915
rect 1081 -3923 1085 -3915
rect 1093 -3923 1097 -3915
rect 1105 -3923 1109 -3915
rect 1114 -3923 1118 -3915
rect 1123 -3923 1127 -3915
rect 1135 -3923 1139 -3915
rect 1147 -3923 1151 -3915
rect 1155 -3923 1159 -3915
rect 1321 -3923 1325 -3915
rect 1330 -3923 1334 -3915
rect 1339 -3923 1343 -3915
rect 1347 -3923 1351 -3915
rect 1355 -3923 1359 -3915
rect 1367 -3923 1371 -3915
rect 1379 -3923 1383 -3915
rect 1388 -3923 1392 -3915
rect 1397 -3923 1401 -3915
rect 1409 -3923 1413 -3915
rect 1421 -3923 1425 -3915
rect 1430 -3923 1434 -3915
rect 1439 -3923 1443 -3915
rect 1451 -3923 1455 -3915
rect 1463 -3923 1467 -3915
rect 1472 -3923 1476 -3915
rect 1481 -3923 1485 -3915
rect 1493 -3923 1497 -3915
rect 1505 -3923 1509 -3915
rect 1513 -3923 1517 -3915
rect -1264 -4048 -1260 -4040
rect -1255 -4048 -1251 -4040
rect -1246 -4048 -1242 -4040
rect -1238 -4048 -1234 -4040
rect -1230 -4048 -1226 -4040
rect -1218 -4048 -1214 -4040
rect -1206 -4048 -1202 -4040
rect -1197 -4048 -1193 -4040
rect -1188 -4048 -1184 -4040
rect -1176 -4048 -1172 -4040
rect -1164 -4048 -1160 -4040
rect -1155 -4048 -1151 -4040
rect -1146 -4048 -1142 -4040
rect -1134 -4048 -1130 -4040
rect -1122 -4048 -1118 -4040
rect -1113 -4048 -1109 -4040
rect -1104 -4048 -1100 -4040
rect -1092 -4048 -1088 -4040
rect -1080 -4048 -1076 -4040
rect -1072 -4048 -1068 -4040
rect -935 -4048 -931 -4040
rect -926 -4048 -922 -4040
rect -917 -4048 -913 -4040
rect -909 -4048 -905 -4040
rect -901 -4048 -897 -4040
rect -889 -4048 -885 -4040
rect -877 -4048 -873 -4040
rect -868 -4048 -864 -4040
rect -859 -4048 -855 -4040
rect -847 -4048 -843 -4040
rect -835 -4048 -831 -4040
rect -826 -4048 -822 -4040
rect -817 -4048 -813 -4040
rect -805 -4048 -801 -4040
rect -793 -4048 -789 -4040
rect -784 -4048 -780 -4040
rect -775 -4048 -771 -4040
rect -763 -4048 -759 -4040
rect -751 -4048 -747 -4040
rect -743 -4048 -739 -4040
rect -577 -4048 -573 -4040
rect -568 -4048 -564 -4040
rect -559 -4048 -555 -4040
rect -551 -4048 -547 -4040
rect -543 -4048 -539 -4040
rect -531 -4048 -527 -4040
rect -519 -4048 -515 -4040
rect -510 -4048 -506 -4040
rect -501 -4048 -497 -4040
rect -489 -4048 -485 -4040
rect -477 -4048 -473 -4040
rect -468 -4048 -464 -4040
rect -459 -4048 -455 -4040
rect -447 -4048 -443 -4040
rect -435 -4048 -431 -4040
rect -426 -4048 -422 -4040
rect -417 -4048 -413 -4040
rect -405 -4048 -401 -4040
rect -393 -4048 -389 -4040
rect -385 -4048 -381 -4040
rect -219 -4048 -215 -4040
rect -210 -4048 -206 -4040
rect -201 -4048 -197 -4040
rect -193 -4048 -189 -4040
rect -185 -4048 -181 -4040
rect -173 -4048 -169 -4040
rect -161 -4048 -157 -4040
rect -152 -4048 -148 -4040
rect -143 -4048 -139 -4040
rect -131 -4048 -127 -4040
rect -119 -4048 -115 -4040
rect -110 -4048 -106 -4040
rect -101 -4048 -97 -4040
rect -89 -4048 -85 -4040
rect -77 -4048 -73 -4040
rect -68 -4048 -64 -4040
rect -59 -4048 -55 -4040
rect -47 -4048 -43 -4040
rect -35 -4048 -31 -4040
rect -27 -4048 -23 -4040
rect 209 -4048 213 -4040
rect 218 -4048 222 -4040
rect 227 -4048 231 -4040
rect 235 -4048 239 -4040
rect 243 -4048 247 -4040
rect 255 -4048 259 -4040
rect 267 -4048 271 -4040
rect 276 -4048 280 -4040
rect 285 -4048 289 -4040
rect 297 -4048 301 -4040
rect 309 -4048 313 -4040
rect 318 -4048 322 -4040
rect 327 -4048 331 -4040
rect 339 -4048 343 -4040
rect 351 -4048 355 -4040
rect 360 -4048 364 -4040
rect 369 -4048 373 -4040
rect 381 -4048 385 -4040
rect 393 -4048 397 -4040
rect 401 -4048 405 -4040
rect 565 -4048 569 -4040
rect 574 -4048 578 -4040
rect 583 -4048 587 -4040
rect 591 -4048 595 -4040
rect 599 -4048 603 -4040
rect 611 -4048 615 -4040
rect 623 -4048 627 -4040
rect 632 -4048 636 -4040
rect 641 -4048 645 -4040
rect 653 -4048 657 -4040
rect 665 -4048 669 -4040
rect 674 -4048 678 -4040
rect 683 -4048 687 -4040
rect 695 -4048 699 -4040
rect 707 -4048 711 -4040
rect 716 -4048 720 -4040
rect 725 -4048 729 -4040
rect 737 -4048 741 -4040
rect 749 -4048 753 -4040
rect 757 -4048 761 -4040
rect 963 -4048 967 -4040
rect 972 -4048 976 -4040
rect 981 -4048 985 -4040
rect 989 -4048 993 -4040
rect 997 -4048 1001 -4040
rect 1009 -4048 1013 -4040
rect 1021 -4048 1025 -4040
rect 1030 -4048 1034 -4040
rect 1039 -4048 1043 -4040
rect 1051 -4048 1055 -4040
rect 1063 -4048 1067 -4040
rect 1072 -4048 1076 -4040
rect 1081 -4048 1085 -4040
rect 1093 -4048 1097 -4040
rect 1105 -4048 1109 -4040
rect 1114 -4048 1118 -4040
rect 1123 -4048 1127 -4040
rect 1135 -4048 1139 -4040
rect 1147 -4048 1151 -4040
rect 1155 -4048 1159 -4040
rect 1321 -4048 1325 -4040
rect 1330 -4048 1334 -4040
rect 1339 -4048 1343 -4040
rect 1347 -4048 1351 -4040
rect 1355 -4048 1359 -4040
rect 1367 -4048 1371 -4040
rect 1379 -4048 1383 -4040
rect 1388 -4048 1392 -4040
rect 1397 -4048 1401 -4040
rect 1409 -4048 1413 -4040
rect 1421 -4048 1425 -4040
rect 1430 -4048 1434 -4040
rect 1439 -4048 1443 -4040
rect 1451 -4048 1455 -4040
rect 1463 -4048 1467 -4040
rect 1472 -4048 1476 -4040
rect 1481 -4048 1485 -4040
rect 1493 -4048 1497 -4040
rect 1505 -4048 1509 -4040
rect 1513 -4048 1517 -4040
rect -1264 -4172 -1260 -4164
rect -1255 -4172 -1251 -4164
rect -1246 -4172 -1242 -4164
rect -1238 -4172 -1234 -4164
rect -1230 -4172 -1226 -4164
rect -1218 -4172 -1214 -4164
rect -1206 -4172 -1202 -4164
rect -1197 -4172 -1193 -4164
rect -1188 -4172 -1184 -4164
rect -1176 -4172 -1172 -4164
rect -1164 -4172 -1160 -4164
rect -1155 -4172 -1151 -4164
rect -1146 -4172 -1142 -4164
rect -1134 -4172 -1130 -4164
rect -1122 -4172 -1118 -4164
rect -1113 -4172 -1109 -4164
rect -1104 -4172 -1100 -4164
rect -1092 -4172 -1088 -4164
rect -1080 -4172 -1076 -4164
rect -1072 -4172 -1068 -4164
rect -1029 -4172 -1025 -4164
rect -1021 -4172 -1017 -4164
rect -935 -4172 -931 -4164
rect -926 -4172 -922 -4164
rect -917 -4172 -913 -4164
rect -909 -4172 -905 -4164
rect -901 -4172 -897 -4164
rect -889 -4172 -885 -4164
rect -877 -4172 -873 -4164
rect -868 -4172 -864 -4164
rect -859 -4172 -855 -4164
rect -847 -4172 -843 -4164
rect -835 -4172 -831 -4164
rect -826 -4172 -822 -4164
rect -817 -4172 -813 -4164
rect -805 -4172 -801 -4164
rect -793 -4172 -789 -4164
rect -784 -4172 -780 -4164
rect -775 -4172 -771 -4164
rect -763 -4172 -759 -4164
rect -751 -4172 -747 -4164
rect -743 -4172 -739 -4164
rect -577 -4172 -573 -4164
rect -568 -4172 -564 -4164
rect -559 -4172 -555 -4164
rect -551 -4172 -547 -4164
rect -543 -4172 -539 -4164
rect -531 -4172 -527 -4164
rect -519 -4172 -515 -4164
rect -510 -4172 -506 -4164
rect -501 -4172 -497 -4164
rect -489 -4172 -485 -4164
rect -477 -4172 -473 -4164
rect -468 -4172 -464 -4164
rect -459 -4172 -455 -4164
rect -447 -4172 -443 -4164
rect -435 -4172 -431 -4164
rect -426 -4172 -422 -4164
rect -417 -4172 -413 -4164
rect -405 -4172 -401 -4164
rect -393 -4172 -389 -4164
rect -385 -4172 -381 -4164
rect -332 -4172 -328 -4164
rect -324 -4172 -320 -4164
rect -219 -4172 -215 -4164
rect -210 -4172 -206 -4164
rect -201 -4172 -197 -4164
rect -193 -4172 -189 -4164
rect -185 -4172 -181 -4164
rect -173 -4172 -169 -4164
rect -161 -4172 -157 -4164
rect -152 -4172 -148 -4164
rect -143 -4172 -139 -4164
rect -131 -4172 -127 -4164
rect -119 -4172 -115 -4164
rect -110 -4172 -106 -4164
rect -101 -4172 -97 -4164
rect -89 -4172 -85 -4164
rect -77 -4172 -73 -4164
rect -68 -4172 -64 -4164
rect -59 -4172 -55 -4164
rect -47 -4172 -43 -4164
rect -35 -4172 -31 -4164
rect -27 -4172 -23 -4164
rect 456 -4172 460 -4164
rect 464 -4172 468 -4164
rect 1201 -4172 1205 -4164
rect 1209 -4172 1213 -4164
rect -1339 -4283 -1335 -4275
rect -1331 -4283 -1327 -4275
rect -1322 -4283 -1318 -4275
rect -1313 -4283 -1309 -4275
rect -1029 -4283 -1025 -4275
rect -1021 -4283 -1017 -4275
rect -935 -4283 -931 -4275
rect -927 -4283 -923 -4275
rect -918 -4283 -914 -4275
rect -909 -4283 -905 -4275
rect -673 -4291 -669 -4275
rect -665 -4291 -661 -4275
rect -577 -4283 -573 -4275
rect -569 -4283 -565 -4275
rect -560 -4283 -556 -4275
rect -551 -4283 -547 -4275
rect -332 -4283 -328 -4275
rect -324 -4283 -320 -4275
rect -219 -4283 -215 -4275
rect -211 -4283 -207 -4275
rect -202 -4283 -198 -4275
rect -193 -4283 -189 -4275
rect 209 -4283 213 -4275
rect 217 -4283 221 -4275
rect 226 -4283 230 -4275
rect 235 -4283 239 -4275
rect 456 -4283 460 -4275
rect 464 -4283 468 -4275
rect 565 -4283 569 -4275
rect 573 -4283 577 -4275
rect 582 -4283 586 -4275
rect 591 -4283 595 -4275
rect 860 -4291 864 -4275
rect 868 -4291 872 -4275
rect 963 -4283 967 -4275
rect 971 -4283 975 -4275
rect 980 -4283 984 -4275
rect 989 -4283 993 -4275
rect 1201 -4283 1205 -4275
rect 1209 -4283 1213 -4275
rect 1321 -4283 1325 -4275
rect 1329 -4283 1333 -4275
rect 1338 -4283 1342 -4275
rect 1347 -4283 1351 -4275
rect -1264 -4402 -1260 -4394
rect -1255 -4402 -1251 -4394
rect -1246 -4402 -1242 -4394
rect -1238 -4402 -1234 -4394
rect -1220 -4402 -1216 -4394
rect -1198 -4402 -1194 -4394
rect -1186 -4402 -1182 -4394
rect -1177 -4402 -1173 -4394
rect -1168 -4402 -1164 -4394
rect -935 -4402 -931 -4394
rect -926 -4402 -922 -4394
rect -917 -4402 -913 -4394
rect -909 -4402 -905 -4394
rect -900 -4402 -896 -4394
rect -891 -4402 -887 -4394
rect -883 -4402 -879 -4394
rect -865 -4402 -861 -4394
rect -843 -4402 -839 -4394
rect -831 -4402 -827 -4394
rect -822 -4402 -818 -4394
rect -813 -4402 -809 -4394
rect -805 -4402 -801 -4394
rect -787 -4402 -783 -4394
rect -765 -4402 -761 -4394
rect -753 -4402 -749 -4394
rect -741 -4402 -737 -4394
rect -729 -4402 -725 -4394
rect -721 -4402 -717 -4394
rect -704 -4402 -700 -4394
rect -695 -4402 -691 -4394
rect -577 -4402 -573 -4394
rect -568 -4402 -564 -4394
rect -559 -4402 -555 -4394
rect -551 -4402 -547 -4394
rect -542 -4402 -538 -4394
rect -533 -4402 -529 -4394
rect -525 -4402 -521 -4394
rect -507 -4402 -503 -4394
rect -485 -4402 -481 -4394
rect -473 -4402 -469 -4394
rect -464 -4402 -460 -4394
rect -455 -4402 -451 -4394
rect -447 -4402 -443 -4394
rect -429 -4402 -425 -4394
rect -407 -4402 -403 -4394
rect -395 -4402 -391 -4394
rect -383 -4402 -379 -4394
rect -371 -4402 -367 -4394
rect -363 -4402 -359 -4394
rect -346 -4402 -342 -4394
rect -337 -4402 -333 -4394
rect -219 -4402 -215 -4394
rect -210 -4402 -206 -4394
rect -201 -4402 -197 -4394
rect -193 -4402 -189 -4394
rect -184 -4402 -180 -4394
rect -175 -4402 -171 -4394
rect -167 -4402 -163 -4394
rect -149 -4402 -145 -4394
rect -127 -4402 -123 -4394
rect -115 -4402 -111 -4394
rect -106 -4402 -102 -4394
rect -97 -4402 -93 -4394
rect -89 -4402 -85 -4394
rect -71 -4402 -67 -4394
rect -49 -4402 -45 -4394
rect -37 -4402 -33 -4394
rect -25 -4402 -21 -4394
rect -13 -4402 -9 -4394
rect -5 -4402 -1 -4394
rect 12 -4402 16 -4394
rect 21 -4402 25 -4394
rect 209 -4402 213 -4394
rect 218 -4402 222 -4394
rect 227 -4402 231 -4394
rect 235 -4402 239 -4394
rect 244 -4402 248 -4394
rect 253 -4402 257 -4394
rect 261 -4402 265 -4394
rect 279 -4402 283 -4394
rect 301 -4402 305 -4394
rect 313 -4402 317 -4394
rect 322 -4402 326 -4394
rect 331 -4402 335 -4394
rect 339 -4402 343 -4394
rect 357 -4402 361 -4394
rect 379 -4402 383 -4394
rect 391 -4402 395 -4394
rect 403 -4402 407 -4394
rect 415 -4402 419 -4394
rect 423 -4402 427 -4394
rect 440 -4402 444 -4394
rect 449 -4402 453 -4394
rect 565 -4402 569 -4394
rect 574 -4402 578 -4394
rect 583 -4402 587 -4394
rect 591 -4402 595 -4394
rect 600 -4402 604 -4394
rect 609 -4402 613 -4394
rect 617 -4402 621 -4394
rect 635 -4402 639 -4394
rect 657 -4402 661 -4394
rect 669 -4402 673 -4394
rect 678 -4402 682 -4394
rect 687 -4402 691 -4394
rect 695 -4402 699 -4394
rect 713 -4402 717 -4394
rect 735 -4402 739 -4394
rect 747 -4402 751 -4394
rect 759 -4402 763 -4394
rect 771 -4402 775 -4394
rect 779 -4402 783 -4394
rect 796 -4402 800 -4394
rect 805 -4402 809 -4394
rect 963 -4402 967 -4394
rect 972 -4402 976 -4394
rect 981 -4402 985 -4394
rect 989 -4402 993 -4394
rect 998 -4402 1002 -4394
rect 1007 -4402 1011 -4394
rect 1015 -4402 1019 -4394
rect 1033 -4402 1037 -4394
rect 1055 -4402 1059 -4394
rect 1067 -4402 1071 -4394
rect 1076 -4402 1080 -4394
rect 1085 -4402 1089 -4394
rect 1093 -4402 1097 -4394
rect 1111 -4402 1115 -4394
rect 1133 -4402 1137 -4394
rect 1145 -4402 1149 -4394
rect 1157 -4402 1161 -4394
rect 1169 -4402 1173 -4394
rect 1177 -4402 1181 -4394
rect 1194 -4402 1198 -4394
rect 1203 -4402 1207 -4394
rect 1321 -4402 1325 -4394
rect 1330 -4402 1334 -4394
rect 1339 -4402 1343 -4394
rect 1347 -4402 1351 -4394
rect 1356 -4402 1360 -4394
rect 1365 -4402 1369 -4394
rect 1373 -4402 1377 -4394
rect 1391 -4402 1395 -4394
rect 1413 -4402 1417 -4394
rect 1425 -4402 1429 -4394
rect 1434 -4402 1438 -4394
rect 1443 -4402 1447 -4394
rect 1451 -4402 1455 -4394
rect 1469 -4402 1473 -4394
rect 1491 -4402 1495 -4394
rect 1503 -4402 1507 -4394
rect 1515 -4402 1519 -4394
rect 1527 -4402 1531 -4394
rect 1535 -4402 1539 -4394
rect 1552 -4402 1556 -4394
rect 1561 -4402 1565 -4394
rect -1264 -4525 -1260 -4517
rect -1255 -4525 -1251 -4517
rect -1246 -4525 -1242 -4517
rect -1238 -4525 -1234 -4517
rect -1230 -4525 -1226 -4517
rect -1218 -4525 -1214 -4517
rect -1206 -4525 -1202 -4517
rect -1197 -4525 -1193 -4517
rect -1188 -4525 -1184 -4517
rect -1176 -4525 -1172 -4517
rect -1164 -4525 -1160 -4517
rect -1155 -4525 -1151 -4517
rect -1146 -4525 -1142 -4517
rect -1134 -4525 -1130 -4517
rect -1122 -4525 -1118 -4517
rect -1113 -4525 -1109 -4517
rect -1104 -4525 -1100 -4517
rect -1092 -4525 -1088 -4517
rect -1080 -4525 -1076 -4517
rect -1072 -4525 -1068 -4517
rect -935 -4525 -931 -4517
rect -926 -4525 -922 -4517
rect -917 -4525 -913 -4517
rect -909 -4525 -905 -4517
rect -901 -4525 -897 -4517
rect -889 -4525 -885 -4517
rect -877 -4525 -873 -4517
rect -868 -4525 -864 -4517
rect -859 -4525 -855 -4517
rect -847 -4525 -843 -4517
rect -835 -4525 -831 -4517
rect -826 -4525 -822 -4517
rect -817 -4525 -813 -4517
rect -805 -4525 -801 -4517
rect -793 -4525 -789 -4517
rect -784 -4525 -780 -4517
rect -775 -4525 -771 -4517
rect -763 -4525 -759 -4517
rect -751 -4525 -747 -4517
rect -743 -4525 -739 -4517
rect -577 -4525 -573 -4517
rect -568 -4525 -564 -4517
rect -559 -4525 -555 -4517
rect -551 -4525 -547 -4517
rect -543 -4525 -539 -4517
rect -531 -4525 -527 -4517
rect -519 -4525 -515 -4517
rect -510 -4525 -506 -4517
rect -501 -4525 -497 -4517
rect -489 -4525 -485 -4517
rect -477 -4525 -473 -4517
rect -468 -4525 -464 -4517
rect -459 -4525 -455 -4517
rect -447 -4525 -443 -4517
rect -435 -4525 -431 -4517
rect -426 -4525 -422 -4517
rect -417 -4525 -413 -4517
rect -405 -4525 -401 -4517
rect -393 -4525 -389 -4517
rect -385 -4525 -381 -4517
rect -1264 -4646 -1260 -4638
rect -1255 -4646 -1251 -4638
rect -1246 -4646 -1242 -4638
rect -1238 -4646 -1234 -4638
rect -1230 -4646 -1226 -4638
rect -1218 -4646 -1214 -4638
rect -1206 -4646 -1202 -4638
rect -1197 -4646 -1193 -4638
rect -1188 -4646 -1184 -4638
rect -1176 -4646 -1172 -4638
rect -1164 -4646 -1160 -4638
rect -1155 -4646 -1151 -4638
rect -1146 -4646 -1142 -4638
rect -1134 -4646 -1130 -4638
rect -1122 -4646 -1118 -4638
rect -1113 -4646 -1109 -4638
rect -1104 -4646 -1100 -4638
rect -1092 -4646 -1088 -4638
rect -1080 -4646 -1076 -4638
rect -1072 -4646 -1068 -4638
rect -935 -4646 -931 -4638
rect -926 -4646 -922 -4638
rect -917 -4646 -913 -4638
rect -909 -4646 -905 -4638
rect -901 -4646 -897 -4638
rect -889 -4646 -885 -4638
rect -877 -4646 -873 -4638
rect -868 -4646 -864 -4638
rect -859 -4646 -855 -4638
rect -847 -4646 -843 -4638
rect -835 -4646 -831 -4638
rect -826 -4646 -822 -4638
rect -817 -4646 -813 -4638
rect -805 -4646 -801 -4638
rect -793 -4646 -789 -4638
rect -784 -4646 -780 -4638
rect -775 -4646 -771 -4638
rect -763 -4646 -759 -4638
rect -751 -4646 -747 -4638
rect -743 -4646 -739 -4638
rect -577 -4646 -573 -4638
rect -568 -4646 -564 -4638
rect -559 -4646 -555 -4638
rect -551 -4646 -547 -4638
rect -543 -4646 -539 -4638
rect -531 -4646 -527 -4638
rect -519 -4646 -515 -4638
rect -510 -4646 -506 -4638
rect -501 -4646 -497 -4638
rect -489 -4646 -485 -4638
rect -477 -4646 -473 -4638
rect -468 -4646 -464 -4638
rect -459 -4646 -455 -4638
rect -447 -4646 -443 -4638
rect -435 -4646 -431 -4638
rect -426 -4646 -422 -4638
rect -417 -4646 -413 -4638
rect -405 -4646 -401 -4638
rect -393 -4646 -389 -4638
rect -385 -4646 -381 -4638
rect -219 -4646 -215 -4638
rect -210 -4646 -206 -4638
rect -201 -4646 -197 -4638
rect -193 -4646 -189 -4638
rect -185 -4646 -181 -4638
rect -173 -4646 -169 -4638
rect -161 -4646 -157 -4638
rect -152 -4646 -148 -4638
rect -143 -4646 -139 -4638
rect -131 -4646 -127 -4638
rect -119 -4646 -115 -4638
rect -110 -4646 -106 -4638
rect -101 -4646 -97 -4638
rect -89 -4646 -85 -4638
rect -77 -4646 -73 -4638
rect -68 -4646 -64 -4638
rect -59 -4646 -55 -4638
rect -47 -4646 -43 -4638
rect -35 -4646 -31 -4638
rect -27 -4646 -23 -4638
rect 209 -4646 213 -4638
rect 218 -4646 222 -4638
rect 227 -4646 231 -4638
rect 235 -4646 239 -4638
rect 243 -4646 247 -4638
rect 255 -4646 259 -4638
rect 267 -4646 271 -4638
rect 276 -4646 280 -4638
rect 285 -4646 289 -4638
rect 297 -4646 301 -4638
rect 309 -4646 313 -4638
rect 318 -4646 322 -4638
rect 327 -4646 331 -4638
rect 339 -4646 343 -4638
rect 351 -4646 355 -4638
rect 360 -4646 364 -4638
rect 369 -4646 373 -4638
rect 381 -4646 385 -4638
rect 393 -4646 397 -4638
rect 401 -4646 405 -4638
rect 565 -4646 569 -4638
rect 574 -4646 578 -4638
rect 583 -4646 587 -4638
rect 591 -4646 595 -4638
rect 599 -4646 603 -4638
rect 611 -4646 615 -4638
rect 623 -4646 627 -4638
rect 632 -4646 636 -4638
rect 641 -4646 645 -4638
rect 653 -4646 657 -4638
rect 665 -4646 669 -4638
rect 674 -4646 678 -4638
rect 683 -4646 687 -4638
rect 695 -4646 699 -4638
rect 707 -4646 711 -4638
rect 716 -4646 720 -4638
rect 725 -4646 729 -4638
rect 737 -4646 741 -4638
rect 749 -4646 753 -4638
rect 757 -4646 761 -4638
rect 963 -4646 967 -4638
rect 972 -4646 976 -4638
rect 981 -4646 985 -4638
rect 989 -4646 993 -4638
rect 997 -4646 1001 -4638
rect 1009 -4646 1013 -4638
rect 1021 -4646 1025 -4638
rect 1030 -4646 1034 -4638
rect 1039 -4646 1043 -4638
rect 1051 -4646 1055 -4638
rect 1063 -4646 1067 -4638
rect 1072 -4646 1076 -4638
rect 1081 -4646 1085 -4638
rect 1093 -4646 1097 -4638
rect 1105 -4646 1109 -4638
rect 1114 -4646 1118 -4638
rect 1123 -4646 1127 -4638
rect 1135 -4646 1139 -4638
rect 1147 -4646 1151 -4638
rect 1155 -4646 1159 -4638
rect 1321 -4646 1325 -4638
rect 1330 -4646 1334 -4638
rect 1339 -4646 1343 -4638
rect 1347 -4646 1351 -4638
rect 1355 -4646 1359 -4638
rect 1367 -4646 1371 -4638
rect 1379 -4646 1383 -4638
rect 1388 -4646 1392 -4638
rect 1397 -4646 1401 -4638
rect 1409 -4646 1413 -4638
rect 1421 -4646 1425 -4638
rect 1430 -4646 1434 -4638
rect 1439 -4646 1443 -4638
rect 1451 -4646 1455 -4638
rect 1463 -4646 1467 -4638
rect 1472 -4646 1476 -4638
rect 1481 -4646 1485 -4638
rect 1493 -4646 1497 -4638
rect 1505 -4646 1509 -4638
rect 1513 -4646 1517 -4638
rect -1264 -4767 -1260 -4759
rect -1255 -4767 -1251 -4759
rect -1246 -4767 -1242 -4759
rect -1238 -4767 -1234 -4759
rect -1230 -4767 -1226 -4759
rect -1218 -4767 -1214 -4759
rect -1206 -4767 -1202 -4759
rect -1197 -4767 -1193 -4759
rect -1188 -4767 -1184 -4759
rect -1176 -4767 -1172 -4759
rect -1164 -4767 -1160 -4759
rect -1155 -4767 -1151 -4759
rect -1146 -4767 -1142 -4759
rect -1134 -4767 -1130 -4759
rect -1122 -4767 -1118 -4759
rect -1113 -4767 -1109 -4759
rect -1104 -4767 -1100 -4759
rect -1092 -4767 -1088 -4759
rect -1080 -4767 -1076 -4759
rect -1072 -4767 -1068 -4759
rect -935 -4767 -931 -4759
rect -926 -4767 -922 -4759
rect -917 -4767 -913 -4759
rect -909 -4767 -905 -4759
rect -901 -4767 -897 -4759
rect -889 -4767 -885 -4759
rect -877 -4767 -873 -4759
rect -868 -4767 -864 -4759
rect -859 -4767 -855 -4759
rect -847 -4767 -843 -4759
rect -835 -4767 -831 -4759
rect -826 -4767 -822 -4759
rect -817 -4767 -813 -4759
rect -805 -4767 -801 -4759
rect -793 -4767 -789 -4759
rect -784 -4767 -780 -4759
rect -775 -4767 -771 -4759
rect -763 -4767 -759 -4759
rect -751 -4767 -747 -4759
rect -743 -4767 -739 -4759
rect -577 -4767 -573 -4759
rect -568 -4767 -564 -4759
rect -559 -4767 -555 -4759
rect -551 -4767 -547 -4759
rect -543 -4767 -539 -4759
rect -531 -4767 -527 -4759
rect -519 -4767 -515 -4759
rect -510 -4767 -506 -4759
rect -501 -4767 -497 -4759
rect -489 -4767 -485 -4759
rect -477 -4767 -473 -4759
rect -468 -4767 -464 -4759
rect -459 -4767 -455 -4759
rect -447 -4767 -443 -4759
rect -435 -4767 -431 -4759
rect -426 -4767 -422 -4759
rect -417 -4767 -413 -4759
rect -405 -4767 -401 -4759
rect -393 -4767 -389 -4759
rect -385 -4767 -381 -4759
rect -219 -4767 -215 -4759
rect -210 -4767 -206 -4759
rect -201 -4767 -197 -4759
rect -193 -4767 -189 -4759
rect -185 -4767 -181 -4759
rect -173 -4767 -169 -4759
rect -161 -4767 -157 -4759
rect -152 -4767 -148 -4759
rect -143 -4767 -139 -4759
rect -131 -4767 -127 -4759
rect -119 -4767 -115 -4759
rect -110 -4767 -106 -4759
rect -101 -4767 -97 -4759
rect -89 -4767 -85 -4759
rect -77 -4767 -73 -4759
rect -68 -4767 -64 -4759
rect -59 -4767 -55 -4759
rect -47 -4767 -43 -4759
rect -35 -4767 -31 -4759
rect -27 -4767 -23 -4759
rect 90 -4791 94 -4759
rect 98 -4791 102 -4759
rect 209 -4767 213 -4759
rect 218 -4767 222 -4759
rect 227 -4767 231 -4759
rect 235 -4767 239 -4759
rect 243 -4767 247 -4759
rect 255 -4767 259 -4759
rect 267 -4767 271 -4759
rect 276 -4767 280 -4759
rect 285 -4767 289 -4759
rect 297 -4767 301 -4759
rect 309 -4767 313 -4759
rect 318 -4767 322 -4759
rect 327 -4767 331 -4759
rect 339 -4767 343 -4759
rect 351 -4767 355 -4759
rect 360 -4767 364 -4759
rect 369 -4767 373 -4759
rect 381 -4767 385 -4759
rect 393 -4767 397 -4759
rect 401 -4767 405 -4759
rect 565 -4767 569 -4759
rect 574 -4767 578 -4759
rect 583 -4767 587 -4759
rect 591 -4767 595 -4759
rect 599 -4767 603 -4759
rect 611 -4767 615 -4759
rect 623 -4767 627 -4759
rect 632 -4767 636 -4759
rect 641 -4767 645 -4759
rect 653 -4767 657 -4759
rect 665 -4767 669 -4759
rect 674 -4767 678 -4759
rect 683 -4767 687 -4759
rect 695 -4767 699 -4759
rect 707 -4767 711 -4759
rect 716 -4767 720 -4759
rect 725 -4767 729 -4759
rect 737 -4767 741 -4759
rect 749 -4767 753 -4759
rect 757 -4767 761 -4759
rect 963 -4767 967 -4759
rect 972 -4767 976 -4759
rect 981 -4767 985 -4759
rect 989 -4767 993 -4759
rect 997 -4767 1001 -4759
rect 1009 -4767 1013 -4759
rect 1021 -4767 1025 -4759
rect 1030 -4767 1034 -4759
rect 1039 -4767 1043 -4759
rect 1051 -4767 1055 -4759
rect 1063 -4767 1067 -4759
rect 1072 -4767 1076 -4759
rect 1081 -4767 1085 -4759
rect 1093 -4767 1097 -4759
rect 1105 -4767 1109 -4759
rect 1114 -4767 1118 -4759
rect 1123 -4767 1127 -4759
rect 1135 -4767 1139 -4759
rect 1147 -4767 1151 -4759
rect 1155 -4767 1159 -4759
rect 1321 -4767 1325 -4759
rect 1330 -4767 1334 -4759
rect 1339 -4767 1343 -4759
rect 1347 -4767 1351 -4759
rect 1355 -4767 1359 -4759
rect 1367 -4767 1371 -4759
rect 1379 -4767 1383 -4759
rect 1388 -4767 1392 -4759
rect 1397 -4767 1401 -4759
rect 1409 -4767 1413 -4759
rect 1421 -4767 1425 -4759
rect 1430 -4767 1434 -4759
rect 1439 -4767 1443 -4759
rect 1451 -4767 1455 -4759
rect 1463 -4767 1467 -4759
rect 1472 -4767 1476 -4759
rect 1481 -4767 1485 -4759
rect 1493 -4767 1497 -4759
rect 1505 -4767 1509 -4759
rect 1513 -4767 1517 -4759
rect -1264 -4885 -1260 -4877
rect -1255 -4885 -1251 -4877
rect -1246 -4885 -1242 -4877
rect -1238 -4885 -1234 -4877
rect -1230 -4885 -1226 -4877
rect -1218 -4885 -1214 -4877
rect -1206 -4885 -1202 -4877
rect -1197 -4885 -1193 -4877
rect -1188 -4885 -1184 -4877
rect -1176 -4885 -1172 -4877
rect -1164 -4885 -1160 -4877
rect -1155 -4885 -1151 -4877
rect -1146 -4885 -1142 -4877
rect -1134 -4885 -1130 -4877
rect -1122 -4885 -1118 -4877
rect -1113 -4885 -1109 -4877
rect -1104 -4885 -1100 -4877
rect -1092 -4885 -1088 -4877
rect -1080 -4885 -1076 -4877
rect -1072 -4885 -1068 -4877
rect -935 -4885 -931 -4877
rect -926 -4885 -922 -4877
rect -917 -4885 -913 -4877
rect -909 -4885 -905 -4877
rect -901 -4885 -897 -4877
rect -889 -4885 -885 -4877
rect -877 -4885 -873 -4877
rect -868 -4885 -864 -4877
rect -859 -4885 -855 -4877
rect -847 -4885 -843 -4877
rect -835 -4885 -831 -4877
rect -826 -4885 -822 -4877
rect -817 -4885 -813 -4877
rect -805 -4885 -801 -4877
rect -793 -4885 -789 -4877
rect -784 -4885 -780 -4877
rect -775 -4885 -771 -4877
rect -763 -4885 -759 -4877
rect -751 -4885 -747 -4877
rect -743 -4885 -739 -4877
rect -577 -4885 -573 -4877
rect -568 -4885 -564 -4877
rect -559 -4885 -555 -4877
rect -551 -4885 -547 -4877
rect -543 -4885 -539 -4877
rect -531 -4885 -527 -4877
rect -519 -4885 -515 -4877
rect -510 -4885 -506 -4877
rect -501 -4885 -497 -4877
rect -489 -4885 -485 -4877
rect -477 -4885 -473 -4877
rect -468 -4885 -464 -4877
rect -459 -4885 -455 -4877
rect -447 -4885 -443 -4877
rect -435 -4885 -431 -4877
rect -426 -4885 -422 -4877
rect -417 -4885 -413 -4877
rect -405 -4885 -401 -4877
rect -393 -4885 -389 -4877
rect -385 -4885 -381 -4877
rect -219 -4885 -215 -4877
rect -210 -4885 -206 -4877
rect -201 -4885 -197 -4877
rect -193 -4885 -189 -4877
rect -185 -4885 -181 -4877
rect -173 -4885 -169 -4877
rect -161 -4885 -157 -4877
rect -152 -4885 -148 -4877
rect -143 -4885 -139 -4877
rect -131 -4885 -127 -4877
rect -119 -4885 -115 -4877
rect -110 -4885 -106 -4877
rect -101 -4885 -97 -4877
rect -89 -4885 -85 -4877
rect -77 -4885 -73 -4877
rect -68 -4885 -64 -4877
rect -59 -4885 -55 -4877
rect -47 -4885 -43 -4877
rect -35 -4885 -31 -4877
rect -27 -4885 -23 -4877
rect 209 -4885 213 -4877
rect 218 -4885 222 -4877
rect 227 -4885 231 -4877
rect 235 -4885 239 -4877
rect 243 -4885 247 -4877
rect 255 -4885 259 -4877
rect 267 -4885 271 -4877
rect 276 -4885 280 -4877
rect 285 -4885 289 -4877
rect 297 -4885 301 -4877
rect 309 -4885 313 -4877
rect 318 -4885 322 -4877
rect 327 -4885 331 -4877
rect 339 -4885 343 -4877
rect 351 -4885 355 -4877
rect 360 -4885 364 -4877
rect 369 -4885 373 -4877
rect 381 -4885 385 -4877
rect 393 -4885 397 -4877
rect 401 -4885 405 -4877
rect -1339 -5002 -1335 -4994
rect -1331 -5002 -1327 -4994
rect -1322 -5002 -1318 -4994
rect -1313 -5002 -1309 -4994
rect -935 -5002 -931 -4994
rect -927 -5002 -923 -4994
rect -918 -5002 -914 -4994
rect -909 -5002 -905 -4994
rect -577 -5002 -573 -4994
rect -569 -5002 -565 -4994
rect -560 -5002 -556 -4994
rect -551 -5002 -547 -4994
rect -219 -5002 -215 -4994
rect -211 -5002 -207 -4994
rect -202 -5002 -198 -4994
rect -193 -5002 -189 -4994
rect 209 -5002 213 -4994
rect 217 -5002 221 -4994
rect 226 -5002 230 -4994
rect 235 -5002 239 -4994
rect 565 -5002 569 -4994
rect 573 -5002 577 -4994
rect 582 -5002 586 -4994
rect 591 -5002 595 -4994
rect 963 -5002 967 -4994
rect 971 -5002 975 -4994
rect 980 -5002 984 -4994
rect 989 -5002 993 -4994
rect 1321 -5002 1325 -4994
rect 1329 -5002 1333 -4994
rect 1338 -5002 1342 -4994
rect 1347 -5002 1351 -4994
rect -1264 -5121 -1260 -5113
rect -1255 -5121 -1251 -5113
rect -1246 -5121 -1242 -5113
rect -1238 -5121 -1234 -5113
rect -1220 -5121 -1216 -5113
rect -1198 -5121 -1194 -5113
rect -1186 -5121 -1182 -5113
rect -1177 -5121 -1173 -5113
rect -1168 -5121 -1164 -5113
rect -935 -5121 -931 -5113
rect -926 -5121 -922 -5113
rect -917 -5121 -913 -5113
rect -909 -5121 -905 -5113
rect -900 -5121 -896 -5113
rect -891 -5121 -887 -5113
rect -883 -5121 -879 -5113
rect -865 -5121 -861 -5113
rect -843 -5121 -839 -5113
rect -831 -5121 -827 -5113
rect -822 -5121 -818 -5113
rect -813 -5121 -809 -5113
rect -805 -5121 -801 -5113
rect -787 -5121 -783 -5113
rect -765 -5121 -761 -5113
rect -753 -5121 -749 -5113
rect -741 -5121 -737 -5113
rect -729 -5121 -725 -5113
rect -721 -5121 -717 -5113
rect -704 -5121 -700 -5113
rect -695 -5121 -691 -5113
rect -577 -5121 -573 -5113
rect -568 -5121 -564 -5113
rect -559 -5121 -555 -5113
rect -551 -5121 -547 -5113
rect -542 -5121 -538 -5113
rect -533 -5121 -529 -5113
rect -525 -5121 -521 -5113
rect -507 -5121 -503 -5113
rect -485 -5121 -481 -5113
rect -473 -5121 -469 -5113
rect -464 -5121 -460 -5113
rect -455 -5121 -451 -5113
rect -447 -5121 -443 -5113
rect -429 -5121 -425 -5113
rect -407 -5121 -403 -5113
rect -395 -5121 -391 -5113
rect -383 -5121 -379 -5113
rect -371 -5121 -367 -5113
rect -363 -5121 -359 -5113
rect -346 -5121 -342 -5113
rect -337 -5121 -333 -5113
rect -219 -5121 -215 -5113
rect -210 -5121 -206 -5113
rect -201 -5121 -197 -5113
rect -193 -5121 -189 -5113
rect -184 -5121 -180 -5113
rect -175 -5121 -171 -5113
rect -167 -5121 -163 -5113
rect -149 -5121 -145 -5113
rect -127 -5121 -123 -5113
rect -115 -5121 -111 -5113
rect -106 -5121 -102 -5113
rect -97 -5121 -93 -5113
rect -89 -5121 -85 -5113
rect -71 -5121 -67 -5113
rect -49 -5121 -45 -5113
rect -37 -5121 -33 -5113
rect -25 -5121 -21 -5113
rect -13 -5121 -9 -5113
rect -5 -5121 -1 -5113
rect 12 -5121 16 -5113
rect 21 -5121 25 -5113
rect 209 -5121 213 -5113
rect 218 -5121 222 -5113
rect 227 -5121 231 -5113
rect 235 -5121 239 -5113
rect 244 -5121 248 -5113
rect 253 -5121 257 -5113
rect 261 -5121 265 -5113
rect 279 -5121 283 -5113
rect 301 -5121 305 -5113
rect 313 -5121 317 -5113
rect 322 -5121 326 -5113
rect 331 -5121 335 -5113
rect 339 -5121 343 -5113
rect 357 -5121 361 -5113
rect 379 -5121 383 -5113
rect 391 -5121 395 -5113
rect 403 -5121 407 -5113
rect 415 -5121 419 -5113
rect 423 -5121 427 -5113
rect 440 -5121 444 -5113
rect 449 -5121 453 -5113
rect 565 -5121 569 -5113
rect 574 -5121 578 -5113
rect 583 -5121 587 -5113
rect 591 -5121 595 -5113
rect 600 -5121 604 -5113
rect 609 -5121 613 -5113
rect 617 -5121 621 -5113
rect 635 -5121 639 -5113
rect 657 -5121 661 -5113
rect 669 -5121 673 -5113
rect 678 -5121 682 -5113
rect 687 -5121 691 -5113
rect 695 -5121 699 -5113
rect 713 -5121 717 -5113
rect 735 -5121 739 -5113
rect 747 -5121 751 -5113
rect 759 -5121 763 -5113
rect 771 -5121 775 -5113
rect 779 -5121 783 -5113
rect 796 -5121 800 -5113
rect 805 -5121 809 -5113
rect 963 -5121 967 -5113
rect 972 -5121 976 -5113
rect 981 -5121 985 -5113
rect 989 -5121 993 -5113
rect 998 -5121 1002 -5113
rect 1007 -5121 1011 -5113
rect 1015 -5121 1019 -5113
rect 1033 -5121 1037 -5113
rect 1055 -5121 1059 -5113
rect 1067 -5121 1071 -5113
rect 1076 -5121 1080 -5113
rect 1085 -5121 1089 -5113
rect 1093 -5121 1097 -5113
rect 1111 -5121 1115 -5113
rect 1133 -5121 1137 -5113
rect 1145 -5121 1149 -5113
rect 1157 -5121 1161 -5113
rect 1169 -5121 1173 -5113
rect 1177 -5121 1181 -5113
rect 1194 -5121 1198 -5113
rect 1203 -5121 1207 -5113
rect 1321 -5121 1325 -5113
rect 1330 -5121 1334 -5113
rect 1339 -5121 1343 -5113
rect 1347 -5121 1351 -5113
rect 1356 -5121 1360 -5113
rect 1365 -5121 1369 -5113
rect 1373 -5121 1377 -5113
rect 1391 -5121 1395 -5113
rect 1413 -5121 1417 -5113
rect 1425 -5121 1429 -5113
rect 1434 -5121 1438 -5113
rect 1443 -5121 1447 -5113
rect 1451 -5121 1455 -5113
rect 1469 -5121 1473 -5113
rect 1491 -5121 1495 -5113
rect 1503 -5121 1507 -5113
rect 1515 -5121 1519 -5113
rect 1527 -5121 1531 -5113
rect 1535 -5121 1539 -5113
rect 1552 -5121 1556 -5113
rect 1561 -5121 1565 -5113
rect -1264 -5240 -1260 -5232
rect -1255 -5240 -1251 -5232
rect -1246 -5240 -1242 -5232
rect -1238 -5240 -1234 -5232
rect -1230 -5240 -1226 -5232
rect -1218 -5240 -1214 -5232
rect -1206 -5240 -1202 -5232
rect -1197 -5240 -1193 -5232
rect -1188 -5240 -1184 -5232
rect -1176 -5240 -1172 -5232
rect -1164 -5240 -1160 -5232
rect -1155 -5240 -1151 -5232
rect -1146 -5240 -1142 -5232
rect -1134 -5240 -1130 -5232
rect -1122 -5240 -1118 -5232
rect -1113 -5240 -1109 -5232
rect -1104 -5240 -1100 -5232
rect -1092 -5240 -1088 -5232
rect -1080 -5240 -1076 -5232
rect -1072 -5240 -1068 -5232
rect -935 -5240 -931 -5232
rect -926 -5240 -922 -5232
rect -917 -5240 -913 -5232
rect -909 -5240 -905 -5232
rect -901 -5240 -897 -5232
rect -889 -5240 -885 -5232
rect -877 -5240 -873 -5232
rect -868 -5240 -864 -5232
rect -859 -5240 -855 -5232
rect -847 -5240 -843 -5232
rect -835 -5240 -831 -5232
rect -826 -5240 -822 -5232
rect -817 -5240 -813 -5232
rect -805 -5240 -801 -5232
rect -793 -5240 -789 -5232
rect -784 -5240 -780 -5232
rect -775 -5240 -771 -5232
rect -763 -5240 -759 -5232
rect -751 -5240 -747 -5232
rect -743 -5240 -739 -5232
rect -1264 -5361 -1260 -5353
rect -1255 -5361 -1251 -5353
rect -1246 -5361 -1242 -5353
rect -1238 -5361 -1234 -5353
rect -1230 -5361 -1226 -5353
rect -1218 -5361 -1214 -5353
rect -1206 -5361 -1202 -5353
rect -1197 -5361 -1193 -5353
rect -1188 -5361 -1184 -5353
rect -1176 -5361 -1172 -5353
rect -1164 -5361 -1160 -5353
rect -1155 -5361 -1151 -5353
rect -1146 -5361 -1142 -5353
rect -1134 -5361 -1130 -5353
rect -1122 -5361 -1118 -5353
rect -1113 -5361 -1109 -5353
rect -1104 -5361 -1100 -5353
rect -1092 -5361 -1088 -5353
rect -1080 -5361 -1076 -5353
rect -1072 -5361 -1068 -5353
rect -1026 -5361 -1022 -5353
rect -1018 -5361 -1014 -5353
rect -935 -5361 -931 -5353
rect -926 -5361 -922 -5353
rect -917 -5361 -913 -5353
rect -909 -5361 -905 -5353
rect -901 -5361 -897 -5353
rect -889 -5361 -885 -5353
rect -877 -5361 -873 -5353
rect -868 -5361 -864 -5353
rect -859 -5361 -855 -5353
rect -847 -5361 -843 -5353
rect -835 -5361 -831 -5353
rect -826 -5361 -822 -5353
rect -817 -5361 -813 -5353
rect -805 -5361 -801 -5353
rect -793 -5361 -789 -5353
rect -784 -5361 -780 -5353
rect -775 -5361 -771 -5353
rect -763 -5361 -759 -5353
rect -751 -5361 -747 -5353
rect -743 -5361 -739 -5353
rect -673 -5369 -669 -5353
rect -665 -5369 -661 -5353
rect -577 -5361 -573 -5353
rect -568 -5361 -564 -5353
rect -559 -5361 -555 -5353
rect -551 -5361 -547 -5353
rect -543 -5361 -539 -5353
rect -531 -5361 -527 -5353
rect -519 -5361 -515 -5353
rect -510 -5361 -506 -5353
rect -501 -5361 -497 -5353
rect -489 -5361 -485 -5353
rect -477 -5361 -473 -5353
rect -468 -5361 -464 -5353
rect -459 -5361 -455 -5353
rect -447 -5361 -443 -5353
rect -435 -5361 -431 -5353
rect -426 -5361 -422 -5353
rect -417 -5361 -413 -5353
rect -405 -5361 -401 -5353
rect -393 -5361 -389 -5353
rect -385 -5361 -381 -5353
rect -327 -5361 -323 -5353
rect -319 -5361 -315 -5353
rect -219 -5361 -215 -5353
rect -210 -5361 -206 -5353
rect -201 -5361 -197 -5353
rect -193 -5361 -189 -5353
rect -185 -5361 -181 -5353
rect -173 -5361 -169 -5353
rect -161 -5361 -157 -5353
rect -152 -5361 -148 -5353
rect -143 -5361 -139 -5353
rect -131 -5361 -127 -5353
rect -119 -5361 -115 -5353
rect -110 -5361 -106 -5353
rect -101 -5361 -97 -5353
rect -89 -5361 -85 -5353
rect -77 -5361 -73 -5353
rect -68 -5361 -64 -5353
rect -59 -5361 -55 -5353
rect -47 -5361 -43 -5353
rect -35 -5361 -31 -5353
rect -27 -5361 -23 -5353
rect 209 -5361 213 -5353
rect 218 -5361 222 -5353
rect 227 -5361 231 -5353
rect 235 -5361 239 -5353
rect 243 -5361 247 -5353
rect 255 -5361 259 -5353
rect 267 -5361 271 -5353
rect 276 -5361 280 -5353
rect 285 -5361 289 -5353
rect 297 -5361 301 -5353
rect 309 -5361 313 -5353
rect 318 -5361 322 -5353
rect 327 -5361 331 -5353
rect 339 -5361 343 -5353
rect 351 -5361 355 -5353
rect 360 -5361 364 -5353
rect 369 -5361 373 -5353
rect 381 -5361 385 -5353
rect 393 -5361 397 -5353
rect 401 -5361 405 -5353
rect 466 -5361 470 -5353
rect 474 -5361 478 -5353
rect 565 -5361 569 -5353
rect 574 -5361 578 -5353
rect 583 -5361 587 -5353
rect 591 -5361 595 -5353
rect 599 -5361 603 -5353
rect 611 -5361 615 -5353
rect 623 -5361 627 -5353
rect 632 -5361 636 -5353
rect 641 -5361 645 -5353
rect 653 -5361 657 -5353
rect 665 -5361 669 -5353
rect 674 -5361 678 -5353
rect 683 -5361 687 -5353
rect 695 -5361 699 -5353
rect 707 -5361 711 -5353
rect 716 -5361 720 -5353
rect 725 -5361 729 -5353
rect 737 -5361 741 -5353
rect 749 -5361 753 -5353
rect 757 -5361 761 -5353
rect 867 -5369 871 -5353
rect 875 -5369 879 -5353
rect 963 -5361 967 -5353
rect 972 -5361 976 -5353
rect 981 -5361 985 -5353
rect 989 -5361 993 -5353
rect 997 -5361 1001 -5353
rect 1009 -5361 1013 -5353
rect 1021 -5361 1025 -5353
rect 1030 -5361 1034 -5353
rect 1039 -5361 1043 -5353
rect 1051 -5361 1055 -5353
rect 1063 -5361 1067 -5353
rect 1072 -5361 1076 -5353
rect 1081 -5361 1085 -5353
rect 1093 -5361 1097 -5353
rect 1105 -5361 1109 -5353
rect 1114 -5361 1118 -5353
rect 1123 -5361 1127 -5353
rect 1135 -5361 1139 -5353
rect 1147 -5361 1151 -5353
rect 1155 -5361 1159 -5353
rect 1210 -5361 1214 -5353
rect 1218 -5361 1222 -5353
rect 1321 -5361 1325 -5353
rect 1330 -5361 1334 -5353
rect 1339 -5361 1343 -5353
rect 1347 -5361 1351 -5353
rect 1355 -5361 1359 -5353
rect 1367 -5361 1371 -5353
rect 1379 -5361 1383 -5353
rect 1388 -5361 1392 -5353
rect 1397 -5361 1401 -5353
rect 1409 -5361 1413 -5353
rect 1421 -5361 1425 -5353
rect 1430 -5361 1434 -5353
rect 1439 -5361 1443 -5353
rect 1451 -5361 1455 -5353
rect 1463 -5361 1467 -5353
rect 1472 -5361 1476 -5353
rect 1481 -5361 1485 -5353
rect 1493 -5361 1497 -5353
rect 1505 -5361 1509 -5353
rect 1513 -5361 1517 -5353
rect -1264 -5481 -1260 -5473
rect -1255 -5481 -1251 -5473
rect -1246 -5481 -1242 -5473
rect -1238 -5481 -1234 -5473
rect -1230 -5481 -1226 -5473
rect -1218 -5481 -1214 -5473
rect -1206 -5481 -1202 -5473
rect -1197 -5481 -1193 -5473
rect -1188 -5481 -1184 -5473
rect -1176 -5481 -1172 -5473
rect -1164 -5481 -1160 -5473
rect -1155 -5481 -1151 -5473
rect -1146 -5481 -1142 -5473
rect -1134 -5481 -1130 -5473
rect -1122 -5481 -1118 -5473
rect -1113 -5481 -1109 -5473
rect -1104 -5481 -1100 -5473
rect -1092 -5481 -1088 -5473
rect -1080 -5481 -1076 -5473
rect -1072 -5481 -1068 -5473
rect -1026 -5481 -1022 -5473
rect -1018 -5481 -1014 -5473
rect -935 -5481 -931 -5473
rect -926 -5481 -922 -5473
rect -917 -5481 -913 -5473
rect -909 -5481 -905 -5473
rect -901 -5481 -897 -5473
rect -889 -5481 -885 -5473
rect -877 -5481 -873 -5473
rect -868 -5481 -864 -5473
rect -859 -5481 -855 -5473
rect -847 -5481 -843 -5473
rect -835 -5481 -831 -5473
rect -826 -5481 -822 -5473
rect -817 -5481 -813 -5473
rect -805 -5481 -801 -5473
rect -793 -5481 -789 -5473
rect -784 -5481 -780 -5473
rect -775 -5481 -771 -5473
rect -763 -5481 -759 -5473
rect -751 -5481 -747 -5473
rect -743 -5481 -739 -5473
rect -577 -5481 -573 -5473
rect -568 -5481 -564 -5473
rect -559 -5481 -555 -5473
rect -551 -5481 -547 -5473
rect -543 -5481 -539 -5473
rect -531 -5481 -527 -5473
rect -519 -5481 -515 -5473
rect -510 -5481 -506 -5473
rect -501 -5481 -497 -5473
rect -489 -5481 -485 -5473
rect -477 -5481 -473 -5473
rect -468 -5481 -464 -5473
rect -459 -5481 -455 -5473
rect -447 -5481 -443 -5473
rect -435 -5481 -431 -5473
rect -426 -5481 -422 -5473
rect -417 -5481 -413 -5473
rect -405 -5481 -401 -5473
rect -393 -5481 -389 -5473
rect -385 -5481 -381 -5473
rect -327 -5481 -323 -5473
rect -319 -5481 -315 -5473
rect -219 -5481 -215 -5473
rect -210 -5481 -206 -5473
rect -201 -5481 -197 -5473
rect -193 -5481 -189 -5473
rect -185 -5481 -181 -5473
rect -173 -5481 -169 -5473
rect -161 -5481 -157 -5473
rect -152 -5481 -148 -5473
rect -143 -5481 -139 -5473
rect -131 -5481 -127 -5473
rect -119 -5481 -115 -5473
rect -110 -5481 -106 -5473
rect -101 -5481 -97 -5473
rect -89 -5481 -85 -5473
rect -77 -5481 -73 -5473
rect -68 -5481 -64 -5473
rect -59 -5481 -55 -5473
rect -47 -5481 -43 -5473
rect -35 -5481 -31 -5473
rect -27 -5481 -23 -5473
rect 209 -5481 213 -5473
rect 218 -5481 222 -5473
rect 227 -5481 231 -5473
rect 235 -5481 239 -5473
rect 243 -5481 247 -5473
rect 255 -5481 259 -5473
rect 267 -5481 271 -5473
rect 276 -5481 280 -5473
rect 285 -5481 289 -5473
rect 297 -5481 301 -5473
rect 309 -5481 313 -5473
rect 318 -5481 322 -5473
rect 327 -5481 331 -5473
rect 339 -5481 343 -5473
rect 351 -5481 355 -5473
rect 360 -5481 364 -5473
rect 369 -5481 373 -5473
rect 381 -5481 385 -5473
rect 393 -5481 397 -5473
rect 401 -5481 405 -5473
rect 466 -5481 470 -5473
rect 474 -5481 478 -5473
rect 565 -5481 569 -5473
rect 574 -5481 578 -5473
rect 583 -5481 587 -5473
rect 591 -5481 595 -5473
rect 599 -5481 603 -5473
rect 611 -5481 615 -5473
rect 623 -5481 627 -5473
rect 632 -5481 636 -5473
rect 641 -5481 645 -5473
rect 653 -5481 657 -5473
rect 665 -5481 669 -5473
rect 674 -5481 678 -5473
rect 683 -5481 687 -5473
rect 695 -5481 699 -5473
rect 707 -5481 711 -5473
rect 716 -5481 720 -5473
rect 725 -5481 729 -5473
rect 737 -5481 741 -5473
rect 749 -5481 753 -5473
rect 757 -5481 761 -5473
rect 963 -5481 967 -5473
rect 972 -5481 976 -5473
rect 981 -5481 985 -5473
rect 989 -5481 993 -5473
rect 997 -5481 1001 -5473
rect 1009 -5481 1013 -5473
rect 1021 -5481 1025 -5473
rect 1030 -5481 1034 -5473
rect 1039 -5481 1043 -5473
rect 1051 -5481 1055 -5473
rect 1063 -5481 1067 -5473
rect 1072 -5481 1076 -5473
rect 1081 -5481 1085 -5473
rect 1093 -5481 1097 -5473
rect 1105 -5481 1109 -5473
rect 1114 -5481 1118 -5473
rect 1123 -5481 1127 -5473
rect 1135 -5481 1139 -5473
rect 1147 -5481 1151 -5473
rect 1155 -5481 1159 -5473
rect 1210 -5481 1214 -5473
rect 1218 -5481 1222 -5473
rect 1321 -5481 1325 -5473
rect 1330 -5481 1334 -5473
rect 1339 -5481 1343 -5473
rect 1347 -5481 1351 -5473
rect 1355 -5481 1359 -5473
rect 1367 -5481 1371 -5473
rect 1379 -5481 1383 -5473
rect 1388 -5481 1392 -5473
rect 1397 -5481 1401 -5473
rect 1409 -5481 1413 -5473
rect 1421 -5481 1425 -5473
rect 1430 -5481 1434 -5473
rect 1439 -5481 1443 -5473
rect 1451 -5481 1455 -5473
rect 1463 -5481 1467 -5473
rect 1472 -5481 1476 -5473
rect 1481 -5481 1485 -5473
rect 1493 -5481 1497 -5473
rect 1505 -5481 1509 -5473
rect 1513 -5481 1517 -5473
rect -1264 -5598 -1260 -5590
rect -1255 -5598 -1251 -5590
rect -1246 -5598 -1242 -5590
rect -1238 -5598 -1234 -5590
rect -1230 -5598 -1226 -5590
rect -1218 -5598 -1214 -5590
rect -1206 -5598 -1202 -5590
rect -1197 -5598 -1193 -5590
rect -1188 -5598 -1184 -5590
rect -1176 -5598 -1172 -5590
rect -1164 -5598 -1160 -5590
rect -1155 -5598 -1151 -5590
rect -1146 -5598 -1142 -5590
rect -1134 -5598 -1130 -5590
rect -1122 -5598 -1118 -5590
rect -1113 -5598 -1109 -5590
rect -1104 -5598 -1100 -5590
rect -1092 -5598 -1088 -5590
rect -1080 -5598 -1076 -5590
rect -1072 -5598 -1068 -5590
rect -935 -5598 -931 -5590
rect -926 -5598 -922 -5590
rect -917 -5598 -913 -5590
rect -909 -5598 -905 -5590
rect -901 -5598 -897 -5590
rect -889 -5598 -885 -5590
rect -877 -5598 -873 -5590
rect -868 -5598 -864 -5590
rect -859 -5598 -855 -5590
rect -847 -5598 -843 -5590
rect -835 -5598 -831 -5590
rect -826 -5598 -822 -5590
rect -817 -5598 -813 -5590
rect -805 -5598 -801 -5590
rect -793 -5598 -789 -5590
rect -784 -5598 -780 -5590
rect -775 -5598 -771 -5590
rect -763 -5598 -759 -5590
rect -751 -5598 -747 -5590
rect -743 -5598 -739 -5590
rect -577 -5598 -573 -5590
rect -568 -5598 -564 -5590
rect -559 -5598 -555 -5590
rect -551 -5598 -547 -5590
rect -543 -5598 -539 -5590
rect -531 -5598 -527 -5590
rect -519 -5598 -515 -5590
rect -510 -5598 -506 -5590
rect -501 -5598 -497 -5590
rect -489 -5598 -485 -5590
rect -477 -5598 -473 -5590
rect -468 -5598 -464 -5590
rect -459 -5598 -455 -5590
rect -447 -5598 -443 -5590
rect -435 -5598 -431 -5590
rect -426 -5598 -422 -5590
rect -417 -5598 -413 -5590
rect -405 -5598 -401 -5590
rect -393 -5598 -389 -5590
rect -385 -5598 -381 -5590
rect -219 -5598 -215 -5590
rect -210 -5598 -206 -5590
rect -201 -5598 -197 -5590
rect -193 -5598 -189 -5590
rect -185 -5598 -181 -5590
rect -173 -5598 -169 -5590
rect -161 -5598 -157 -5590
rect -152 -5598 -148 -5590
rect -143 -5598 -139 -5590
rect -131 -5598 -127 -5590
rect -119 -5598 -115 -5590
rect -110 -5598 -106 -5590
rect -101 -5598 -97 -5590
rect -89 -5598 -85 -5590
rect -77 -5598 -73 -5590
rect -68 -5598 -64 -5590
rect -59 -5598 -55 -5590
rect -47 -5598 -43 -5590
rect -35 -5598 -31 -5590
rect -27 -5598 -23 -5590
rect 209 -5598 213 -5590
rect 218 -5598 222 -5590
rect 227 -5598 231 -5590
rect 235 -5598 239 -5590
rect 243 -5598 247 -5590
rect 255 -5598 259 -5590
rect 267 -5598 271 -5590
rect 276 -5598 280 -5590
rect 285 -5598 289 -5590
rect 297 -5598 301 -5590
rect 309 -5598 313 -5590
rect 318 -5598 322 -5590
rect 327 -5598 331 -5590
rect 339 -5598 343 -5590
rect 351 -5598 355 -5590
rect 360 -5598 364 -5590
rect 369 -5598 373 -5590
rect 381 -5598 385 -5590
rect 393 -5598 397 -5590
rect 401 -5598 405 -5590
rect 565 -5598 569 -5590
rect 574 -5598 578 -5590
rect 583 -5598 587 -5590
rect 591 -5598 595 -5590
rect 599 -5598 603 -5590
rect 611 -5598 615 -5590
rect 623 -5598 627 -5590
rect 632 -5598 636 -5590
rect 641 -5598 645 -5590
rect 653 -5598 657 -5590
rect 665 -5598 669 -5590
rect 674 -5598 678 -5590
rect 683 -5598 687 -5590
rect 695 -5598 699 -5590
rect 707 -5598 711 -5590
rect 716 -5598 720 -5590
rect 725 -5598 729 -5590
rect 737 -5598 741 -5590
rect 749 -5598 753 -5590
rect 757 -5598 761 -5590
rect -1339 -5715 -1335 -5707
rect -1331 -5715 -1327 -5707
rect -1322 -5715 -1318 -5707
rect -1313 -5715 -1309 -5707
rect -935 -5715 -931 -5707
rect -927 -5715 -923 -5707
rect -918 -5715 -914 -5707
rect -909 -5715 -905 -5707
rect -577 -5715 -573 -5707
rect -569 -5715 -565 -5707
rect -560 -5715 -556 -5707
rect -551 -5715 -547 -5707
rect -219 -5715 -215 -5707
rect -211 -5715 -207 -5707
rect -202 -5715 -198 -5707
rect -193 -5715 -189 -5707
rect 209 -5715 213 -5707
rect 217 -5715 221 -5707
rect 226 -5715 230 -5707
rect 235 -5715 239 -5707
rect 565 -5715 569 -5707
rect 573 -5715 577 -5707
rect 582 -5715 586 -5707
rect 591 -5715 595 -5707
rect 963 -5715 967 -5707
rect 971 -5715 975 -5707
rect 980 -5715 984 -5707
rect 989 -5715 993 -5707
rect 1321 -5715 1325 -5707
rect 1329 -5715 1333 -5707
rect 1338 -5715 1342 -5707
rect 1347 -5715 1351 -5707
rect -1264 -5834 -1260 -5826
rect -1255 -5834 -1251 -5826
rect -1246 -5834 -1242 -5826
rect -1238 -5834 -1234 -5826
rect -1220 -5834 -1216 -5826
rect -1198 -5834 -1194 -5826
rect -1186 -5834 -1182 -5826
rect -1177 -5834 -1173 -5826
rect -1168 -5834 -1164 -5826
rect -935 -5834 -931 -5826
rect -926 -5834 -922 -5826
rect -917 -5834 -913 -5826
rect -909 -5834 -905 -5826
rect -900 -5834 -896 -5826
rect -891 -5834 -887 -5826
rect -883 -5834 -879 -5826
rect -865 -5834 -861 -5826
rect -843 -5834 -839 -5826
rect -831 -5834 -827 -5826
rect -822 -5834 -818 -5826
rect -813 -5834 -809 -5826
rect -805 -5834 -801 -5826
rect -787 -5834 -783 -5826
rect -765 -5834 -761 -5826
rect -753 -5834 -749 -5826
rect -741 -5834 -737 -5826
rect -729 -5834 -725 -5826
rect -721 -5834 -717 -5826
rect -704 -5834 -700 -5826
rect -695 -5834 -691 -5826
rect -577 -5834 -573 -5826
rect -568 -5834 -564 -5826
rect -559 -5834 -555 -5826
rect -551 -5834 -547 -5826
rect -542 -5834 -538 -5826
rect -533 -5834 -529 -5826
rect -525 -5834 -521 -5826
rect -507 -5834 -503 -5826
rect -485 -5834 -481 -5826
rect -473 -5834 -469 -5826
rect -464 -5834 -460 -5826
rect -455 -5834 -451 -5826
rect -447 -5834 -443 -5826
rect -429 -5834 -425 -5826
rect -407 -5834 -403 -5826
rect -395 -5834 -391 -5826
rect -383 -5834 -379 -5826
rect -371 -5834 -367 -5826
rect -363 -5834 -359 -5826
rect -346 -5834 -342 -5826
rect -337 -5834 -333 -5826
rect -219 -5834 -215 -5826
rect -210 -5834 -206 -5826
rect -201 -5834 -197 -5826
rect -193 -5834 -189 -5826
rect -184 -5834 -180 -5826
rect -175 -5834 -171 -5826
rect -167 -5834 -163 -5826
rect -149 -5834 -145 -5826
rect -127 -5834 -123 -5826
rect -115 -5834 -111 -5826
rect -106 -5834 -102 -5826
rect -97 -5834 -93 -5826
rect -89 -5834 -85 -5826
rect -71 -5834 -67 -5826
rect -49 -5834 -45 -5826
rect -37 -5834 -33 -5826
rect -25 -5834 -21 -5826
rect -13 -5834 -9 -5826
rect -5 -5834 -1 -5826
rect 12 -5834 16 -5826
rect 21 -5834 25 -5826
rect 209 -5834 213 -5826
rect 218 -5834 222 -5826
rect 227 -5834 231 -5826
rect 235 -5834 239 -5826
rect 244 -5834 248 -5826
rect 253 -5834 257 -5826
rect 261 -5834 265 -5826
rect 279 -5834 283 -5826
rect 301 -5834 305 -5826
rect 313 -5834 317 -5826
rect 322 -5834 326 -5826
rect 331 -5834 335 -5826
rect 339 -5834 343 -5826
rect 357 -5834 361 -5826
rect 379 -5834 383 -5826
rect 391 -5834 395 -5826
rect 403 -5834 407 -5826
rect 415 -5834 419 -5826
rect 423 -5834 427 -5826
rect 440 -5834 444 -5826
rect 449 -5834 453 -5826
rect 565 -5834 569 -5826
rect 574 -5834 578 -5826
rect 583 -5834 587 -5826
rect 591 -5834 595 -5826
rect 600 -5834 604 -5826
rect 609 -5834 613 -5826
rect 617 -5834 621 -5826
rect 635 -5834 639 -5826
rect 657 -5834 661 -5826
rect 669 -5834 673 -5826
rect 678 -5834 682 -5826
rect 687 -5834 691 -5826
rect 695 -5834 699 -5826
rect 713 -5834 717 -5826
rect 735 -5834 739 -5826
rect 747 -5834 751 -5826
rect 759 -5834 763 -5826
rect 771 -5834 775 -5826
rect 779 -5834 783 -5826
rect 796 -5834 800 -5826
rect 805 -5834 809 -5826
rect 963 -5834 967 -5826
rect 972 -5834 976 -5826
rect 981 -5834 985 -5826
rect 989 -5834 993 -5826
rect 998 -5834 1002 -5826
rect 1007 -5834 1011 -5826
rect 1015 -5834 1019 -5826
rect 1033 -5834 1037 -5826
rect 1055 -5834 1059 -5826
rect 1067 -5834 1071 -5826
rect 1076 -5834 1080 -5826
rect 1085 -5834 1089 -5826
rect 1093 -5834 1097 -5826
rect 1111 -5834 1115 -5826
rect 1133 -5834 1137 -5826
rect 1145 -5834 1149 -5826
rect 1157 -5834 1161 -5826
rect 1169 -5834 1173 -5826
rect 1177 -5834 1181 -5826
rect 1194 -5834 1198 -5826
rect 1203 -5834 1207 -5826
rect 1321 -5834 1325 -5826
rect 1330 -5834 1334 -5826
rect 1339 -5834 1343 -5826
rect 1347 -5834 1351 -5826
rect 1356 -5834 1360 -5826
rect 1365 -5834 1369 -5826
rect 1373 -5834 1377 -5826
rect 1391 -5834 1395 -5826
rect 1413 -5834 1417 -5826
rect 1425 -5834 1429 -5826
rect 1434 -5834 1438 -5826
rect 1443 -5834 1447 -5826
rect 1451 -5834 1455 -5826
rect 1469 -5834 1473 -5826
rect 1491 -5834 1495 -5826
rect 1503 -5834 1507 -5826
rect 1515 -5834 1519 -5826
rect 1527 -5834 1531 -5826
rect 1535 -5834 1539 -5826
rect 1552 -5834 1556 -5826
rect 1561 -5834 1565 -5826
rect -1264 -5957 -1260 -5949
rect -1255 -5957 -1251 -5949
rect -1246 -5957 -1242 -5949
rect -1238 -5957 -1234 -5949
rect -1230 -5957 -1226 -5949
rect -1218 -5957 -1214 -5949
rect -1206 -5957 -1202 -5949
rect -1197 -5957 -1193 -5949
rect -1188 -5957 -1184 -5949
rect -1176 -5957 -1172 -5949
rect -1164 -5957 -1160 -5949
rect -1155 -5957 -1151 -5949
rect -1146 -5957 -1142 -5949
rect -1134 -5957 -1130 -5949
rect -1122 -5957 -1118 -5949
rect -1113 -5957 -1109 -5949
rect -1104 -5957 -1100 -5949
rect -1092 -5957 -1088 -5949
rect -1080 -5957 -1076 -5949
rect -1072 -5957 -1068 -5949
rect -935 -5957 -931 -5949
rect -926 -5957 -922 -5949
rect -917 -5957 -913 -5949
rect -909 -5957 -905 -5949
rect -901 -5957 -897 -5949
rect -889 -5957 -885 -5949
rect -877 -5957 -873 -5949
rect -868 -5957 -864 -5949
rect -859 -5957 -855 -5949
rect -847 -5957 -843 -5949
rect -835 -5957 -831 -5949
rect -826 -5957 -822 -5949
rect -817 -5957 -813 -5949
rect -805 -5957 -801 -5949
rect -793 -5957 -789 -5949
rect -784 -5957 -780 -5949
rect -775 -5957 -771 -5949
rect -763 -5957 -759 -5949
rect -751 -5957 -747 -5949
rect -743 -5957 -739 -5949
rect -577 -5957 -573 -5949
rect -568 -5957 -564 -5949
rect -559 -5957 -555 -5949
rect -551 -5957 -547 -5949
rect -543 -5957 -539 -5949
rect -531 -5957 -527 -5949
rect -519 -5957 -515 -5949
rect -510 -5957 -506 -5949
rect -501 -5957 -497 -5949
rect -489 -5957 -485 -5949
rect -477 -5957 -473 -5949
rect -468 -5957 -464 -5949
rect -459 -5957 -455 -5949
rect -447 -5957 -443 -5949
rect -435 -5957 -431 -5949
rect -426 -5957 -422 -5949
rect -417 -5957 -413 -5949
rect -405 -5957 -401 -5949
rect -393 -5957 -389 -5949
rect -385 -5957 -381 -5949
rect -219 -5957 -215 -5949
rect -210 -5957 -206 -5949
rect -201 -5957 -197 -5949
rect -193 -5957 -189 -5949
rect -185 -5957 -181 -5949
rect -173 -5957 -169 -5949
rect -161 -5957 -157 -5949
rect -152 -5957 -148 -5949
rect -143 -5957 -139 -5949
rect -131 -5957 -127 -5949
rect -119 -5957 -115 -5949
rect -110 -5957 -106 -5949
rect -101 -5957 -97 -5949
rect -89 -5957 -85 -5949
rect -77 -5957 -73 -5949
rect -68 -5957 -64 -5949
rect -59 -5957 -55 -5949
rect -47 -5957 -43 -5949
rect -35 -5957 -31 -5949
rect -27 -5957 -23 -5949
rect 209 -5957 213 -5949
rect 218 -5957 222 -5949
rect 227 -5957 231 -5949
rect 235 -5957 239 -5949
rect 243 -5957 247 -5949
rect 255 -5957 259 -5949
rect 267 -5957 271 -5949
rect 276 -5957 280 -5949
rect 285 -5957 289 -5949
rect 297 -5957 301 -5949
rect 309 -5957 313 -5949
rect 318 -5957 322 -5949
rect 327 -5957 331 -5949
rect 339 -5957 343 -5949
rect 351 -5957 355 -5949
rect 360 -5957 364 -5949
rect 369 -5957 373 -5949
rect 381 -5957 385 -5949
rect 393 -5957 397 -5949
rect 401 -5957 405 -5949
rect 565 -5957 569 -5949
rect 574 -5957 578 -5949
rect 583 -5957 587 -5949
rect 591 -5957 595 -5949
rect 599 -5957 603 -5949
rect 611 -5957 615 -5949
rect 623 -5957 627 -5949
rect 632 -5957 636 -5949
rect 641 -5957 645 -5949
rect 653 -5957 657 -5949
rect 665 -5957 669 -5949
rect 674 -5957 678 -5949
rect 683 -5957 687 -5949
rect 695 -5957 699 -5949
rect 707 -5957 711 -5949
rect 716 -5957 720 -5949
rect 725 -5957 729 -5949
rect 737 -5957 741 -5949
rect 749 -5957 753 -5949
rect 757 -5957 761 -5949
rect 963 -5957 967 -5949
rect 972 -5957 976 -5949
rect 981 -5957 985 -5949
rect 989 -5957 993 -5949
rect 997 -5957 1001 -5949
rect 1009 -5957 1013 -5949
rect 1021 -5957 1025 -5949
rect 1030 -5957 1034 -5949
rect 1039 -5957 1043 -5949
rect 1051 -5957 1055 -5949
rect 1063 -5957 1067 -5949
rect 1072 -5957 1076 -5949
rect 1081 -5957 1085 -5949
rect 1093 -5957 1097 -5949
rect 1105 -5957 1109 -5949
rect 1114 -5957 1118 -5949
rect 1123 -5957 1127 -5949
rect 1135 -5957 1139 -5949
rect 1147 -5957 1151 -5949
rect 1155 -5957 1159 -5949
rect 1321 -5957 1325 -5949
rect 1330 -5957 1334 -5949
rect 1339 -5957 1343 -5949
rect 1347 -5957 1351 -5949
rect 1355 -5957 1359 -5949
rect 1367 -5957 1371 -5949
rect 1379 -5957 1383 -5949
rect 1388 -5957 1392 -5949
rect 1397 -5957 1401 -5949
rect 1409 -5957 1413 -5949
rect 1421 -5957 1425 -5949
rect 1430 -5957 1434 -5949
rect 1439 -5957 1443 -5949
rect 1451 -5957 1455 -5949
rect 1463 -5957 1467 -5949
rect 1472 -5957 1476 -5949
rect 1481 -5957 1485 -5949
rect 1493 -5957 1497 -5949
rect 1505 -5957 1509 -5949
rect 1513 -5957 1517 -5949
rect 1321 -6075 1325 -6067
rect 1330 -6075 1334 -6067
rect 1339 -6075 1343 -6067
rect 1347 -6075 1351 -6067
rect 1355 -6075 1359 -6067
rect 1367 -6075 1371 -6067
rect 1379 -6075 1383 -6067
rect 1388 -6075 1392 -6067
rect 1397 -6075 1401 -6067
rect 1409 -6075 1413 -6067
rect 1421 -6075 1425 -6067
rect 1430 -6075 1434 -6067
rect 1439 -6075 1443 -6067
rect 1451 -6075 1455 -6067
rect 1463 -6075 1467 -6067
rect 1472 -6075 1476 -6067
rect 1481 -6075 1485 -6067
rect 1493 -6075 1497 -6067
rect 1505 -6075 1509 -6067
rect 1513 -6075 1517 -6067
<< m2contact >>
rect -1337 -1034 -1333 -1030
rect -1320 -1034 -1316 -1030
rect -936 -1034 -932 -1030
rect -919 -1034 -915 -1030
rect -948 -1082 -944 -1078
rect -1320 -1126 -1316 -1122
rect -1311 -1204 -1307 -1200
rect -1266 -1090 -1262 -1086
rect -1339 -1264 -1335 -1260
rect -1322 -1264 -1318 -1260
rect -1322 -1356 -1318 -1352
rect -1251 -1148 -1247 -1144
rect -1234 -1148 -1230 -1144
rect -1214 -1148 -1210 -1144
rect -1193 -1148 -1189 -1144
rect -1172 -1148 -1168 -1144
rect -1151 -1148 -1147 -1144
rect -1130 -1148 -1126 -1144
rect -1109 -1148 -1105 -1144
rect -1088 -1148 -1084 -1144
rect -1068 -1148 -1064 -1144
rect -1260 -1211 -1256 -1207
rect -1202 -1204 -1198 -1200
rect -1160 -1211 -1156 -1207
rect -1142 -1204 -1138 -1200
rect -1100 -1196 -1096 -1192
rect -1100 -1204 -1096 -1200
rect -1118 -1218 -1114 -1214
rect -1218 -1225 -1214 -1221
rect -1176 -1225 -1172 -1221
rect -1076 -1211 -1072 -1207
rect -1251 -1240 -1247 -1236
rect -1234 -1240 -1230 -1236
rect -1193 -1240 -1189 -1236
rect -1151 -1240 -1147 -1236
rect -1109 -1240 -1105 -1236
rect -1068 -1240 -1064 -1236
rect -954 -1317 -950 -1313
rect -1251 -1378 -1247 -1374
rect -1234 -1378 -1230 -1374
rect -1194 -1378 -1190 -1374
rect -1173 -1378 -1169 -1374
rect -1266 -1434 -1262 -1430
rect -1260 -1427 -1256 -1423
rect -1313 -1441 -1309 -1437
rect -1216 -1448 -1212 -1444
rect -1164 -1426 -1160 -1422
rect -1234 -1455 -1230 -1451
rect -1198 -1455 -1194 -1451
rect -948 -1418 -944 -1414
rect -577 -1034 -573 -1030
rect -560 -1034 -556 -1030
rect -910 -1090 -906 -1086
rect -589 -1090 -585 -1086
rect -919 -1126 -915 -1122
rect -926 -1148 -922 -1144
rect -909 -1148 -905 -1144
rect -889 -1148 -885 -1144
rect -868 -1148 -864 -1144
rect -847 -1148 -843 -1144
rect -826 -1148 -822 -1144
rect -805 -1148 -801 -1144
rect -784 -1148 -780 -1144
rect -763 -1148 -759 -1144
rect -743 -1148 -739 -1144
rect -935 -1211 -931 -1207
rect -877 -1204 -873 -1200
rect -835 -1211 -831 -1207
rect -817 -1204 -813 -1200
rect -775 -1196 -771 -1192
rect -775 -1204 -771 -1200
rect -793 -1218 -789 -1214
rect -893 -1225 -889 -1221
rect -851 -1225 -847 -1221
rect -751 -1211 -747 -1207
rect -926 -1240 -922 -1236
rect -909 -1240 -905 -1236
rect -868 -1240 -864 -1236
rect -826 -1240 -822 -1236
rect -784 -1240 -780 -1236
rect -743 -1240 -739 -1236
rect -935 -1264 -931 -1260
rect -918 -1264 -914 -1260
rect -954 -1433 -950 -1429
rect -1158 -1448 -1154 -1444
rect -1251 -1470 -1247 -1466
rect -1207 -1470 -1203 -1466
rect -1173 -1470 -1169 -1466
rect -1272 -1477 -1268 -1473
rect -1266 -1484 -1262 -1480
rect -1158 -1484 -1154 -1480
rect -948 -1484 -944 -1480
rect -1251 -1501 -1247 -1497
rect -1234 -1501 -1230 -1497
rect -1214 -1501 -1210 -1497
rect -1193 -1501 -1189 -1497
rect -1172 -1501 -1168 -1497
rect -1151 -1501 -1147 -1497
rect -1130 -1501 -1126 -1497
rect -1109 -1501 -1105 -1497
rect -1088 -1501 -1084 -1497
rect -1068 -1501 -1064 -1497
rect -1266 -1557 -1262 -1553
rect -1260 -1564 -1256 -1560
rect -1202 -1557 -1198 -1553
rect -1160 -1564 -1156 -1560
rect -1142 -1557 -1138 -1553
rect -1100 -1549 -1096 -1545
rect -1100 -1557 -1096 -1553
rect -1118 -1571 -1114 -1567
rect -1218 -1578 -1214 -1574
rect -1176 -1578 -1172 -1574
rect -1076 -1564 -1072 -1560
rect -1251 -1593 -1247 -1589
rect -1234 -1593 -1230 -1589
rect -1193 -1593 -1189 -1589
rect -1151 -1593 -1147 -1589
rect -1109 -1593 -1105 -1589
rect -1068 -1593 -1064 -1589
rect -1251 -1622 -1247 -1618
rect -1234 -1622 -1230 -1618
rect -1214 -1622 -1210 -1618
rect -1193 -1622 -1189 -1618
rect -1172 -1622 -1168 -1618
rect -1151 -1622 -1147 -1618
rect -1130 -1622 -1126 -1618
rect -1109 -1622 -1105 -1618
rect -1088 -1622 -1084 -1618
rect -1068 -1622 -1064 -1618
rect -1272 -1678 -1268 -1674
rect -1260 -1685 -1256 -1681
rect -1202 -1678 -1198 -1674
rect -1160 -1685 -1156 -1681
rect -1142 -1678 -1138 -1674
rect -1100 -1670 -1096 -1666
rect -1100 -1678 -1096 -1674
rect -1118 -1692 -1114 -1688
rect -1218 -1699 -1214 -1695
rect -1176 -1699 -1172 -1695
rect -1062 -1670 -1058 -1666
rect -1076 -1685 -1072 -1681
rect -1251 -1714 -1247 -1710
rect -1234 -1714 -1230 -1710
rect -1193 -1714 -1189 -1710
rect -1151 -1714 -1147 -1710
rect -1109 -1714 -1105 -1710
rect -1068 -1714 -1064 -1710
rect -948 -1678 -944 -1674
rect -1349 -1799 -1345 -1795
rect -1266 -1721 -1262 -1717
rect -1062 -1721 -1058 -1717
rect -1339 -1970 -1335 -1966
rect -1322 -1970 -1318 -1966
rect -1322 -2062 -1318 -2058
rect -953 -1722 -949 -1718
rect -1251 -1743 -1247 -1739
rect -1234 -1743 -1230 -1739
rect -1214 -1743 -1210 -1739
rect -1193 -1743 -1189 -1739
rect -1172 -1743 -1168 -1739
rect -1151 -1743 -1147 -1739
rect -1130 -1743 -1126 -1739
rect -1109 -1743 -1105 -1739
rect -1088 -1743 -1084 -1739
rect -1068 -1743 -1064 -1739
rect -1029 -1743 -1025 -1739
rect -1260 -1806 -1256 -1802
rect -1202 -1799 -1198 -1795
rect -1160 -1806 -1156 -1802
rect -1142 -1799 -1138 -1795
rect -1100 -1791 -1096 -1787
rect -1100 -1799 -1096 -1795
rect -1118 -1813 -1114 -1809
rect -1218 -1820 -1214 -1816
rect -1176 -1820 -1172 -1816
rect -1056 -1791 -1052 -1787
rect -1076 -1806 -1072 -1802
rect -1251 -1835 -1247 -1831
rect -1234 -1835 -1230 -1831
rect -1193 -1835 -1189 -1831
rect -1151 -1835 -1147 -1831
rect -1109 -1835 -1105 -1831
rect -1068 -1835 -1064 -1831
rect -1251 -1858 -1247 -1854
rect -1234 -1858 -1230 -1854
rect -1214 -1858 -1210 -1854
rect -1193 -1858 -1189 -1854
rect -1172 -1858 -1168 -1854
rect -1151 -1858 -1147 -1854
rect -1130 -1858 -1126 -1854
rect -1109 -1858 -1105 -1854
rect -1088 -1858 -1084 -1854
rect -1068 -1858 -1064 -1854
rect -1260 -1921 -1256 -1917
rect -1202 -1914 -1198 -1910
rect -1160 -1921 -1156 -1917
rect -1142 -1914 -1138 -1910
rect -1100 -1898 -1096 -1894
rect -1100 -1914 -1096 -1910
rect -1118 -1928 -1114 -1924
rect -1218 -1935 -1214 -1931
rect -1176 -1935 -1172 -1931
rect -1062 -1898 -1058 -1894
rect -1076 -1921 -1072 -1917
rect -1251 -1950 -1247 -1946
rect -1234 -1950 -1230 -1946
rect -1193 -1950 -1189 -1946
rect -1151 -1950 -1147 -1946
rect -1109 -1950 -1105 -1946
rect -1068 -1950 -1064 -1946
rect -1021 -1792 -1017 -1788
rect -1029 -1835 -1025 -1831
rect -1029 -1858 -1025 -1854
rect -1021 -1907 -1017 -1903
rect -1029 -1950 -1025 -1946
rect -1056 -2002 -1052 -1998
rect -1062 -2010 -1058 -2006
rect -1251 -2089 -1247 -2085
rect -1234 -2089 -1230 -2085
rect -1194 -2089 -1190 -2085
rect -1173 -2089 -1169 -2085
rect -1266 -2145 -1262 -2141
rect -1260 -2138 -1256 -2134
rect -1313 -2152 -1309 -2148
rect -1216 -2159 -1212 -2155
rect -909 -1317 -905 -1313
rect -595 -1317 -591 -1313
rect -918 -1356 -914 -1352
rect -926 -1378 -922 -1374
rect -900 -1378 -896 -1374
rect -883 -1378 -879 -1374
rect -843 -1378 -839 -1374
rect -822 -1378 -818 -1374
rect -805 -1378 -801 -1374
rect -765 -1378 -761 -1374
rect -741 -1378 -737 -1374
rect -704 -1378 -700 -1374
rect -935 -1411 -931 -1407
rect -917 -1404 -913 -1400
rect -891 -1426 -887 -1422
rect -909 -1433 -905 -1429
rect -865 -1418 -861 -1414
rect -813 -1411 -809 -1407
rect -883 -1455 -879 -1451
rect -847 -1455 -843 -1451
rect -787 -1426 -783 -1422
rect -805 -1455 -801 -1451
rect -769 -1455 -765 -1451
rect -695 -1418 -691 -1414
rect -689 -1426 -685 -1422
rect -926 -1470 -922 -1466
rect -900 -1470 -896 -1466
rect -857 -1470 -853 -1466
rect -822 -1470 -818 -1466
rect -778 -1470 -774 -1466
rect -761 -1470 -757 -1466
rect -725 -1470 -721 -1466
rect -704 -1470 -700 -1466
rect -589 -1418 -585 -1414
rect -219 -1034 -215 -1030
rect -202 -1034 -198 -1030
rect -551 -1082 -547 -1078
rect -231 -1082 -227 -1078
rect -560 -1126 -556 -1122
rect -568 -1148 -564 -1144
rect -551 -1148 -547 -1144
rect -531 -1148 -527 -1144
rect -510 -1148 -506 -1144
rect -489 -1148 -485 -1144
rect -468 -1148 -464 -1144
rect -447 -1148 -443 -1144
rect -426 -1148 -422 -1144
rect -405 -1148 -401 -1144
rect -385 -1148 -381 -1144
rect -577 -1211 -573 -1207
rect -519 -1204 -515 -1200
rect -477 -1211 -473 -1207
rect -459 -1204 -455 -1200
rect -417 -1196 -413 -1192
rect -417 -1204 -413 -1200
rect -435 -1218 -431 -1214
rect -535 -1225 -531 -1221
rect -493 -1225 -489 -1221
rect -393 -1211 -389 -1207
rect -568 -1240 -564 -1236
rect -551 -1240 -547 -1236
rect -510 -1240 -506 -1236
rect -468 -1240 -464 -1236
rect -426 -1240 -422 -1236
rect -385 -1240 -381 -1236
rect -577 -1264 -573 -1260
rect -560 -1264 -556 -1260
rect -595 -1433 -591 -1429
rect -689 -1477 -685 -1473
rect -589 -1491 -585 -1487
rect -926 -1501 -922 -1497
rect -909 -1501 -905 -1497
rect -889 -1501 -885 -1497
rect -868 -1501 -864 -1497
rect -847 -1501 -843 -1497
rect -826 -1501 -822 -1497
rect -805 -1501 -801 -1497
rect -784 -1501 -780 -1497
rect -763 -1501 -759 -1497
rect -743 -1501 -739 -1497
rect -935 -1564 -931 -1560
rect -877 -1557 -873 -1553
rect -835 -1564 -831 -1560
rect -817 -1557 -813 -1553
rect -775 -1549 -771 -1545
rect -775 -1557 -771 -1553
rect -793 -1571 -789 -1567
rect -893 -1578 -889 -1574
rect -851 -1578 -847 -1574
rect -751 -1564 -747 -1560
rect -926 -1593 -922 -1589
rect -909 -1593 -905 -1589
rect -868 -1593 -864 -1589
rect -826 -1593 -822 -1589
rect -784 -1593 -780 -1589
rect -743 -1593 -739 -1589
rect -926 -1622 -922 -1618
rect -909 -1622 -905 -1618
rect -889 -1622 -885 -1618
rect -868 -1622 -864 -1618
rect -847 -1622 -843 -1618
rect -826 -1622 -822 -1618
rect -805 -1622 -801 -1618
rect -784 -1622 -780 -1618
rect -763 -1622 -759 -1618
rect -743 -1622 -739 -1618
rect -935 -1685 -931 -1681
rect -877 -1678 -873 -1674
rect -835 -1685 -831 -1681
rect -817 -1678 -813 -1674
rect -775 -1670 -771 -1666
rect -775 -1678 -771 -1674
rect -793 -1692 -789 -1688
rect -893 -1699 -889 -1695
rect -851 -1699 -847 -1695
rect -737 -1670 -733 -1666
rect -751 -1685 -747 -1681
rect -926 -1714 -922 -1710
rect -909 -1714 -905 -1710
rect -868 -1714 -864 -1710
rect -826 -1714 -822 -1710
rect -784 -1714 -780 -1710
rect -743 -1714 -739 -1710
rect -589 -1678 -585 -1674
rect -737 -1722 -733 -1718
rect -589 -1722 -585 -1718
rect -926 -1743 -922 -1739
rect -909 -1743 -905 -1739
rect -889 -1743 -885 -1739
rect -868 -1743 -864 -1739
rect -847 -1743 -843 -1739
rect -826 -1743 -822 -1739
rect -805 -1743 -801 -1739
rect -784 -1743 -780 -1739
rect -763 -1743 -759 -1739
rect -743 -1743 -739 -1739
rect -942 -1799 -938 -1795
rect -935 -1806 -931 -1802
rect -877 -1799 -873 -1795
rect -835 -1806 -831 -1802
rect -817 -1799 -813 -1795
rect -775 -1791 -771 -1787
rect -775 -1799 -771 -1795
rect -793 -1813 -789 -1809
rect -893 -1820 -889 -1816
rect -851 -1820 -847 -1816
rect -737 -1791 -733 -1787
rect -751 -1806 -747 -1802
rect -926 -1835 -922 -1831
rect -909 -1835 -905 -1831
rect -868 -1835 -864 -1831
rect -826 -1835 -822 -1831
rect -784 -1835 -780 -1831
rect -743 -1835 -739 -1831
rect -935 -1970 -931 -1966
rect -918 -1970 -914 -1966
rect -953 -2129 -949 -2125
rect -947 -2023 -943 -2019
rect -1164 -2137 -1160 -2133
rect -1234 -2166 -1230 -2162
rect -1198 -2166 -1194 -2162
rect -947 -2144 -943 -2140
rect -1158 -2159 -1154 -2155
rect -1251 -2181 -1247 -2177
rect -1207 -2181 -1203 -2177
rect -1173 -2181 -1169 -2177
rect -1276 -2188 -1272 -2184
rect -1270 -2195 -1266 -2191
rect -1158 -2195 -1154 -2191
rect -947 -2195 -943 -2191
rect -1255 -2233 -1251 -2229
rect -1238 -2233 -1234 -2229
rect -1218 -2233 -1214 -2229
rect -1197 -2233 -1193 -2229
rect -1176 -2233 -1172 -2229
rect -1155 -2233 -1151 -2229
rect -1134 -2233 -1130 -2229
rect -1113 -2233 -1109 -2229
rect -1092 -2233 -1088 -2229
rect -1072 -2233 -1068 -2229
rect -1270 -2289 -1266 -2285
rect -1264 -2296 -1260 -2292
rect -1206 -2289 -1202 -2285
rect -1164 -2296 -1160 -2292
rect -1146 -2289 -1142 -2285
rect -1104 -2281 -1100 -2277
rect -1104 -2289 -1100 -2285
rect -1122 -2303 -1118 -2299
rect -1222 -2310 -1218 -2306
rect -1180 -2310 -1176 -2306
rect -1080 -2296 -1076 -2292
rect -1255 -2325 -1251 -2321
rect -1238 -2325 -1234 -2321
rect -1197 -2325 -1193 -2321
rect -1155 -2325 -1151 -2321
rect -1113 -2325 -1109 -2321
rect -1072 -2325 -1068 -2321
rect -1255 -2364 -1251 -2360
rect -1238 -2364 -1234 -2360
rect -1218 -2364 -1214 -2360
rect -1197 -2364 -1193 -2360
rect -1176 -2364 -1172 -2360
rect -1155 -2364 -1151 -2360
rect -1134 -2364 -1130 -2360
rect -1113 -2364 -1109 -2360
rect -1092 -2364 -1088 -2360
rect -1072 -2364 -1068 -2360
rect -1276 -2420 -1272 -2416
rect -1264 -2427 -1260 -2423
rect -1206 -2420 -1202 -2416
rect -1164 -2427 -1160 -2423
rect -1146 -2420 -1142 -2416
rect -1104 -2412 -1100 -2408
rect -1104 -2420 -1100 -2416
rect -1122 -2434 -1118 -2430
rect -1222 -2441 -1218 -2437
rect -1180 -2441 -1176 -2437
rect -1066 -2412 -1062 -2408
rect -1080 -2427 -1076 -2423
rect -1255 -2456 -1251 -2452
rect -1238 -2456 -1234 -2452
rect -1197 -2456 -1193 -2452
rect -1155 -2456 -1151 -2452
rect -1113 -2456 -1109 -2452
rect -1072 -2456 -1068 -2452
rect -947 -2420 -943 -2416
rect -1349 -2551 -1345 -2547
rect -1270 -2464 -1266 -2460
rect -1066 -2464 -1062 -2460
rect -947 -2463 -943 -2459
rect -1339 -2720 -1335 -2716
rect -1322 -2720 -1318 -2716
rect -1322 -2812 -1318 -2808
rect -1255 -2495 -1251 -2491
rect -1238 -2495 -1234 -2491
rect -1218 -2495 -1214 -2491
rect -1197 -2495 -1193 -2491
rect -1176 -2495 -1172 -2491
rect -1155 -2495 -1151 -2491
rect -1134 -2495 -1130 -2491
rect -1113 -2495 -1109 -2491
rect -1092 -2495 -1088 -2491
rect -1072 -2495 -1068 -2491
rect -1264 -2558 -1260 -2554
rect -1206 -2551 -1202 -2547
rect -1164 -2558 -1160 -2554
rect -1146 -2551 -1142 -2547
rect -1104 -2543 -1100 -2539
rect -1104 -2551 -1100 -2547
rect -1122 -2565 -1118 -2561
rect -1222 -2572 -1218 -2568
rect -1180 -2572 -1176 -2568
rect -1066 -2543 -1062 -2539
rect -1080 -2558 -1076 -2554
rect -1255 -2587 -1251 -2583
rect -1238 -2587 -1234 -2583
rect -1197 -2587 -1193 -2583
rect -1155 -2587 -1151 -2583
rect -1113 -2587 -1109 -2583
rect -1072 -2587 -1068 -2583
rect -1255 -2607 -1251 -2603
rect -1238 -2607 -1234 -2603
rect -1218 -2607 -1214 -2603
rect -1197 -2607 -1193 -2603
rect -1176 -2607 -1172 -2603
rect -1155 -2607 -1151 -2603
rect -1134 -2607 -1130 -2603
rect -1113 -2607 -1109 -2603
rect -1092 -2607 -1088 -2603
rect -1072 -2607 -1068 -2603
rect -1264 -2670 -1260 -2666
rect -1206 -2663 -1202 -2659
rect -1164 -2670 -1160 -2666
rect -1146 -2663 -1142 -2659
rect -1104 -2655 -1100 -2651
rect -1104 -2663 -1100 -2659
rect -1122 -2677 -1118 -2673
rect -1222 -2684 -1218 -2680
rect -1180 -2684 -1176 -2680
rect -1080 -2670 -1076 -2666
rect -1255 -2699 -1251 -2695
rect -1238 -2699 -1234 -2695
rect -1197 -2699 -1193 -2695
rect -1155 -2699 -1151 -2695
rect -1113 -2699 -1109 -2695
rect -1072 -2699 -1068 -2695
rect -1066 -2752 -1062 -2748
rect -953 -2773 -949 -2769
rect -1255 -2839 -1251 -2835
rect -1238 -2839 -1234 -2835
rect -1198 -2839 -1194 -2835
rect -1177 -2839 -1173 -2835
rect -1270 -2895 -1266 -2891
rect -1264 -2888 -1260 -2884
rect -1313 -2902 -1309 -2898
rect -1220 -2909 -1216 -2905
rect -953 -2879 -949 -2875
rect -1168 -2887 -1164 -2883
rect -1238 -2916 -1234 -2912
rect -1202 -2916 -1198 -2912
rect -673 -1858 -669 -1854
rect -665 -1907 -661 -1903
rect -673 -1950 -669 -1946
rect -737 -2002 -733 -1998
rect -909 -2023 -905 -2019
rect -595 -2023 -591 -2019
rect -918 -2062 -914 -2058
rect -926 -2089 -922 -2085
rect -900 -2089 -896 -2085
rect -883 -2089 -879 -2085
rect -843 -2089 -839 -2085
rect -822 -2089 -818 -2085
rect -805 -2089 -801 -2085
rect -765 -2089 -761 -2085
rect -741 -2089 -737 -2085
rect -704 -2089 -700 -2085
rect -935 -2122 -931 -2118
rect -917 -2115 -913 -2111
rect -891 -2137 -887 -2133
rect -909 -2144 -905 -2140
rect -865 -2129 -861 -2125
rect -813 -2122 -809 -2118
rect -883 -2166 -879 -2162
rect -847 -2166 -843 -2162
rect -787 -2137 -783 -2133
rect -805 -2166 -801 -2162
rect -769 -2166 -765 -2162
rect -695 -2129 -691 -2125
rect -689 -2137 -685 -2133
rect -926 -2181 -922 -2177
rect -900 -2181 -896 -2177
rect -857 -2181 -853 -2177
rect -822 -2181 -818 -2177
rect -778 -2181 -774 -2177
rect -761 -2181 -757 -2177
rect -725 -2181 -721 -2177
rect -704 -2181 -700 -2177
rect -551 -1317 -547 -1313
rect -237 -1317 -233 -1313
rect -560 -1356 -556 -1352
rect -568 -1378 -564 -1374
rect -542 -1378 -538 -1374
rect -525 -1378 -521 -1374
rect -485 -1378 -481 -1374
rect -464 -1378 -460 -1374
rect -447 -1378 -443 -1374
rect -407 -1378 -403 -1374
rect -383 -1378 -379 -1374
rect -346 -1378 -342 -1374
rect -577 -1411 -573 -1407
rect -559 -1404 -555 -1400
rect -533 -1426 -529 -1422
rect -551 -1433 -547 -1429
rect -507 -1418 -503 -1414
rect -455 -1411 -451 -1407
rect -525 -1455 -521 -1451
rect -489 -1455 -485 -1451
rect -429 -1426 -425 -1422
rect -447 -1455 -443 -1451
rect -411 -1455 -407 -1451
rect -337 -1418 -333 -1414
rect -331 -1426 -327 -1422
rect -568 -1470 -564 -1466
rect -542 -1470 -538 -1466
rect -499 -1470 -495 -1466
rect -464 -1470 -460 -1466
rect -420 -1470 -416 -1466
rect -403 -1470 -399 -1466
rect -367 -1470 -363 -1466
rect -346 -1470 -342 -1466
rect -231 -1418 -227 -1414
rect 209 -1034 213 -1030
rect 226 -1034 230 -1030
rect -193 -1090 -189 -1086
rect 197 -1090 201 -1086
rect -202 -1126 -198 -1122
rect -210 -1148 -206 -1144
rect -193 -1148 -189 -1144
rect -173 -1148 -169 -1144
rect -152 -1148 -148 -1144
rect -131 -1148 -127 -1144
rect -110 -1148 -106 -1144
rect -89 -1148 -85 -1144
rect -68 -1148 -64 -1144
rect -47 -1148 -43 -1144
rect -27 -1148 -23 -1144
rect -219 -1211 -215 -1207
rect -161 -1204 -157 -1200
rect -119 -1211 -115 -1207
rect -101 -1204 -97 -1200
rect -59 -1196 -55 -1192
rect -59 -1204 -55 -1200
rect -77 -1218 -73 -1214
rect -177 -1225 -173 -1221
rect -135 -1225 -131 -1221
rect -35 -1211 -31 -1207
rect -210 -1240 -206 -1236
rect -193 -1240 -189 -1236
rect -152 -1240 -148 -1236
rect -110 -1240 -106 -1236
rect -68 -1240 -64 -1236
rect -27 -1240 -23 -1236
rect -219 -1264 -215 -1260
rect -202 -1264 -198 -1260
rect -237 -1433 -233 -1429
rect -331 -1484 -327 -1480
rect -231 -1484 -227 -1480
rect -568 -1501 -564 -1497
rect -551 -1501 -547 -1497
rect -531 -1501 -527 -1497
rect -510 -1501 -506 -1497
rect -489 -1501 -485 -1497
rect -468 -1501 -464 -1497
rect -447 -1501 -443 -1497
rect -426 -1501 -422 -1497
rect -405 -1501 -401 -1497
rect -385 -1501 -381 -1497
rect -577 -1564 -573 -1560
rect -519 -1557 -515 -1553
rect -477 -1564 -473 -1560
rect -459 -1557 -455 -1553
rect -417 -1549 -413 -1545
rect -417 -1557 -413 -1553
rect -435 -1571 -431 -1567
rect -535 -1578 -531 -1574
rect -493 -1578 -489 -1574
rect -393 -1564 -389 -1560
rect -568 -1593 -564 -1589
rect -551 -1593 -547 -1589
rect -510 -1593 -506 -1589
rect -468 -1593 -464 -1589
rect -426 -1593 -422 -1589
rect -385 -1593 -381 -1589
rect -568 -1622 -564 -1618
rect -551 -1622 -547 -1618
rect -531 -1622 -527 -1618
rect -510 -1622 -506 -1618
rect -489 -1622 -485 -1618
rect -468 -1622 -464 -1618
rect -447 -1622 -443 -1618
rect -426 -1622 -422 -1618
rect -405 -1622 -401 -1618
rect -385 -1622 -381 -1618
rect -577 -1685 -573 -1681
rect -519 -1678 -515 -1674
rect -477 -1685 -473 -1681
rect -459 -1678 -455 -1674
rect -417 -1670 -413 -1666
rect -417 -1678 -413 -1674
rect -435 -1692 -431 -1688
rect -535 -1699 -531 -1695
rect -493 -1699 -489 -1695
rect -379 -1670 -375 -1666
rect -393 -1685 -389 -1681
rect -568 -1714 -564 -1710
rect -551 -1714 -547 -1710
rect -510 -1714 -506 -1710
rect -468 -1714 -464 -1710
rect -426 -1714 -422 -1710
rect -385 -1714 -381 -1710
rect -231 -1678 -227 -1674
rect -379 -1722 -375 -1718
rect -231 -1721 -227 -1717
rect -568 -1743 -564 -1739
rect -551 -1743 -547 -1739
rect -531 -1743 -527 -1739
rect -510 -1743 -506 -1739
rect -489 -1743 -485 -1739
rect -468 -1743 -464 -1739
rect -447 -1743 -443 -1739
rect -426 -1743 -422 -1739
rect -405 -1743 -401 -1739
rect -385 -1743 -381 -1739
rect -583 -1799 -579 -1795
rect -332 -1743 -328 -1739
rect -577 -1806 -573 -1802
rect -519 -1799 -515 -1795
rect -477 -1806 -473 -1802
rect -459 -1799 -455 -1795
rect -417 -1791 -413 -1787
rect -417 -1799 -413 -1795
rect -435 -1813 -431 -1809
rect -535 -1820 -531 -1816
rect -493 -1820 -489 -1816
rect -379 -1791 -375 -1787
rect -393 -1806 -389 -1802
rect -568 -1835 -564 -1831
rect -551 -1835 -547 -1831
rect -510 -1835 -506 -1831
rect -468 -1835 -464 -1831
rect -426 -1835 -422 -1831
rect -385 -1835 -381 -1831
rect -577 -1970 -573 -1966
rect -560 -1970 -556 -1966
rect -589 -2129 -585 -2125
rect -595 -2144 -591 -2140
rect -689 -2188 -685 -2184
rect -589 -2188 -585 -2184
rect -926 -2233 -922 -2229
rect -909 -2233 -905 -2229
rect -889 -2233 -885 -2229
rect -868 -2233 -864 -2229
rect -847 -2233 -843 -2229
rect -826 -2233 -822 -2229
rect -805 -2233 -801 -2229
rect -784 -2233 -780 -2229
rect -763 -2233 -759 -2229
rect -743 -2233 -739 -2229
rect -935 -2296 -931 -2292
rect -877 -2289 -873 -2285
rect -835 -2296 -831 -2292
rect -817 -2289 -813 -2285
rect -775 -2281 -771 -2277
rect -775 -2289 -771 -2285
rect -793 -2303 -789 -2299
rect -893 -2310 -889 -2306
rect -851 -2310 -847 -2306
rect -751 -2296 -747 -2292
rect -926 -2325 -922 -2321
rect -909 -2325 -905 -2321
rect -868 -2325 -864 -2321
rect -826 -2325 -822 -2321
rect -784 -2325 -780 -2321
rect -743 -2325 -739 -2321
rect -926 -2364 -922 -2360
rect -909 -2364 -905 -2360
rect -889 -2364 -885 -2360
rect -868 -2364 -864 -2360
rect -847 -2364 -843 -2360
rect -826 -2364 -822 -2360
rect -805 -2364 -801 -2360
rect -784 -2364 -780 -2360
rect -763 -2364 -759 -2360
rect -743 -2364 -739 -2360
rect -935 -2427 -931 -2423
rect -877 -2420 -873 -2416
rect -835 -2427 -831 -2423
rect -817 -2420 -813 -2416
rect -775 -2412 -771 -2408
rect -775 -2420 -771 -2416
rect -793 -2434 -789 -2430
rect -893 -2441 -889 -2437
rect -851 -2441 -847 -2437
rect -737 -2412 -733 -2408
rect -751 -2427 -747 -2423
rect -926 -2456 -922 -2452
rect -909 -2456 -905 -2452
rect -868 -2456 -864 -2452
rect -826 -2456 -822 -2452
rect -784 -2456 -780 -2452
rect -743 -2456 -739 -2452
rect -589 -2420 -585 -2416
rect -737 -2463 -733 -2459
rect -589 -2464 -585 -2460
rect -926 -2495 -922 -2491
rect -909 -2495 -905 -2491
rect -889 -2495 -885 -2491
rect -868 -2495 -864 -2491
rect -847 -2495 -843 -2491
rect -826 -2495 -822 -2491
rect -805 -2495 -801 -2491
rect -784 -2495 -780 -2491
rect -763 -2495 -759 -2491
rect -743 -2495 -739 -2491
rect -941 -2551 -937 -2547
rect -935 -2558 -931 -2554
rect -877 -2551 -873 -2547
rect -835 -2558 -831 -2554
rect -817 -2551 -813 -2547
rect -775 -2543 -771 -2539
rect -775 -2551 -771 -2547
rect -793 -2565 -789 -2561
rect -893 -2572 -889 -2568
rect -851 -2572 -847 -2568
rect -731 -2543 -727 -2539
rect -751 -2558 -747 -2554
rect -926 -2587 -922 -2583
rect -909 -2587 -905 -2583
rect -868 -2587 -864 -2583
rect -826 -2587 -822 -2583
rect -784 -2587 -780 -2583
rect -743 -2587 -739 -2583
rect -926 -2607 -922 -2603
rect -909 -2607 -905 -2603
rect -889 -2607 -885 -2603
rect -868 -2607 -864 -2603
rect -847 -2607 -843 -2603
rect -826 -2607 -822 -2603
rect -805 -2607 -801 -2603
rect -784 -2607 -780 -2603
rect -763 -2607 -759 -2603
rect -743 -2607 -739 -2603
rect -935 -2670 -931 -2666
rect -877 -2663 -873 -2659
rect -835 -2670 -831 -2666
rect -817 -2663 -813 -2659
rect -775 -2655 -771 -2651
rect -775 -2663 -771 -2659
rect -793 -2677 -789 -2673
rect -893 -2684 -889 -2680
rect -851 -2684 -847 -2680
rect -737 -2655 -733 -2651
rect -751 -2670 -747 -2666
rect -926 -2699 -922 -2695
rect -909 -2699 -905 -2695
rect -868 -2699 -864 -2695
rect -826 -2699 -822 -2695
rect -784 -2699 -780 -2695
rect -743 -2699 -739 -2695
rect -935 -2720 -931 -2716
rect -918 -2720 -914 -2716
rect -947 -2894 -943 -2890
rect -1162 -2909 -1158 -2905
rect -1255 -2931 -1251 -2927
rect -1211 -2931 -1207 -2927
rect -1177 -2931 -1173 -2927
rect -1276 -2938 -1272 -2934
rect -1270 -2946 -1266 -2942
rect -1162 -2946 -1158 -2942
rect -947 -2945 -943 -2941
rect -1255 -2958 -1251 -2954
rect -1238 -2958 -1234 -2954
rect -1218 -2958 -1214 -2954
rect -1197 -2958 -1193 -2954
rect -1176 -2958 -1172 -2954
rect -1155 -2958 -1151 -2954
rect -1134 -2958 -1130 -2954
rect -1113 -2958 -1109 -2954
rect -1092 -2958 -1088 -2954
rect -1072 -2958 -1068 -2954
rect -1270 -3014 -1266 -3010
rect -1026 -2958 -1022 -2954
rect -1264 -3021 -1260 -3017
rect -1206 -3014 -1202 -3010
rect -1164 -3021 -1160 -3017
rect -1146 -3014 -1142 -3010
rect -1104 -2979 -1100 -2975
rect -1104 -3014 -1100 -3010
rect -1122 -3028 -1118 -3024
rect -1222 -3035 -1218 -3031
rect -1180 -3035 -1176 -3031
rect -1018 -3008 -1014 -3004
rect -1080 -3021 -1076 -3017
rect -1255 -3050 -1251 -3046
rect -1238 -3050 -1234 -3046
rect -1197 -3050 -1193 -3046
rect -1155 -3050 -1151 -3046
rect -1113 -3050 -1109 -3046
rect -1072 -3050 -1068 -3046
rect -1026 -3050 -1022 -3046
rect -1255 -3074 -1251 -3070
rect -1238 -3074 -1234 -3070
rect -1218 -3074 -1214 -3070
rect -1197 -3074 -1193 -3070
rect -1176 -3074 -1172 -3070
rect -1155 -3074 -1151 -3070
rect -1134 -3074 -1130 -3070
rect -1113 -3074 -1109 -3070
rect -1092 -3074 -1088 -3070
rect -1072 -3074 -1068 -3070
rect -1276 -3130 -1272 -3126
rect -1026 -3074 -1022 -3070
rect -1264 -3137 -1260 -3133
rect -1206 -3130 -1202 -3126
rect -1164 -3137 -1160 -3133
rect -1146 -3130 -1142 -3126
rect -1104 -3122 -1100 -3118
rect -1104 -3130 -1100 -3126
rect -1122 -3144 -1118 -3140
rect -1222 -3151 -1218 -3147
rect -1180 -3151 -1176 -3147
rect -1066 -3122 -1062 -3118
rect -1080 -3137 -1076 -3133
rect -1255 -3166 -1251 -3162
rect -1238 -3166 -1234 -3162
rect -1197 -3166 -1193 -3162
rect -1155 -3166 -1151 -3162
rect -1113 -3166 -1109 -3162
rect -1072 -3166 -1068 -3162
rect -1018 -3123 -1014 -3119
rect -947 -3130 -943 -3126
rect -1026 -3166 -1022 -3162
rect -1349 -3251 -1345 -3247
rect -1270 -3174 -1266 -3170
rect -1066 -3174 -1062 -3170
rect -947 -3174 -943 -3170
rect -1339 -3426 -1335 -3422
rect -1322 -3426 -1318 -3422
rect -1621 -3851 -1607 -3837
rect -1322 -3518 -1318 -3514
rect -1255 -3195 -1251 -3191
rect -1238 -3195 -1234 -3191
rect -1218 -3195 -1214 -3191
rect -1197 -3195 -1193 -3191
rect -1176 -3195 -1172 -3191
rect -1155 -3195 -1151 -3191
rect -1134 -3195 -1130 -3191
rect -1113 -3195 -1109 -3191
rect -1092 -3195 -1088 -3191
rect -1072 -3195 -1068 -3191
rect -1264 -3258 -1260 -3254
rect -1206 -3251 -1202 -3247
rect -1164 -3258 -1160 -3254
rect -1146 -3251 -1142 -3247
rect -1104 -3243 -1100 -3239
rect -1104 -3251 -1100 -3247
rect -1122 -3265 -1118 -3261
rect -1222 -3272 -1218 -3268
rect -1180 -3272 -1176 -3268
rect -1066 -3243 -1062 -3239
rect -1080 -3258 -1076 -3254
rect -1255 -3287 -1251 -3283
rect -1238 -3287 -1234 -3283
rect -1197 -3287 -1193 -3283
rect -1155 -3287 -1151 -3283
rect -1113 -3287 -1109 -3283
rect -1072 -3287 -1068 -3283
rect -1255 -3309 -1251 -3305
rect -1238 -3309 -1234 -3305
rect -1218 -3309 -1214 -3305
rect -1197 -3309 -1193 -3305
rect -1176 -3309 -1172 -3305
rect -1155 -3309 -1151 -3305
rect -1134 -3309 -1130 -3305
rect -1113 -3309 -1109 -3305
rect -1092 -3309 -1088 -3305
rect -1072 -3309 -1068 -3305
rect -1264 -3372 -1260 -3368
rect -1206 -3365 -1202 -3361
rect -1164 -3372 -1160 -3368
rect -1146 -3365 -1142 -3361
rect -1104 -3357 -1100 -3353
rect -1104 -3365 -1100 -3361
rect -1122 -3379 -1118 -3375
rect -1222 -3386 -1218 -3382
rect -1180 -3386 -1176 -3382
rect -1080 -3372 -1076 -3368
rect -1255 -3401 -1251 -3397
rect -1238 -3401 -1234 -3397
rect -1197 -3401 -1193 -3397
rect -1155 -3401 -1151 -3397
rect -1113 -3401 -1109 -3397
rect -1072 -3401 -1068 -3397
rect -1066 -3458 -1062 -3454
rect -953 -3479 -949 -3475
rect -1255 -3550 -1251 -3546
rect -1238 -3550 -1234 -3546
rect -1198 -3550 -1194 -3546
rect -1177 -3550 -1173 -3546
rect -1270 -3606 -1266 -3602
rect -1264 -3599 -1260 -3595
rect -1313 -3613 -1309 -3609
rect -1220 -3620 -1216 -3616
rect -953 -3590 -949 -3586
rect -1168 -3598 -1164 -3594
rect -1238 -3627 -1234 -3623
rect -1202 -3627 -1198 -3623
rect -731 -2752 -727 -2748
rect -737 -2760 -733 -2756
rect -909 -2773 -905 -2769
rect -595 -2773 -591 -2769
rect -918 -2812 -914 -2808
rect -926 -2839 -922 -2835
rect -900 -2839 -896 -2835
rect -883 -2839 -879 -2835
rect -843 -2839 -839 -2835
rect -822 -2839 -818 -2835
rect -805 -2839 -801 -2835
rect -765 -2839 -761 -2835
rect -741 -2839 -737 -2835
rect -704 -2839 -700 -2835
rect -935 -2872 -931 -2868
rect -917 -2865 -913 -2861
rect -891 -2887 -887 -2883
rect -909 -2894 -905 -2890
rect -865 -2879 -861 -2875
rect -813 -2872 -809 -2868
rect -883 -2916 -879 -2912
rect -847 -2916 -843 -2912
rect -787 -2887 -783 -2883
rect -805 -2916 -801 -2912
rect -769 -2916 -765 -2912
rect -695 -2879 -691 -2875
rect -689 -2887 -685 -2883
rect -926 -2931 -922 -2927
rect -900 -2931 -896 -2927
rect -857 -2931 -853 -2927
rect -822 -2931 -818 -2927
rect -778 -2931 -774 -2927
rect -761 -2931 -757 -2927
rect -725 -2931 -721 -2927
rect -704 -2931 -700 -2927
rect -324 -1792 -320 -1788
rect -332 -1835 -328 -1831
rect -332 -1858 -328 -1854
rect -324 -1907 -320 -1903
rect -332 -1950 -328 -1946
rect -379 -2002 -375 -1998
rect -551 -2023 -547 -2019
rect -237 -2023 -233 -2019
rect -560 -2062 -556 -2058
rect -568 -2089 -564 -2085
rect -542 -2089 -538 -2085
rect -525 -2089 -521 -2085
rect -485 -2089 -481 -2085
rect -464 -2089 -460 -2085
rect -447 -2089 -443 -2085
rect -407 -2089 -403 -2085
rect -383 -2089 -379 -2085
rect -346 -2089 -342 -2085
rect -577 -2122 -573 -2118
rect -559 -2115 -555 -2111
rect -533 -2137 -529 -2133
rect -551 -2144 -547 -2140
rect -507 -2129 -503 -2125
rect -455 -2122 -451 -2118
rect -525 -2166 -521 -2162
rect -489 -2166 -485 -2162
rect -429 -2137 -425 -2133
rect -447 -2166 -443 -2162
rect -411 -2166 -407 -2162
rect -337 -2126 -333 -2122
rect -331 -2137 -327 -2133
rect -568 -2181 -564 -2177
rect -542 -2181 -538 -2177
rect -499 -2181 -495 -2177
rect -464 -2181 -460 -2177
rect -420 -2181 -416 -2177
rect -403 -2181 -399 -2177
rect -367 -2181 -363 -2177
rect -346 -2181 -342 -2177
rect -193 -1317 -189 -1313
rect 191 -1317 195 -1313
rect -202 -1356 -198 -1352
rect -210 -1378 -206 -1374
rect -184 -1378 -180 -1374
rect -167 -1378 -163 -1374
rect -127 -1378 -123 -1374
rect -106 -1378 -102 -1374
rect -89 -1378 -85 -1374
rect -49 -1378 -45 -1374
rect -25 -1378 -21 -1374
rect 12 -1378 16 -1374
rect -219 -1411 -215 -1407
rect -201 -1404 -197 -1400
rect -175 -1426 -171 -1422
rect -193 -1433 -189 -1429
rect -149 -1418 -145 -1414
rect -97 -1411 -93 -1407
rect -167 -1455 -163 -1451
rect -131 -1455 -127 -1451
rect -71 -1426 -67 -1422
rect -89 -1455 -85 -1451
rect -53 -1455 -49 -1451
rect 21 -1418 25 -1414
rect 27 -1426 31 -1422
rect -210 -1470 -206 -1466
rect -184 -1470 -180 -1466
rect -141 -1470 -137 -1466
rect -106 -1470 -102 -1466
rect -62 -1470 -58 -1466
rect -45 -1470 -41 -1466
rect -9 -1470 -5 -1466
rect 12 -1470 16 -1466
rect 197 -1418 201 -1414
rect 565 -1034 569 -1030
rect 582 -1034 586 -1030
rect 235 -1082 239 -1078
rect 553 -1082 557 -1078
rect 226 -1126 230 -1122
rect 218 -1148 222 -1144
rect 235 -1148 239 -1144
rect 255 -1148 259 -1144
rect 276 -1148 280 -1144
rect 297 -1148 301 -1144
rect 318 -1148 322 -1144
rect 339 -1148 343 -1144
rect 360 -1148 364 -1144
rect 381 -1148 385 -1144
rect 401 -1148 405 -1144
rect 209 -1211 213 -1207
rect 267 -1204 271 -1200
rect 309 -1211 313 -1207
rect 327 -1204 331 -1200
rect 369 -1196 373 -1192
rect 369 -1204 373 -1200
rect 351 -1218 355 -1214
rect 251 -1225 255 -1221
rect 293 -1225 297 -1221
rect 393 -1211 397 -1207
rect 218 -1240 222 -1236
rect 235 -1240 239 -1236
rect 276 -1240 280 -1236
rect 318 -1240 322 -1236
rect 360 -1240 364 -1236
rect 401 -1240 405 -1236
rect 209 -1264 213 -1260
rect 226 -1264 230 -1260
rect 191 -1433 195 -1429
rect 27 -1491 31 -1487
rect 197 -1491 201 -1487
rect -210 -1501 -206 -1497
rect -193 -1501 -189 -1497
rect -173 -1501 -169 -1497
rect -152 -1501 -148 -1497
rect -131 -1501 -127 -1497
rect -110 -1501 -106 -1497
rect -89 -1501 -85 -1497
rect -68 -1501 -64 -1497
rect -47 -1501 -43 -1497
rect -27 -1501 -23 -1497
rect -219 -1564 -215 -1560
rect -161 -1557 -157 -1553
rect -119 -1564 -115 -1560
rect -101 -1557 -97 -1553
rect -59 -1549 -55 -1545
rect -59 -1557 -55 -1553
rect -77 -1571 -73 -1567
rect -177 -1578 -173 -1574
rect -135 -1578 -131 -1574
rect -35 -1564 -31 -1560
rect -210 -1593 -206 -1589
rect -193 -1593 -189 -1589
rect -152 -1593 -148 -1589
rect -110 -1593 -106 -1589
rect -68 -1593 -64 -1589
rect -27 -1593 -23 -1589
rect -210 -1622 -206 -1618
rect -193 -1622 -189 -1618
rect -173 -1622 -169 -1618
rect -152 -1622 -148 -1618
rect -131 -1622 -127 -1618
rect -110 -1622 -106 -1618
rect -89 -1622 -85 -1618
rect -68 -1622 -64 -1618
rect -47 -1622 -43 -1618
rect -27 -1622 -23 -1618
rect -219 -1685 -215 -1681
rect -161 -1678 -157 -1674
rect -119 -1685 -115 -1681
rect -101 -1678 -97 -1674
rect -59 -1670 -55 -1666
rect -59 -1678 -55 -1674
rect -77 -1692 -73 -1688
rect -177 -1699 -173 -1695
rect -135 -1699 -131 -1695
rect -21 -1670 -17 -1666
rect -35 -1685 -31 -1681
rect -210 -1714 -206 -1710
rect -193 -1714 -189 -1710
rect -152 -1714 -148 -1710
rect -110 -1714 -106 -1710
rect -68 -1714 -64 -1710
rect -27 -1714 -23 -1710
rect 197 -1678 201 -1674
rect -21 -1721 -17 -1717
rect 197 -1722 201 -1718
rect -210 -1743 -206 -1739
rect -193 -1743 -189 -1739
rect -173 -1743 -169 -1739
rect -152 -1743 -148 -1739
rect -131 -1743 -127 -1739
rect -110 -1743 -106 -1739
rect -89 -1743 -85 -1739
rect -68 -1743 -64 -1739
rect -47 -1743 -43 -1739
rect -27 -1743 -23 -1739
rect -225 -1799 -221 -1795
rect -219 -1806 -215 -1802
rect -161 -1799 -157 -1795
rect -119 -1806 -115 -1802
rect -101 -1799 -97 -1795
rect -59 -1791 -55 -1787
rect -59 -1799 -55 -1795
rect -77 -1813 -73 -1809
rect -177 -1820 -173 -1816
rect -135 -1820 -131 -1816
rect -21 -1791 -17 -1787
rect -35 -1806 -31 -1802
rect -210 -1835 -206 -1831
rect -193 -1835 -189 -1831
rect -152 -1835 -148 -1831
rect -110 -1835 -106 -1831
rect -68 -1835 -64 -1831
rect -27 -1835 -23 -1831
rect -219 -1970 -215 -1966
rect -202 -1970 -198 -1966
rect -231 -2129 -227 -2125
rect -237 -2144 -233 -2140
rect -331 -2195 -327 -2191
rect -231 -2195 -227 -2191
rect -568 -2233 -564 -2229
rect -551 -2233 -547 -2229
rect -531 -2233 -527 -2229
rect -510 -2233 -506 -2229
rect -489 -2233 -485 -2229
rect -468 -2233 -464 -2229
rect -447 -2233 -443 -2229
rect -426 -2233 -422 -2229
rect -405 -2233 -401 -2229
rect -385 -2233 -381 -2229
rect -577 -2296 -573 -2292
rect -519 -2289 -515 -2285
rect -477 -2296 -473 -2292
rect -459 -2289 -455 -2285
rect -417 -2281 -413 -2277
rect -417 -2289 -413 -2285
rect -435 -2303 -431 -2299
rect -535 -2310 -531 -2306
rect -493 -2310 -489 -2306
rect -393 -2296 -389 -2292
rect -568 -2325 -564 -2321
rect -551 -2325 -547 -2321
rect -510 -2325 -506 -2321
rect -468 -2325 -464 -2321
rect -426 -2325 -422 -2321
rect -385 -2325 -381 -2321
rect -568 -2364 -564 -2360
rect -551 -2364 -547 -2360
rect -531 -2364 -527 -2360
rect -510 -2364 -506 -2360
rect -489 -2364 -485 -2360
rect -468 -2364 -464 -2360
rect -447 -2364 -443 -2360
rect -426 -2364 -422 -2360
rect -405 -2364 -401 -2360
rect -385 -2364 -381 -2360
rect -577 -2427 -573 -2423
rect -519 -2420 -515 -2416
rect -477 -2427 -473 -2423
rect -459 -2420 -455 -2416
rect -417 -2412 -413 -2408
rect -417 -2420 -413 -2416
rect -435 -2434 -431 -2430
rect -535 -2441 -531 -2437
rect -493 -2441 -489 -2437
rect -379 -2412 -375 -2408
rect -393 -2427 -389 -2423
rect -568 -2456 -564 -2452
rect -551 -2456 -547 -2452
rect -510 -2456 -506 -2452
rect -468 -2456 -464 -2452
rect -426 -2456 -422 -2452
rect -385 -2456 -381 -2452
rect -231 -2420 -227 -2416
rect -379 -2464 -375 -2460
rect -231 -2464 -227 -2460
rect -568 -2495 -564 -2491
rect -551 -2495 -547 -2491
rect -531 -2495 -527 -2491
rect -510 -2495 -506 -2491
rect -489 -2495 -485 -2491
rect -468 -2495 -464 -2491
rect -447 -2495 -443 -2491
rect -426 -2495 -422 -2491
rect -405 -2495 -401 -2491
rect -385 -2495 -381 -2491
rect -583 -2551 -579 -2547
rect -577 -2558 -573 -2554
rect -519 -2551 -515 -2547
rect -477 -2558 -473 -2554
rect -459 -2551 -455 -2547
rect -417 -2543 -413 -2539
rect -417 -2551 -413 -2547
rect -435 -2565 -431 -2561
rect -535 -2572 -531 -2568
rect -493 -2572 -489 -2568
rect -379 -2543 -375 -2539
rect -393 -2558 -389 -2554
rect -568 -2587 -564 -2583
rect -551 -2587 -547 -2583
rect -510 -2587 -506 -2583
rect -468 -2587 -464 -2583
rect -426 -2587 -422 -2583
rect -385 -2587 -381 -2583
rect -577 -2720 -573 -2716
rect -560 -2720 -556 -2716
rect -589 -2879 -585 -2875
rect -595 -2894 -591 -2890
rect -689 -2938 -685 -2934
rect -589 -2938 -585 -2934
rect -926 -2958 -922 -2954
rect -909 -2958 -905 -2954
rect -889 -2958 -885 -2954
rect -868 -2958 -864 -2954
rect -847 -2958 -843 -2954
rect -826 -2958 -822 -2954
rect -805 -2958 -801 -2954
rect -784 -2958 -780 -2954
rect -763 -2958 -759 -2954
rect -743 -2958 -739 -2954
rect -672 -2958 -668 -2954
rect -935 -3021 -931 -3017
rect -877 -3014 -873 -3010
rect -835 -3021 -831 -3017
rect -817 -3014 -813 -3010
rect -775 -2996 -771 -2992
rect -775 -3014 -771 -3010
rect -793 -3028 -789 -3024
rect -893 -3035 -889 -3031
rect -851 -3035 -847 -3031
rect -664 -3007 -660 -3003
rect -751 -3021 -747 -3017
rect -926 -3050 -922 -3046
rect -909 -3050 -905 -3046
rect -868 -3050 -864 -3046
rect -826 -3050 -822 -3046
rect -784 -3050 -780 -3046
rect -743 -3050 -739 -3046
rect -672 -3050 -668 -3046
rect -926 -3074 -922 -3070
rect -909 -3074 -905 -3070
rect -889 -3074 -885 -3070
rect -868 -3074 -864 -3070
rect -847 -3074 -843 -3070
rect -826 -3074 -822 -3070
rect -805 -3074 -801 -3070
rect -784 -3074 -780 -3070
rect -763 -3074 -759 -3070
rect -743 -3074 -739 -3070
rect -935 -3137 -931 -3133
rect -877 -3130 -873 -3126
rect -835 -3137 -831 -3133
rect -817 -3130 -813 -3126
rect -775 -3122 -771 -3118
rect -775 -3130 -771 -3126
rect -793 -3144 -789 -3140
rect -893 -3151 -889 -3147
rect -851 -3151 -847 -3147
rect -737 -3122 -733 -3118
rect -751 -3137 -747 -3133
rect -926 -3166 -922 -3162
rect -909 -3166 -905 -3162
rect -868 -3166 -864 -3162
rect -826 -3166 -822 -3162
rect -784 -3166 -780 -3162
rect -743 -3166 -739 -3162
rect -589 -3130 -585 -3126
rect -737 -3174 -733 -3170
rect -589 -3173 -585 -3169
rect -926 -3195 -922 -3191
rect -909 -3195 -905 -3191
rect -889 -3195 -885 -3191
rect -868 -3195 -864 -3191
rect -847 -3195 -843 -3191
rect -826 -3195 -822 -3191
rect -805 -3195 -801 -3191
rect -784 -3195 -780 -3191
rect -763 -3195 -759 -3191
rect -743 -3195 -739 -3191
rect -941 -3251 -937 -3247
rect -935 -3258 -931 -3254
rect -877 -3251 -873 -3247
rect -835 -3258 -831 -3254
rect -817 -3251 -813 -3247
rect -775 -3243 -771 -3239
rect -775 -3251 -771 -3247
rect -793 -3265 -789 -3261
rect -893 -3272 -889 -3268
rect -851 -3272 -847 -3268
rect -737 -3243 -733 -3239
rect -751 -3258 -747 -3254
rect -926 -3287 -922 -3283
rect -909 -3287 -905 -3283
rect -868 -3287 -864 -3283
rect -826 -3287 -822 -3283
rect -784 -3287 -780 -3283
rect -743 -3287 -739 -3283
rect -926 -3309 -922 -3305
rect -909 -3309 -905 -3305
rect -889 -3309 -885 -3305
rect -868 -3309 -864 -3305
rect -847 -3309 -843 -3305
rect -826 -3309 -822 -3305
rect -805 -3309 -801 -3305
rect -784 -3309 -780 -3305
rect -763 -3309 -759 -3305
rect -743 -3309 -739 -3305
rect -935 -3372 -931 -3368
rect -877 -3365 -873 -3361
rect -835 -3372 -831 -3368
rect -817 -3365 -813 -3361
rect -775 -3357 -771 -3353
rect -775 -3365 -771 -3361
rect -793 -3379 -789 -3375
rect -893 -3386 -889 -3382
rect -851 -3386 -847 -3382
rect -751 -3372 -747 -3368
rect -926 -3401 -922 -3397
rect -909 -3401 -905 -3397
rect -868 -3401 -864 -3397
rect -826 -3401 -822 -3397
rect -784 -3401 -780 -3397
rect -743 -3401 -739 -3397
rect -935 -3426 -931 -3422
rect -918 -3426 -914 -3422
rect -947 -3605 -943 -3601
rect -1162 -3620 -1158 -3616
rect -1255 -3642 -1251 -3638
rect -1211 -3642 -1207 -3638
rect -1177 -3642 -1173 -3638
rect -1276 -3649 -1272 -3645
rect -1270 -3656 -1266 -3652
rect -1162 -3656 -1158 -3652
rect -947 -3656 -943 -3652
rect -1255 -3680 -1251 -3676
rect -1238 -3680 -1234 -3676
rect -1218 -3680 -1214 -3676
rect -1197 -3680 -1193 -3676
rect -1176 -3680 -1172 -3676
rect -1155 -3680 -1151 -3676
rect -1134 -3680 -1130 -3676
rect -1113 -3680 -1109 -3676
rect -1092 -3680 -1088 -3676
rect -1072 -3680 -1068 -3676
rect -1270 -3736 -1266 -3732
rect -1264 -3743 -1260 -3739
rect -1206 -3736 -1202 -3732
rect -1164 -3743 -1160 -3739
rect -1146 -3736 -1142 -3732
rect -1104 -3728 -1100 -3724
rect -1104 -3736 -1100 -3732
rect -1122 -3750 -1118 -3746
rect -1222 -3757 -1218 -3753
rect -1180 -3757 -1176 -3753
rect -1080 -3743 -1076 -3739
rect -1255 -3772 -1251 -3768
rect -1238 -3772 -1234 -3768
rect -1197 -3772 -1193 -3768
rect -1155 -3772 -1151 -3768
rect -1113 -3772 -1109 -3768
rect -1072 -3772 -1068 -3768
rect -1255 -3911 -1251 -3907
rect -1238 -3911 -1234 -3907
rect -1218 -3911 -1214 -3907
rect -1197 -3911 -1193 -3907
rect -1176 -3911 -1172 -3907
rect -1155 -3911 -1151 -3907
rect -1134 -3911 -1130 -3907
rect -1113 -3911 -1109 -3907
rect -1092 -3911 -1088 -3907
rect -1072 -3911 -1068 -3907
rect -1276 -3967 -1272 -3963
rect -1264 -3974 -1260 -3970
rect -1206 -3967 -1202 -3963
rect -1164 -3974 -1160 -3970
rect -1146 -3967 -1142 -3963
rect -1104 -3959 -1100 -3955
rect -1104 -3967 -1100 -3963
rect -1122 -3981 -1118 -3977
rect -1222 -3988 -1218 -3984
rect -1180 -3988 -1176 -3984
rect -1066 -3959 -1062 -3955
rect -1080 -3974 -1076 -3970
rect -1255 -4003 -1251 -3999
rect -1238 -4003 -1234 -3999
rect -1197 -4003 -1193 -3999
rect -1155 -4003 -1151 -3999
rect -1113 -4003 -1109 -3999
rect -1072 -4003 -1068 -3999
rect -947 -3967 -943 -3963
rect -1349 -4092 -1345 -4088
rect -1270 -4010 -1266 -4006
rect -1066 -4010 -1062 -4006
rect -1339 -4271 -1335 -4267
rect -1322 -4271 -1318 -4267
rect -1322 -4363 -1318 -4359
rect -947 -4011 -943 -4007
rect -1255 -4036 -1251 -4032
rect -1238 -4036 -1234 -4032
rect -1218 -4036 -1214 -4032
rect -1197 -4036 -1193 -4032
rect -1176 -4036 -1172 -4032
rect -1155 -4036 -1151 -4032
rect -1134 -4036 -1130 -4032
rect -1113 -4036 -1109 -4032
rect -1092 -4036 -1088 -4032
rect -1072 -4036 -1068 -4032
rect -1264 -4099 -1260 -4095
rect -1206 -4092 -1202 -4088
rect -1164 -4099 -1160 -4095
rect -1146 -4092 -1142 -4088
rect -1104 -4084 -1100 -4080
rect -1104 -4092 -1100 -4088
rect -1122 -4106 -1118 -4102
rect -1222 -4113 -1218 -4109
rect -1180 -4113 -1176 -4109
rect -1066 -4084 -1062 -4080
rect -1080 -4099 -1076 -4095
rect -1255 -4128 -1251 -4124
rect -1238 -4128 -1234 -4124
rect -1197 -4128 -1193 -4124
rect -1155 -4128 -1151 -4124
rect -1113 -4128 -1109 -4124
rect -1072 -4128 -1068 -4124
rect -1255 -4160 -1251 -4156
rect -1238 -4160 -1234 -4156
rect -1218 -4160 -1214 -4156
rect -1197 -4160 -1193 -4156
rect -1176 -4160 -1172 -4156
rect -1155 -4160 -1151 -4156
rect -1134 -4160 -1130 -4156
rect -1113 -4160 -1109 -4156
rect -1092 -4160 -1088 -4156
rect -1072 -4160 -1068 -4156
rect -1264 -4223 -1260 -4219
rect -1206 -4216 -1202 -4212
rect -1164 -4223 -1160 -4219
rect -1146 -4216 -1142 -4212
rect -1104 -4183 -1100 -4179
rect -1104 -4216 -1100 -4212
rect -1122 -4230 -1118 -4226
rect -1222 -4237 -1218 -4233
rect -1180 -4237 -1176 -4233
rect -1080 -4223 -1076 -4219
rect -1255 -4252 -1251 -4248
rect -1238 -4252 -1234 -4248
rect -1197 -4252 -1193 -4248
rect -1155 -4252 -1151 -4248
rect -1113 -4252 -1109 -4248
rect -1072 -4252 -1068 -4248
rect -1029 -4160 -1025 -4156
rect -1021 -4205 -1017 -4201
rect -1029 -4252 -1025 -4248
rect -1029 -4271 -1025 -4267
rect -1066 -4303 -1062 -4299
rect -1021 -4320 -1017 -4316
rect -953 -4324 -949 -4320
rect -1029 -4363 -1025 -4359
rect -1255 -4390 -1251 -4386
rect -1238 -4390 -1234 -4386
rect -1198 -4390 -1194 -4386
rect -1177 -4390 -1173 -4386
rect -1270 -4446 -1266 -4442
rect -1264 -4439 -1260 -4435
rect -1313 -4453 -1309 -4449
rect -1220 -4460 -1216 -4456
rect -953 -4430 -949 -4426
rect -1168 -4438 -1164 -4434
rect -1238 -4467 -1234 -4463
rect -1202 -4467 -1198 -4463
rect -737 -3458 -733 -3454
rect -909 -3479 -905 -3475
rect -595 -3479 -591 -3475
rect -918 -3518 -914 -3514
rect -926 -3550 -922 -3546
rect -900 -3550 -896 -3546
rect -883 -3550 -879 -3546
rect -843 -3550 -839 -3546
rect -822 -3550 -818 -3546
rect -805 -3550 -801 -3546
rect -765 -3550 -761 -3546
rect -741 -3550 -737 -3546
rect -704 -3550 -700 -3546
rect -935 -3583 -931 -3579
rect -917 -3576 -913 -3572
rect -891 -3598 -887 -3594
rect -909 -3605 -905 -3601
rect -865 -3590 -861 -3586
rect -813 -3583 -809 -3579
rect -883 -3627 -879 -3623
rect -847 -3627 -843 -3623
rect -787 -3598 -783 -3594
rect -805 -3627 -801 -3623
rect -769 -3627 -765 -3623
rect -695 -3590 -691 -3586
rect -689 -3598 -685 -3594
rect -926 -3642 -922 -3638
rect -900 -3642 -896 -3638
rect -857 -3642 -853 -3638
rect -822 -3642 -818 -3638
rect -778 -3642 -774 -3638
rect -761 -3642 -757 -3638
rect -725 -3642 -721 -3638
rect -704 -3642 -700 -3638
rect -379 -2752 -375 -2748
rect -551 -2773 -547 -2769
rect -237 -2773 -233 -2769
rect -560 -2812 -556 -2808
rect -568 -2839 -564 -2835
rect -542 -2839 -538 -2835
rect -525 -2839 -521 -2835
rect -485 -2839 -481 -2835
rect -464 -2839 -460 -2835
rect -447 -2839 -443 -2835
rect -407 -2839 -403 -2835
rect -383 -2839 -379 -2835
rect -346 -2839 -342 -2835
rect -577 -2872 -573 -2868
rect -559 -2865 -555 -2861
rect -533 -2887 -529 -2883
rect -551 -2894 -547 -2890
rect -507 -2879 -503 -2875
rect -455 -2872 -451 -2868
rect -525 -2916 -521 -2912
rect -489 -2916 -485 -2912
rect -429 -2887 -425 -2883
rect -447 -2916 -443 -2912
rect -411 -2916 -407 -2912
rect -337 -2878 -333 -2874
rect -331 -2887 -327 -2883
rect -568 -2931 -564 -2927
rect -542 -2931 -538 -2927
rect -499 -2931 -495 -2927
rect -464 -2931 -460 -2927
rect -420 -2931 -416 -2927
rect -403 -2931 -399 -2927
rect -367 -2931 -363 -2927
rect -346 -2931 -342 -2927
rect -21 -2002 -17 -1998
rect -193 -2023 -189 -2019
rect 191 -2023 195 -2019
rect -202 -2062 -198 -2058
rect -210 -2089 -206 -2085
rect -184 -2089 -180 -2085
rect -167 -2089 -163 -2085
rect -127 -2089 -123 -2085
rect -106 -2089 -102 -2085
rect -89 -2089 -85 -2085
rect -49 -2089 -45 -2085
rect -25 -2089 -21 -2085
rect 12 -2089 16 -2085
rect -219 -2122 -215 -2118
rect -201 -2115 -197 -2111
rect -175 -2137 -171 -2133
rect -193 -2144 -189 -2140
rect -149 -2129 -145 -2125
rect -97 -2122 -93 -2118
rect -167 -2166 -163 -2162
rect -131 -2166 -127 -2162
rect -71 -2137 -67 -2133
rect -89 -2166 -85 -2162
rect -53 -2166 -49 -2162
rect 21 -2129 25 -2125
rect 27 -2137 31 -2133
rect -210 -2181 -206 -2177
rect -184 -2181 -180 -2177
rect -141 -2181 -137 -2177
rect -106 -2181 -102 -2177
rect -62 -2181 -58 -2177
rect -45 -2181 -41 -2177
rect -9 -2181 -5 -2177
rect 12 -2181 16 -2177
rect 235 -1317 239 -1313
rect 547 -1317 551 -1313
rect 226 -1356 230 -1352
rect 218 -1378 222 -1374
rect 244 -1378 248 -1374
rect 261 -1378 265 -1374
rect 301 -1378 305 -1374
rect 322 -1378 326 -1374
rect 339 -1378 343 -1374
rect 379 -1378 383 -1374
rect 403 -1378 407 -1374
rect 440 -1378 444 -1374
rect 209 -1411 213 -1407
rect 227 -1404 231 -1400
rect 253 -1426 257 -1422
rect 235 -1433 239 -1429
rect 279 -1418 283 -1414
rect 331 -1411 335 -1407
rect 261 -1455 265 -1451
rect 297 -1455 301 -1451
rect 357 -1426 361 -1422
rect 339 -1455 343 -1451
rect 375 -1455 379 -1451
rect 449 -1418 453 -1414
rect 455 -1426 459 -1422
rect 218 -1470 222 -1466
rect 244 -1470 248 -1466
rect 287 -1470 291 -1466
rect 322 -1470 326 -1466
rect 366 -1470 370 -1466
rect 383 -1470 387 -1466
rect 419 -1470 423 -1466
rect 440 -1470 444 -1466
rect 553 -1418 557 -1414
rect 963 -1034 967 -1030
rect 980 -1034 984 -1030
rect 591 -1090 595 -1086
rect 951 -1090 955 -1086
rect 582 -1126 586 -1122
rect 574 -1148 578 -1144
rect 591 -1148 595 -1144
rect 611 -1148 615 -1144
rect 632 -1148 636 -1144
rect 653 -1148 657 -1144
rect 674 -1148 678 -1144
rect 695 -1148 699 -1144
rect 716 -1148 720 -1144
rect 737 -1148 741 -1144
rect 757 -1148 761 -1144
rect 565 -1211 569 -1207
rect 623 -1204 627 -1200
rect 665 -1211 669 -1207
rect 683 -1204 687 -1200
rect 725 -1196 729 -1192
rect 725 -1204 729 -1200
rect 707 -1218 711 -1214
rect 607 -1225 611 -1221
rect 649 -1225 653 -1221
rect 749 -1211 753 -1207
rect 574 -1240 578 -1236
rect 591 -1240 595 -1236
rect 632 -1240 636 -1236
rect 674 -1240 678 -1236
rect 716 -1240 720 -1236
rect 757 -1240 761 -1236
rect 565 -1264 569 -1260
rect 582 -1264 586 -1260
rect 547 -1433 551 -1429
rect 455 -1484 459 -1480
rect 553 -1484 557 -1480
rect 218 -1501 222 -1497
rect 235 -1501 239 -1497
rect 255 -1501 259 -1497
rect 276 -1501 280 -1497
rect 297 -1501 301 -1497
rect 318 -1501 322 -1497
rect 339 -1501 343 -1497
rect 360 -1501 364 -1497
rect 381 -1501 385 -1497
rect 401 -1501 405 -1497
rect 209 -1564 213 -1560
rect 267 -1557 271 -1553
rect 309 -1564 313 -1560
rect 327 -1557 331 -1553
rect 369 -1549 373 -1545
rect 369 -1557 373 -1553
rect 351 -1571 355 -1567
rect 251 -1578 255 -1574
rect 293 -1578 297 -1574
rect 393 -1564 397 -1560
rect 218 -1593 222 -1589
rect 235 -1593 239 -1589
rect 276 -1593 280 -1589
rect 318 -1593 322 -1589
rect 360 -1593 364 -1589
rect 401 -1593 405 -1589
rect 218 -1622 222 -1618
rect 235 -1622 239 -1618
rect 255 -1622 259 -1618
rect 276 -1622 280 -1618
rect 297 -1622 301 -1618
rect 318 -1622 322 -1618
rect 339 -1622 343 -1618
rect 360 -1622 364 -1618
rect 381 -1622 385 -1618
rect 401 -1622 405 -1618
rect 209 -1685 213 -1681
rect 267 -1678 271 -1674
rect 309 -1685 313 -1681
rect 327 -1678 331 -1674
rect 369 -1670 373 -1666
rect 369 -1678 373 -1674
rect 351 -1692 355 -1688
rect 251 -1699 255 -1695
rect 293 -1699 297 -1695
rect 407 -1670 411 -1666
rect 393 -1685 397 -1681
rect 218 -1714 222 -1710
rect 235 -1714 239 -1710
rect 276 -1714 280 -1710
rect 318 -1714 322 -1710
rect 360 -1714 364 -1710
rect 401 -1714 405 -1710
rect 553 -1678 557 -1674
rect 407 -1722 411 -1718
rect 553 -1721 557 -1717
rect 218 -1743 222 -1739
rect 235 -1743 239 -1739
rect 255 -1743 259 -1739
rect 276 -1743 280 -1739
rect 297 -1743 301 -1739
rect 318 -1743 322 -1739
rect 339 -1743 343 -1739
rect 360 -1743 364 -1739
rect 381 -1743 385 -1739
rect 401 -1743 405 -1739
rect 203 -1799 207 -1795
rect 464 -1743 468 -1739
rect 209 -1806 213 -1802
rect 267 -1799 271 -1795
rect 309 -1806 313 -1802
rect 327 -1799 331 -1795
rect 369 -1791 373 -1787
rect 369 -1799 373 -1795
rect 351 -1813 355 -1809
rect 251 -1820 255 -1816
rect 293 -1820 297 -1816
rect 407 -1791 411 -1787
rect 393 -1806 397 -1802
rect 218 -1835 222 -1831
rect 235 -1835 239 -1831
rect 276 -1835 280 -1831
rect 318 -1835 322 -1831
rect 360 -1835 364 -1831
rect 401 -1835 405 -1831
rect 209 -1970 213 -1966
rect 226 -1970 230 -1966
rect 197 -2129 201 -2125
rect 191 -2144 195 -2140
rect 27 -2188 31 -2184
rect 197 -2188 201 -2184
rect -210 -2233 -206 -2229
rect -193 -2233 -189 -2229
rect -173 -2233 -169 -2229
rect -152 -2233 -148 -2229
rect -131 -2233 -127 -2229
rect -110 -2233 -106 -2229
rect -89 -2233 -85 -2229
rect -68 -2233 -64 -2229
rect -47 -2233 -43 -2229
rect -27 -2233 -23 -2229
rect -219 -2296 -215 -2292
rect -161 -2289 -157 -2285
rect -119 -2296 -115 -2292
rect -101 -2289 -97 -2285
rect -59 -2281 -55 -2277
rect -59 -2289 -55 -2285
rect -77 -2303 -73 -2299
rect -177 -2310 -173 -2306
rect -135 -2310 -131 -2306
rect -35 -2296 -31 -2292
rect -210 -2325 -206 -2321
rect -193 -2325 -189 -2321
rect -152 -2325 -148 -2321
rect -110 -2325 -106 -2321
rect -68 -2325 -64 -2321
rect -27 -2325 -23 -2321
rect -210 -2364 -206 -2360
rect -193 -2364 -189 -2360
rect -173 -2364 -169 -2360
rect -152 -2364 -148 -2360
rect -131 -2364 -127 -2360
rect -110 -2364 -106 -2360
rect -89 -2364 -85 -2360
rect -68 -2364 -64 -2360
rect -47 -2364 -43 -2360
rect -27 -2364 -23 -2360
rect -219 -2427 -215 -2423
rect -161 -2420 -157 -2416
rect -119 -2427 -115 -2423
rect -101 -2420 -97 -2416
rect -59 -2412 -55 -2408
rect -59 -2420 -55 -2416
rect -77 -2434 -73 -2430
rect -177 -2441 -173 -2437
rect -135 -2441 -131 -2437
rect -21 -2412 -17 -2408
rect -35 -2427 -31 -2423
rect -210 -2456 -206 -2452
rect -193 -2456 -189 -2452
rect -152 -2456 -148 -2452
rect -110 -2456 -106 -2452
rect -68 -2456 -64 -2452
rect -27 -2456 -23 -2452
rect 197 -2420 201 -2416
rect -21 -2464 -17 -2460
rect 197 -2463 201 -2459
rect -210 -2495 -206 -2491
rect -193 -2495 -189 -2491
rect -173 -2495 -169 -2491
rect -152 -2495 -148 -2491
rect -131 -2495 -127 -2491
rect -110 -2495 -106 -2491
rect -89 -2495 -85 -2491
rect -68 -2495 -64 -2491
rect -47 -2495 -43 -2491
rect -27 -2495 -23 -2491
rect -225 -2551 -221 -2547
rect 90 -2495 94 -2491
rect -219 -2558 -215 -2554
rect -161 -2551 -157 -2547
rect -119 -2558 -115 -2554
rect -101 -2551 -97 -2547
rect -59 -2543 -55 -2539
rect -59 -2551 -55 -2547
rect -77 -2565 -73 -2561
rect -177 -2572 -173 -2568
rect -135 -2572 -131 -2568
rect -21 -2543 -17 -2539
rect -35 -2558 -31 -2554
rect -210 -2587 -206 -2583
rect -193 -2587 -189 -2583
rect -152 -2587 -148 -2583
rect -110 -2587 -106 -2583
rect -68 -2587 -64 -2583
rect -27 -2587 -23 -2583
rect -219 -2720 -215 -2716
rect -202 -2720 -198 -2716
rect -231 -2879 -227 -2875
rect -237 -2894 -233 -2890
rect -331 -2945 -327 -2941
rect -231 -2945 -227 -2941
rect -568 -2958 -564 -2954
rect -551 -2958 -547 -2954
rect -531 -2958 -527 -2954
rect -510 -2958 -506 -2954
rect -489 -2958 -485 -2954
rect -468 -2958 -464 -2954
rect -447 -2958 -443 -2954
rect -426 -2958 -422 -2954
rect -405 -2958 -401 -2954
rect -385 -2958 -381 -2954
rect -329 -2958 -325 -2954
rect -577 -3021 -573 -3017
rect -519 -3014 -515 -3010
rect -477 -3021 -473 -3017
rect -459 -3014 -455 -3010
rect -417 -2980 -413 -2976
rect -417 -3014 -413 -3010
rect -435 -3028 -431 -3024
rect -535 -3035 -531 -3031
rect -493 -3035 -489 -3031
rect -321 -3009 -317 -3005
rect -393 -3021 -389 -3017
rect -568 -3050 -564 -3046
rect -551 -3050 -547 -3046
rect -510 -3050 -506 -3046
rect -468 -3050 -464 -3046
rect -426 -3050 -422 -3046
rect -385 -3050 -381 -3046
rect -329 -3050 -325 -3046
rect -568 -3074 -564 -3070
rect -551 -3074 -547 -3070
rect -531 -3074 -527 -3070
rect -510 -3074 -506 -3070
rect -489 -3074 -485 -3070
rect -468 -3074 -464 -3070
rect -447 -3074 -443 -3070
rect -426 -3074 -422 -3070
rect -405 -3074 -401 -3070
rect -385 -3074 -381 -3070
rect -329 -3074 -325 -3070
rect -577 -3137 -573 -3133
rect -519 -3130 -515 -3126
rect -477 -3137 -473 -3133
rect -459 -3130 -455 -3126
rect -417 -3122 -413 -3118
rect -417 -3130 -413 -3126
rect -435 -3144 -431 -3140
rect -535 -3151 -531 -3147
rect -493 -3151 -489 -3147
rect -379 -3122 -375 -3118
rect -393 -3137 -389 -3133
rect -568 -3166 -564 -3162
rect -551 -3166 -547 -3162
rect -510 -3166 -506 -3162
rect -468 -3166 -464 -3162
rect -426 -3166 -422 -3162
rect -385 -3166 -381 -3162
rect -321 -3124 -317 -3120
rect -231 -3130 -227 -3126
rect -329 -3166 -325 -3162
rect -379 -3173 -375 -3169
rect -231 -3174 -227 -3170
rect -568 -3195 -564 -3191
rect -551 -3195 -547 -3191
rect -531 -3195 -527 -3191
rect -510 -3195 -506 -3191
rect -489 -3195 -485 -3191
rect -468 -3195 -464 -3191
rect -447 -3195 -443 -3191
rect -426 -3195 -422 -3191
rect -405 -3195 -401 -3191
rect -385 -3195 -381 -3191
rect -583 -3251 -579 -3247
rect -577 -3258 -573 -3254
rect -519 -3251 -515 -3247
rect -477 -3258 -473 -3254
rect -459 -3251 -455 -3247
rect -417 -3243 -413 -3239
rect -417 -3251 -413 -3247
rect -435 -3265 -431 -3261
rect -535 -3272 -531 -3268
rect -493 -3272 -489 -3268
rect -373 -3243 -369 -3239
rect -393 -3258 -389 -3254
rect -568 -3287 -564 -3283
rect -551 -3287 -547 -3283
rect -510 -3287 -506 -3283
rect -468 -3287 -464 -3283
rect -426 -3287 -422 -3283
rect -385 -3287 -381 -3283
rect -568 -3309 -564 -3305
rect -551 -3309 -547 -3305
rect -531 -3309 -527 -3305
rect -510 -3309 -506 -3305
rect -489 -3309 -485 -3305
rect -468 -3309 -464 -3305
rect -447 -3309 -443 -3305
rect -426 -3309 -422 -3305
rect -405 -3309 -401 -3305
rect -385 -3309 -381 -3305
rect -577 -3372 -573 -3368
rect -519 -3365 -515 -3361
rect -477 -3372 -473 -3368
rect -459 -3365 -455 -3361
rect -417 -3357 -413 -3353
rect -417 -3365 -413 -3361
rect -435 -3379 -431 -3375
rect -535 -3386 -531 -3382
rect -493 -3386 -489 -3382
rect -379 -3357 -375 -3353
rect -393 -3372 -389 -3368
rect -568 -3401 -564 -3397
rect -551 -3401 -547 -3397
rect -510 -3401 -506 -3397
rect -468 -3401 -464 -3397
rect -426 -3401 -422 -3397
rect -385 -3401 -381 -3397
rect -577 -3426 -573 -3422
rect -560 -3426 -556 -3422
rect -589 -3590 -585 -3586
rect -595 -3605 -591 -3601
rect -689 -3649 -685 -3645
rect -589 -3649 -585 -3645
rect -926 -3680 -922 -3676
rect -909 -3680 -905 -3676
rect -889 -3680 -885 -3676
rect -868 -3680 -864 -3676
rect -847 -3680 -843 -3676
rect -826 -3680 -822 -3676
rect -805 -3680 -801 -3676
rect -784 -3680 -780 -3676
rect -763 -3680 -759 -3676
rect -743 -3680 -739 -3676
rect -935 -3743 -931 -3739
rect -877 -3736 -873 -3732
rect -835 -3743 -831 -3739
rect -817 -3736 -813 -3732
rect -775 -3728 -771 -3724
rect -775 -3736 -771 -3732
rect -793 -3750 -789 -3746
rect -893 -3757 -889 -3753
rect -851 -3757 -847 -3753
rect -751 -3743 -747 -3739
rect -926 -3772 -922 -3768
rect -909 -3772 -905 -3768
rect -868 -3772 -864 -3768
rect -826 -3772 -822 -3768
rect -784 -3772 -780 -3768
rect -743 -3772 -739 -3768
rect -926 -3911 -922 -3907
rect -909 -3911 -905 -3907
rect -889 -3911 -885 -3907
rect -868 -3911 -864 -3907
rect -847 -3911 -843 -3907
rect -826 -3911 -822 -3907
rect -805 -3911 -801 -3907
rect -784 -3911 -780 -3907
rect -763 -3911 -759 -3907
rect -743 -3911 -739 -3907
rect -935 -3974 -931 -3970
rect -877 -3967 -873 -3963
rect -835 -3974 -831 -3970
rect -817 -3967 -813 -3963
rect -775 -3959 -771 -3955
rect -775 -3967 -771 -3963
rect -793 -3981 -789 -3977
rect -893 -3988 -889 -3984
rect -851 -3988 -847 -3984
rect -737 -3959 -733 -3955
rect -751 -3974 -747 -3970
rect -926 -4003 -922 -3999
rect -909 -4003 -905 -3999
rect -868 -4003 -864 -3999
rect -826 -4003 -822 -3999
rect -784 -4003 -780 -3999
rect -743 -4003 -739 -3999
rect -589 -3967 -585 -3963
rect -737 -4011 -733 -4007
rect -589 -4010 -585 -4006
rect -926 -4036 -922 -4032
rect -909 -4036 -905 -4032
rect -889 -4036 -885 -4032
rect -868 -4036 -864 -4032
rect -847 -4036 -843 -4032
rect -826 -4036 -822 -4032
rect -805 -4036 -801 -4032
rect -784 -4036 -780 -4032
rect -763 -4036 -759 -4032
rect -743 -4036 -739 -4032
rect -941 -4092 -937 -4088
rect -935 -4099 -931 -4095
rect -877 -4092 -873 -4088
rect -835 -4099 -831 -4095
rect -817 -4092 -813 -4088
rect -775 -4084 -771 -4080
rect -775 -4092 -771 -4088
rect -793 -4106 -789 -4102
rect -893 -4113 -889 -4109
rect -851 -4113 -847 -4109
rect -737 -4084 -733 -4080
rect -751 -4099 -747 -4095
rect -926 -4128 -922 -4124
rect -909 -4128 -905 -4124
rect -868 -4128 -864 -4124
rect -826 -4128 -822 -4124
rect -784 -4128 -780 -4124
rect -743 -4128 -739 -4124
rect -926 -4160 -922 -4156
rect -909 -4160 -905 -4156
rect -889 -4160 -885 -4156
rect -868 -4160 -864 -4156
rect -847 -4160 -843 -4156
rect -826 -4160 -822 -4156
rect -805 -4160 -801 -4156
rect -784 -4160 -780 -4156
rect -763 -4160 -759 -4156
rect -743 -4160 -739 -4156
rect -935 -4223 -931 -4219
rect -877 -4216 -873 -4212
rect -835 -4223 -831 -4219
rect -817 -4216 -813 -4212
rect -775 -4208 -771 -4204
rect -775 -4216 -771 -4212
rect -793 -4230 -789 -4226
rect -893 -4237 -889 -4233
rect -851 -4237 -847 -4233
rect -751 -4223 -747 -4219
rect -926 -4252 -922 -4248
rect -909 -4252 -905 -4248
rect -868 -4252 -864 -4248
rect -826 -4252 -822 -4248
rect -784 -4252 -780 -4248
rect -743 -4252 -739 -4248
rect -935 -4271 -931 -4267
rect -918 -4271 -914 -4267
rect -947 -4445 -943 -4441
rect -1162 -4460 -1158 -4456
rect -1255 -4482 -1251 -4478
rect -1211 -4482 -1207 -4478
rect -1177 -4482 -1173 -4478
rect -1276 -4489 -1272 -4485
rect -1270 -4496 -1266 -4492
rect -1162 -4496 -1158 -4492
rect -947 -4496 -943 -4492
rect -1255 -4513 -1251 -4509
rect -1238 -4513 -1234 -4509
rect -1218 -4513 -1214 -4509
rect -1197 -4513 -1193 -4509
rect -1176 -4513 -1172 -4509
rect -1155 -4513 -1151 -4509
rect -1134 -4513 -1130 -4509
rect -1113 -4513 -1109 -4509
rect -1092 -4513 -1088 -4509
rect -1072 -4513 -1068 -4509
rect -1270 -4569 -1266 -4565
rect -1264 -4576 -1260 -4572
rect -1206 -4569 -1202 -4565
rect -1164 -4576 -1160 -4572
rect -1146 -4569 -1142 -4565
rect -1104 -4561 -1100 -4557
rect -1104 -4569 -1100 -4565
rect -1122 -4583 -1118 -4579
rect -1222 -4590 -1218 -4586
rect -1180 -4590 -1176 -4586
rect -1080 -4576 -1076 -4572
rect -1255 -4605 -1251 -4601
rect -1238 -4605 -1234 -4601
rect -1197 -4605 -1193 -4601
rect -1155 -4605 -1151 -4601
rect -1113 -4605 -1109 -4601
rect -1072 -4605 -1068 -4601
rect -1255 -4634 -1251 -4630
rect -1238 -4634 -1234 -4630
rect -1218 -4634 -1214 -4630
rect -1197 -4634 -1193 -4630
rect -1176 -4634 -1172 -4630
rect -1155 -4634 -1151 -4630
rect -1134 -4634 -1130 -4630
rect -1113 -4634 -1109 -4630
rect -1092 -4634 -1088 -4630
rect -1072 -4634 -1068 -4630
rect -1276 -4690 -1272 -4686
rect -1264 -4697 -1260 -4693
rect -1206 -4690 -1202 -4686
rect -1164 -4697 -1160 -4693
rect -1146 -4690 -1142 -4686
rect -1104 -4682 -1100 -4678
rect -1104 -4690 -1100 -4686
rect -1122 -4704 -1118 -4700
rect -1222 -4711 -1218 -4707
rect -1180 -4711 -1176 -4707
rect -1066 -4682 -1062 -4678
rect -1080 -4697 -1076 -4693
rect -1255 -4726 -1251 -4722
rect -1238 -4726 -1234 -4722
rect -1197 -4726 -1193 -4722
rect -1155 -4726 -1151 -4722
rect -1113 -4726 -1109 -4722
rect -1072 -4726 -1068 -4722
rect -947 -4690 -943 -4686
rect -1349 -4811 -1345 -4807
rect -1270 -4734 -1266 -4730
rect -1066 -4734 -1062 -4730
rect -947 -4733 -943 -4729
rect -1339 -4990 -1335 -4986
rect -1322 -4990 -1318 -4986
rect -1322 -5082 -1318 -5078
rect -1255 -4755 -1251 -4751
rect -1238 -4755 -1234 -4751
rect -1218 -4755 -1214 -4751
rect -1197 -4755 -1193 -4751
rect -1176 -4755 -1172 -4751
rect -1155 -4755 -1151 -4751
rect -1134 -4755 -1130 -4751
rect -1113 -4755 -1109 -4751
rect -1092 -4755 -1088 -4751
rect -1072 -4755 -1068 -4751
rect -1264 -4818 -1260 -4814
rect -1206 -4811 -1202 -4807
rect -1164 -4818 -1160 -4814
rect -1146 -4811 -1142 -4807
rect -1104 -4803 -1100 -4799
rect -1104 -4811 -1100 -4807
rect -1122 -4825 -1118 -4821
rect -1222 -4832 -1218 -4828
rect -1180 -4832 -1176 -4828
rect -1066 -4803 -1062 -4799
rect -1080 -4818 -1076 -4814
rect -1255 -4847 -1251 -4843
rect -1238 -4847 -1234 -4843
rect -1197 -4847 -1193 -4843
rect -1155 -4847 -1151 -4843
rect -1113 -4847 -1109 -4843
rect -1072 -4847 -1068 -4843
rect -1255 -4873 -1251 -4869
rect -1238 -4873 -1234 -4869
rect -1218 -4873 -1214 -4869
rect -1197 -4873 -1193 -4869
rect -1176 -4873 -1172 -4869
rect -1155 -4873 -1151 -4869
rect -1134 -4873 -1130 -4869
rect -1113 -4873 -1109 -4869
rect -1092 -4873 -1088 -4869
rect -1072 -4873 -1068 -4869
rect -1264 -4936 -1260 -4932
rect -1206 -4929 -1202 -4925
rect -1164 -4936 -1160 -4932
rect -1146 -4929 -1142 -4925
rect -1104 -4921 -1100 -4917
rect -1104 -4929 -1100 -4925
rect -1122 -4943 -1118 -4939
rect -1222 -4950 -1218 -4946
rect -1180 -4950 -1176 -4946
rect -1080 -4936 -1076 -4932
rect -1255 -4965 -1251 -4961
rect -1238 -4965 -1234 -4961
rect -1197 -4965 -1193 -4961
rect -1155 -4965 -1151 -4961
rect -1113 -4965 -1109 -4961
rect -1072 -4965 -1068 -4961
rect -1066 -5022 -1062 -5018
rect -953 -5043 -949 -5039
rect -1255 -5109 -1251 -5105
rect -1238 -5109 -1234 -5105
rect -1198 -5109 -1194 -5105
rect -1177 -5109 -1173 -5105
rect -1270 -5165 -1266 -5161
rect -1264 -5158 -1260 -5154
rect -1313 -5172 -1309 -5168
rect -1220 -5179 -1216 -5175
rect -953 -5149 -949 -5145
rect -1168 -5157 -1164 -5153
rect -1238 -5186 -1234 -5182
rect -1202 -5186 -1198 -5182
rect -673 -4271 -669 -4267
rect -737 -4303 -733 -4299
rect -909 -4324 -905 -4320
rect -665 -4321 -661 -4317
rect -595 -4324 -591 -4320
rect -918 -4363 -914 -4359
rect -673 -4363 -669 -4359
rect -926 -4390 -922 -4386
rect -900 -4390 -896 -4386
rect -883 -4390 -879 -4386
rect -843 -4390 -839 -4386
rect -822 -4390 -818 -4386
rect -805 -4390 -801 -4386
rect -765 -4390 -761 -4386
rect -741 -4390 -737 -4386
rect -704 -4390 -700 -4386
rect -935 -4423 -931 -4419
rect -917 -4416 -913 -4412
rect -891 -4438 -887 -4434
rect -909 -4445 -905 -4441
rect -865 -4430 -861 -4426
rect -813 -4423 -809 -4419
rect -883 -4467 -879 -4463
rect -847 -4467 -843 -4463
rect -787 -4438 -783 -4434
rect -805 -4467 -801 -4463
rect -769 -4467 -765 -4463
rect -695 -4430 -691 -4426
rect -689 -4438 -685 -4434
rect -926 -4482 -922 -4478
rect -900 -4482 -896 -4478
rect -857 -4482 -853 -4478
rect -822 -4482 -818 -4478
rect -778 -4482 -774 -4478
rect -761 -4482 -757 -4478
rect -725 -4482 -721 -4478
rect -704 -4482 -700 -4478
rect -373 -3458 -369 -3454
rect -379 -3466 -375 -3462
rect -551 -3479 -547 -3475
rect -237 -3479 -233 -3475
rect -560 -3518 -556 -3514
rect -568 -3550 -564 -3546
rect -542 -3550 -538 -3546
rect -525 -3550 -521 -3546
rect -485 -3550 -481 -3546
rect -464 -3550 -460 -3546
rect -447 -3550 -443 -3546
rect -407 -3550 -403 -3546
rect -383 -3550 -379 -3546
rect -346 -3550 -342 -3546
rect -577 -3583 -573 -3579
rect -559 -3576 -555 -3572
rect -533 -3598 -529 -3594
rect -551 -3605 -547 -3601
rect -507 -3590 -503 -3586
rect -455 -3583 -451 -3579
rect -525 -3627 -521 -3623
rect -489 -3627 -485 -3623
rect -429 -3598 -425 -3594
rect -447 -3627 -443 -3623
rect -411 -3627 -407 -3623
rect -337 -3589 -333 -3585
rect -331 -3598 -327 -3594
rect -568 -3642 -564 -3638
rect -542 -3642 -538 -3638
rect -499 -3642 -495 -3638
rect -464 -3642 -460 -3638
rect -420 -3642 -416 -3638
rect -403 -3642 -399 -3638
rect -367 -3642 -363 -3638
rect -346 -3642 -342 -3638
rect 98 -2546 102 -2542
rect 90 -2587 94 -2583
rect -21 -2752 -17 -2748
rect -193 -2773 -189 -2769
rect 191 -2773 195 -2769
rect -202 -2812 -198 -2808
rect -210 -2839 -206 -2835
rect -184 -2839 -180 -2835
rect -167 -2839 -163 -2835
rect -127 -2839 -123 -2835
rect -106 -2839 -102 -2835
rect -89 -2839 -85 -2835
rect -49 -2839 -45 -2835
rect -25 -2839 -21 -2835
rect 12 -2839 16 -2835
rect -219 -2872 -215 -2868
rect -201 -2865 -197 -2861
rect -175 -2887 -171 -2883
rect -193 -2894 -189 -2890
rect -149 -2879 -145 -2875
rect -97 -2872 -93 -2868
rect -167 -2916 -163 -2912
rect -131 -2916 -127 -2912
rect -71 -2887 -67 -2883
rect -89 -2916 -85 -2912
rect -53 -2916 -49 -2912
rect 21 -2879 25 -2875
rect 27 -2887 31 -2883
rect -210 -2931 -206 -2927
rect -184 -2931 -180 -2927
rect -141 -2931 -137 -2927
rect -106 -2931 -102 -2927
rect -62 -2931 -58 -2927
rect -45 -2931 -41 -2927
rect -9 -2931 -5 -2927
rect 12 -2931 16 -2927
rect 472 -1792 476 -1788
rect 464 -1835 468 -1831
rect 464 -1858 468 -1854
rect 472 -1907 476 -1903
rect 464 -1950 468 -1946
rect 407 -2002 411 -1998
rect 235 -2023 239 -2019
rect 547 -2023 551 -2019
rect 226 -2062 230 -2058
rect 218 -2089 222 -2085
rect 244 -2089 248 -2085
rect 261 -2089 265 -2085
rect 301 -2089 305 -2085
rect 322 -2089 326 -2085
rect 339 -2089 343 -2085
rect 379 -2089 383 -2085
rect 403 -2089 407 -2085
rect 440 -2089 444 -2085
rect 209 -2122 213 -2118
rect 227 -2115 231 -2111
rect 253 -2137 257 -2133
rect 235 -2144 239 -2140
rect 279 -2129 283 -2125
rect 331 -2122 335 -2118
rect 261 -2166 265 -2162
rect 297 -2166 301 -2162
rect 357 -2137 361 -2133
rect 339 -2166 343 -2162
rect 375 -2166 379 -2162
rect 449 -2129 453 -2125
rect 455 -2137 459 -2133
rect 218 -2181 222 -2177
rect 244 -2181 248 -2177
rect 287 -2181 291 -2177
rect 322 -2181 326 -2177
rect 366 -2181 370 -2177
rect 383 -2181 387 -2177
rect 419 -2181 423 -2177
rect 440 -2181 444 -2177
rect 591 -1317 595 -1313
rect 945 -1317 949 -1313
rect 582 -1356 586 -1352
rect 574 -1378 578 -1374
rect 600 -1378 604 -1374
rect 617 -1378 621 -1374
rect 657 -1378 661 -1374
rect 678 -1378 682 -1374
rect 695 -1378 699 -1374
rect 735 -1378 739 -1374
rect 759 -1378 763 -1374
rect 796 -1378 800 -1374
rect 565 -1411 569 -1407
rect 583 -1404 587 -1400
rect 609 -1426 613 -1422
rect 591 -1433 595 -1429
rect 635 -1418 639 -1414
rect 687 -1411 691 -1407
rect 617 -1455 621 -1451
rect 653 -1455 657 -1451
rect 713 -1426 717 -1422
rect 695 -1455 699 -1451
rect 731 -1455 735 -1451
rect 805 -1418 809 -1414
rect 811 -1426 815 -1422
rect 574 -1470 578 -1466
rect 600 -1470 604 -1466
rect 643 -1470 647 -1466
rect 678 -1470 682 -1466
rect 722 -1470 726 -1466
rect 739 -1470 743 -1466
rect 775 -1470 779 -1466
rect 796 -1470 800 -1466
rect 951 -1418 955 -1414
rect 989 -1082 993 -1078
rect 1321 -1034 1325 -1030
rect 1338 -1034 1342 -1030
rect 980 -1126 984 -1122
rect 972 -1148 976 -1144
rect 989 -1148 993 -1144
rect 1009 -1148 1013 -1144
rect 1030 -1148 1034 -1144
rect 1051 -1148 1055 -1144
rect 1072 -1148 1076 -1144
rect 1093 -1148 1097 -1144
rect 1114 -1148 1118 -1144
rect 1135 -1148 1139 -1144
rect 1155 -1148 1159 -1144
rect 963 -1211 967 -1207
rect 1021 -1204 1025 -1200
rect 1063 -1211 1067 -1207
rect 1081 -1204 1085 -1200
rect 1123 -1196 1127 -1192
rect 1123 -1204 1127 -1200
rect 1105 -1218 1109 -1214
rect 1005 -1225 1009 -1221
rect 1047 -1225 1051 -1221
rect 1147 -1211 1151 -1207
rect 972 -1240 976 -1236
rect 989 -1240 993 -1236
rect 1030 -1240 1034 -1236
rect 1072 -1240 1076 -1236
rect 1114 -1240 1118 -1236
rect 1155 -1240 1159 -1236
rect 963 -1264 967 -1260
rect 980 -1264 984 -1260
rect 945 -1433 949 -1429
rect 811 -1491 815 -1487
rect 951 -1491 955 -1487
rect 574 -1501 578 -1497
rect 591 -1501 595 -1497
rect 611 -1501 615 -1497
rect 632 -1501 636 -1497
rect 653 -1501 657 -1497
rect 674 -1501 678 -1497
rect 695 -1501 699 -1497
rect 716 -1501 720 -1497
rect 737 -1501 741 -1497
rect 757 -1501 761 -1497
rect 565 -1564 569 -1560
rect 623 -1557 627 -1553
rect 665 -1564 669 -1560
rect 683 -1557 687 -1553
rect 725 -1549 729 -1545
rect 725 -1557 729 -1553
rect 707 -1571 711 -1567
rect 607 -1578 611 -1574
rect 649 -1578 653 -1574
rect 749 -1564 753 -1560
rect 574 -1593 578 -1589
rect 591 -1593 595 -1589
rect 632 -1593 636 -1589
rect 674 -1593 678 -1589
rect 716 -1593 720 -1589
rect 757 -1593 761 -1589
rect 574 -1622 578 -1618
rect 591 -1622 595 -1618
rect 611 -1622 615 -1618
rect 632 -1622 636 -1618
rect 653 -1622 657 -1618
rect 674 -1622 678 -1618
rect 695 -1622 699 -1618
rect 716 -1622 720 -1618
rect 737 -1622 741 -1618
rect 757 -1622 761 -1618
rect 565 -1685 569 -1681
rect 623 -1678 627 -1674
rect 665 -1685 669 -1681
rect 683 -1678 687 -1674
rect 725 -1670 729 -1666
rect 725 -1678 729 -1674
rect 707 -1692 711 -1688
rect 607 -1699 611 -1695
rect 649 -1699 653 -1695
rect 763 -1670 767 -1666
rect 749 -1685 753 -1681
rect 574 -1714 578 -1710
rect 591 -1714 595 -1710
rect 632 -1714 636 -1710
rect 674 -1714 678 -1710
rect 716 -1714 720 -1710
rect 757 -1714 761 -1710
rect 951 -1678 955 -1674
rect 763 -1721 767 -1717
rect 951 -1721 955 -1717
rect 574 -1743 578 -1739
rect 591 -1743 595 -1739
rect 611 -1743 615 -1739
rect 632 -1743 636 -1739
rect 653 -1743 657 -1739
rect 674 -1743 678 -1739
rect 695 -1743 699 -1739
rect 716 -1743 720 -1739
rect 737 -1743 741 -1739
rect 757 -1743 761 -1739
rect 559 -1799 563 -1795
rect 565 -1806 569 -1802
rect 623 -1799 627 -1795
rect 665 -1806 669 -1802
rect 683 -1799 687 -1795
rect 725 -1791 729 -1787
rect 725 -1799 729 -1795
rect 707 -1813 711 -1809
rect 607 -1820 611 -1816
rect 649 -1820 653 -1816
rect 763 -1791 767 -1787
rect 749 -1806 753 -1802
rect 574 -1835 578 -1831
rect 591 -1835 595 -1831
rect 632 -1835 636 -1831
rect 674 -1835 678 -1831
rect 716 -1835 720 -1831
rect 757 -1835 761 -1831
rect 565 -1970 569 -1966
rect 582 -1970 586 -1966
rect 553 -2129 557 -2125
rect 547 -2144 551 -2140
rect 455 -2195 459 -2191
rect 553 -2195 557 -2191
rect 218 -2233 222 -2229
rect 235 -2233 239 -2229
rect 255 -2233 259 -2229
rect 276 -2233 280 -2229
rect 297 -2233 301 -2229
rect 318 -2233 322 -2229
rect 339 -2233 343 -2229
rect 360 -2233 364 -2229
rect 381 -2233 385 -2229
rect 401 -2233 405 -2229
rect 209 -2296 213 -2292
rect 267 -2289 271 -2285
rect 309 -2296 313 -2292
rect 327 -2289 331 -2285
rect 369 -2281 373 -2277
rect 369 -2289 373 -2285
rect 351 -2303 355 -2299
rect 251 -2310 255 -2306
rect 293 -2310 297 -2306
rect 393 -2296 397 -2292
rect 218 -2325 222 -2321
rect 235 -2325 239 -2321
rect 276 -2325 280 -2321
rect 318 -2325 322 -2321
rect 360 -2325 364 -2321
rect 401 -2325 405 -2321
rect 218 -2364 222 -2360
rect 235 -2364 239 -2360
rect 255 -2364 259 -2360
rect 276 -2364 280 -2360
rect 297 -2364 301 -2360
rect 318 -2364 322 -2360
rect 339 -2364 343 -2360
rect 360 -2364 364 -2360
rect 381 -2364 385 -2360
rect 401 -2364 405 -2360
rect 209 -2427 213 -2423
rect 267 -2420 271 -2416
rect 309 -2427 313 -2423
rect 327 -2420 331 -2416
rect 369 -2412 373 -2408
rect 369 -2420 373 -2416
rect 351 -2434 355 -2430
rect 251 -2441 255 -2437
rect 293 -2441 297 -2437
rect 407 -2412 411 -2408
rect 393 -2427 397 -2423
rect 218 -2456 222 -2452
rect 235 -2456 239 -2452
rect 276 -2456 280 -2452
rect 318 -2456 322 -2452
rect 360 -2456 364 -2452
rect 401 -2456 405 -2452
rect 553 -2420 557 -2416
rect 407 -2463 411 -2459
rect 553 -2463 557 -2459
rect 218 -2495 222 -2491
rect 235 -2495 239 -2491
rect 255 -2495 259 -2491
rect 276 -2495 280 -2491
rect 297 -2495 301 -2491
rect 318 -2495 322 -2491
rect 339 -2495 343 -2491
rect 360 -2495 364 -2491
rect 381 -2495 385 -2491
rect 401 -2495 405 -2491
rect 203 -2551 207 -2547
rect 209 -2558 213 -2554
rect 267 -2551 271 -2547
rect 309 -2558 313 -2554
rect 327 -2551 331 -2547
rect 369 -2543 373 -2539
rect 369 -2551 373 -2547
rect 351 -2565 355 -2561
rect 251 -2572 255 -2568
rect 293 -2572 297 -2568
rect 407 -2543 411 -2539
rect 393 -2558 397 -2554
rect 218 -2587 222 -2583
rect 235 -2587 239 -2583
rect 276 -2587 280 -2583
rect 318 -2587 322 -2583
rect 360 -2587 364 -2583
rect 401 -2587 405 -2583
rect 209 -2720 213 -2716
rect 226 -2720 230 -2716
rect 197 -2879 201 -2875
rect 191 -2894 195 -2890
rect 27 -2938 31 -2934
rect 197 -2938 201 -2934
rect -210 -2958 -206 -2954
rect -193 -2958 -189 -2954
rect -173 -2958 -169 -2954
rect -152 -2958 -148 -2954
rect -131 -2958 -127 -2954
rect -110 -2958 -106 -2954
rect -89 -2958 -85 -2954
rect -68 -2958 -64 -2954
rect -47 -2958 -43 -2954
rect -27 -2958 -23 -2954
rect -219 -3021 -215 -3017
rect -161 -3014 -157 -3010
rect -119 -3021 -115 -3017
rect -101 -3014 -97 -3010
rect -59 -3006 -55 -3002
rect -59 -3014 -55 -3010
rect -77 -3028 -73 -3024
rect -177 -3035 -173 -3031
rect -135 -3035 -131 -3031
rect -35 -3021 -31 -3017
rect -210 -3050 -206 -3046
rect -193 -3050 -189 -3046
rect -152 -3050 -148 -3046
rect -110 -3050 -106 -3046
rect -68 -3050 -64 -3046
rect -27 -3050 -23 -3046
rect -210 -3074 -206 -3070
rect -193 -3074 -189 -3070
rect -173 -3074 -169 -3070
rect -152 -3074 -148 -3070
rect -131 -3074 -127 -3070
rect -110 -3074 -106 -3070
rect -89 -3074 -85 -3070
rect -68 -3074 -64 -3070
rect -47 -3074 -43 -3070
rect -27 -3074 -23 -3070
rect -219 -3137 -215 -3133
rect -161 -3130 -157 -3126
rect -119 -3137 -115 -3133
rect -101 -3130 -97 -3126
rect -59 -3122 -55 -3118
rect -59 -3130 -55 -3126
rect -77 -3144 -73 -3140
rect -177 -3151 -173 -3147
rect -135 -3151 -131 -3147
rect -21 -3122 -17 -3118
rect -35 -3137 -31 -3133
rect -210 -3166 -206 -3162
rect -193 -3166 -189 -3162
rect -152 -3166 -148 -3162
rect -110 -3166 -106 -3162
rect -68 -3166 -64 -3162
rect -27 -3166 -23 -3162
rect 197 -3130 201 -3126
rect -21 -3174 -17 -3170
rect 197 -3173 201 -3169
rect -210 -3195 -206 -3191
rect -193 -3195 -189 -3191
rect -173 -3195 -169 -3191
rect -152 -3195 -148 -3191
rect -131 -3195 -127 -3191
rect -110 -3195 -106 -3191
rect -89 -3195 -85 -3191
rect -68 -3195 -64 -3191
rect -47 -3195 -43 -3191
rect -27 -3195 -23 -3191
rect -225 -3251 -221 -3247
rect -219 -3258 -215 -3254
rect -161 -3251 -157 -3247
rect -119 -3258 -115 -3254
rect -101 -3251 -97 -3247
rect -59 -3243 -55 -3239
rect -59 -3251 -55 -3247
rect -77 -3265 -73 -3261
rect -177 -3272 -173 -3268
rect -135 -3272 -131 -3268
rect -21 -3243 -17 -3239
rect -35 -3258 -31 -3254
rect -210 -3287 -206 -3283
rect -193 -3287 -189 -3283
rect -152 -3287 -148 -3283
rect -110 -3287 -106 -3283
rect -68 -3287 -64 -3283
rect -27 -3287 -23 -3283
rect -219 -3426 -215 -3422
rect -202 -3426 -198 -3422
rect -231 -3590 -227 -3586
rect -237 -3605 -233 -3601
rect -331 -3656 -327 -3652
rect -231 -3656 -227 -3652
rect -568 -3680 -564 -3676
rect -551 -3680 -547 -3676
rect -531 -3680 -527 -3676
rect -510 -3680 -506 -3676
rect -489 -3680 -485 -3676
rect -468 -3680 -464 -3676
rect -447 -3680 -443 -3676
rect -426 -3680 -422 -3676
rect -405 -3680 -401 -3676
rect -385 -3680 -381 -3676
rect -577 -3743 -573 -3739
rect -519 -3736 -515 -3732
rect -477 -3743 -473 -3739
rect -459 -3736 -455 -3732
rect -417 -3728 -413 -3724
rect -417 -3736 -413 -3732
rect -435 -3750 -431 -3746
rect -535 -3757 -531 -3753
rect -493 -3757 -489 -3753
rect -393 -3743 -389 -3739
rect -568 -3772 -564 -3768
rect -551 -3772 -547 -3768
rect -510 -3772 -506 -3768
rect -468 -3772 -464 -3768
rect -426 -3772 -422 -3768
rect -385 -3772 -381 -3768
rect -568 -3911 -564 -3907
rect -551 -3911 -547 -3907
rect -531 -3911 -527 -3907
rect -510 -3911 -506 -3907
rect -489 -3911 -485 -3907
rect -468 -3911 -464 -3907
rect -447 -3911 -443 -3907
rect -426 -3911 -422 -3907
rect -405 -3911 -401 -3907
rect -385 -3911 -381 -3907
rect -577 -3974 -573 -3970
rect -519 -3967 -515 -3963
rect -477 -3974 -473 -3970
rect -459 -3967 -455 -3963
rect -417 -3959 -413 -3955
rect -417 -3967 -413 -3963
rect -435 -3981 -431 -3977
rect -535 -3988 -531 -3984
rect -493 -3988 -489 -3984
rect -379 -3959 -375 -3955
rect -393 -3974 -389 -3970
rect -568 -4003 -564 -3999
rect -551 -4003 -547 -3999
rect -510 -4003 -506 -3999
rect -468 -4003 -464 -3999
rect -426 -4003 -422 -3999
rect -385 -4003 -381 -3999
rect -231 -3967 -227 -3963
rect -379 -4010 -375 -4006
rect -231 -4010 -227 -4006
rect -568 -4036 -564 -4032
rect -551 -4036 -547 -4032
rect -531 -4036 -527 -4032
rect -510 -4036 -506 -4032
rect -489 -4036 -485 -4032
rect -468 -4036 -464 -4032
rect -447 -4036 -443 -4032
rect -426 -4036 -422 -4032
rect -405 -4036 -401 -4032
rect -385 -4036 -381 -4032
rect -583 -4092 -579 -4088
rect -577 -4099 -573 -4095
rect -519 -4092 -515 -4088
rect -477 -4099 -473 -4095
rect -459 -4092 -455 -4088
rect -417 -4084 -413 -4080
rect -417 -4092 -413 -4088
rect -435 -4106 -431 -4102
rect -535 -4113 -531 -4109
rect -493 -4113 -489 -4109
rect -379 -4084 -375 -4080
rect -393 -4099 -389 -4095
rect -568 -4128 -564 -4124
rect -551 -4128 -547 -4124
rect -510 -4128 -506 -4124
rect -468 -4128 -464 -4124
rect -426 -4128 -422 -4124
rect -385 -4128 -381 -4124
rect -568 -4160 -564 -4156
rect -551 -4160 -547 -4156
rect -531 -4160 -527 -4156
rect -510 -4160 -506 -4156
rect -489 -4160 -485 -4156
rect -468 -4160 -464 -4156
rect -447 -4160 -443 -4156
rect -426 -4160 -422 -4156
rect -405 -4160 -401 -4156
rect -385 -4160 -381 -4156
rect -577 -4223 -573 -4219
rect -519 -4216 -515 -4212
rect -477 -4223 -473 -4219
rect -459 -4216 -455 -4212
rect -417 -4186 -413 -4182
rect -417 -4216 -413 -4212
rect -435 -4230 -431 -4226
rect -535 -4237 -531 -4233
rect -493 -4237 -489 -4233
rect -393 -4223 -389 -4219
rect -568 -4252 -564 -4248
rect -551 -4252 -547 -4248
rect -510 -4252 -506 -4248
rect -468 -4252 -464 -4248
rect -426 -4252 -422 -4248
rect -385 -4252 -381 -4248
rect -577 -4271 -573 -4267
rect -560 -4271 -556 -4267
rect -589 -4430 -585 -4426
rect -595 -4445 -591 -4441
rect -689 -4489 -685 -4485
rect -589 -4489 -585 -4485
rect -926 -4513 -922 -4509
rect -909 -4513 -905 -4509
rect -889 -4513 -885 -4509
rect -868 -4513 -864 -4509
rect -847 -4513 -843 -4509
rect -826 -4513 -822 -4509
rect -805 -4513 -801 -4509
rect -784 -4513 -780 -4509
rect -763 -4513 -759 -4509
rect -743 -4513 -739 -4509
rect -935 -4576 -931 -4572
rect -877 -4569 -873 -4565
rect -835 -4576 -831 -4572
rect -817 -4569 -813 -4565
rect -775 -4561 -771 -4557
rect -775 -4569 -771 -4565
rect -793 -4583 -789 -4579
rect -893 -4590 -889 -4586
rect -851 -4590 -847 -4586
rect -751 -4576 -747 -4572
rect -926 -4605 -922 -4601
rect -909 -4605 -905 -4601
rect -868 -4605 -864 -4601
rect -826 -4605 -822 -4601
rect -784 -4605 -780 -4601
rect -743 -4605 -739 -4601
rect -926 -4634 -922 -4630
rect -909 -4634 -905 -4630
rect -889 -4634 -885 -4630
rect -868 -4634 -864 -4630
rect -847 -4634 -843 -4630
rect -826 -4634 -822 -4630
rect -805 -4634 -801 -4630
rect -784 -4634 -780 -4630
rect -763 -4634 -759 -4630
rect -743 -4634 -739 -4630
rect -935 -4697 -931 -4693
rect -877 -4690 -873 -4686
rect -835 -4697 -831 -4693
rect -817 -4690 -813 -4686
rect -775 -4682 -771 -4678
rect -775 -4690 -771 -4686
rect -793 -4704 -789 -4700
rect -893 -4711 -889 -4707
rect -851 -4711 -847 -4707
rect -737 -4682 -733 -4678
rect -751 -4697 -747 -4693
rect -926 -4726 -922 -4722
rect -909 -4726 -905 -4722
rect -868 -4726 -864 -4722
rect -826 -4726 -822 -4722
rect -784 -4726 -780 -4722
rect -743 -4726 -739 -4722
rect -589 -4690 -585 -4686
rect -737 -4733 -733 -4729
rect -589 -4733 -585 -4729
rect -926 -4755 -922 -4751
rect -909 -4755 -905 -4751
rect -889 -4755 -885 -4751
rect -868 -4755 -864 -4751
rect -847 -4755 -843 -4751
rect -826 -4755 -822 -4751
rect -805 -4755 -801 -4751
rect -784 -4755 -780 -4751
rect -763 -4755 -759 -4751
rect -743 -4755 -739 -4751
rect -941 -4811 -937 -4807
rect -935 -4818 -931 -4814
rect -877 -4811 -873 -4807
rect -835 -4818 -831 -4814
rect -817 -4811 -813 -4807
rect -775 -4803 -771 -4799
rect -775 -4811 -771 -4807
rect -793 -4825 -789 -4821
rect -893 -4832 -889 -4828
rect -851 -4832 -847 -4828
rect -737 -4803 -733 -4799
rect -751 -4818 -747 -4814
rect -926 -4847 -922 -4843
rect -909 -4847 -905 -4843
rect -868 -4847 -864 -4843
rect -826 -4847 -822 -4843
rect -784 -4847 -780 -4843
rect -743 -4847 -739 -4843
rect -926 -4873 -922 -4869
rect -909 -4873 -905 -4869
rect -889 -4873 -885 -4869
rect -868 -4873 -864 -4869
rect -847 -4873 -843 -4869
rect -826 -4873 -822 -4869
rect -805 -4873 -801 -4869
rect -784 -4873 -780 -4869
rect -763 -4873 -759 -4869
rect -743 -4873 -739 -4869
rect -935 -4936 -931 -4932
rect -877 -4929 -873 -4925
rect -835 -4936 -831 -4932
rect -817 -4929 -813 -4925
rect -775 -4921 -771 -4917
rect -775 -4929 -771 -4925
rect -793 -4943 -789 -4939
rect -893 -4950 -889 -4946
rect -851 -4950 -847 -4946
rect -751 -4936 -747 -4932
rect -926 -4965 -922 -4961
rect -909 -4965 -905 -4961
rect -868 -4965 -864 -4961
rect -826 -4965 -822 -4961
rect -784 -4965 -780 -4961
rect -743 -4965 -739 -4961
rect -935 -4990 -931 -4986
rect -918 -4990 -914 -4986
rect -947 -5164 -943 -5160
rect -1162 -5179 -1158 -5175
rect -1255 -5201 -1251 -5197
rect -1211 -5201 -1207 -5197
rect -1177 -5201 -1173 -5197
rect -1276 -5208 -1272 -5204
rect -1270 -5216 -1266 -5212
rect -1162 -5216 -1158 -5212
rect -947 -5215 -943 -5211
rect -1255 -5228 -1251 -5224
rect -1238 -5228 -1234 -5224
rect -1218 -5228 -1214 -5224
rect -1197 -5228 -1193 -5224
rect -1176 -5228 -1172 -5224
rect -1155 -5228 -1151 -5224
rect -1134 -5228 -1130 -5224
rect -1113 -5228 -1109 -5224
rect -1092 -5228 -1088 -5224
rect -1072 -5228 -1068 -5224
rect -1270 -5284 -1266 -5280
rect -1264 -5291 -1260 -5287
rect -1206 -5284 -1202 -5280
rect -1164 -5291 -1160 -5287
rect -1146 -5284 -1142 -5280
rect -1104 -5276 -1100 -5272
rect -1104 -5284 -1100 -5280
rect -1122 -5298 -1118 -5294
rect -1222 -5305 -1218 -5301
rect -1180 -5305 -1176 -5301
rect -1080 -5291 -1076 -5287
rect -1255 -5320 -1251 -5316
rect -1238 -5320 -1234 -5316
rect -1197 -5320 -1193 -5316
rect -1155 -5320 -1151 -5316
rect -1113 -5320 -1109 -5316
rect -1072 -5320 -1068 -5316
rect -1255 -5349 -1251 -5345
rect -1238 -5349 -1234 -5345
rect -1218 -5349 -1214 -5345
rect -1197 -5349 -1193 -5345
rect -1176 -5349 -1172 -5345
rect -1155 -5349 -1151 -5345
rect -1134 -5349 -1130 -5345
rect -1113 -5349 -1109 -5345
rect -1092 -5349 -1088 -5345
rect -1072 -5349 -1068 -5345
rect -1276 -5405 -1272 -5401
rect -1026 -5349 -1022 -5345
rect -1264 -5412 -1260 -5408
rect -1206 -5405 -1202 -5401
rect -1164 -5412 -1160 -5408
rect -1146 -5405 -1142 -5401
rect -1104 -5397 -1100 -5393
rect -1104 -5405 -1100 -5401
rect -1122 -5419 -1118 -5415
rect -1222 -5426 -1218 -5422
rect -1180 -5426 -1176 -5422
rect -1066 -5397 -1062 -5393
rect -1018 -5394 -1014 -5390
rect -1080 -5412 -1076 -5408
rect -1255 -5441 -1251 -5437
rect -1238 -5441 -1234 -5437
rect -1197 -5441 -1193 -5437
rect -1155 -5441 -1151 -5437
rect -1113 -5441 -1109 -5437
rect -1072 -5441 -1068 -5437
rect -947 -5405 -943 -5401
rect -1026 -5441 -1022 -5437
rect -1349 -5525 -1345 -5521
rect -1270 -5448 -1266 -5444
rect -1066 -5448 -1062 -5444
rect -947 -5448 -943 -5444
rect -1339 -5703 -1335 -5699
rect -1322 -5703 -1318 -5699
rect -1322 -5795 -1318 -5791
rect -1255 -5469 -1251 -5465
rect -1238 -5469 -1234 -5465
rect -1218 -5469 -1214 -5465
rect -1197 -5469 -1193 -5465
rect -1176 -5469 -1172 -5465
rect -1155 -5469 -1151 -5465
rect -1134 -5469 -1130 -5465
rect -1113 -5469 -1109 -5465
rect -1092 -5469 -1088 -5465
rect -1072 -5469 -1068 -5465
rect -1026 -5469 -1022 -5465
rect -1264 -5532 -1260 -5528
rect -1206 -5525 -1202 -5521
rect -1164 -5532 -1160 -5528
rect -1146 -5525 -1142 -5521
rect -1104 -5517 -1100 -5513
rect -1104 -5525 -1100 -5521
rect -1122 -5539 -1118 -5535
rect -1222 -5546 -1218 -5542
rect -1180 -5546 -1176 -5542
rect -1066 -5517 -1062 -5513
rect -1080 -5532 -1076 -5528
rect -1255 -5561 -1251 -5557
rect -1238 -5561 -1234 -5557
rect -1197 -5561 -1193 -5557
rect -1155 -5561 -1151 -5557
rect -1113 -5561 -1109 -5557
rect -1072 -5561 -1068 -5557
rect -1255 -5586 -1251 -5582
rect -1238 -5586 -1234 -5582
rect -1218 -5586 -1214 -5582
rect -1197 -5586 -1193 -5582
rect -1176 -5586 -1172 -5582
rect -1155 -5586 -1151 -5582
rect -1134 -5586 -1130 -5582
rect -1113 -5586 -1109 -5582
rect -1092 -5586 -1088 -5582
rect -1072 -5586 -1068 -5582
rect -1264 -5649 -1260 -5645
rect -1206 -5642 -1202 -5638
rect -1164 -5649 -1160 -5645
rect -1146 -5642 -1142 -5638
rect -1104 -5634 -1100 -5630
rect -1104 -5642 -1100 -5638
rect -1122 -5656 -1118 -5652
rect -1222 -5663 -1218 -5659
rect -1180 -5663 -1176 -5659
rect -1080 -5649 -1076 -5645
rect -1255 -5678 -1251 -5674
rect -1238 -5678 -1234 -5674
rect -1197 -5678 -1193 -5674
rect -1155 -5678 -1151 -5674
rect -1113 -5678 -1109 -5674
rect -1072 -5678 -1068 -5674
rect -1018 -5518 -1014 -5514
rect -1026 -5561 -1022 -5557
rect -1066 -5735 -1062 -5731
rect -953 -5756 -949 -5752
rect -1255 -5822 -1251 -5818
rect -1238 -5822 -1234 -5818
rect -1198 -5822 -1194 -5818
rect -1177 -5822 -1173 -5818
rect -1270 -5878 -1266 -5874
rect -1264 -5871 -1260 -5867
rect -1313 -5885 -1309 -5881
rect -1220 -5892 -1216 -5888
rect -953 -5862 -949 -5858
rect -1168 -5870 -1164 -5866
rect -1238 -5899 -1234 -5895
rect -1202 -5899 -1198 -5895
rect -737 -5022 -733 -5018
rect -909 -5043 -905 -5039
rect -595 -5043 -591 -5039
rect -918 -5082 -914 -5078
rect -926 -5109 -922 -5105
rect -900 -5109 -896 -5105
rect -883 -5109 -879 -5105
rect -843 -5109 -839 -5105
rect -822 -5109 -818 -5105
rect -805 -5109 -801 -5105
rect -765 -5109 -761 -5105
rect -741 -5109 -737 -5105
rect -704 -5109 -700 -5105
rect -935 -5142 -931 -5138
rect -917 -5135 -913 -5131
rect -891 -5157 -887 -5153
rect -909 -5164 -905 -5160
rect -865 -5149 -861 -5145
rect -813 -5142 -809 -5138
rect -883 -5186 -879 -5182
rect -847 -5186 -843 -5182
rect -787 -5157 -783 -5153
rect -805 -5186 -801 -5182
rect -769 -5186 -765 -5182
rect -695 -5149 -691 -5145
rect -689 -5157 -685 -5153
rect -926 -5201 -922 -5197
rect -900 -5201 -896 -5197
rect -857 -5201 -853 -5197
rect -822 -5201 -818 -5197
rect -778 -5201 -774 -5197
rect -761 -5201 -757 -5197
rect -725 -5201 -721 -5197
rect -704 -5201 -700 -5197
rect -332 -4160 -328 -4156
rect -324 -4207 -320 -4203
rect -332 -4252 -328 -4248
rect -332 -4271 -328 -4267
rect -379 -4303 -375 -4299
rect -551 -4324 -547 -4320
rect -324 -4322 -320 -4318
rect -237 -4324 -233 -4320
rect -560 -4363 -556 -4359
rect -332 -4363 -328 -4359
rect -568 -4390 -564 -4386
rect -542 -4390 -538 -4386
rect -525 -4390 -521 -4386
rect -485 -4390 -481 -4386
rect -464 -4390 -460 -4386
rect -447 -4390 -443 -4386
rect -407 -4390 -403 -4386
rect -383 -4390 -379 -4386
rect -346 -4390 -342 -4386
rect -577 -4423 -573 -4419
rect -559 -4416 -555 -4412
rect -533 -4438 -529 -4434
rect -551 -4445 -547 -4441
rect -507 -4430 -503 -4426
rect -455 -4423 -451 -4419
rect -525 -4467 -521 -4463
rect -489 -4467 -485 -4463
rect -429 -4438 -425 -4434
rect -447 -4467 -443 -4463
rect -411 -4467 -407 -4463
rect -337 -4429 -333 -4425
rect -331 -4438 -327 -4434
rect -568 -4482 -564 -4478
rect -542 -4482 -538 -4478
rect -499 -4482 -495 -4478
rect -464 -4482 -460 -4478
rect -420 -4482 -416 -4478
rect -403 -4482 -399 -4478
rect -367 -4482 -363 -4478
rect -346 -4482 -342 -4478
rect -21 -3458 -17 -3454
rect -193 -3479 -189 -3475
rect 191 -3479 195 -3475
rect -202 -3518 -198 -3514
rect -210 -3550 -206 -3546
rect -184 -3550 -180 -3546
rect -167 -3550 -163 -3546
rect -127 -3550 -123 -3546
rect -106 -3550 -102 -3546
rect -89 -3550 -85 -3546
rect -49 -3550 -45 -3546
rect -25 -3550 -21 -3546
rect 12 -3550 16 -3546
rect -219 -3583 -215 -3579
rect -201 -3576 -197 -3572
rect -175 -3598 -171 -3594
rect -193 -3605 -189 -3601
rect -149 -3590 -145 -3586
rect -97 -3583 -93 -3579
rect -167 -3627 -163 -3623
rect -131 -3627 -127 -3623
rect -71 -3598 -67 -3594
rect -89 -3627 -85 -3623
rect -53 -3627 -49 -3623
rect 21 -3590 25 -3586
rect 27 -3598 31 -3594
rect -210 -3642 -206 -3638
rect -184 -3642 -180 -3638
rect -141 -3642 -137 -3638
rect -106 -3642 -102 -3638
rect -62 -3642 -58 -3638
rect -45 -3642 -41 -3638
rect -9 -3642 -5 -3638
rect 12 -3642 16 -3638
rect 407 -2752 411 -2748
rect 235 -2773 239 -2769
rect 547 -2773 551 -2769
rect 226 -2812 230 -2808
rect 218 -2839 222 -2835
rect 244 -2839 248 -2835
rect 261 -2839 265 -2835
rect 301 -2839 305 -2835
rect 322 -2839 326 -2835
rect 339 -2839 343 -2835
rect 379 -2839 383 -2835
rect 403 -2839 407 -2835
rect 440 -2839 444 -2835
rect 209 -2872 213 -2868
rect 227 -2865 231 -2861
rect 253 -2887 257 -2883
rect 235 -2894 239 -2890
rect 279 -2879 283 -2875
rect 331 -2872 335 -2868
rect 261 -2916 265 -2912
rect 297 -2916 301 -2912
rect 357 -2887 361 -2883
rect 339 -2916 343 -2912
rect 375 -2916 379 -2912
rect 449 -2879 453 -2875
rect 455 -2887 459 -2883
rect 218 -2931 222 -2927
rect 244 -2931 248 -2927
rect 287 -2931 291 -2927
rect 322 -2931 326 -2927
rect 366 -2931 370 -2927
rect 383 -2931 387 -2927
rect 419 -2931 423 -2927
rect 440 -2931 444 -2927
rect 841 -1858 845 -1854
rect 849 -1907 853 -1903
rect 841 -1950 845 -1946
rect 763 -2002 767 -1998
rect 591 -2023 595 -2019
rect 945 -2023 949 -2019
rect 582 -2062 586 -2058
rect 574 -2089 578 -2085
rect 600 -2089 604 -2085
rect 617 -2089 621 -2085
rect 657 -2089 661 -2085
rect 678 -2089 682 -2085
rect 695 -2089 699 -2085
rect 735 -2089 739 -2085
rect 759 -2089 763 -2085
rect 796 -2089 800 -2085
rect 565 -2122 569 -2118
rect 583 -2115 587 -2111
rect 609 -2137 613 -2133
rect 591 -2144 595 -2140
rect 635 -2129 639 -2125
rect 687 -2122 691 -2118
rect 617 -2166 621 -2162
rect 653 -2166 657 -2162
rect 713 -2137 717 -2133
rect 695 -2166 699 -2162
rect 731 -2166 735 -2162
rect 805 -2129 809 -2125
rect 811 -2137 815 -2133
rect 574 -2181 578 -2177
rect 600 -2181 604 -2177
rect 643 -2181 647 -2177
rect 678 -2181 682 -2177
rect 722 -2181 726 -2177
rect 739 -2181 743 -2177
rect 775 -2181 779 -2177
rect 796 -2181 800 -2177
rect 1347 -1090 1351 -1086
rect 1338 -1126 1342 -1122
rect 1321 -1264 1325 -1260
rect 1338 -1264 1342 -1260
rect 989 -1317 993 -1313
rect 1309 -1317 1313 -1313
rect 980 -1356 984 -1352
rect 972 -1378 976 -1374
rect 998 -1378 1002 -1374
rect 1015 -1378 1019 -1374
rect 1055 -1378 1059 -1374
rect 1076 -1378 1080 -1374
rect 1093 -1378 1097 -1374
rect 1133 -1378 1137 -1374
rect 1157 -1378 1161 -1374
rect 1194 -1378 1198 -1374
rect 963 -1411 967 -1407
rect 981 -1404 985 -1400
rect 1007 -1426 1011 -1422
rect 989 -1433 993 -1429
rect 1033 -1418 1037 -1414
rect 1085 -1411 1089 -1407
rect 1015 -1455 1019 -1451
rect 1051 -1455 1055 -1451
rect 1111 -1426 1115 -1422
rect 1093 -1455 1097 -1451
rect 1129 -1455 1133 -1451
rect 1203 -1434 1207 -1430
rect 1209 -1426 1213 -1422
rect 972 -1470 976 -1466
rect 998 -1470 1002 -1466
rect 1041 -1470 1045 -1466
rect 1076 -1470 1080 -1466
rect 1120 -1470 1124 -1466
rect 1137 -1470 1141 -1466
rect 1173 -1470 1177 -1466
rect 1194 -1470 1198 -1466
rect 1309 -1441 1313 -1437
rect 1209 -1484 1213 -1480
rect 1309 -1484 1313 -1480
rect 972 -1501 976 -1497
rect 989 -1501 993 -1497
rect 1009 -1501 1013 -1497
rect 1030 -1501 1034 -1497
rect 1051 -1501 1055 -1497
rect 1072 -1501 1076 -1497
rect 1093 -1501 1097 -1497
rect 1114 -1501 1118 -1497
rect 1135 -1501 1139 -1497
rect 1155 -1501 1159 -1497
rect 963 -1564 967 -1560
rect 1021 -1557 1025 -1553
rect 1063 -1564 1067 -1560
rect 1081 -1557 1085 -1553
rect 1123 -1549 1127 -1545
rect 1123 -1557 1127 -1553
rect 1105 -1571 1109 -1567
rect 1005 -1578 1009 -1574
rect 1047 -1578 1051 -1574
rect 1147 -1564 1151 -1560
rect 972 -1593 976 -1589
rect 989 -1593 993 -1589
rect 1030 -1593 1034 -1589
rect 1072 -1593 1076 -1589
rect 1114 -1593 1118 -1589
rect 1155 -1593 1159 -1589
rect 972 -1622 976 -1618
rect 989 -1622 993 -1618
rect 1009 -1622 1013 -1618
rect 1030 -1622 1034 -1618
rect 1051 -1622 1055 -1618
rect 1072 -1622 1076 -1618
rect 1093 -1622 1097 -1618
rect 1114 -1622 1118 -1618
rect 1135 -1622 1139 -1618
rect 1155 -1622 1159 -1618
rect 963 -1685 967 -1681
rect 1021 -1678 1025 -1674
rect 1063 -1685 1067 -1681
rect 1081 -1678 1085 -1674
rect 1123 -1670 1127 -1666
rect 1123 -1678 1127 -1674
rect 1105 -1692 1109 -1688
rect 1005 -1699 1009 -1695
rect 1047 -1699 1051 -1695
rect 1161 -1670 1165 -1666
rect 1147 -1685 1151 -1681
rect 972 -1714 976 -1710
rect 989 -1714 993 -1710
rect 1030 -1714 1034 -1710
rect 1072 -1714 1076 -1710
rect 1114 -1714 1118 -1710
rect 1155 -1714 1159 -1710
rect 1309 -1678 1313 -1674
rect 1161 -1721 1165 -1717
rect 1309 -1722 1313 -1718
rect 972 -1743 976 -1739
rect 989 -1743 993 -1739
rect 1009 -1743 1013 -1739
rect 1030 -1743 1034 -1739
rect 1051 -1743 1055 -1739
rect 1072 -1743 1076 -1739
rect 1093 -1743 1097 -1739
rect 1114 -1743 1118 -1739
rect 1135 -1743 1139 -1739
rect 1155 -1743 1159 -1739
rect 957 -1799 961 -1795
rect 1203 -1743 1207 -1739
rect 963 -1806 967 -1802
rect 1021 -1799 1025 -1795
rect 1063 -1806 1067 -1802
rect 1081 -1799 1085 -1795
rect 1123 -1791 1127 -1787
rect 1123 -1799 1127 -1795
rect 1105 -1813 1109 -1809
rect 1005 -1820 1009 -1816
rect 1047 -1820 1051 -1816
rect 1161 -1791 1165 -1787
rect 1147 -1806 1151 -1802
rect 972 -1835 976 -1831
rect 989 -1835 993 -1831
rect 1030 -1835 1034 -1831
rect 1072 -1835 1076 -1831
rect 1114 -1835 1118 -1831
rect 1155 -1835 1159 -1831
rect 963 -1970 967 -1966
rect 980 -1970 984 -1966
rect 951 -2129 955 -2125
rect 945 -2144 949 -2140
rect 811 -2188 815 -2184
rect 951 -2188 955 -2184
rect 574 -2233 578 -2229
rect 591 -2233 595 -2229
rect 611 -2233 615 -2229
rect 632 -2233 636 -2229
rect 653 -2233 657 -2229
rect 674 -2233 678 -2229
rect 695 -2233 699 -2229
rect 716 -2233 720 -2229
rect 737 -2233 741 -2229
rect 757 -2233 761 -2229
rect 565 -2296 569 -2292
rect 623 -2289 627 -2285
rect 665 -2296 669 -2292
rect 683 -2289 687 -2285
rect 725 -2281 729 -2277
rect 725 -2289 729 -2285
rect 707 -2303 711 -2299
rect 607 -2310 611 -2306
rect 649 -2310 653 -2306
rect 749 -2296 753 -2292
rect 574 -2325 578 -2321
rect 591 -2325 595 -2321
rect 632 -2325 636 -2321
rect 674 -2325 678 -2321
rect 716 -2325 720 -2321
rect 757 -2325 761 -2321
rect 574 -2364 578 -2360
rect 591 -2364 595 -2360
rect 611 -2364 615 -2360
rect 632 -2364 636 -2360
rect 653 -2364 657 -2360
rect 674 -2364 678 -2360
rect 695 -2364 699 -2360
rect 716 -2364 720 -2360
rect 737 -2364 741 -2360
rect 757 -2364 761 -2360
rect 565 -2427 569 -2423
rect 623 -2420 627 -2416
rect 665 -2427 669 -2423
rect 683 -2420 687 -2416
rect 725 -2412 729 -2408
rect 725 -2420 729 -2416
rect 707 -2434 711 -2430
rect 607 -2441 611 -2437
rect 649 -2441 653 -2437
rect 763 -2412 767 -2408
rect 749 -2427 753 -2423
rect 574 -2456 578 -2452
rect 591 -2456 595 -2452
rect 632 -2456 636 -2452
rect 674 -2456 678 -2452
rect 716 -2456 720 -2452
rect 757 -2456 761 -2452
rect 951 -2420 955 -2416
rect 763 -2463 767 -2459
rect 951 -2464 955 -2460
rect 574 -2495 578 -2491
rect 591 -2495 595 -2491
rect 611 -2495 615 -2491
rect 632 -2495 636 -2491
rect 653 -2495 657 -2491
rect 674 -2495 678 -2491
rect 695 -2495 699 -2491
rect 716 -2495 720 -2491
rect 737 -2495 741 -2491
rect 757 -2495 761 -2491
rect 559 -2551 563 -2547
rect 565 -2558 569 -2554
rect 623 -2551 627 -2547
rect 665 -2558 669 -2554
rect 683 -2551 687 -2547
rect 725 -2543 729 -2539
rect 725 -2551 729 -2547
rect 707 -2565 711 -2561
rect 607 -2572 611 -2568
rect 649 -2572 653 -2568
rect 763 -2543 767 -2539
rect 749 -2558 753 -2554
rect 574 -2587 578 -2583
rect 591 -2587 595 -2583
rect 632 -2587 636 -2583
rect 674 -2587 678 -2583
rect 716 -2587 720 -2583
rect 757 -2587 761 -2583
rect 565 -2720 569 -2716
rect 582 -2720 586 -2716
rect 553 -2879 557 -2875
rect 547 -2894 551 -2890
rect 455 -2945 459 -2941
rect 553 -2945 557 -2941
rect 218 -2958 222 -2954
rect 235 -2958 239 -2954
rect 255 -2958 259 -2954
rect 276 -2958 280 -2954
rect 297 -2958 301 -2954
rect 318 -2958 322 -2954
rect 339 -2958 343 -2954
rect 360 -2958 364 -2954
rect 381 -2958 385 -2954
rect 401 -2958 405 -2954
rect 472 -2958 476 -2954
rect 209 -3021 213 -3017
rect 267 -3014 271 -3010
rect 309 -3021 313 -3017
rect 327 -3014 331 -3010
rect 369 -3006 373 -3002
rect 369 -3014 373 -3010
rect 351 -3028 355 -3024
rect 251 -3035 255 -3031
rect 293 -3035 297 -3031
rect 480 -3007 484 -3003
rect 393 -3021 397 -3017
rect 218 -3050 222 -3046
rect 235 -3050 239 -3046
rect 276 -3050 280 -3046
rect 318 -3050 322 -3046
rect 360 -3050 364 -3046
rect 401 -3050 405 -3046
rect 472 -3050 476 -3046
rect 218 -3074 222 -3070
rect 235 -3074 239 -3070
rect 255 -3074 259 -3070
rect 276 -3074 280 -3070
rect 297 -3074 301 -3070
rect 318 -3074 322 -3070
rect 339 -3074 343 -3070
rect 360 -3074 364 -3070
rect 381 -3074 385 -3070
rect 401 -3074 405 -3070
rect 472 -3074 476 -3070
rect 209 -3137 213 -3133
rect 267 -3130 271 -3126
rect 309 -3137 313 -3133
rect 327 -3130 331 -3126
rect 369 -3122 373 -3118
rect 369 -3130 373 -3126
rect 351 -3144 355 -3140
rect 251 -3151 255 -3147
rect 293 -3151 297 -3147
rect 407 -3122 411 -3118
rect 393 -3137 397 -3133
rect 218 -3166 222 -3162
rect 235 -3166 239 -3162
rect 276 -3166 280 -3162
rect 318 -3166 322 -3162
rect 360 -3166 364 -3162
rect 401 -3166 405 -3162
rect 480 -3123 484 -3119
rect 553 -3130 557 -3126
rect 472 -3166 476 -3162
rect 407 -3173 411 -3169
rect 553 -3173 557 -3169
rect 218 -3195 222 -3191
rect 235 -3195 239 -3191
rect 255 -3195 259 -3191
rect 276 -3195 280 -3191
rect 297 -3195 301 -3191
rect 318 -3195 322 -3191
rect 339 -3195 343 -3191
rect 360 -3195 364 -3191
rect 381 -3195 385 -3191
rect 401 -3195 405 -3191
rect 203 -3251 207 -3247
rect 209 -3258 213 -3254
rect 267 -3251 271 -3247
rect 309 -3258 313 -3254
rect 327 -3251 331 -3247
rect 369 -3243 373 -3239
rect 369 -3251 373 -3247
rect 351 -3265 355 -3261
rect 251 -3272 255 -3268
rect 293 -3272 297 -3268
rect 407 -3243 411 -3239
rect 393 -3258 397 -3254
rect 218 -3287 222 -3283
rect 235 -3287 239 -3283
rect 276 -3287 280 -3283
rect 318 -3287 322 -3283
rect 360 -3287 364 -3283
rect 401 -3287 405 -3283
rect 209 -3426 213 -3422
rect 226 -3426 230 -3422
rect 197 -3590 201 -3586
rect 191 -3605 195 -3601
rect 27 -3649 31 -3645
rect 197 -3649 201 -3645
rect -210 -3680 -206 -3676
rect -193 -3680 -189 -3676
rect -173 -3680 -169 -3676
rect -152 -3680 -148 -3676
rect -131 -3680 -127 -3676
rect -110 -3680 -106 -3676
rect -89 -3680 -85 -3676
rect -68 -3680 -64 -3676
rect -47 -3680 -43 -3676
rect -27 -3680 -23 -3676
rect -219 -3743 -215 -3739
rect -161 -3736 -157 -3732
rect -119 -3743 -115 -3739
rect -101 -3736 -97 -3732
rect -59 -3728 -55 -3724
rect -59 -3736 -55 -3732
rect -77 -3750 -73 -3746
rect -177 -3757 -173 -3753
rect -135 -3757 -131 -3753
rect -35 -3743 -31 -3739
rect -210 -3772 -206 -3768
rect -193 -3772 -189 -3768
rect -152 -3772 -148 -3768
rect -110 -3772 -106 -3768
rect -68 -3772 -64 -3768
rect -27 -3772 -23 -3768
rect 68 -3795 72 -3791
rect 76 -3846 80 -3842
rect 68 -3887 72 -3883
rect -210 -3911 -206 -3907
rect -193 -3911 -189 -3907
rect -173 -3911 -169 -3907
rect -152 -3911 -148 -3907
rect -131 -3911 -127 -3907
rect -110 -3911 -106 -3907
rect -89 -3911 -85 -3907
rect -68 -3911 -64 -3907
rect -47 -3911 -43 -3907
rect -27 -3911 -23 -3907
rect -219 -3974 -215 -3970
rect -161 -3967 -157 -3963
rect -119 -3974 -115 -3970
rect -101 -3967 -97 -3963
rect -59 -3959 -55 -3955
rect -59 -3967 -55 -3963
rect -77 -3981 -73 -3977
rect -177 -3988 -173 -3984
rect -135 -3988 -131 -3984
rect -21 -3959 -17 -3955
rect -35 -3974 -31 -3970
rect -210 -4003 -206 -3999
rect -193 -4003 -189 -3999
rect -152 -4003 -148 -3999
rect -110 -4003 -106 -3999
rect -68 -4003 -64 -3999
rect -27 -4003 -23 -3999
rect 197 -3967 201 -3963
rect -21 -4010 -17 -4006
rect 197 -4010 201 -4006
rect -210 -4036 -206 -4032
rect -193 -4036 -189 -4032
rect -173 -4036 -169 -4032
rect -152 -4036 -148 -4032
rect -131 -4036 -127 -4032
rect -110 -4036 -106 -4032
rect -89 -4036 -85 -4032
rect -68 -4036 -64 -4032
rect -47 -4036 -43 -4032
rect -27 -4036 -23 -4032
rect -225 -4092 -221 -4088
rect -219 -4099 -215 -4095
rect -161 -4092 -157 -4088
rect -119 -4099 -115 -4095
rect -101 -4092 -97 -4088
rect -59 -4084 -55 -4080
rect -59 -4092 -55 -4088
rect -77 -4106 -73 -4102
rect -177 -4113 -173 -4109
rect -135 -4113 -131 -4109
rect -15 -4084 -11 -4080
rect -35 -4099 -31 -4095
rect -210 -4128 -206 -4124
rect -193 -4128 -189 -4124
rect -152 -4128 -148 -4124
rect -110 -4128 -106 -4124
rect -68 -4128 -64 -4124
rect -27 -4128 -23 -4124
rect -210 -4160 -206 -4156
rect -193 -4160 -189 -4156
rect -173 -4160 -169 -4156
rect -152 -4160 -148 -4156
rect -131 -4160 -127 -4156
rect -110 -4160 -106 -4156
rect -89 -4160 -85 -4156
rect -68 -4160 -64 -4156
rect -47 -4160 -43 -4156
rect -27 -4160 -23 -4156
rect -219 -4223 -215 -4219
rect -161 -4216 -157 -4212
rect -119 -4223 -115 -4219
rect -101 -4216 -97 -4212
rect -59 -4208 -55 -4204
rect -59 -4216 -55 -4212
rect -77 -4230 -73 -4226
rect -177 -4237 -173 -4233
rect -135 -4237 -131 -4233
rect -21 -4208 -17 -4204
rect -35 -4223 -31 -4219
rect -210 -4252 -206 -4248
rect -193 -4252 -189 -4248
rect -152 -4252 -148 -4248
rect -110 -4252 -106 -4248
rect -68 -4252 -64 -4248
rect -27 -4252 -23 -4248
rect -219 -4271 -215 -4267
rect -202 -4271 -198 -4267
rect -231 -4430 -227 -4426
rect -237 -4445 -233 -4441
rect -331 -4496 -327 -4492
rect -231 -4496 -227 -4492
rect -568 -4513 -564 -4509
rect -551 -4513 -547 -4509
rect -531 -4513 -527 -4509
rect -510 -4513 -506 -4509
rect -489 -4513 -485 -4509
rect -468 -4513 -464 -4509
rect -447 -4513 -443 -4509
rect -426 -4513 -422 -4509
rect -405 -4513 -401 -4509
rect -385 -4513 -381 -4509
rect -577 -4576 -573 -4572
rect -519 -4569 -515 -4565
rect -477 -4576 -473 -4572
rect -459 -4569 -455 -4565
rect -417 -4561 -413 -4557
rect -417 -4569 -413 -4565
rect -435 -4583 -431 -4579
rect -535 -4590 -531 -4586
rect -493 -4590 -489 -4586
rect -393 -4576 -389 -4572
rect -568 -4605 -564 -4601
rect -551 -4605 -547 -4601
rect -510 -4605 -506 -4601
rect -468 -4605 -464 -4601
rect -426 -4605 -422 -4601
rect -385 -4605 -381 -4601
rect -568 -4634 -564 -4630
rect -551 -4634 -547 -4630
rect -531 -4634 -527 -4630
rect -510 -4634 -506 -4630
rect -489 -4634 -485 -4630
rect -468 -4634 -464 -4630
rect -447 -4634 -443 -4630
rect -426 -4634 -422 -4630
rect -405 -4634 -401 -4630
rect -385 -4634 -381 -4630
rect -577 -4697 -573 -4693
rect -519 -4690 -515 -4686
rect -477 -4697 -473 -4693
rect -459 -4690 -455 -4686
rect -417 -4682 -413 -4678
rect -417 -4690 -413 -4686
rect -435 -4704 -431 -4700
rect -535 -4711 -531 -4707
rect -493 -4711 -489 -4707
rect -379 -4682 -375 -4678
rect -393 -4697 -389 -4693
rect -568 -4726 -564 -4722
rect -551 -4726 -547 -4722
rect -510 -4726 -506 -4722
rect -468 -4726 -464 -4722
rect -426 -4726 -422 -4722
rect -385 -4726 -381 -4722
rect -231 -4690 -227 -4686
rect -379 -4733 -375 -4729
rect -231 -4733 -227 -4729
rect -568 -4755 -564 -4751
rect -551 -4755 -547 -4751
rect -531 -4755 -527 -4751
rect -510 -4755 -506 -4751
rect -489 -4755 -485 -4751
rect -468 -4755 -464 -4751
rect -447 -4755 -443 -4751
rect -426 -4755 -422 -4751
rect -405 -4755 -401 -4751
rect -385 -4755 -381 -4751
rect -583 -4811 -579 -4807
rect -577 -4818 -573 -4814
rect -519 -4811 -515 -4807
rect -477 -4818 -473 -4814
rect -459 -4811 -455 -4807
rect -417 -4803 -413 -4799
rect -417 -4811 -413 -4807
rect -435 -4825 -431 -4821
rect -535 -4832 -531 -4828
rect -493 -4832 -489 -4828
rect -379 -4803 -375 -4799
rect -393 -4818 -389 -4814
rect -568 -4847 -564 -4843
rect -551 -4847 -547 -4843
rect -510 -4847 -506 -4843
rect -468 -4847 -464 -4843
rect -426 -4847 -422 -4843
rect -385 -4847 -381 -4843
rect -568 -4873 -564 -4869
rect -551 -4873 -547 -4869
rect -531 -4873 -527 -4869
rect -510 -4873 -506 -4869
rect -489 -4873 -485 -4869
rect -468 -4873 -464 -4869
rect -447 -4873 -443 -4869
rect -426 -4873 -422 -4869
rect -405 -4873 -401 -4869
rect -385 -4873 -381 -4869
rect -577 -4936 -573 -4932
rect -519 -4929 -515 -4925
rect -477 -4936 -473 -4932
rect -459 -4929 -455 -4925
rect -417 -4921 -413 -4917
rect -417 -4929 -413 -4925
rect -435 -4943 -431 -4939
rect -535 -4950 -531 -4946
rect -493 -4950 -489 -4946
rect -393 -4936 -389 -4932
rect -568 -4965 -564 -4961
rect -551 -4965 -547 -4961
rect -510 -4965 -506 -4961
rect -468 -4965 -464 -4961
rect -426 -4965 -422 -4961
rect -385 -4965 -381 -4961
rect -577 -4990 -573 -4986
rect -560 -4990 -556 -4986
rect -589 -5149 -585 -5145
rect -595 -5164 -591 -5160
rect -689 -5208 -685 -5204
rect -589 -5208 -585 -5204
rect -926 -5228 -922 -5224
rect -909 -5228 -905 -5224
rect -889 -5228 -885 -5224
rect -868 -5228 -864 -5224
rect -847 -5228 -843 -5224
rect -826 -5228 -822 -5224
rect -805 -5228 -801 -5224
rect -784 -5228 -780 -5224
rect -763 -5228 -759 -5224
rect -743 -5228 -739 -5224
rect -935 -5291 -931 -5287
rect -877 -5284 -873 -5280
rect -835 -5291 -831 -5287
rect -817 -5284 -813 -5280
rect -775 -5276 -771 -5272
rect -775 -5284 -771 -5280
rect -793 -5298 -789 -5294
rect -893 -5305 -889 -5301
rect -851 -5305 -847 -5301
rect -751 -5291 -747 -5287
rect -926 -5320 -922 -5316
rect -909 -5320 -905 -5316
rect -868 -5320 -864 -5316
rect -826 -5320 -822 -5316
rect -784 -5320 -780 -5316
rect -743 -5320 -739 -5316
rect -926 -5349 -922 -5345
rect -909 -5349 -905 -5345
rect -889 -5349 -885 -5345
rect -868 -5349 -864 -5345
rect -847 -5349 -843 -5345
rect -826 -5349 -822 -5345
rect -805 -5349 -801 -5345
rect -784 -5349 -780 -5345
rect -763 -5349 -759 -5345
rect -743 -5349 -739 -5345
rect -673 -5349 -669 -5345
rect -935 -5412 -931 -5408
rect -877 -5405 -873 -5401
rect -835 -5412 -831 -5408
rect -817 -5405 -813 -5401
rect -775 -5397 -771 -5393
rect -775 -5405 -771 -5401
rect -793 -5419 -789 -5415
rect -893 -5426 -889 -5422
rect -851 -5426 -847 -5422
rect -737 -5397 -733 -5393
rect -751 -5412 -747 -5408
rect -926 -5441 -922 -5437
rect -909 -5441 -905 -5437
rect -868 -5441 -864 -5437
rect -826 -5441 -822 -5437
rect -784 -5441 -780 -5437
rect -743 -5441 -739 -5437
rect -665 -5399 -661 -5395
rect -589 -5405 -585 -5401
rect -673 -5441 -669 -5437
rect -737 -5448 -733 -5444
rect -589 -5449 -585 -5445
rect -926 -5469 -922 -5465
rect -909 -5469 -905 -5465
rect -889 -5469 -885 -5465
rect -868 -5469 -864 -5465
rect -847 -5469 -843 -5465
rect -826 -5469 -822 -5465
rect -805 -5469 -801 -5465
rect -784 -5469 -780 -5465
rect -763 -5469 -759 -5465
rect -743 -5469 -739 -5465
rect -941 -5525 -937 -5521
rect -935 -5532 -931 -5528
rect -877 -5525 -873 -5521
rect -835 -5532 -831 -5528
rect -817 -5525 -813 -5521
rect -775 -5517 -771 -5513
rect -775 -5525 -771 -5521
rect -793 -5539 -789 -5535
rect -893 -5546 -889 -5542
rect -851 -5546 -847 -5542
rect -737 -5517 -733 -5513
rect -751 -5532 -747 -5528
rect -926 -5561 -922 -5557
rect -909 -5561 -905 -5557
rect -868 -5561 -864 -5557
rect -826 -5561 -822 -5557
rect -784 -5561 -780 -5557
rect -743 -5561 -739 -5557
rect -926 -5586 -922 -5582
rect -909 -5586 -905 -5582
rect -889 -5586 -885 -5582
rect -868 -5586 -864 -5582
rect -847 -5586 -843 -5582
rect -826 -5586 -822 -5582
rect -805 -5586 -801 -5582
rect -784 -5586 -780 -5582
rect -763 -5586 -759 -5582
rect -743 -5586 -739 -5582
rect -935 -5649 -931 -5645
rect -877 -5642 -873 -5638
rect -835 -5649 -831 -5645
rect -817 -5642 -813 -5638
rect -775 -5634 -771 -5630
rect -775 -5642 -771 -5638
rect -793 -5656 -789 -5652
rect -893 -5663 -889 -5659
rect -851 -5663 -847 -5659
rect -751 -5649 -747 -5645
rect -926 -5678 -922 -5674
rect -909 -5678 -905 -5674
rect -868 -5678 -864 -5674
rect -826 -5678 -822 -5674
rect -784 -5678 -780 -5674
rect -743 -5678 -739 -5674
rect -935 -5703 -931 -5699
rect -918 -5703 -914 -5699
rect -737 -5735 -733 -5731
rect -909 -5756 -905 -5752
rect -595 -5756 -591 -5752
rect -918 -5795 -914 -5791
rect -926 -5822 -922 -5818
rect -900 -5822 -896 -5818
rect -883 -5822 -879 -5818
rect -843 -5822 -839 -5818
rect -822 -5822 -818 -5818
rect -805 -5822 -801 -5818
rect -765 -5822 -761 -5818
rect -741 -5822 -737 -5818
rect -704 -5822 -700 -5818
rect -947 -5877 -943 -5873
rect -935 -5855 -931 -5851
rect -1162 -5892 -1158 -5888
rect -1255 -5914 -1251 -5910
rect -1211 -5914 -1207 -5910
rect -1177 -5914 -1173 -5910
rect -917 -5848 -913 -5844
rect -891 -5870 -887 -5866
rect -909 -5877 -905 -5873
rect -865 -5862 -861 -5858
rect -813 -5855 -809 -5851
rect -883 -5899 -879 -5895
rect -847 -5899 -843 -5895
rect -787 -5870 -783 -5866
rect -805 -5899 -801 -5895
rect -769 -5899 -765 -5895
rect -695 -5862 -691 -5858
rect -689 -5870 -685 -5866
rect -926 -5914 -922 -5910
rect -900 -5914 -896 -5910
rect -857 -5914 -853 -5910
rect -822 -5914 -818 -5910
rect -778 -5914 -774 -5910
rect -761 -5914 -757 -5910
rect -725 -5914 -721 -5910
rect -704 -5914 -700 -5910
rect -379 -5022 -375 -5018
rect -551 -5043 -547 -5039
rect -237 -5043 -233 -5039
rect -560 -5082 -556 -5078
rect -568 -5109 -564 -5105
rect -542 -5109 -538 -5105
rect -525 -5109 -521 -5105
rect -485 -5109 -481 -5105
rect -464 -5109 -460 -5105
rect -447 -5109 -443 -5105
rect -407 -5109 -403 -5105
rect -383 -5109 -379 -5105
rect -346 -5109 -342 -5105
rect -577 -5142 -573 -5138
rect -559 -5135 -555 -5131
rect -533 -5157 -529 -5153
rect -551 -5164 -547 -5160
rect -507 -5149 -503 -5145
rect -455 -5142 -451 -5138
rect -525 -5186 -521 -5182
rect -489 -5186 -485 -5182
rect -429 -5157 -425 -5153
rect -447 -5186 -443 -5182
rect -411 -5186 -407 -5182
rect -337 -5148 -333 -5144
rect -331 -5157 -327 -5153
rect -568 -5201 -564 -5197
rect -542 -5201 -538 -5197
rect -499 -5201 -495 -5197
rect -464 -5201 -460 -5197
rect -420 -5201 -416 -5197
rect -403 -5201 -399 -5197
rect -367 -5201 -363 -5197
rect -346 -5201 -342 -5197
rect -15 -4303 -11 -4299
rect -21 -4311 -17 -4307
rect -193 -4324 -189 -4320
rect 191 -4324 195 -4320
rect -202 -4363 -198 -4359
rect -210 -4390 -206 -4386
rect -184 -4390 -180 -4386
rect -167 -4390 -163 -4386
rect -127 -4390 -123 -4386
rect -106 -4390 -102 -4386
rect -89 -4390 -85 -4386
rect -49 -4390 -45 -4386
rect -25 -4390 -21 -4386
rect 12 -4390 16 -4386
rect -219 -4423 -215 -4419
rect -201 -4416 -197 -4412
rect -175 -4438 -171 -4434
rect -193 -4445 -189 -4441
rect -149 -4430 -145 -4426
rect -97 -4423 -93 -4419
rect -167 -4467 -163 -4463
rect -131 -4467 -127 -4463
rect -71 -4438 -67 -4434
rect -89 -4467 -85 -4463
rect -53 -4467 -49 -4463
rect 21 -4430 25 -4426
rect 27 -4438 31 -4434
rect -210 -4482 -206 -4478
rect -184 -4482 -180 -4478
rect -141 -4482 -137 -4478
rect -106 -4482 -102 -4478
rect -62 -4482 -58 -4478
rect -45 -4482 -41 -4478
rect -9 -4482 -5 -4478
rect 12 -4482 16 -4478
rect 407 -3458 411 -3454
rect 235 -3479 239 -3475
rect 547 -3479 551 -3475
rect 226 -3518 230 -3514
rect 218 -3550 222 -3546
rect 244 -3550 248 -3546
rect 261 -3550 265 -3546
rect 301 -3550 305 -3546
rect 322 -3550 326 -3546
rect 339 -3550 343 -3546
rect 379 -3550 383 -3546
rect 403 -3550 407 -3546
rect 440 -3550 444 -3546
rect 209 -3583 213 -3579
rect 227 -3576 231 -3572
rect 253 -3598 257 -3594
rect 235 -3605 239 -3601
rect 279 -3590 283 -3586
rect 331 -3583 335 -3579
rect 261 -3627 265 -3623
rect 297 -3627 301 -3623
rect 357 -3598 361 -3594
rect 339 -3627 343 -3623
rect 375 -3627 379 -3623
rect 449 -3590 453 -3586
rect 455 -3598 459 -3594
rect 218 -3642 222 -3638
rect 244 -3642 248 -3638
rect 287 -3642 291 -3638
rect 322 -3642 326 -3638
rect 366 -3642 370 -3638
rect 383 -3642 387 -3638
rect 419 -3642 423 -3638
rect 440 -3642 444 -3638
rect 763 -2752 767 -2748
rect 591 -2773 595 -2769
rect 945 -2773 949 -2769
rect 582 -2812 586 -2808
rect 574 -2839 578 -2835
rect 600 -2839 604 -2835
rect 617 -2839 621 -2835
rect 657 -2839 661 -2835
rect 678 -2839 682 -2835
rect 695 -2839 699 -2835
rect 735 -2839 739 -2835
rect 759 -2839 763 -2835
rect 796 -2839 800 -2835
rect 565 -2872 569 -2868
rect 583 -2865 587 -2861
rect 609 -2887 613 -2883
rect 591 -2894 595 -2890
rect 635 -2879 639 -2875
rect 687 -2872 691 -2868
rect 617 -2916 621 -2912
rect 653 -2916 657 -2912
rect 713 -2887 717 -2883
rect 695 -2916 699 -2912
rect 731 -2916 735 -2912
rect 805 -2879 809 -2875
rect 811 -2887 815 -2883
rect 574 -2931 578 -2927
rect 600 -2931 604 -2927
rect 643 -2931 647 -2927
rect 678 -2931 682 -2927
rect 722 -2931 726 -2927
rect 739 -2931 743 -2927
rect 775 -2931 779 -2927
rect 796 -2931 800 -2927
rect 1211 -1792 1215 -1788
rect 1203 -1835 1207 -1831
rect 1203 -1858 1207 -1854
rect 1211 -1907 1215 -1903
rect 1203 -1950 1207 -1946
rect 1161 -2002 1165 -1998
rect 989 -2023 993 -2019
rect 1303 -2023 1307 -2019
rect 980 -2062 984 -2058
rect 972 -2089 976 -2085
rect 998 -2089 1002 -2085
rect 1015 -2089 1019 -2085
rect 1055 -2089 1059 -2085
rect 1076 -2089 1080 -2085
rect 1093 -2089 1097 -2085
rect 1133 -2089 1137 -2085
rect 1157 -2089 1161 -2085
rect 1194 -2089 1198 -2085
rect 963 -2122 967 -2118
rect 981 -2115 985 -2111
rect 1007 -2137 1011 -2133
rect 989 -2144 993 -2140
rect 1033 -2129 1037 -2125
rect 1085 -2122 1089 -2118
rect 1015 -2166 1019 -2162
rect 1051 -2166 1055 -2162
rect 1111 -2137 1115 -2133
rect 1093 -2166 1097 -2162
rect 1129 -2166 1133 -2162
rect 1203 -2127 1207 -2123
rect 1303 -2129 1307 -2125
rect 1209 -2137 1213 -2133
rect 972 -2181 976 -2177
rect 998 -2181 1002 -2177
rect 1041 -2181 1045 -2177
rect 1076 -2181 1080 -2177
rect 1120 -2181 1124 -2177
rect 1137 -2181 1141 -2177
rect 1173 -2181 1177 -2177
rect 1194 -2181 1198 -2177
rect 1347 -1317 1351 -1313
rect 1338 -1356 1342 -1352
rect 1330 -1378 1334 -1374
rect 1347 -1378 1351 -1374
rect 1387 -1378 1391 -1374
rect 1408 -1378 1412 -1374
rect 1321 -1427 1325 -1423
rect 1365 -1448 1369 -1444
rect 1347 -1455 1351 -1451
rect 1383 -1455 1387 -1451
rect 1330 -1470 1334 -1466
rect 1374 -1470 1378 -1466
rect 1408 -1470 1412 -1466
rect 1417 -1484 1421 -1480
rect 1423 -1448 1427 -1444
rect 1423 -1491 1427 -1487
rect 1330 -1622 1334 -1618
rect 1347 -1622 1351 -1618
rect 1367 -1622 1371 -1618
rect 1388 -1622 1392 -1618
rect 1409 -1622 1413 -1618
rect 1430 -1622 1434 -1618
rect 1451 -1622 1455 -1618
rect 1472 -1622 1476 -1618
rect 1493 -1622 1497 -1618
rect 1513 -1622 1517 -1618
rect 1321 -1685 1325 -1681
rect 1379 -1678 1383 -1674
rect 1421 -1685 1425 -1681
rect 1439 -1678 1443 -1674
rect 1481 -1670 1485 -1666
rect 1481 -1678 1485 -1674
rect 1463 -1692 1467 -1688
rect 1363 -1699 1367 -1695
rect 1405 -1699 1409 -1695
rect 1519 -1670 1523 -1666
rect 1505 -1685 1509 -1681
rect 1330 -1714 1334 -1710
rect 1347 -1714 1351 -1710
rect 1388 -1714 1392 -1710
rect 1430 -1714 1434 -1710
rect 1472 -1714 1476 -1710
rect 1513 -1714 1517 -1710
rect 1519 -1722 1523 -1718
rect 1330 -1743 1334 -1739
rect 1347 -1743 1351 -1739
rect 1367 -1743 1371 -1739
rect 1388 -1743 1392 -1739
rect 1409 -1743 1413 -1739
rect 1430 -1743 1434 -1739
rect 1451 -1743 1455 -1739
rect 1472 -1743 1476 -1739
rect 1493 -1743 1497 -1739
rect 1513 -1743 1517 -1739
rect 1315 -1799 1319 -1795
rect 1321 -1806 1325 -1802
rect 1379 -1799 1383 -1795
rect 1421 -1806 1425 -1802
rect 1439 -1799 1443 -1795
rect 1481 -1791 1485 -1787
rect 1481 -1799 1485 -1795
rect 1463 -1813 1467 -1809
rect 1363 -1820 1367 -1816
rect 1405 -1820 1409 -1816
rect 1519 -1791 1523 -1787
rect 1505 -1806 1509 -1802
rect 1330 -1835 1334 -1831
rect 1347 -1835 1351 -1831
rect 1388 -1835 1392 -1831
rect 1430 -1835 1434 -1831
rect 1472 -1835 1476 -1831
rect 1513 -1835 1517 -1831
rect 1321 -1970 1325 -1966
rect 1338 -1970 1342 -1966
rect 1309 -2144 1313 -2140
rect 1209 -2195 1213 -2191
rect 1309 -2195 1313 -2191
rect 972 -2364 976 -2360
rect 989 -2364 993 -2360
rect 1009 -2364 1013 -2360
rect 1030 -2364 1034 -2360
rect 1051 -2364 1055 -2360
rect 1072 -2364 1076 -2360
rect 1093 -2364 1097 -2360
rect 1114 -2364 1118 -2360
rect 1135 -2364 1139 -2360
rect 1155 -2364 1159 -2360
rect 963 -2427 967 -2423
rect 1021 -2420 1025 -2416
rect 1063 -2427 1067 -2423
rect 1081 -2420 1085 -2416
rect 1123 -2412 1127 -2408
rect 1123 -2420 1127 -2416
rect 1105 -2434 1109 -2430
rect 1005 -2441 1009 -2437
rect 1047 -2441 1051 -2437
rect 1161 -2412 1165 -2408
rect 1147 -2427 1151 -2423
rect 972 -2456 976 -2452
rect 989 -2456 993 -2452
rect 1030 -2456 1034 -2452
rect 1072 -2456 1076 -2452
rect 1114 -2456 1118 -2452
rect 1155 -2456 1159 -2452
rect 1309 -2420 1313 -2416
rect 1161 -2464 1165 -2460
rect 1309 -2464 1313 -2460
rect 972 -2495 976 -2491
rect 989 -2495 993 -2491
rect 1009 -2495 1013 -2491
rect 1030 -2495 1034 -2491
rect 1051 -2495 1055 -2491
rect 1072 -2495 1076 -2491
rect 1093 -2495 1097 -2491
rect 1114 -2495 1118 -2491
rect 1135 -2495 1139 -2491
rect 1155 -2495 1159 -2491
rect 957 -2551 961 -2547
rect 963 -2558 967 -2554
rect 1021 -2551 1025 -2547
rect 1063 -2558 1067 -2554
rect 1081 -2551 1085 -2547
rect 1123 -2543 1127 -2539
rect 1123 -2551 1127 -2547
rect 1105 -2565 1109 -2561
rect 1005 -2572 1009 -2568
rect 1047 -2572 1051 -2568
rect 1161 -2543 1165 -2539
rect 1147 -2558 1151 -2554
rect 972 -2587 976 -2583
rect 989 -2587 993 -2583
rect 1030 -2587 1034 -2583
rect 1072 -2587 1076 -2583
rect 1114 -2587 1118 -2583
rect 1155 -2587 1159 -2583
rect 963 -2720 967 -2716
rect 980 -2720 984 -2716
rect 951 -2879 955 -2875
rect 945 -2894 949 -2890
rect 811 -2938 815 -2934
rect 951 -2938 955 -2934
rect 841 -2958 845 -2954
rect 849 -3007 853 -3003
rect 841 -3050 845 -3046
rect 574 -3074 578 -3070
rect 591 -3074 595 -3070
rect 611 -3074 615 -3070
rect 632 -3074 636 -3070
rect 653 -3074 657 -3070
rect 674 -3074 678 -3070
rect 695 -3074 699 -3070
rect 716 -3074 720 -3070
rect 737 -3074 741 -3070
rect 757 -3074 761 -3070
rect 565 -3137 569 -3133
rect 623 -3130 627 -3126
rect 665 -3137 669 -3133
rect 683 -3130 687 -3126
rect 725 -3122 729 -3118
rect 725 -3130 729 -3126
rect 707 -3144 711 -3140
rect 607 -3151 611 -3147
rect 649 -3151 653 -3147
rect 763 -3122 767 -3118
rect 749 -3137 753 -3133
rect 574 -3166 578 -3162
rect 591 -3166 595 -3162
rect 632 -3166 636 -3162
rect 674 -3166 678 -3162
rect 716 -3166 720 -3162
rect 757 -3166 761 -3162
rect 951 -3130 955 -3126
rect 763 -3173 767 -3169
rect 951 -3173 955 -3169
rect 574 -3195 578 -3191
rect 591 -3195 595 -3191
rect 611 -3195 615 -3191
rect 632 -3195 636 -3191
rect 653 -3195 657 -3191
rect 674 -3195 678 -3191
rect 695 -3195 699 -3191
rect 716 -3195 720 -3191
rect 737 -3195 741 -3191
rect 757 -3195 761 -3191
rect 559 -3251 563 -3247
rect 565 -3258 569 -3254
rect 623 -3251 627 -3247
rect 665 -3258 669 -3254
rect 683 -3251 687 -3247
rect 725 -3243 729 -3239
rect 725 -3251 729 -3247
rect 707 -3265 711 -3261
rect 607 -3272 611 -3268
rect 649 -3272 653 -3268
rect 763 -3243 767 -3239
rect 749 -3258 753 -3254
rect 574 -3287 578 -3283
rect 591 -3287 595 -3283
rect 632 -3287 636 -3283
rect 674 -3287 678 -3283
rect 716 -3287 720 -3283
rect 757 -3287 761 -3283
rect 565 -3426 569 -3422
rect 582 -3426 586 -3422
rect 553 -3590 557 -3586
rect 547 -3605 551 -3601
rect 455 -3656 459 -3652
rect 553 -3656 557 -3652
rect 218 -3911 222 -3907
rect 235 -3911 239 -3907
rect 255 -3911 259 -3907
rect 276 -3911 280 -3907
rect 297 -3911 301 -3907
rect 318 -3911 322 -3907
rect 339 -3911 343 -3907
rect 360 -3911 364 -3907
rect 381 -3911 385 -3907
rect 401 -3911 405 -3907
rect 209 -3974 213 -3970
rect 267 -3967 271 -3963
rect 309 -3974 313 -3970
rect 327 -3967 331 -3963
rect 369 -3959 373 -3955
rect 369 -3967 373 -3963
rect 351 -3981 355 -3977
rect 251 -3988 255 -3984
rect 293 -3988 297 -3984
rect 407 -3959 411 -3955
rect 393 -3974 397 -3970
rect 218 -4003 222 -3999
rect 235 -4003 239 -3999
rect 276 -4003 280 -3999
rect 318 -4003 322 -3999
rect 360 -4003 364 -3999
rect 401 -4003 405 -3999
rect 553 -3967 557 -3963
rect 407 -4010 411 -4006
rect 553 -4011 557 -4007
rect 218 -4036 222 -4032
rect 235 -4036 239 -4032
rect 255 -4036 259 -4032
rect 276 -4036 280 -4032
rect 297 -4036 301 -4032
rect 318 -4036 322 -4032
rect 339 -4036 343 -4032
rect 360 -4036 364 -4032
rect 381 -4036 385 -4032
rect 401 -4036 405 -4032
rect 203 -4092 207 -4088
rect 209 -4099 213 -4095
rect 267 -4092 271 -4088
rect 309 -4099 313 -4095
rect 327 -4092 331 -4088
rect 369 -4084 373 -4080
rect 369 -4092 373 -4088
rect 351 -4106 355 -4102
rect 251 -4113 255 -4109
rect 293 -4113 297 -4109
rect 407 -4084 411 -4080
rect 393 -4099 397 -4095
rect 218 -4128 222 -4124
rect 235 -4128 239 -4124
rect 276 -4128 280 -4124
rect 318 -4128 322 -4124
rect 360 -4128 364 -4124
rect 401 -4128 405 -4124
rect 209 -4271 213 -4267
rect 226 -4271 230 -4267
rect 197 -4430 201 -4426
rect 191 -4445 195 -4441
rect 27 -4489 31 -4485
rect 197 -4489 201 -4485
rect -210 -4634 -206 -4630
rect -193 -4634 -189 -4630
rect -173 -4634 -169 -4630
rect -152 -4634 -148 -4630
rect -131 -4634 -127 -4630
rect -110 -4634 -106 -4630
rect -89 -4634 -85 -4630
rect -68 -4634 -64 -4630
rect -47 -4634 -43 -4630
rect -27 -4634 -23 -4630
rect -219 -4697 -215 -4693
rect -161 -4690 -157 -4686
rect -119 -4697 -115 -4693
rect -101 -4690 -97 -4686
rect -59 -4682 -55 -4678
rect -59 -4690 -55 -4686
rect -77 -4704 -73 -4700
rect -177 -4711 -173 -4707
rect -135 -4711 -131 -4707
rect -21 -4682 -17 -4678
rect -35 -4697 -31 -4693
rect -210 -4726 -206 -4722
rect -193 -4726 -189 -4722
rect -152 -4726 -148 -4722
rect -110 -4726 -106 -4722
rect -68 -4726 -64 -4722
rect -27 -4726 -23 -4722
rect 197 -4690 201 -4686
rect -21 -4733 -17 -4729
rect 197 -4735 201 -4731
rect -210 -4755 -206 -4751
rect -193 -4755 -189 -4751
rect -173 -4755 -169 -4751
rect -152 -4755 -148 -4751
rect -131 -4755 -127 -4751
rect -110 -4755 -106 -4751
rect -89 -4755 -85 -4751
rect -68 -4755 -64 -4751
rect -47 -4755 -43 -4751
rect -27 -4755 -23 -4751
rect -225 -4811 -221 -4807
rect 90 -4755 94 -4751
rect -219 -4818 -215 -4814
rect -161 -4811 -157 -4807
rect -119 -4818 -115 -4814
rect -101 -4811 -97 -4807
rect -59 -4803 -55 -4799
rect -59 -4811 -55 -4807
rect -77 -4825 -73 -4821
rect -177 -4832 -173 -4828
rect -135 -4832 -131 -4828
rect -21 -4803 -17 -4799
rect -35 -4818 -31 -4814
rect -210 -4847 -206 -4843
rect -193 -4847 -189 -4843
rect -152 -4847 -148 -4843
rect -110 -4847 -106 -4843
rect -68 -4847 -64 -4843
rect -27 -4847 -23 -4843
rect -210 -4873 -206 -4869
rect -193 -4873 -189 -4869
rect -173 -4873 -169 -4869
rect -152 -4873 -148 -4869
rect -131 -4873 -127 -4869
rect -110 -4873 -106 -4869
rect -89 -4873 -85 -4869
rect -68 -4873 -64 -4869
rect -47 -4873 -43 -4869
rect -27 -4873 -23 -4869
rect -219 -4936 -215 -4932
rect -161 -4929 -157 -4925
rect -119 -4936 -115 -4932
rect -101 -4929 -97 -4925
rect -59 -4921 -55 -4917
rect -59 -4929 -55 -4925
rect -77 -4943 -73 -4939
rect -177 -4950 -173 -4946
rect -135 -4950 -131 -4946
rect -35 -4936 -31 -4932
rect -210 -4965 -206 -4961
rect -193 -4965 -189 -4961
rect -152 -4965 -148 -4961
rect -110 -4965 -106 -4961
rect -68 -4965 -64 -4961
rect -27 -4965 -23 -4961
rect -219 -4990 -215 -4986
rect -202 -4990 -198 -4986
rect -231 -5149 -227 -5145
rect -237 -5164 -233 -5160
rect -331 -5215 -327 -5211
rect -231 -5215 -227 -5211
rect -568 -5349 -564 -5345
rect -551 -5349 -547 -5345
rect -531 -5349 -527 -5345
rect -510 -5349 -506 -5345
rect -489 -5349 -485 -5345
rect -468 -5349 -464 -5345
rect -447 -5349 -443 -5345
rect -426 -5349 -422 -5345
rect -405 -5349 -401 -5345
rect -385 -5349 -381 -5345
rect -327 -5349 -323 -5345
rect -577 -5412 -573 -5408
rect -519 -5405 -515 -5401
rect -477 -5412 -473 -5408
rect -459 -5405 -455 -5401
rect -417 -5397 -413 -5393
rect -417 -5405 -413 -5401
rect -435 -5419 -431 -5415
rect -535 -5426 -531 -5422
rect -493 -5426 -489 -5422
rect -379 -5397 -375 -5393
rect -393 -5412 -389 -5408
rect -568 -5441 -564 -5437
rect -551 -5441 -547 -5437
rect -510 -5441 -506 -5437
rect -468 -5441 -464 -5437
rect -426 -5441 -422 -5437
rect -385 -5441 -381 -5437
rect -319 -5400 -315 -5396
rect -231 -5405 -227 -5401
rect -327 -5441 -323 -5437
rect -379 -5449 -375 -5445
rect -231 -5448 -227 -5444
rect -568 -5469 -564 -5465
rect -551 -5469 -547 -5465
rect -531 -5469 -527 -5465
rect -510 -5469 -506 -5465
rect -489 -5469 -485 -5465
rect -468 -5469 -464 -5465
rect -447 -5469 -443 -5465
rect -426 -5469 -422 -5465
rect -405 -5469 -401 -5465
rect -385 -5469 -381 -5465
rect -583 -5525 -579 -5521
rect -327 -5469 -323 -5465
rect -577 -5532 -573 -5528
rect -519 -5525 -515 -5521
rect -477 -5532 -473 -5528
rect -459 -5525 -455 -5521
rect -417 -5517 -413 -5513
rect -417 -5525 -413 -5521
rect -435 -5539 -431 -5535
rect -535 -5546 -531 -5542
rect -493 -5546 -489 -5542
rect -379 -5517 -375 -5513
rect -393 -5532 -389 -5528
rect -568 -5561 -564 -5557
rect -551 -5561 -547 -5557
rect -510 -5561 -506 -5557
rect -468 -5561 -464 -5557
rect -426 -5561 -422 -5557
rect -385 -5561 -381 -5557
rect -568 -5586 -564 -5582
rect -551 -5586 -547 -5582
rect -531 -5586 -527 -5582
rect -510 -5586 -506 -5582
rect -489 -5586 -485 -5582
rect -468 -5586 -464 -5582
rect -447 -5586 -443 -5582
rect -426 -5586 -422 -5582
rect -405 -5586 -401 -5582
rect -385 -5586 -381 -5582
rect -577 -5649 -573 -5645
rect -519 -5642 -515 -5638
rect -477 -5649 -473 -5645
rect -459 -5642 -455 -5638
rect -417 -5634 -413 -5630
rect -417 -5642 -413 -5638
rect -435 -5656 -431 -5652
rect -535 -5663 -531 -5659
rect -493 -5663 -489 -5659
rect -393 -5649 -389 -5645
rect -568 -5678 -564 -5674
rect -551 -5678 -547 -5674
rect -510 -5678 -506 -5674
rect -468 -5678 -464 -5674
rect -426 -5678 -422 -5674
rect -385 -5678 -381 -5674
rect -577 -5703 -573 -5699
rect -560 -5703 -556 -5699
rect -319 -5515 -315 -5511
rect -327 -5561 -323 -5557
rect -379 -5735 -375 -5731
rect -551 -5756 -547 -5752
rect -237 -5756 -233 -5752
rect -560 -5795 -556 -5791
rect -568 -5822 -564 -5818
rect -542 -5822 -538 -5818
rect -525 -5822 -521 -5818
rect -485 -5822 -481 -5818
rect -464 -5822 -460 -5818
rect -447 -5822 -443 -5818
rect -407 -5822 -403 -5818
rect -383 -5822 -379 -5818
rect -346 -5822 -342 -5818
rect -589 -5862 -585 -5858
rect -577 -5855 -573 -5851
rect -595 -5877 -591 -5873
rect -559 -5848 -555 -5844
rect -533 -5870 -529 -5866
rect -551 -5877 -547 -5873
rect -507 -5862 -503 -5858
rect -455 -5855 -451 -5851
rect -525 -5899 -521 -5895
rect -489 -5899 -485 -5895
rect -429 -5870 -425 -5866
rect -447 -5899 -443 -5895
rect -411 -5899 -407 -5895
rect -337 -5861 -333 -5857
rect -331 -5870 -327 -5866
rect -568 -5914 -564 -5910
rect -542 -5914 -538 -5910
rect -499 -5914 -495 -5910
rect -464 -5914 -460 -5910
rect -420 -5914 -416 -5910
rect -403 -5914 -399 -5910
rect -367 -5914 -363 -5910
rect -346 -5914 -342 -5910
rect 98 -4806 102 -4802
rect 90 -4847 94 -4843
rect -21 -5022 -17 -5018
rect -193 -5043 -189 -5039
rect 191 -5043 195 -5039
rect -202 -5082 -198 -5078
rect -210 -5109 -206 -5105
rect -184 -5109 -180 -5105
rect -167 -5109 -163 -5105
rect -127 -5109 -123 -5105
rect -106 -5109 -102 -5105
rect -89 -5109 -85 -5105
rect -49 -5109 -45 -5105
rect -25 -5109 -21 -5105
rect 12 -5109 16 -5105
rect -219 -5142 -215 -5138
rect -201 -5135 -197 -5131
rect -175 -5157 -171 -5153
rect -193 -5164 -189 -5160
rect -149 -5149 -145 -5145
rect -97 -5142 -93 -5138
rect -167 -5186 -163 -5182
rect -131 -5186 -127 -5182
rect -71 -5157 -67 -5153
rect -89 -5186 -85 -5182
rect -53 -5186 -49 -5182
rect 21 -5149 25 -5145
rect 27 -5157 31 -5153
rect -210 -5201 -206 -5197
rect -184 -5201 -180 -5197
rect -141 -5201 -137 -5197
rect -106 -5201 -102 -5197
rect -62 -5201 -58 -5197
rect -45 -5201 -41 -5197
rect -9 -5201 -5 -5197
rect 12 -5201 16 -5197
rect 456 -4160 460 -4156
rect 464 -4205 468 -4201
rect 456 -4252 460 -4248
rect 456 -4271 460 -4267
rect 407 -4303 411 -4299
rect 235 -4324 239 -4320
rect 464 -4320 468 -4316
rect 547 -4324 551 -4320
rect 226 -4363 230 -4359
rect 456 -4363 460 -4359
rect 218 -4390 222 -4386
rect 244 -4390 248 -4386
rect 261 -4390 265 -4386
rect 301 -4390 305 -4386
rect 322 -4390 326 -4386
rect 339 -4390 343 -4386
rect 379 -4390 383 -4386
rect 403 -4390 407 -4386
rect 440 -4390 444 -4386
rect 209 -4423 213 -4419
rect 227 -4416 231 -4412
rect 253 -4438 257 -4434
rect 235 -4445 239 -4441
rect 279 -4430 283 -4426
rect 331 -4423 335 -4419
rect 261 -4467 265 -4463
rect 297 -4467 301 -4463
rect 357 -4438 361 -4434
rect 339 -4467 343 -4463
rect 375 -4467 379 -4463
rect 449 -4430 453 -4426
rect 455 -4438 459 -4434
rect 218 -4482 222 -4478
rect 244 -4482 248 -4478
rect 287 -4482 291 -4478
rect 322 -4482 326 -4478
rect 366 -4482 370 -4478
rect 383 -4482 387 -4478
rect 419 -4482 423 -4478
rect 440 -4482 444 -4478
rect 763 -3458 767 -3454
rect 591 -3479 595 -3475
rect 945 -3479 949 -3475
rect 582 -3518 586 -3514
rect 574 -3550 578 -3546
rect 600 -3550 604 -3546
rect 617 -3550 621 -3546
rect 657 -3550 661 -3546
rect 678 -3550 682 -3546
rect 695 -3550 699 -3546
rect 735 -3550 739 -3546
rect 759 -3550 763 -3546
rect 796 -3550 800 -3546
rect 565 -3583 569 -3579
rect 583 -3576 587 -3572
rect 609 -3598 613 -3594
rect 591 -3605 595 -3601
rect 635 -3590 639 -3586
rect 687 -3583 691 -3579
rect 617 -3627 621 -3623
rect 653 -3627 657 -3623
rect 713 -3598 717 -3594
rect 695 -3627 699 -3623
rect 731 -3627 735 -3623
rect 805 -3590 809 -3586
rect 811 -3598 815 -3594
rect 574 -3642 578 -3638
rect 600 -3642 604 -3638
rect 643 -3642 647 -3638
rect 678 -3642 682 -3638
rect 722 -3642 726 -3638
rect 739 -3642 743 -3638
rect 775 -3642 779 -3638
rect 796 -3642 800 -3638
rect 1161 -2752 1165 -2748
rect 989 -2773 993 -2769
rect 1303 -2773 1307 -2769
rect 980 -2812 984 -2808
rect 972 -2839 976 -2835
rect 998 -2839 1002 -2835
rect 1015 -2839 1019 -2835
rect 1055 -2839 1059 -2835
rect 1076 -2839 1080 -2835
rect 1093 -2839 1097 -2835
rect 1133 -2839 1137 -2835
rect 1157 -2839 1161 -2835
rect 1194 -2839 1198 -2835
rect 963 -2872 967 -2868
rect 981 -2865 985 -2861
rect 1007 -2887 1011 -2883
rect 989 -2894 993 -2890
rect 1033 -2879 1037 -2875
rect 1085 -2872 1089 -2868
rect 1015 -2916 1019 -2912
rect 1051 -2916 1055 -2912
rect 1111 -2887 1115 -2883
rect 1093 -2916 1097 -2912
rect 1129 -2916 1133 -2912
rect 1203 -2877 1207 -2873
rect 1303 -2879 1307 -2875
rect 1209 -2887 1213 -2883
rect 972 -2931 976 -2927
rect 998 -2931 1002 -2927
rect 1041 -2931 1045 -2927
rect 1076 -2931 1080 -2927
rect 1120 -2931 1124 -2927
rect 1137 -2931 1141 -2927
rect 1173 -2931 1177 -2927
rect 1194 -2931 1198 -2927
rect 1519 -2002 1523 -1998
rect 1347 -2023 1351 -2019
rect 1338 -2062 1342 -2058
rect 1330 -2089 1334 -2085
rect 1356 -2089 1360 -2085
rect 1373 -2089 1377 -2085
rect 1413 -2089 1417 -2085
rect 1434 -2089 1438 -2085
rect 1451 -2089 1455 -2085
rect 1491 -2089 1495 -2085
rect 1515 -2089 1519 -2085
rect 1552 -2089 1556 -2085
rect 1321 -2122 1325 -2118
rect 1339 -2115 1343 -2111
rect 1365 -2137 1369 -2133
rect 1347 -2144 1351 -2140
rect 1391 -2129 1395 -2125
rect 1443 -2122 1447 -2118
rect 1373 -2166 1377 -2162
rect 1409 -2166 1413 -2162
rect 1469 -2137 1473 -2133
rect 1451 -2166 1455 -2162
rect 1487 -2166 1491 -2162
rect 1330 -2181 1334 -2177
rect 1356 -2181 1360 -2177
rect 1399 -2181 1403 -2177
rect 1434 -2181 1438 -2177
rect 1478 -2181 1482 -2177
rect 1495 -2181 1499 -2177
rect 1531 -2181 1535 -2177
rect 1552 -2181 1556 -2177
rect 1567 -2137 1571 -2133
rect 1567 -2188 1571 -2184
rect 1561 -2195 1565 -2191
rect 1330 -2364 1334 -2360
rect 1347 -2364 1351 -2360
rect 1367 -2364 1371 -2360
rect 1388 -2364 1392 -2360
rect 1409 -2364 1413 -2360
rect 1430 -2364 1434 -2360
rect 1451 -2364 1455 -2360
rect 1472 -2364 1476 -2360
rect 1493 -2364 1497 -2360
rect 1513 -2364 1517 -2360
rect 1321 -2427 1325 -2423
rect 1379 -2420 1383 -2416
rect 1421 -2427 1425 -2423
rect 1439 -2420 1443 -2416
rect 1481 -2412 1485 -2408
rect 1481 -2420 1485 -2416
rect 1463 -2434 1467 -2430
rect 1363 -2441 1367 -2437
rect 1405 -2441 1409 -2437
rect 1519 -2412 1523 -2408
rect 1505 -2427 1509 -2423
rect 1330 -2456 1334 -2452
rect 1347 -2456 1351 -2452
rect 1388 -2456 1392 -2452
rect 1430 -2456 1434 -2452
rect 1472 -2456 1476 -2452
rect 1513 -2456 1517 -2452
rect 1519 -2464 1523 -2460
rect 1330 -2495 1334 -2491
rect 1347 -2495 1351 -2491
rect 1367 -2495 1371 -2491
rect 1388 -2495 1392 -2491
rect 1409 -2495 1413 -2491
rect 1430 -2495 1434 -2491
rect 1451 -2495 1455 -2491
rect 1472 -2495 1476 -2491
rect 1493 -2495 1497 -2491
rect 1513 -2495 1517 -2491
rect 1315 -2551 1319 -2547
rect 1321 -2558 1325 -2554
rect 1379 -2551 1383 -2547
rect 1421 -2558 1425 -2554
rect 1439 -2551 1443 -2547
rect 1481 -2543 1485 -2539
rect 1481 -2551 1485 -2547
rect 1463 -2565 1467 -2561
rect 1363 -2572 1367 -2568
rect 1405 -2572 1409 -2568
rect 1519 -2543 1523 -2539
rect 1505 -2558 1509 -2554
rect 1330 -2587 1334 -2583
rect 1347 -2587 1351 -2583
rect 1388 -2587 1392 -2583
rect 1430 -2587 1434 -2583
rect 1472 -2587 1476 -2583
rect 1513 -2587 1517 -2583
rect 1321 -2720 1325 -2716
rect 1338 -2720 1342 -2716
rect 1309 -2894 1313 -2890
rect 1209 -2945 1213 -2941
rect 1309 -2945 1313 -2941
rect 1199 -2958 1203 -2954
rect 1207 -3008 1211 -3004
rect 1199 -3050 1203 -3046
rect 972 -3074 976 -3070
rect 989 -3074 993 -3070
rect 1009 -3074 1013 -3070
rect 1030 -3074 1034 -3070
rect 1051 -3074 1055 -3070
rect 1072 -3074 1076 -3070
rect 1093 -3074 1097 -3070
rect 1114 -3074 1118 -3070
rect 1135 -3074 1139 -3070
rect 1155 -3074 1159 -3070
rect 1199 -3074 1203 -3070
rect 963 -3137 967 -3133
rect 1021 -3130 1025 -3126
rect 1063 -3137 1067 -3133
rect 1081 -3130 1085 -3126
rect 1123 -3122 1127 -3118
rect 1123 -3130 1127 -3126
rect 1105 -3144 1109 -3140
rect 1005 -3151 1009 -3147
rect 1047 -3151 1051 -3147
rect 1161 -3122 1165 -3118
rect 1147 -3137 1151 -3133
rect 972 -3166 976 -3162
rect 989 -3166 993 -3162
rect 1030 -3166 1034 -3162
rect 1072 -3166 1076 -3162
rect 1114 -3166 1118 -3162
rect 1155 -3166 1159 -3162
rect 1207 -3123 1211 -3119
rect 1309 -3130 1313 -3126
rect 1199 -3166 1203 -3162
rect 1161 -3173 1165 -3169
rect 1309 -3174 1313 -3170
rect 972 -3195 976 -3191
rect 989 -3195 993 -3191
rect 1009 -3195 1013 -3191
rect 1030 -3195 1034 -3191
rect 1051 -3195 1055 -3191
rect 1072 -3195 1076 -3191
rect 1093 -3195 1097 -3191
rect 1114 -3195 1118 -3191
rect 1135 -3195 1139 -3191
rect 1155 -3195 1159 -3191
rect 957 -3251 961 -3247
rect 963 -3258 967 -3254
rect 1021 -3251 1025 -3247
rect 1063 -3258 1067 -3254
rect 1081 -3251 1085 -3247
rect 1123 -3243 1127 -3239
rect 1123 -3251 1127 -3247
rect 1105 -3265 1109 -3261
rect 1005 -3272 1009 -3268
rect 1047 -3272 1051 -3268
rect 1161 -3243 1165 -3239
rect 1147 -3258 1151 -3254
rect 972 -3287 976 -3283
rect 989 -3287 993 -3283
rect 1030 -3287 1034 -3283
rect 1072 -3287 1076 -3283
rect 1114 -3287 1118 -3283
rect 1155 -3287 1159 -3283
rect 963 -3426 967 -3422
rect 980 -3426 984 -3422
rect 951 -3590 955 -3586
rect 945 -3605 949 -3601
rect 811 -3649 815 -3645
rect 951 -3649 955 -3645
rect 574 -3911 578 -3907
rect 591 -3911 595 -3907
rect 611 -3911 615 -3907
rect 632 -3911 636 -3907
rect 653 -3911 657 -3907
rect 674 -3911 678 -3907
rect 695 -3911 699 -3907
rect 716 -3911 720 -3907
rect 737 -3911 741 -3907
rect 757 -3911 761 -3907
rect 565 -3974 569 -3970
rect 623 -3967 627 -3963
rect 665 -3974 669 -3970
rect 683 -3967 687 -3963
rect 725 -3959 729 -3955
rect 725 -3967 729 -3963
rect 707 -3981 711 -3977
rect 607 -3988 611 -3984
rect 649 -3988 653 -3984
rect 763 -3959 767 -3955
rect 749 -3974 753 -3970
rect 574 -4003 578 -3999
rect 591 -4003 595 -3999
rect 632 -4003 636 -3999
rect 674 -4003 678 -3999
rect 716 -4003 720 -3999
rect 757 -4003 761 -3999
rect 951 -3967 955 -3963
rect 763 -4011 767 -4007
rect 951 -4010 955 -4006
rect 574 -4036 578 -4032
rect 591 -4036 595 -4032
rect 611 -4036 615 -4032
rect 632 -4036 636 -4032
rect 653 -4036 657 -4032
rect 674 -4036 678 -4032
rect 695 -4036 699 -4032
rect 716 -4036 720 -4032
rect 737 -4036 741 -4032
rect 757 -4036 761 -4032
rect 559 -4092 563 -4088
rect 565 -4099 569 -4095
rect 623 -4092 627 -4088
rect 665 -4099 669 -4095
rect 683 -4092 687 -4088
rect 725 -4084 729 -4080
rect 725 -4092 729 -4088
rect 707 -4106 711 -4102
rect 607 -4113 611 -4109
rect 649 -4113 653 -4109
rect 763 -4084 767 -4080
rect 749 -4099 753 -4095
rect 574 -4128 578 -4124
rect 591 -4128 595 -4124
rect 632 -4128 636 -4124
rect 674 -4128 678 -4124
rect 716 -4128 720 -4124
rect 757 -4128 761 -4124
rect 565 -4271 569 -4267
rect 582 -4271 586 -4267
rect 553 -4430 557 -4426
rect 547 -4445 551 -4441
rect 455 -4496 459 -4492
rect 553 -4496 557 -4492
rect 218 -4634 222 -4630
rect 235 -4634 239 -4630
rect 255 -4634 259 -4630
rect 276 -4634 280 -4630
rect 297 -4634 301 -4630
rect 318 -4634 322 -4630
rect 339 -4634 343 -4630
rect 360 -4634 364 -4630
rect 381 -4634 385 -4630
rect 401 -4634 405 -4630
rect 209 -4697 213 -4693
rect 267 -4690 271 -4686
rect 309 -4697 313 -4693
rect 327 -4690 331 -4686
rect 369 -4682 373 -4678
rect 369 -4690 373 -4686
rect 351 -4704 355 -4700
rect 251 -4711 255 -4707
rect 293 -4711 297 -4707
rect 407 -4682 411 -4678
rect 393 -4697 397 -4693
rect 218 -4726 222 -4722
rect 235 -4726 239 -4722
rect 276 -4726 280 -4722
rect 318 -4726 322 -4722
rect 360 -4726 364 -4722
rect 401 -4726 405 -4722
rect 553 -4690 557 -4686
rect 407 -4735 411 -4731
rect 553 -4734 557 -4730
rect 218 -4755 222 -4751
rect 235 -4755 239 -4751
rect 255 -4755 259 -4751
rect 276 -4755 280 -4751
rect 297 -4755 301 -4751
rect 318 -4755 322 -4751
rect 339 -4755 343 -4751
rect 360 -4755 364 -4751
rect 381 -4755 385 -4751
rect 401 -4755 405 -4751
rect 203 -4811 207 -4807
rect 209 -4818 213 -4814
rect 267 -4811 271 -4807
rect 309 -4818 313 -4814
rect 327 -4811 331 -4807
rect 369 -4803 373 -4799
rect 369 -4811 373 -4807
rect 351 -4825 355 -4821
rect 251 -4832 255 -4828
rect 293 -4832 297 -4828
rect 413 -4803 417 -4799
rect 393 -4818 397 -4814
rect 218 -4847 222 -4843
rect 235 -4847 239 -4843
rect 276 -4847 280 -4843
rect 318 -4847 322 -4843
rect 360 -4847 364 -4843
rect 401 -4847 405 -4843
rect 218 -4873 222 -4869
rect 235 -4873 239 -4869
rect 255 -4873 259 -4869
rect 276 -4873 280 -4869
rect 297 -4873 301 -4869
rect 318 -4873 322 -4869
rect 339 -4873 343 -4869
rect 360 -4873 364 -4869
rect 381 -4873 385 -4869
rect 401 -4873 405 -4869
rect 209 -4936 213 -4932
rect 267 -4929 271 -4925
rect 309 -4936 313 -4932
rect 327 -4929 331 -4925
rect 369 -4921 373 -4917
rect 369 -4929 373 -4925
rect 351 -4943 355 -4939
rect 251 -4950 255 -4946
rect 293 -4950 297 -4946
rect 407 -4921 411 -4917
rect 393 -4936 397 -4932
rect 218 -4965 222 -4961
rect 235 -4965 239 -4961
rect 276 -4965 280 -4961
rect 318 -4965 322 -4961
rect 360 -4965 364 -4961
rect 401 -4965 405 -4961
rect 209 -4990 213 -4986
rect 226 -4990 230 -4986
rect 197 -5149 201 -5145
rect 191 -5164 195 -5160
rect 27 -5208 31 -5204
rect 197 -5208 201 -5204
rect -210 -5349 -206 -5345
rect -193 -5349 -189 -5345
rect -173 -5349 -169 -5345
rect -152 -5349 -148 -5345
rect -131 -5349 -127 -5345
rect -110 -5349 -106 -5345
rect -89 -5349 -85 -5345
rect -68 -5349 -64 -5345
rect -47 -5349 -43 -5345
rect -27 -5349 -23 -5345
rect -219 -5412 -215 -5408
rect -161 -5405 -157 -5401
rect -119 -5412 -115 -5408
rect -101 -5405 -97 -5401
rect -59 -5397 -55 -5393
rect -59 -5405 -55 -5401
rect -77 -5419 -73 -5415
rect -177 -5426 -173 -5422
rect -135 -5426 -131 -5422
rect -21 -5397 -17 -5393
rect -35 -5412 -31 -5408
rect -210 -5441 -206 -5437
rect -193 -5441 -189 -5437
rect -152 -5441 -148 -5437
rect -110 -5441 -106 -5437
rect -68 -5441 -64 -5437
rect -27 -5441 -23 -5437
rect 197 -5405 201 -5401
rect -21 -5448 -17 -5444
rect 197 -5448 201 -5444
rect -210 -5469 -206 -5465
rect -193 -5469 -189 -5465
rect -173 -5469 -169 -5465
rect -152 -5469 -148 -5465
rect -131 -5469 -127 -5465
rect -110 -5469 -106 -5465
rect -89 -5469 -85 -5465
rect -68 -5469 -64 -5465
rect -47 -5469 -43 -5465
rect -27 -5469 -23 -5465
rect -225 -5525 -221 -5521
rect -219 -5532 -215 -5528
rect -161 -5525 -157 -5521
rect -119 -5532 -115 -5528
rect -101 -5525 -97 -5521
rect -59 -5517 -55 -5513
rect -59 -5525 -55 -5521
rect -77 -5539 -73 -5535
rect -177 -5546 -173 -5542
rect -135 -5546 -131 -5542
rect -21 -5517 -17 -5513
rect -35 -5532 -31 -5528
rect -210 -5561 -206 -5557
rect -193 -5561 -189 -5557
rect -152 -5561 -148 -5557
rect -110 -5561 -106 -5557
rect -68 -5561 -64 -5557
rect -27 -5561 -23 -5557
rect -210 -5586 -206 -5582
rect -193 -5586 -189 -5582
rect -173 -5586 -169 -5582
rect -152 -5586 -148 -5582
rect -131 -5586 -127 -5582
rect -110 -5586 -106 -5582
rect -89 -5586 -85 -5582
rect -68 -5586 -64 -5582
rect -47 -5586 -43 -5582
rect -27 -5586 -23 -5582
rect -219 -5649 -215 -5645
rect -161 -5642 -157 -5638
rect -119 -5649 -115 -5645
rect -101 -5642 -97 -5638
rect -59 -5634 -55 -5630
rect -59 -5642 -55 -5638
rect -77 -5656 -73 -5652
rect -177 -5663 -173 -5659
rect -135 -5663 -131 -5659
rect -35 -5649 -31 -5645
rect -210 -5678 -206 -5674
rect -193 -5678 -189 -5674
rect -152 -5678 -148 -5674
rect -110 -5678 -106 -5674
rect -68 -5678 -64 -5674
rect -27 -5678 -23 -5674
rect -219 -5703 -215 -5699
rect -202 -5703 -198 -5699
rect -21 -5735 -17 -5731
rect -193 -5756 -189 -5752
rect 191 -5756 195 -5752
rect -202 -5795 -198 -5791
rect -210 -5822 -206 -5818
rect -184 -5822 -180 -5818
rect -167 -5822 -163 -5818
rect -127 -5822 -123 -5818
rect -106 -5822 -102 -5818
rect -89 -5822 -85 -5818
rect -49 -5822 -45 -5818
rect -25 -5822 -21 -5818
rect 12 -5822 16 -5818
rect -231 -5862 -227 -5858
rect -219 -5855 -215 -5851
rect -237 -5877 -233 -5873
rect -201 -5848 -197 -5844
rect -175 -5870 -171 -5866
rect -193 -5877 -189 -5873
rect -149 -5862 -145 -5858
rect -97 -5855 -93 -5851
rect -167 -5899 -163 -5895
rect -131 -5899 -127 -5895
rect -71 -5870 -67 -5866
rect -89 -5899 -85 -5895
rect -53 -5899 -49 -5895
rect 21 -5862 25 -5858
rect 27 -5870 31 -5866
rect -210 -5914 -206 -5910
rect -184 -5914 -180 -5910
rect -141 -5914 -137 -5910
rect -106 -5914 -102 -5910
rect -62 -5914 -58 -5910
rect -45 -5914 -41 -5910
rect -9 -5914 -5 -5910
rect 12 -5914 16 -5910
rect 413 -5022 417 -5018
rect 407 -5030 411 -5026
rect 235 -5043 239 -5039
rect 547 -5043 551 -5039
rect 226 -5082 230 -5078
rect 218 -5109 222 -5105
rect 244 -5109 248 -5105
rect 261 -5109 265 -5105
rect 301 -5109 305 -5105
rect 322 -5109 326 -5105
rect 339 -5109 343 -5105
rect 379 -5109 383 -5105
rect 403 -5109 407 -5105
rect 440 -5109 444 -5105
rect 209 -5142 213 -5138
rect 227 -5135 231 -5131
rect 253 -5157 257 -5153
rect 235 -5164 239 -5160
rect 279 -5149 283 -5145
rect 331 -5142 335 -5138
rect 261 -5186 265 -5182
rect 297 -5186 301 -5182
rect 357 -5157 361 -5153
rect 339 -5186 343 -5182
rect 375 -5186 379 -5182
rect 449 -5149 453 -5145
rect 455 -5157 459 -5153
rect 218 -5201 222 -5197
rect 244 -5201 248 -5197
rect 287 -5201 291 -5197
rect 322 -5201 326 -5197
rect 366 -5201 370 -5197
rect 383 -5201 387 -5197
rect 419 -5201 423 -5197
rect 440 -5201 444 -5197
rect 860 -4271 864 -4267
rect 763 -4303 767 -4299
rect 591 -4324 595 -4320
rect 868 -4321 872 -4317
rect 945 -4324 949 -4320
rect 582 -4363 586 -4359
rect 860 -4363 864 -4359
rect 574 -4390 578 -4386
rect 600 -4390 604 -4386
rect 617 -4390 621 -4386
rect 657 -4390 661 -4386
rect 678 -4390 682 -4386
rect 695 -4390 699 -4386
rect 735 -4390 739 -4386
rect 759 -4390 763 -4386
rect 796 -4390 800 -4386
rect 565 -4423 569 -4419
rect 583 -4416 587 -4412
rect 609 -4438 613 -4434
rect 591 -4445 595 -4441
rect 635 -4430 639 -4426
rect 687 -4423 691 -4419
rect 617 -4467 621 -4463
rect 653 -4467 657 -4463
rect 713 -4438 717 -4434
rect 695 -4467 699 -4463
rect 731 -4467 735 -4463
rect 805 -4430 809 -4426
rect 811 -4438 815 -4434
rect 574 -4482 578 -4478
rect 600 -4482 604 -4478
rect 643 -4482 647 -4478
rect 678 -4482 682 -4478
rect 722 -4482 726 -4478
rect 739 -4482 743 -4478
rect 775 -4482 779 -4478
rect 796 -4482 800 -4478
rect 1161 -3458 1165 -3454
rect 989 -3479 993 -3475
rect 1303 -3479 1307 -3475
rect 980 -3518 984 -3514
rect 972 -3550 976 -3546
rect 998 -3550 1002 -3546
rect 1015 -3550 1019 -3546
rect 1055 -3550 1059 -3546
rect 1076 -3550 1080 -3546
rect 1093 -3550 1097 -3546
rect 1133 -3550 1137 -3546
rect 1157 -3550 1161 -3546
rect 1194 -3550 1198 -3546
rect 963 -3583 967 -3579
rect 981 -3576 985 -3572
rect 1007 -3598 1011 -3594
rect 989 -3605 993 -3601
rect 1033 -3590 1037 -3586
rect 1085 -3583 1089 -3579
rect 1015 -3627 1019 -3623
rect 1051 -3627 1055 -3623
rect 1111 -3598 1115 -3594
rect 1093 -3627 1097 -3623
rect 1129 -3627 1133 -3623
rect 1203 -3588 1207 -3584
rect 1303 -3590 1307 -3586
rect 1209 -3598 1213 -3594
rect 972 -3642 976 -3638
rect 998 -3642 1002 -3638
rect 1041 -3642 1045 -3638
rect 1076 -3642 1080 -3638
rect 1120 -3642 1124 -3638
rect 1137 -3642 1141 -3638
rect 1173 -3642 1177 -3638
rect 1194 -3642 1198 -3638
rect 1519 -2752 1523 -2748
rect 1347 -2773 1351 -2769
rect 1338 -2812 1342 -2808
rect 1330 -2839 1334 -2835
rect 1356 -2839 1360 -2835
rect 1373 -2839 1377 -2835
rect 1413 -2839 1417 -2835
rect 1434 -2839 1438 -2835
rect 1451 -2839 1455 -2835
rect 1491 -2839 1495 -2835
rect 1515 -2839 1519 -2835
rect 1552 -2839 1556 -2835
rect 1321 -2872 1325 -2868
rect 1339 -2865 1343 -2861
rect 1365 -2887 1369 -2883
rect 1347 -2894 1351 -2890
rect 1391 -2879 1395 -2875
rect 1443 -2872 1447 -2868
rect 1373 -2916 1377 -2912
rect 1409 -2916 1413 -2912
rect 1469 -2887 1473 -2883
rect 1451 -2916 1455 -2912
rect 1487 -2916 1491 -2912
rect 1330 -2931 1334 -2927
rect 1356 -2931 1360 -2927
rect 1399 -2931 1403 -2927
rect 1434 -2931 1438 -2927
rect 1478 -2931 1482 -2927
rect 1495 -2931 1499 -2927
rect 1531 -2931 1535 -2927
rect 1552 -2931 1556 -2927
rect 1567 -2887 1571 -2883
rect 1567 -2938 1571 -2934
rect 1561 -2945 1565 -2941
rect 1330 -3074 1334 -3070
rect 1347 -3074 1351 -3070
rect 1367 -3074 1371 -3070
rect 1388 -3074 1392 -3070
rect 1409 -3074 1413 -3070
rect 1430 -3074 1434 -3070
rect 1451 -3074 1455 -3070
rect 1472 -3074 1476 -3070
rect 1493 -3074 1497 -3070
rect 1513 -3074 1517 -3070
rect 1321 -3137 1325 -3133
rect 1379 -3130 1383 -3126
rect 1421 -3137 1425 -3133
rect 1439 -3130 1443 -3126
rect 1481 -3122 1485 -3118
rect 1481 -3130 1485 -3126
rect 1463 -3144 1467 -3140
rect 1363 -3151 1367 -3147
rect 1405 -3151 1409 -3147
rect 1519 -3122 1523 -3118
rect 1505 -3137 1509 -3133
rect 1330 -3166 1334 -3162
rect 1347 -3166 1351 -3162
rect 1388 -3166 1392 -3162
rect 1430 -3166 1434 -3162
rect 1472 -3166 1476 -3162
rect 1513 -3166 1517 -3162
rect 1519 -3174 1523 -3170
rect 1330 -3195 1334 -3191
rect 1347 -3195 1351 -3191
rect 1367 -3195 1371 -3191
rect 1388 -3195 1392 -3191
rect 1409 -3195 1413 -3191
rect 1430 -3195 1434 -3191
rect 1451 -3195 1455 -3191
rect 1472 -3195 1476 -3191
rect 1493 -3195 1497 -3191
rect 1513 -3195 1517 -3191
rect 1315 -3251 1319 -3247
rect 1321 -3258 1325 -3254
rect 1379 -3251 1383 -3247
rect 1421 -3258 1425 -3254
rect 1439 -3251 1443 -3247
rect 1481 -3243 1485 -3239
rect 1481 -3251 1485 -3247
rect 1463 -3265 1467 -3261
rect 1363 -3272 1367 -3268
rect 1405 -3272 1409 -3268
rect 1519 -3243 1523 -3239
rect 1505 -3258 1509 -3254
rect 1330 -3287 1334 -3283
rect 1347 -3287 1351 -3283
rect 1388 -3287 1392 -3283
rect 1430 -3287 1434 -3283
rect 1472 -3287 1476 -3283
rect 1513 -3287 1517 -3283
rect 1321 -3426 1325 -3422
rect 1338 -3426 1342 -3422
rect 1309 -3605 1313 -3601
rect 1209 -3656 1213 -3652
rect 1309 -3656 1313 -3652
rect 972 -3911 976 -3907
rect 989 -3911 993 -3907
rect 1009 -3911 1013 -3907
rect 1030 -3911 1034 -3907
rect 1051 -3911 1055 -3907
rect 1072 -3911 1076 -3907
rect 1093 -3911 1097 -3907
rect 1114 -3911 1118 -3907
rect 1135 -3911 1139 -3907
rect 1155 -3911 1159 -3907
rect 963 -3974 967 -3970
rect 1021 -3967 1025 -3963
rect 1063 -3974 1067 -3970
rect 1081 -3967 1085 -3963
rect 1123 -3959 1127 -3955
rect 1123 -3967 1127 -3963
rect 1105 -3981 1109 -3977
rect 1005 -3988 1009 -3984
rect 1047 -3988 1051 -3984
rect 1161 -3959 1165 -3955
rect 1147 -3974 1151 -3970
rect 972 -4003 976 -3999
rect 989 -4003 993 -3999
rect 1030 -4003 1034 -3999
rect 1072 -4003 1076 -3999
rect 1114 -4003 1118 -3999
rect 1155 -4003 1159 -3999
rect 1309 -3967 1313 -3963
rect 1161 -4010 1165 -4006
rect 1309 -4010 1313 -4006
rect 972 -4036 976 -4032
rect 989 -4036 993 -4032
rect 1009 -4036 1013 -4032
rect 1030 -4036 1034 -4032
rect 1051 -4036 1055 -4032
rect 1072 -4036 1076 -4032
rect 1093 -4036 1097 -4032
rect 1114 -4036 1118 -4032
rect 1135 -4036 1139 -4032
rect 1155 -4036 1159 -4032
rect 957 -4092 961 -4088
rect 963 -4099 967 -4095
rect 1021 -4092 1025 -4088
rect 1063 -4099 1067 -4095
rect 1081 -4092 1085 -4088
rect 1123 -4084 1127 -4080
rect 1123 -4092 1127 -4088
rect 1105 -4106 1109 -4102
rect 1005 -4113 1009 -4109
rect 1047 -4113 1051 -4109
rect 1161 -4084 1165 -4080
rect 1147 -4099 1151 -4095
rect 972 -4128 976 -4124
rect 989 -4128 993 -4124
rect 1030 -4128 1034 -4124
rect 1072 -4128 1076 -4124
rect 1114 -4128 1118 -4124
rect 1155 -4128 1159 -4124
rect 963 -4271 967 -4267
rect 980 -4271 984 -4267
rect 951 -4430 955 -4426
rect 945 -4445 949 -4441
rect 811 -4489 815 -4485
rect 951 -4489 955 -4485
rect 574 -4634 578 -4630
rect 591 -4634 595 -4630
rect 611 -4634 615 -4630
rect 632 -4634 636 -4630
rect 653 -4634 657 -4630
rect 674 -4634 678 -4630
rect 695 -4634 699 -4630
rect 716 -4634 720 -4630
rect 737 -4634 741 -4630
rect 757 -4634 761 -4630
rect 565 -4697 569 -4693
rect 623 -4690 627 -4686
rect 665 -4697 669 -4693
rect 683 -4690 687 -4686
rect 725 -4682 729 -4678
rect 725 -4690 729 -4686
rect 707 -4704 711 -4700
rect 607 -4711 611 -4707
rect 649 -4711 653 -4707
rect 763 -4682 767 -4678
rect 749 -4697 753 -4693
rect 574 -4726 578 -4722
rect 591 -4726 595 -4722
rect 632 -4726 636 -4722
rect 674 -4726 678 -4722
rect 716 -4726 720 -4722
rect 757 -4726 761 -4722
rect 951 -4690 955 -4686
rect 763 -4734 767 -4730
rect 951 -4733 955 -4729
rect 574 -4755 578 -4751
rect 591 -4755 595 -4751
rect 611 -4755 615 -4751
rect 632 -4755 636 -4751
rect 653 -4755 657 -4751
rect 674 -4755 678 -4751
rect 695 -4755 699 -4751
rect 716 -4755 720 -4751
rect 737 -4755 741 -4751
rect 757 -4755 761 -4751
rect 559 -4811 563 -4807
rect 565 -4818 569 -4814
rect 623 -4811 627 -4807
rect 665 -4818 669 -4814
rect 683 -4811 687 -4807
rect 725 -4803 729 -4799
rect 725 -4811 729 -4807
rect 707 -4825 711 -4821
rect 607 -4832 611 -4828
rect 649 -4832 653 -4828
rect 763 -4803 767 -4799
rect 749 -4818 753 -4814
rect 574 -4847 578 -4843
rect 591 -4847 595 -4843
rect 632 -4847 636 -4843
rect 674 -4847 678 -4843
rect 716 -4847 720 -4843
rect 757 -4847 761 -4843
rect 565 -4990 569 -4986
rect 582 -4990 586 -4986
rect 553 -5149 557 -5145
rect 547 -5164 551 -5160
rect 455 -5215 459 -5211
rect 553 -5215 557 -5211
rect 218 -5349 222 -5345
rect 235 -5349 239 -5345
rect 255 -5349 259 -5345
rect 276 -5349 280 -5345
rect 297 -5349 301 -5345
rect 318 -5349 322 -5345
rect 339 -5349 343 -5345
rect 360 -5349 364 -5345
rect 381 -5349 385 -5345
rect 401 -5349 405 -5345
rect 466 -5349 470 -5345
rect 209 -5412 213 -5408
rect 267 -5405 271 -5401
rect 309 -5412 313 -5408
rect 327 -5405 331 -5401
rect 369 -5397 373 -5393
rect 369 -5405 373 -5401
rect 351 -5419 355 -5415
rect 251 -5426 255 -5422
rect 293 -5426 297 -5422
rect 407 -5397 411 -5393
rect 474 -5394 478 -5390
rect 393 -5412 397 -5408
rect 218 -5441 222 -5437
rect 235 -5441 239 -5437
rect 276 -5441 280 -5437
rect 318 -5441 322 -5437
rect 360 -5441 364 -5437
rect 401 -5441 405 -5437
rect 553 -5405 557 -5401
rect 466 -5441 470 -5437
rect 407 -5448 411 -5444
rect 553 -5450 557 -5446
rect 218 -5469 222 -5465
rect 235 -5469 239 -5465
rect 255 -5469 259 -5465
rect 276 -5469 280 -5465
rect 297 -5469 301 -5465
rect 318 -5469 322 -5465
rect 339 -5469 343 -5465
rect 360 -5469 364 -5465
rect 381 -5469 385 -5465
rect 401 -5469 405 -5465
rect 203 -5525 207 -5521
rect 466 -5469 470 -5465
rect 209 -5532 213 -5528
rect 267 -5525 271 -5521
rect 309 -5532 313 -5528
rect 327 -5525 331 -5521
rect 369 -5517 373 -5513
rect 369 -5525 373 -5521
rect 351 -5539 355 -5535
rect 251 -5546 255 -5542
rect 293 -5546 297 -5542
rect 407 -5517 411 -5513
rect 393 -5532 397 -5528
rect 218 -5561 222 -5557
rect 235 -5561 239 -5557
rect 276 -5561 280 -5557
rect 318 -5561 322 -5557
rect 360 -5561 364 -5557
rect 401 -5561 405 -5557
rect 218 -5586 222 -5582
rect 235 -5586 239 -5582
rect 255 -5586 259 -5582
rect 276 -5586 280 -5582
rect 297 -5586 301 -5582
rect 318 -5586 322 -5582
rect 339 -5586 343 -5582
rect 360 -5586 364 -5582
rect 381 -5586 385 -5582
rect 401 -5586 405 -5582
rect 209 -5649 213 -5645
rect 267 -5642 271 -5638
rect 309 -5649 313 -5645
rect 327 -5642 331 -5638
rect 369 -5634 373 -5630
rect 369 -5642 373 -5638
rect 351 -5656 355 -5652
rect 251 -5663 255 -5659
rect 293 -5663 297 -5659
rect 393 -5649 397 -5645
rect 218 -5678 222 -5674
rect 235 -5678 239 -5674
rect 276 -5678 280 -5674
rect 318 -5678 322 -5674
rect 360 -5678 364 -5674
rect 401 -5678 405 -5674
rect 209 -5703 213 -5699
rect 226 -5703 230 -5699
rect 474 -5518 478 -5514
rect 466 -5561 470 -5557
rect 407 -5735 411 -5731
rect 235 -5756 239 -5752
rect 547 -5756 551 -5752
rect 226 -5795 230 -5791
rect 218 -5822 222 -5818
rect 244 -5822 248 -5818
rect 261 -5822 265 -5818
rect 301 -5822 305 -5818
rect 322 -5822 326 -5818
rect 339 -5822 343 -5818
rect 379 -5822 383 -5818
rect 403 -5822 407 -5818
rect 440 -5822 444 -5818
rect 197 -5862 201 -5858
rect 209 -5855 213 -5851
rect 191 -5877 195 -5873
rect 227 -5848 231 -5844
rect 253 -5870 257 -5866
rect 235 -5877 239 -5873
rect 279 -5862 283 -5858
rect 331 -5855 335 -5851
rect 261 -5899 265 -5895
rect 297 -5899 301 -5895
rect 357 -5870 361 -5866
rect 339 -5899 343 -5895
rect 375 -5899 379 -5895
rect 449 -5862 453 -5858
rect 455 -5870 459 -5866
rect 218 -5914 222 -5910
rect 244 -5914 248 -5910
rect 287 -5914 291 -5910
rect 322 -5914 326 -5910
rect 366 -5914 370 -5910
rect 383 -5914 387 -5910
rect 419 -5914 423 -5910
rect 440 -5914 444 -5910
rect -1270 -5924 -1266 -5920
rect -1162 -5924 -1158 -5920
rect -941 -5921 -937 -5917
rect -689 -5921 -685 -5917
rect -583 -5921 -579 -5917
rect -331 -5921 -327 -5917
rect -225 -5921 -221 -5917
rect 27 -5921 31 -5917
rect 763 -5022 767 -5018
rect 591 -5043 595 -5039
rect 945 -5043 949 -5039
rect 582 -5082 586 -5078
rect 574 -5109 578 -5105
rect 600 -5109 604 -5105
rect 617 -5109 621 -5105
rect 657 -5109 661 -5105
rect 678 -5109 682 -5105
rect 695 -5109 699 -5105
rect 735 -5109 739 -5105
rect 759 -5109 763 -5105
rect 796 -5109 800 -5105
rect 565 -5142 569 -5138
rect 583 -5135 587 -5131
rect 609 -5157 613 -5153
rect 591 -5164 595 -5160
rect 635 -5149 639 -5145
rect 687 -5142 691 -5138
rect 617 -5186 621 -5182
rect 653 -5186 657 -5182
rect 713 -5157 717 -5153
rect 695 -5186 699 -5182
rect 731 -5186 735 -5182
rect 805 -5149 809 -5145
rect 811 -5157 815 -5153
rect 574 -5201 578 -5197
rect 600 -5201 604 -5197
rect 643 -5201 647 -5197
rect 678 -5201 682 -5197
rect 722 -5201 726 -5197
rect 739 -5201 743 -5197
rect 775 -5201 779 -5197
rect 796 -5201 800 -5197
rect 1201 -4160 1205 -4156
rect 1209 -4205 1213 -4201
rect 1201 -4252 1205 -4248
rect 1201 -4271 1205 -4267
rect 1161 -4303 1165 -4299
rect 989 -4324 993 -4320
rect 1209 -4320 1213 -4316
rect 1303 -4324 1307 -4320
rect 980 -4363 984 -4359
rect 1201 -4363 1205 -4359
rect 972 -4390 976 -4386
rect 998 -4390 1002 -4386
rect 1015 -4390 1019 -4386
rect 1055 -4390 1059 -4386
rect 1076 -4390 1080 -4386
rect 1093 -4390 1097 -4386
rect 1133 -4390 1137 -4386
rect 1157 -4390 1161 -4386
rect 1194 -4390 1198 -4386
rect 963 -4423 967 -4419
rect 981 -4416 985 -4412
rect 1007 -4438 1011 -4434
rect 989 -4445 993 -4441
rect 1033 -4430 1037 -4426
rect 1085 -4423 1089 -4419
rect 1015 -4467 1019 -4463
rect 1051 -4467 1055 -4463
rect 1111 -4438 1115 -4434
rect 1093 -4467 1097 -4463
rect 1129 -4467 1133 -4463
rect 1203 -4428 1207 -4424
rect 1303 -4430 1307 -4426
rect 1209 -4438 1213 -4434
rect 972 -4482 976 -4478
rect 998 -4482 1002 -4478
rect 1041 -4482 1045 -4478
rect 1076 -4482 1080 -4478
rect 1120 -4482 1124 -4478
rect 1137 -4482 1141 -4478
rect 1173 -4482 1177 -4478
rect 1194 -4482 1198 -4478
rect 1519 -3458 1523 -3454
rect 1347 -3479 1351 -3475
rect 1338 -3518 1342 -3514
rect 1330 -3550 1334 -3546
rect 1356 -3550 1360 -3546
rect 1373 -3550 1377 -3546
rect 1413 -3550 1417 -3546
rect 1434 -3550 1438 -3546
rect 1451 -3550 1455 -3546
rect 1491 -3550 1495 -3546
rect 1515 -3550 1519 -3546
rect 1552 -3550 1556 -3546
rect 1321 -3583 1325 -3579
rect 1339 -3576 1343 -3572
rect 1365 -3598 1369 -3594
rect 1347 -3605 1351 -3601
rect 1391 -3590 1395 -3586
rect 1443 -3583 1447 -3579
rect 1373 -3627 1377 -3623
rect 1409 -3627 1413 -3623
rect 1469 -3598 1473 -3594
rect 1451 -3627 1455 -3623
rect 1487 -3627 1491 -3623
rect 1330 -3642 1334 -3638
rect 1356 -3642 1360 -3638
rect 1399 -3642 1403 -3638
rect 1434 -3642 1438 -3638
rect 1478 -3642 1482 -3638
rect 1495 -3642 1499 -3638
rect 1531 -3642 1535 -3638
rect 1552 -3642 1556 -3638
rect 1567 -3598 1571 -3594
rect 1567 -3649 1571 -3645
rect 1561 -3656 1565 -3652
rect 1330 -3911 1334 -3907
rect 1347 -3911 1351 -3907
rect 1367 -3911 1371 -3907
rect 1388 -3911 1392 -3907
rect 1409 -3911 1413 -3907
rect 1430 -3911 1434 -3907
rect 1451 -3911 1455 -3907
rect 1472 -3911 1476 -3907
rect 1493 -3911 1497 -3907
rect 1513 -3911 1517 -3907
rect 1321 -3974 1325 -3970
rect 1379 -3967 1383 -3963
rect 1421 -3974 1425 -3970
rect 1439 -3967 1443 -3963
rect 1481 -3959 1485 -3955
rect 1481 -3967 1485 -3963
rect 1463 -3981 1467 -3977
rect 1363 -3988 1367 -3984
rect 1405 -3988 1409 -3984
rect 1519 -3959 1523 -3955
rect 1505 -3974 1509 -3970
rect 1330 -4003 1334 -3999
rect 1347 -4003 1351 -3999
rect 1388 -4003 1392 -3999
rect 1430 -4003 1434 -3999
rect 1472 -4003 1476 -3999
rect 1513 -4003 1517 -3999
rect 1519 -4010 1523 -4006
rect 1330 -4036 1334 -4032
rect 1347 -4036 1351 -4032
rect 1367 -4036 1371 -4032
rect 1388 -4036 1392 -4032
rect 1409 -4036 1413 -4032
rect 1430 -4036 1434 -4032
rect 1451 -4036 1455 -4032
rect 1472 -4036 1476 -4032
rect 1493 -4036 1497 -4032
rect 1513 -4036 1517 -4032
rect 1315 -4092 1319 -4088
rect 1321 -4099 1325 -4095
rect 1379 -4092 1383 -4088
rect 1421 -4099 1425 -4095
rect 1439 -4092 1443 -4088
rect 1481 -4084 1485 -4080
rect 1481 -4092 1485 -4088
rect 1463 -4106 1467 -4102
rect 1363 -4113 1367 -4109
rect 1405 -4113 1409 -4109
rect 1519 -4084 1523 -4080
rect 1505 -4099 1509 -4095
rect 1330 -4128 1334 -4124
rect 1347 -4128 1351 -4124
rect 1388 -4128 1392 -4124
rect 1430 -4128 1434 -4124
rect 1472 -4128 1476 -4124
rect 1513 -4128 1517 -4124
rect 1321 -4271 1325 -4267
rect 1338 -4271 1342 -4267
rect 1309 -4445 1313 -4441
rect 1209 -4496 1213 -4492
rect 1309 -4496 1313 -4492
rect 972 -4634 976 -4630
rect 989 -4634 993 -4630
rect 1009 -4634 1013 -4630
rect 1030 -4634 1034 -4630
rect 1051 -4634 1055 -4630
rect 1072 -4634 1076 -4630
rect 1093 -4634 1097 -4630
rect 1114 -4634 1118 -4630
rect 1135 -4634 1139 -4630
rect 1155 -4634 1159 -4630
rect 963 -4697 967 -4693
rect 1021 -4690 1025 -4686
rect 1063 -4697 1067 -4693
rect 1081 -4690 1085 -4686
rect 1123 -4682 1127 -4678
rect 1123 -4690 1127 -4686
rect 1105 -4704 1109 -4700
rect 1005 -4711 1009 -4707
rect 1047 -4711 1051 -4707
rect 1161 -4682 1165 -4678
rect 1147 -4697 1151 -4693
rect 972 -4726 976 -4722
rect 989 -4726 993 -4722
rect 1030 -4726 1034 -4722
rect 1072 -4726 1076 -4722
rect 1114 -4726 1118 -4722
rect 1155 -4726 1159 -4722
rect 1309 -4690 1313 -4686
rect 1161 -4733 1165 -4729
rect 1309 -4733 1313 -4729
rect 972 -4755 976 -4751
rect 989 -4755 993 -4751
rect 1009 -4755 1013 -4751
rect 1030 -4755 1034 -4751
rect 1051 -4755 1055 -4751
rect 1072 -4755 1076 -4751
rect 1093 -4755 1097 -4751
rect 1114 -4755 1118 -4751
rect 1135 -4755 1139 -4751
rect 1155 -4755 1159 -4751
rect 957 -4811 961 -4807
rect 963 -4818 967 -4814
rect 1021 -4811 1025 -4807
rect 1063 -4818 1067 -4814
rect 1081 -4811 1085 -4807
rect 1123 -4803 1127 -4799
rect 1123 -4811 1127 -4807
rect 1105 -4825 1109 -4821
rect 1005 -4832 1009 -4828
rect 1047 -4832 1051 -4828
rect 1161 -4803 1165 -4799
rect 1147 -4818 1151 -4814
rect 972 -4847 976 -4843
rect 989 -4847 993 -4843
rect 1030 -4847 1034 -4843
rect 1072 -4847 1076 -4843
rect 1114 -4847 1118 -4843
rect 1155 -4847 1159 -4843
rect 963 -4990 967 -4986
rect 980 -4990 984 -4986
rect 951 -5149 955 -5145
rect 945 -5164 949 -5160
rect 811 -5208 815 -5204
rect 951 -5208 955 -5204
rect 574 -5349 578 -5345
rect 591 -5349 595 -5345
rect 611 -5349 615 -5345
rect 632 -5349 636 -5345
rect 653 -5349 657 -5345
rect 674 -5349 678 -5345
rect 695 -5349 699 -5345
rect 716 -5349 720 -5345
rect 737 -5349 741 -5345
rect 757 -5349 761 -5345
rect 867 -5349 871 -5345
rect 565 -5412 569 -5408
rect 623 -5405 627 -5401
rect 665 -5412 669 -5408
rect 683 -5405 687 -5401
rect 725 -5397 729 -5393
rect 725 -5405 729 -5401
rect 707 -5419 711 -5415
rect 607 -5426 611 -5422
rect 649 -5426 653 -5422
rect 763 -5397 767 -5393
rect 749 -5412 753 -5408
rect 574 -5441 578 -5437
rect 591 -5441 595 -5437
rect 632 -5441 636 -5437
rect 674 -5441 678 -5437
rect 716 -5441 720 -5437
rect 757 -5441 761 -5437
rect 875 -5399 879 -5395
rect 951 -5405 955 -5401
rect 867 -5441 871 -5437
rect 763 -5450 767 -5446
rect 951 -5449 955 -5445
rect 574 -5469 578 -5465
rect 591 -5469 595 -5465
rect 611 -5469 615 -5465
rect 632 -5469 636 -5465
rect 653 -5469 657 -5465
rect 674 -5469 678 -5465
rect 695 -5469 699 -5465
rect 716 -5469 720 -5465
rect 737 -5469 741 -5465
rect 757 -5469 761 -5465
rect 559 -5525 563 -5521
rect 565 -5532 569 -5528
rect 623 -5525 627 -5521
rect 665 -5532 669 -5528
rect 683 -5525 687 -5521
rect 725 -5517 729 -5513
rect 725 -5525 729 -5521
rect 707 -5539 711 -5535
rect 607 -5546 611 -5542
rect 649 -5546 653 -5542
rect 769 -5517 773 -5513
rect 749 -5532 753 -5528
rect 574 -5561 578 -5557
rect 591 -5561 595 -5557
rect 632 -5561 636 -5557
rect 674 -5561 678 -5557
rect 716 -5561 720 -5557
rect 757 -5561 761 -5557
rect 574 -5586 578 -5582
rect 591 -5586 595 -5582
rect 611 -5586 615 -5582
rect 632 -5586 636 -5582
rect 653 -5586 657 -5582
rect 674 -5586 678 -5582
rect 695 -5586 699 -5582
rect 716 -5586 720 -5582
rect 737 -5586 741 -5582
rect 757 -5586 761 -5582
rect 565 -5649 569 -5645
rect 623 -5642 627 -5638
rect 665 -5649 669 -5645
rect 683 -5642 687 -5638
rect 725 -5634 729 -5630
rect 725 -5642 729 -5638
rect 707 -5656 711 -5652
rect 607 -5663 611 -5659
rect 649 -5663 653 -5659
rect 763 -5634 767 -5630
rect 749 -5649 753 -5645
rect 574 -5678 578 -5674
rect 591 -5678 595 -5674
rect 632 -5678 636 -5674
rect 674 -5678 678 -5674
rect 716 -5678 720 -5674
rect 757 -5678 761 -5674
rect 565 -5703 569 -5699
rect 582 -5703 586 -5699
rect 769 -5735 773 -5731
rect 763 -5743 767 -5739
rect 591 -5756 595 -5752
rect 945 -5756 949 -5752
rect 582 -5795 586 -5791
rect 574 -5822 578 -5818
rect 600 -5822 604 -5818
rect 617 -5822 621 -5818
rect 657 -5822 661 -5818
rect 678 -5822 682 -5818
rect 695 -5822 699 -5818
rect 735 -5822 739 -5818
rect 759 -5822 763 -5818
rect 796 -5822 800 -5818
rect 553 -5862 557 -5858
rect 565 -5855 569 -5851
rect 547 -5877 551 -5873
rect 583 -5848 587 -5844
rect 609 -5870 613 -5866
rect 591 -5877 595 -5873
rect 635 -5862 639 -5858
rect 687 -5855 691 -5851
rect 617 -5899 621 -5895
rect 653 -5899 657 -5895
rect 713 -5870 717 -5866
rect 695 -5899 699 -5895
rect 731 -5899 735 -5895
rect 805 -5862 809 -5858
rect 811 -5870 815 -5866
rect 574 -5914 578 -5910
rect 600 -5914 604 -5910
rect 643 -5914 647 -5910
rect 678 -5914 682 -5910
rect 722 -5914 726 -5910
rect 739 -5914 743 -5910
rect 775 -5914 779 -5910
rect 796 -5914 800 -5910
rect 1161 -5022 1165 -5018
rect 989 -5043 993 -5039
rect 1303 -5043 1307 -5039
rect 980 -5082 984 -5078
rect 972 -5109 976 -5105
rect 998 -5109 1002 -5105
rect 1015 -5109 1019 -5105
rect 1055 -5109 1059 -5105
rect 1076 -5109 1080 -5105
rect 1093 -5109 1097 -5105
rect 1133 -5109 1137 -5105
rect 1157 -5109 1161 -5105
rect 1194 -5109 1198 -5105
rect 963 -5142 967 -5138
rect 981 -5135 985 -5131
rect 1007 -5157 1011 -5153
rect 989 -5164 993 -5160
rect 1033 -5149 1037 -5145
rect 1085 -5142 1089 -5138
rect 1015 -5186 1019 -5182
rect 1051 -5186 1055 -5182
rect 1111 -5157 1115 -5153
rect 1093 -5186 1097 -5182
rect 1129 -5186 1133 -5182
rect 1203 -5147 1207 -5143
rect 1303 -5149 1307 -5145
rect 1209 -5157 1213 -5153
rect 972 -5201 976 -5197
rect 998 -5201 1002 -5197
rect 1041 -5201 1045 -5197
rect 1076 -5201 1080 -5197
rect 1120 -5201 1124 -5197
rect 1137 -5201 1141 -5197
rect 1173 -5201 1177 -5197
rect 1194 -5201 1198 -5197
rect 1519 -4303 1523 -4299
rect 1347 -4324 1351 -4320
rect 1338 -4363 1342 -4359
rect 1330 -4390 1334 -4386
rect 1356 -4390 1360 -4386
rect 1373 -4390 1377 -4386
rect 1413 -4390 1417 -4386
rect 1434 -4390 1438 -4386
rect 1451 -4390 1455 -4386
rect 1491 -4390 1495 -4386
rect 1515 -4390 1519 -4386
rect 1552 -4390 1556 -4386
rect 1321 -4423 1325 -4419
rect 1339 -4416 1343 -4412
rect 1365 -4438 1369 -4434
rect 1347 -4445 1351 -4441
rect 1391 -4430 1395 -4426
rect 1443 -4423 1447 -4419
rect 1373 -4467 1377 -4463
rect 1409 -4467 1413 -4463
rect 1469 -4438 1473 -4434
rect 1451 -4467 1455 -4463
rect 1487 -4467 1491 -4463
rect 1330 -4482 1334 -4478
rect 1356 -4482 1360 -4478
rect 1399 -4482 1403 -4478
rect 1434 -4482 1438 -4478
rect 1478 -4482 1482 -4478
rect 1495 -4482 1499 -4478
rect 1531 -4482 1535 -4478
rect 1552 -4482 1556 -4478
rect 1567 -4438 1571 -4434
rect 1567 -4489 1571 -4485
rect 1561 -4496 1565 -4492
rect 1330 -4634 1334 -4630
rect 1347 -4634 1351 -4630
rect 1367 -4634 1371 -4630
rect 1388 -4634 1392 -4630
rect 1409 -4634 1413 -4630
rect 1430 -4634 1434 -4630
rect 1451 -4634 1455 -4630
rect 1472 -4634 1476 -4630
rect 1493 -4634 1497 -4630
rect 1513 -4634 1517 -4630
rect 1321 -4697 1325 -4693
rect 1379 -4690 1383 -4686
rect 1421 -4697 1425 -4693
rect 1439 -4690 1443 -4686
rect 1481 -4682 1485 -4678
rect 1481 -4690 1485 -4686
rect 1463 -4704 1467 -4700
rect 1363 -4711 1367 -4707
rect 1405 -4711 1409 -4707
rect 1519 -4682 1523 -4678
rect 1505 -4697 1509 -4693
rect 1330 -4726 1334 -4722
rect 1347 -4726 1351 -4722
rect 1388 -4726 1392 -4722
rect 1430 -4726 1434 -4722
rect 1472 -4726 1476 -4722
rect 1513 -4726 1517 -4722
rect 1519 -4733 1523 -4729
rect 1330 -4755 1334 -4751
rect 1347 -4755 1351 -4751
rect 1367 -4755 1371 -4751
rect 1388 -4755 1392 -4751
rect 1409 -4755 1413 -4751
rect 1430 -4755 1434 -4751
rect 1451 -4755 1455 -4751
rect 1472 -4755 1476 -4751
rect 1493 -4755 1497 -4751
rect 1513 -4755 1517 -4751
rect 1315 -4811 1319 -4807
rect 1321 -4818 1325 -4814
rect 1379 -4811 1383 -4807
rect 1421 -4818 1425 -4814
rect 1439 -4811 1443 -4807
rect 1481 -4803 1485 -4799
rect 1481 -4811 1485 -4807
rect 1463 -4825 1467 -4821
rect 1363 -4832 1367 -4828
rect 1405 -4832 1409 -4828
rect 1519 -4803 1523 -4799
rect 1505 -4818 1509 -4814
rect 1330 -4847 1334 -4843
rect 1347 -4847 1351 -4843
rect 1388 -4847 1392 -4843
rect 1430 -4847 1434 -4843
rect 1472 -4847 1476 -4843
rect 1513 -4847 1517 -4843
rect 1321 -4990 1325 -4986
rect 1338 -4990 1342 -4986
rect 1309 -5164 1313 -5160
rect 1209 -5215 1213 -5211
rect 1309 -5215 1313 -5211
rect 972 -5349 976 -5345
rect 989 -5349 993 -5345
rect 1009 -5349 1013 -5345
rect 1030 -5349 1034 -5345
rect 1051 -5349 1055 -5345
rect 1072 -5349 1076 -5345
rect 1093 -5349 1097 -5345
rect 1114 -5349 1118 -5345
rect 1135 -5349 1139 -5345
rect 1155 -5349 1159 -5345
rect 1210 -5349 1214 -5345
rect 963 -5412 967 -5408
rect 1021 -5405 1025 -5401
rect 1063 -5412 1067 -5408
rect 1081 -5405 1085 -5401
rect 1123 -5397 1127 -5393
rect 1123 -5405 1127 -5401
rect 1105 -5419 1109 -5415
rect 1005 -5426 1009 -5422
rect 1047 -5426 1051 -5422
rect 1161 -5397 1165 -5393
rect 1147 -5412 1151 -5408
rect 972 -5441 976 -5437
rect 989 -5441 993 -5437
rect 1030 -5441 1034 -5437
rect 1072 -5441 1076 -5437
rect 1114 -5441 1118 -5437
rect 1155 -5441 1159 -5437
rect 1218 -5403 1222 -5399
rect 1309 -5405 1313 -5401
rect 1210 -5441 1214 -5437
rect 1161 -5449 1165 -5445
rect 1309 -5448 1313 -5444
rect 972 -5469 976 -5465
rect 989 -5469 993 -5465
rect 1009 -5469 1013 -5465
rect 1030 -5469 1034 -5465
rect 1051 -5469 1055 -5465
rect 1072 -5469 1076 -5465
rect 1093 -5469 1097 -5465
rect 1114 -5469 1118 -5465
rect 1135 -5469 1139 -5465
rect 1155 -5469 1159 -5465
rect 957 -5525 961 -5521
rect 1210 -5469 1214 -5465
rect 963 -5532 967 -5528
rect 1021 -5525 1025 -5521
rect 1063 -5532 1067 -5528
rect 1081 -5525 1085 -5521
rect 1123 -5517 1127 -5513
rect 1123 -5525 1127 -5521
rect 1105 -5539 1109 -5535
rect 1005 -5546 1009 -5542
rect 1047 -5546 1051 -5542
rect 1161 -5517 1165 -5513
rect 1147 -5532 1151 -5528
rect 972 -5561 976 -5557
rect 989 -5561 993 -5557
rect 1030 -5561 1034 -5557
rect 1072 -5561 1076 -5557
rect 1114 -5561 1118 -5557
rect 1155 -5561 1159 -5557
rect 963 -5703 967 -5699
rect 980 -5703 984 -5699
rect 1218 -5518 1222 -5514
rect 1210 -5561 1214 -5557
rect 1161 -5735 1165 -5731
rect 989 -5756 993 -5752
rect 1303 -5756 1307 -5752
rect 980 -5795 984 -5791
rect 972 -5822 976 -5818
rect 998 -5822 1002 -5818
rect 1015 -5822 1019 -5818
rect 1055 -5822 1059 -5818
rect 1076 -5822 1080 -5818
rect 1093 -5822 1097 -5818
rect 1133 -5822 1137 -5818
rect 1157 -5822 1161 -5818
rect 1194 -5822 1198 -5818
rect 951 -5862 955 -5858
rect 963 -5855 967 -5851
rect 945 -5877 949 -5873
rect 981 -5848 985 -5844
rect 1007 -5870 1011 -5866
rect 989 -5877 993 -5873
rect 1033 -5862 1037 -5858
rect 1085 -5855 1089 -5851
rect 1015 -5899 1019 -5895
rect 1051 -5899 1055 -5895
rect 1111 -5870 1115 -5866
rect 1093 -5899 1097 -5895
rect 1129 -5899 1133 -5895
rect 1203 -5860 1207 -5856
rect 1303 -5862 1307 -5858
rect 1209 -5870 1213 -5866
rect 972 -5914 976 -5910
rect 998 -5914 1002 -5910
rect 1041 -5914 1045 -5910
rect 1076 -5914 1080 -5910
rect 1120 -5914 1124 -5910
rect 1137 -5914 1141 -5910
rect 1173 -5914 1177 -5910
rect 1194 -5914 1198 -5910
rect 1519 -5022 1523 -5018
rect 1347 -5043 1351 -5039
rect 1338 -5082 1342 -5078
rect 1330 -5109 1334 -5105
rect 1356 -5109 1360 -5105
rect 1373 -5109 1377 -5105
rect 1413 -5109 1417 -5105
rect 1434 -5109 1438 -5105
rect 1451 -5109 1455 -5105
rect 1491 -5109 1495 -5105
rect 1515 -5109 1519 -5105
rect 1552 -5109 1556 -5105
rect 1321 -5142 1325 -5138
rect 1339 -5135 1343 -5131
rect 1365 -5157 1369 -5153
rect 1347 -5164 1351 -5160
rect 1391 -5149 1395 -5145
rect 1443 -5142 1447 -5138
rect 1373 -5186 1377 -5182
rect 1409 -5186 1413 -5182
rect 1469 -5157 1473 -5153
rect 1451 -5186 1455 -5182
rect 1487 -5186 1491 -5182
rect 1330 -5201 1334 -5197
rect 1356 -5201 1360 -5197
rect 1399 -5201 1403 -5197
rect 1434 -5201 1438 -5197
rect 1478 -5201 1482 -5197
rect 1495 -5201 1499 -5197
rect 1531 -5201 1535 -5197
rect 1552 -5201 1556 -5197
rect 1567 -5157 1571 -5153
rect 1567 -5208 1571 -5204
rect 1561 -5215 1565 -5211
rect 1330 -5349 1334 -5345
rect 1347 -5349 1351 -5345
rect 1367 -5349 1371 -5345
rect 1388 -5349 1392 -5345
rect 1409 -5349 1413 -5345
rect 1430 -5349 1434 -5345
rect 1451 -5349 1455 -5345
rect 1472 -5349 1476 -5345
rect 1493 -5349 1497 -5345
rect 1513 -5349 1517 -5345
rect 1321 -5412 1325 -5408
rect 1379 -5405 1383 -5401
rect 1421 -5412 1425 -5408
rect 1439 -5405 1443 -5401
rect 1481 -5397 1485 -5393
rect 1481 -5405 1485 -5401
rect 1463 -5419 1467 -5415
rect 1363 -5426 1367 -5422
rect 1405 -5426 1409 -5422
rect 1519 -5397 1523 -5393
rect 1505 -5412 1509 -5408
rect 1330 -5441 1334 -5437
rect 1347 -5441 1351 -5437
rect 1388 -5441 1392 -5437
rect 1430 -5441 1434 -5437
rect 1472 -5441 1476 -5437
rect 1513 -5441 1517 -5437
rect 1519 -5448 1523 -5444
rect 1330 -5469 1334 -5465
rect 1347 -5469 1351 -5465
rect 1367 -5469 1371 -5465
rect 1388 -5469 1392 -5465
rect 1409 -5469 1413 -5465
rect 1430 -5469 1434 -5465
rect 1451 -5469 1455 -5465
rect 1472 -5469 1476 -5465
rect 1493 -5469 1497 -5465
rect 1513 -5469 1517 -5465
rect 1315 -5525 1319 -5521
rect 1321 -5532 1325 -5528
rect 1379 -5525 1383 -5521
rect 1421 -5532 1425 -5528
rect 1439 -5525 1443 -5521
rect 1481 -5517 1485 -5513
rect 1481 -5525 1485 -5521
rect 1463 -5539 1467 -5535
rect 1363 -5546 1367 -5542
rect 1405 -5546 1409 -5542
rect 1519 -5517 1523 -5513
rect 1505 -5532 1509 -5528
rect 1330 -5561 1334 -5557
rect 1347 -5561 1351 -5557
rect 1388 -5561 1392 -5557
rect 1430 -5561 1434 -5557
rect 1472 -5561 1476 -5557
rect 1513 -5561 1517 -5557
rect 1321 -5703 1325 -5699
rect 1338 -5703 1342 -5699
rect 1519 -5735 1523 -5731
rect 1347 -5756 1351 -5752
rect 1338 -5795 1342 -5791
rect 1330 -5822 1334 -5818
rect 1356 -5822 1360 -5818
rect 1373 -5822 1377 -5818
rect 1413 -5822 1417 -5818
rect 1434 -5822 1438 -5818
rect 1451 -5822 1455 -5818
rect 1491 -5822 1495 -5818
rect 1515 -5822 1519 -5818
rect 1552 -5822 1556 -5818
rect 1309 -5877 1313 -5873
rect 1321 -5855 1325 -5851
rect 1339 -5848 1343 -5844
rect 1365 -5870 1369 -5866
rect 1347 -5877 1351 -5873
rect 1391 -5862 1395 -5858
rect 1443 -5855 1447 -5851
rect 1373 -5899 1377 -5895
rect 1409 -5899 1413 -5895
rect 1469 -5870 1473 -5866
rect 1451 -5899 1455 -5895
rect 1487 -5899 1491 -5895
rect 1330 -5914 1334 -5910
rect 1356 -5914 1360 -5910
rect 1399 -5914 1403 -5910
rect 1434 -5914 1438 -5910
rect 1478 -5914 1482 -5910
rect 1495 -5914 1499 -5910
rect 1531 -5914 1535 -5910
rect 1552 -5914 1556 -5910
rect -1255 -5945 -1251 -5941
rect -1238 -5945 -1234 -5941
rect -1218 -5945 -1214 -5941
rect -1197 -5945 -1193 -5941
rect -1176 -5945 -1172 -5941
rect -1155 -5945 -1151 -5941
rect -1134 -5945 -1130 -5941
rect -1113 -5945 -1109 -5941
rect -1092 -5945 -1088 -5941
rect -1072 -5945 -1068 -5941
rect -1270 -6001 -1266 -5997
rect -1264 -6008 -1260 -6004
rect -1206 -6001 -1202 -5997
rect -1164 -6008 -1160 -6004
rect -1146 -6001 -1142 -5997
rect -1104 -5993 -1100 -5989
rect -1104 -6001 -1100 -5997
rect -1122 -6015 -1118 -6011
rect -1222 -6022 -1218 -6018
rect -1180 -6022 -1176 -6018
rect -926 -5945 -922 -5941
rect -909 -5945 -905 -5941
rect -889 -5945 -885 -5941
rect -868 -5945 -864 -5941
rect -847 -5945 -843 -5941
rect -826 -5945 -822 -5941
rect -805 -5945 -801 -5941
rect -784 -5945 -780 -5941
rect -763 -5945 -759 -5941
rect -743 -5945 -739 -5941
rect -941 -6001 -937 -5997
rect -1080 -6008 -1076 -6004
rect -935 -6008 -931 -6004
rect -877 -6001 -873 -5997
rect -835 -6008 -831 -6004
rect -817 -6001 -813 -5997
rect -775 -5993 -771 -5989
rect -775 -6001 -771 -5997
rect -793 -6015 -789 -6011
rect -893 -6022 -889 -6018
rect -851 -6022 -847 -6018
rect -568 -5945 -564 -5941
rect -551 -5945 -547 -5941
rect -531 -5945 -527 -5941
rect -510 -5945 -506 -5941
rect -489 -5945 -485 -5941
rect -468 -5945 -464 -5941
rect -447 -5945 -443 -5941
rect -426 -5945 -422 -5941
rect -405 -5945 -401 -5941
rect -385 -5945 -381 -5941
rect -583 -6001 -579 -5997
rect -751 -6008 -747 -6004
rect -577 -6008 -573 -6004
rect -519 -6001 -515 -5997
rect -477 -6008 -473 -6004
rect -459 -6001 -455 -5997
rect -417 -5993 -413 -5989
rect -417 -6001 -413 -5997
rect -435 -6015 -431 -6011
rect -535 -6022 -531 -6018
rect -493 -6022 -489 -6018
rect 203 -5922 207 -5918
rect 455 -5922 459 -5918
rect 559 -5921 563 -5917
rect 811 -5921 815 -5917
rect 957 -5921 961 -5917
rect 1209 -5921 1213 -5917
rect 1315 -5921 1319 -5917
rect -210 -5945 -206 -5941
rect -193 -5945 -189 -5941
rect -173 -5945 -169 -5941
rect -152 -5945 -148 -5941
rect -131 -5945 -127 -5941
rect -110 -5945 -106 -5941
rect -89 -5945 -85 -5941
rect -68 -5945 -64 -5941
rect -47 -5945 -43 -5941
rect -27 -5945 -23 -5941
rect -225 -6001 -221 -5997
rect -393 -6008 -389 -6004
rect -219 -6008 -215 -6004
rect -161 -6001 -157 -5997
rect -119 -6008 -115 -6004
rect -101 -6001 -97 -5997
rect -59 -5993 -55 -5989
rect -59 -6001 -55 -5997
rect -77 -6015 -73 -6011
rect -177 -6022 -173 -6018
rect -135 -6022 -131 -6018
rect 218 -5945 222 -5941
rect 235 -5945 239 -5941
rect 255 -5945 259 -5941
rect 276 -5945 280 -5941
rect 297 -5945 301 -5941
rect 318 -5945 322 -5941
rect 339 -5945 343 -5941
rect 360 -5945 364 -5941
rect 381 -5945 385 -5941
rect 401 -5945 405 -5941
rect 203 -6001 207 -5997
rect -35 -6008 -31 -6004
rect 209 -6008 213 -6004
rect 267 -6001 271 -5997
rect 309 -6008 313 -6004
rect 327 -6001 331 -5997
rect 369 -5993 373 -5989
rect 369 -6001 373 -5997
rect 351 -6015 355 -6011
rect 251 -6022 255 -6018
rect 293 -6022 297 -6018
rect 574 -5945 578 -5941
rect 591 -5945 595 -5941
rect 611 -5945 615 -5941
rect 632 -5945 636 -5941
rect 653 -5945 657 -5941
rect 674 -5945 678 -5941
rect 695 -5945 699 -5941
rect 716 -5945 720 -5941
rect 737 -5945 741 -5941
rect 757 -5945 761 -5941
rect 559 -6001 563 -5997
rect 393 -6008 397 -6004
rect 565 -6008 569 -6004
rect 623 -6001 627 -5997
rect 665 -6008 669 -6004
rect 683 -6001 687 -5997
rect 725 -5993 729 -5989
rect 725 -6001 729 -5997
rect 707 -6015 711 -6011
rect 607 -6022 611 -6018
rect 649 -6022 653 -6018
rect 972 -5945 976 -5941
rect 989 -5945 993 -5941
rect 1009 -5945 1013 -5941
rect 1030 -5945 1034 -5941
rect 1051 -5945 1055 -5941
rect 1072 -5945 1076 -5941
rect 1093 -5945 1097 -5941
rect 1114 -5945 1118 -5941
rect 1135 -5945 1139 -5941
rect 1155 -5945 1159 -5941
rect 957 -6001 961 -5997
rect 749 -6008 753 -6004
rect 963 -6008 967 -6004
rect 1021 -6001 1025 -5997
rect 1063 -6008 1067 -6004
rect 1081 -6001 1085 -5997
rect 1123 -5993 1127 -5989
rect 1123 -6001 1127 -5997
rect 1105 -6015 1109 -6011
rect 1005 -6022 1009 -6018
rect 1047 -6022 1051 -6018
rect 1330 -5945 1334 -5941
rect 1347 -5945 1351 -5941
rect 1367 -5945 1371 -5941
rect 1388 -5945 1392 -5941
rect 1409 -5945 1413 -5941
rect 1430 -5945 1434 -5941
rect 1451 -5945 1455 -5941
rect 1472 -5945 1476 -5941
rect 1493 -5945 1497 -5941
rect 1513 -5945 1517 -5941
rect 1315 -6001 1319 -5997
rect 1147 -6008 1151 -6004
rect 1321 -6008 1325 -6004
rect 1379 -6001 1383 -5997
rect 1421 -6008 1425 -6004
rect 1439 -6001 1443 -5997
rect 1481 -5993 1485 -5989
rect 1481 -6001 1485 -5997
rect 1463 -6015 1467 -6011
rect 1363 -6022 1367 -6018
rect 1405 -6022 1409 -6018
rect 1505 -6008 1509 -6004
rect -1255 -6037 -1251 -6033
rect -1238 -6037 -1234 -6033
rect -1197 -6037 -1193 -6033
rect -1155 -6037 -1151 -6033
rect -1113 -6037 -1109 -6033
rect -1072 -6037 -1068 -6033
rect -926 -6037 -922 -6033
rect -909 -6037 -905 -6033
rect -868 -6037 -864 -6033
rect -826 -6037 -822 -6033
rect -784 -6037 -780 -6033
rect -743 -6037 -739 -6033
rect -568 -6037 -564 -6033
rect -551 -6037 -547 -6033
rect -510 -6037 -506 -6033
rect -468 -6037 -464 -6033
rect -426 -6037 -422 -6033
rect -385 -6037 -381 -6033
rect -210 -6037 -206 -6033
rect -193 -6037 -189 -6033
rect -152 -6037 -148 -6033
rect -110 -6037 -106 -6033
rect -68 -6037 -64 -6033
rect -27 -6037 -23 -6033
rect 218 -6037 222 -6033
rect 235 -6037 239 -6033
rect 276 -6037 280 -6033
rect 318 -6037 322 -6033
rect 360 -6037 364 -6033
rect 401 -6037 405 -6033
rect 574 -6037 578 -6033
rect 591 -6037 595 -6033
rect 632 -6037 636 -6033
rect 674 -6037 678 -6033
rect 716 -6037 720 -6033
rect 757 -6037 761 -6033
rect 972 -6037 976 -6033
rect 989 -6037 993 -6033
rect 1030 -6037 1034 -6033
rect 1072 -6037 1076 -6033
rect 1114 -6037 1118 -6033
rect 1155 -6037 1159 -6033
rect 1330 -6037 1334 -6033
rect 1347 -6037 1351 -6033
rect 1388 -6037 1392 -6033
rect 1430 -6037 1434 -6033
rect 1472 -6037 1476 -6033
rect 1513 -6037 1517 -6033
rect 1567 -5870 1571 -5866
rect 1567 -5921 1571 -5917
rect 1315 -6044 1319 -6040
rect 1561 -6044 1565 -6040
rect 1330 -6063 1334 -6059
rect 1347 -6063 1351 -6059
rect 1367 -6063 1371 -6059
rect 1388 -6063 1392 -6059
rect 1409 -6063 1413 -6059
rect 1430 -6063 1434 -6059
rect 1451 -6063 1455 -6059
rect 1472 -6063 1476 -6059
rect 1493 -6063 1497 -6059
rect 1513 -6063 1517 -6059
rect 1315 -6119 1319 -6115
rect 1321 -6126 1325 -6122
rect 1379 -6119 1383 -6115
rect 1421 -6126 1425 -6122
rect 1439 -6119 1443 -6115
rect 1481 -6111 1485 -6107
rect 1481 -6119 1485 -6115
rect 1463 -6133 1467 -6129
rect 1363 -6140 1367 -6136
rect 1405 -6140 1409 -6136
rect 1505 -6126 1509 -6122
rect 1330 -6155 1334 -6151
rect 1347 -6155 1351 -6151
rect 1388 -6155 1392 -6151
rect 1430 -6155 1434 -6151
rect 1472 -6155 1476 -6151
rect 1513 -6155 1517 -6151
<< m3contact >>
rect -1274 -1218 -1270 -1214
rect -956 -1218 -952 -1214
rect -587 -1218 -583 -1214
rect -240 -1218 -236 -1214
rect 198 -1218 202 -1214
rect 536 -1218 540 -1214
rect 952 -1218 956 -1214
rect -1265 -1571 -1261 -1567
rect -946 -1571 -942 -1567
rect -588 -1571 -584 -1567
rect -230 -1571 -226 -1567
rect 199 -1571 203 -1567
rect 553 -1571 557 -1567
rect 951 -1571 955 -1567
rect -1270 -1692 -1266 -1688
rect -941 -1692 -937 -1688
rect -588 -1692 -584 -1688
rect -230 -1692 -226 -1688
rect 199 -1692 203 -1688
rect 560 -1692 564 -1688
rect 951 -1692 955 -1688
rect 1311 -1692 1315 -1688
rect -1013 -1792 -1009 -1788
rect -316 -1792 -312 -1788
rect 480 -1792 484 -1788
rect 1219 -1792 1223 -1788
rect -1270 -1813 -1266 -1809
rect -946 -1813 -942 -1809
rect -588 -1813 -584 -1809
rect -230 -1813 -226 -1809
rect 199 -1813 203 -1809
rect 553 -1813 557 -1809
rect 951 -1813 955 -1809
rect 1309 -1813 1313 -1809
rect -1013 -1907 -1009 -1903
rect -657 -1907 -653 -1903
rect -316 -1907 -312 -1903
rect 480 -1907 484 -1903
rect 857 -1907 861 -1903
rect 1219 -1907 1223 -1903
rect -1273 -1928 -1269 -1924
rect -1284 -2303 -1280 -2299
rect -954 -2303 -950 -2299
rect -595 -2303 -591 -2299
rect -239 -2303 -235 -2299
rect 192 -2303 196 -2299
rect 543 -2303 547 -2299
rect -1284 -2434 -1280 -2430
rect -954 -2434 -950 -2430
rect -595 -2434 -591 -2430
rect -239 -2434 -235 -2430
rect 192 -2434 196 -2430
rect 543 -2434 547 -2430
rect 950 -2434 954 -2430
rect 1302 -2434 1306 -2430
rect 106 -2546 110 -2542
rect -1275 -2565 -1271 -2561
rect -942 -2565 -938 -2561
rect -586 -2565 -582 -2561
rect -228 -2565 -224 -2561
rect 198 -2565 202 -2561
rect 556 -2565 560 -2561
rect 944 -2565 948 -2561
rect 1313 -2565 1317 -2561
rect -1275 -2677 -1271 -2673
rect -942 -2677 -938 -2673
rect -1010 -3008 -1006 -3004
rect -656 -3007 -652 -3003
rect -313 -3009 -309 -3005
rect 488 -3007 492 -3003
rect 857 -3007 861 -3003
rect 1215 -3008 1219 -3004
rect -1267 -3028 -1263 -3024
rect -940 -3028 -936 -3024
rect -590 -3028 -586 -3024
rect -227 -3028 -223 -3024
rect 195 -3028 199 -3024
rect -1010 -3123 -1006 -3119
rect -313 -3124 -309 -3120
rect 488 -3123 492 -3119
rect 1215 -3123 1219 -3119
rect -1278 -3144 -1274 -3140
rect -940 -3144 -936 -3140
rect -584 -3144 -580 -3140
rect -225 -3144 -221 -3140
rect 201 -3144 205 -3140
rect 558 -3144 562 -3140
rect 954 -3144 958 -3140
rect 1314 -3144 1318 -3140
rect -1278 -3265 -1274 -3261
rect -940 -3265 -936 -3261
rect -584 -3265 -580 -3261
rect -225 -3265 -221 -3261
rect 201 -3265 205 -3261
rect 558 -3265 562 -3261
rect 954 -3265 958 -3261
rect 1314 -3265 1318 -3261
rect -1278 -3379 -1274 -3375
rect -940 -3379 -936 -3375
rect -584 -3379 -580 -3375
rect -1281 -3750 -1277 -3746
rect -940 -3750 -936 -3746
rect -580 -3750 -576 -3746
rect -225 -3750 -221 -3746
rect -1598 -3851 -1584 -3837
rect 92 -3846 96 -3842
rect -1272 -3981 -1268 -3977
rect -941 -3981 -937 -3977
rect -583 -3981 -579 -3977
rect -226 -3981 -222 -3977
rect 204 -3981 208 -3977
rect 560 -3981 564 -3977
rect 945 -3981 949 -3977
rect 1315 -3981 1319 -3977
rect -1272 -4106 -1268 -4102
rect -941 -4106 -937 -4102
rect -583 -4106 -579 -4102
rect -226 -4106 -222 -4102
rect 204 -4106 208 -4102
rect 560 -4106 564 -4102
rect 945 -4106 949 -4102
rect 1315 -4106 1319 -4102
rect -1013 -4205 -1009 -4201
rect -316 -4207 -312 -4203
rect 472 -4205 476 -4201
rect 1217 -4205 1221 -4201
rect -1272 -4230 -1268 -4226
rect -941 -4230 -937 -4226
rect -583 -4230 -579 -4226
rect -226 -4230 -222 -4226
rect -1013 -4320 -1009 -4316
rect -657 -4321 -653 -4317
rect -316 -4322 -312 -4318
rect 472 -4320 476 -4316
rect 876 -4321 880 -4317
rect 1217 -4320 1221 -4316
rect -1271 -4583 -1267 -4579
rect -942 -4583 -938 -4579
rect -587 -4583 -583 -4579
rect -1272 -4704 -1268 -4700
rect -941 -4704 -937 -4700
rect -587 -4704 -583 -4700
rect -226 -4704 -222 -4700
rect 202 -4704 206 -4700
rect 558 -4704 562 -4700
rect 955 -4704 959 -4700
rect 1315 -4704 1319 -4700
rect 106 -4806 110 -4802
rect -1272 -4825 -1268 -4821
rect -941 -4825 -937 -4821
rect -587 -4825 -583 -4821
rect -226 -4825 -222 -4821
rect 202 -4825 206 -4821
rect 558 -4825 562 -4821
rect 955 -4825 959 -4821
rect 1315 -4825 1319 -4821
rect -1275 -4943 -1271 -4939
rect -940 -4943 -936 -4939
rect -583 -4943 -579 -4939
rect -225 -4943 -221 -4939
rect 202 -4943 206 -4939
rect -1270 -5298 -1266 -5294
rect -942 -5298 -938 -5294
rect -1010 -5394 -1006 -5390
rect -657 -5399 -653 -5395
rect -311 -5400 -307 -5396
rect 482 -5394 486 -5390
rect 883 -5399 887 -5395
rect 1226 -5403 1230 -5399
rect -1270 -5419 -1266 -5415
rect -942 -5419 -938 -5415
rect -585 -5419 -581 -5415
rect -226 -5419 -222 -5415
rect 205 -5419 209 -5415
rect 557 -5419 561 -5415
rect 952 -5419 956 -5415
rect 1313 -5419 1317 -5415
rect -1010 -5518 -1006 -5514
rect -311 -5515 -307 -5511
rect 482 -5518 486 -5514
rect 1226 -5518 1230 -5514
rect -1278 -5539 -1274 -5535
rect -941 -5539 -937 -5535
rect -581 -5539 -577 -5535
rect -227 -5539 -223 -5535
rect 203 -5539 207 -5535
rect 561 -5539 565 -5535
rect 953 -5539 957 -5535
rect 1316 -5539 1320 -5535
rect -1278 -5656 -1274 -5652
rect -941 -5656 -937 -5652
rect -581 -5656 -577 -5652
rect -227 -5656 -223 -5652
rect 203 -5656 207 -5652
rect 561 -5656 565 -5652
rect -1271 -6015 -1267 -6011
rect -940 -6015 -936 -6011
rect -584 -6015 -580 -6011
rect -227 -6015 -223 -6011
rect 201 -6015 205 -6011
rect 559 -6015 563 -6011
rect 957 -6015 961 -6011
rect 1314 -6015 1318 -6011
rect 1316 -6133 1320 -6129
<< pad >>
rect -1325 -1074 -1321 -1070
rect -924 -1074 -920 -1070
rect -565 -1074 -561 -1070
rect -207 -1074 -203 -1070
rect 221 -1074 225 -1070
rect 577 -1074 581 -1070
rect 975 -1074 979 -1070
rect 1333 -1074 1337 -1070
rect -1233 -1196 -1229 -1192
rect -1195 -1196 -1191 -1192
rect -1135 -1196 -1131 -1192
rect -1111 -1196 -1107 -1192
rect -908 -1196 -904 -1192
rect -870 -1196 -866 -1192
rect -810 -1196 -806 -1192
rect -786 -1196 -782 -1192
rect -550 -1196 -546 -1192
rect -512 -1196 -508 -1192
rect -452 -1196 -448 -1192
rect -428 -1196 -424 -1192
rect -192 -1196 -188 -1192
rect -154 -1196 -150 -1192
rect -94 -1196 -90 -1192
rect -70 -1196 -66 -1192
rect 236 -1196 240 -1192
rect 274 -1196 278 -1192
rect 334 -1196 338 -1192
rect 358 -1196 362 -1192
rect 592 -1196 596 -1192
rect 630 -1196 634 -1192
rect 690 -1196 694 -1192
rect 714 -1196 718 -1192
rect 990 -1196 994 -1192
rect 1028 -1196 1032 -1192
rect 1088 -1196 1092 -1192
rect 1112 -1196 1116 -1192
rect -1253 -1204 -1249 -1200
rect -1219 -1204 -1215 -1200
rect -1167 -1204 -1163 -1200
rect -1107 -1204 -1103 -1200
rect -1069 -1204 -1065 -1200
rect -928 -1204 -924 -1200
rect -894 -1204 -890 -1200
rect -842 -1204 -838 -1200
rect -782 -1204 -778 -1200
rect -744 -1204 -740 -1200
rect -570 -1204 -566 -1200
rect -536 -1204 -532 -1200
rect -484 -1204 -480 -1200
rect -424 -1204 -420 -1200
rect -386 -1204 -382 -1200
rect -212 -1204 -208 -1200
rect -178 -1204 -174 -1200
rect -126 -1204 -122 -1200
rect -66 -1204 -62 -1200
rect -28 -1204 -24 -1200
rect 216 -1204 220 -1200
rect 250 -1204 254 -1200
rect 302 -1204 306 -1200
rect 362 -1204 366 -1200
rect 400 -1204 404 -1200
rect 572 -1204 576 -1200
rect 606 -1204 610 -1200
rect 658 -1204 662 -1200
rect 718 -1204 722 -1200
rect 756 -1204 760 -1200
rect 970 -1204 974 -1200
rect 1004 -1204 1008 -1200
rect 1056 -1204 1060 -1200
rect 1116 -1204 1120 -1200
rect 1154 -1204 1158 -1200
rect -1209 -1211 -1205 -1207
rect -1177 -1211 -1173 -1207
rect -1125 -1211 -1121 -1207
rect -1093 -1211 -1089 -1207
rect -884 -1211 -880 -1207
rect -852 -1211 -848 -1207
rect -800 -1211 -796 -1207
rect -768 -1211 -764 -1207
rect -526 -1211 -522 -1207
rect -494 -1211 -490 -1207
rect -442 -1211 -438 -1207
rect -410 -1211 -406 -1207
rect -168 -1211 -164 -1207
rect -136 -1211 -132 -1207
rect -84 -1211 -80 -1207
rect -52 -1211 -48 -1207
rect 260 -1211 264 -1207
rect 292 -1211 296 -1207
rect 344 -1211 348 -1207
rect 376 -1211 380 -1207
rect 616 -1211 620 -1207
rect 648 -1211 652 -1207
rect 700 -1211 704 -1207
rect 732 -1211 736 -1207
rect 1014 -1211 1018 -1207
rect 1046 -1211 1050 -1207
rect 1098 -1211 1102 -1207
rect 1130 -1211 1134 -1207
rect -1249 -1218 -1245 -1214
rect -1135 -1218 -1131 -1214
rect -1083 -1218 -1079 -1214
rect -924 -1218 -920 -1214
rect -810 -1218 -806 -1214
rect -758 -1218 -754 -1214
rect -566 -1218 -562 -1214
rect -452 -1218 -448 -1214
rect -400 -1218 -396 -1214
rect -208 -1218 -204 -1214
rect -94 -1218 -90 -1214
rect -42 -1218 -38 -1214
rect 220 -1218 224 -1214
rect 334 -1218 338 -1214
rect 386 -1218 390 -1214
rect 576 -1218 580 -1214
rect 690 -1218 694 -1214
rect 742 -1218 746 -1214
rect 974 -1218 978 -1214
rect 1088 -1218 1092 -1214
rect 1140 -1218 1144 -1214
rect -1191 -1225 -1187 -1221
rect -1153 -1225 -1149 -1221
rect -866 -1225 -862 -1221
rect -828 -1225 -824 -1221
rect -508 -1225 -504 -1221
rect -470 -1225 -466 -1221
rect -150 -1225 -146 -1221
rect -112 -1225 -108 -1221
rect 278 -1225 282 -1221
rect 316 -1225 320 -1221
rect 634 -1225 638 -1221
rect 672 -1225 676 -1221
rect 1032 -1225 1036 -1221
rect 1070 -1225 1074 -1221
rect -1327 -1304 -1323 -1300
rect -923 -1304 -919 -1300
rect -565 -1304 -561 -1300
rect -207 -1304 -203 -1300
rect 221 -1304 225 -1300
rect 577 -1304 581 -1300
rect 975 -1304 979 -1300
rect 1333 -1304 1337 -1300
rect -924 -1397 -920 -1393
rect -858 -1397 -854 -1393
rect -824 -1397 -820 -1393
rect -780 -1397 -776 -1393
rect -746 -1397 -742 -1393
rect -566 -1397 -562 -1393
rect -500 -1397 -496 -1393
rect -466 -1397 -462 -1393
rect -422 -1397 -418 -1393
rect -388 -1397 -384 -1393
rect -208 -1397 -204 -1393
rect -142 -1397 -138 -1393
rect -108 -1397 -104 -1393
rect -64 -1397 -60 -1393
rect -30 -1397 -26 -1393
rect 220 -1397 224 -1393
rect 286 -1397 290 -1393
rect 320 -1397 324 -1393
rect 364 -1397 368 -1393
rect 398 -1397 402 -1393
rect 576 -1397 580 -1393
rect 642 -1397 646 -1393
rect 676 -1397 680 -1393
rect 720 -1397 724 -1393
rect 754 -1397 758 -1393
rect 974 -1397 978 -1393
rect 1040 -1397 1044 -1393
rect 1074 -1397 1078 -1393
rect 1118 -1397 1122 -1393
rect 1152 -1397 1156 -1393
rect -882 -1404 -878 -1400
rect -524 -1404 -520 -1400
rect -166 -1404 -162 -1400
rect 262 -1404 266 -1400
rect 618 -1404 622 -1400
rect 1016 -1404 1020 -1400
rect -848 -1411 -844 -1407
rect -706 -1411 -702 -1407
rect -490 -1411 -486 -1407
rect -348 -1411 -344 -1407
rect -132 -1411 -128 -1407
rect 10 -1411 14 -1407
rect 296 -1411 300 -1407
rect 438 -1411 442 -1407
rect 652 -1411 656 -1407
rect 794 -1411 798 -1407
rect 1050 -1411 1054 -1407
rect 1192 -1411 1196 -1407
rect -928 -1418 -924 -1414
rect -898 -1418 -894 -1414
rect -780 -1418 -776 -1414
rect -570 -1418 -566 -1414
rect -540 -1418 -536 -1414
rect -422 -1418 -418 -1414
rect -212 -1418 -208 -1414
rect -182 -1418 -178 -1414
rect -64 -1418 -60 -1414
rect 216 -1418 220 -1414
rect 246 -1418 250 -1414
rect 364 -1418 368 -1414
rect 572 -1418 576 -1414
rect 602 -1418 606 -1414
rect 720 -1418 724 -1414
rect 970 -1418 974 -1414
rect 1000 -1418 1004 -1414
rect 1118 -1418 1122 -1414
rect -1199 -1427 -1195 -1423
rect -902 -1426 -898 -1422
rect -804 -1426 -800 -1422
rect -544 -1426 -540 -1422
rect -446 -1426 -442 -1422
rect -186 -1426 -182 -1422
rect -88 -1426 -84 -1422
rect 242 -1426 246 -1422
rect 340 -1426 344 -1422
rect 598 -1426 602 -1422
rect 696 -1426 700 -1422
rect 996 -1426 1000 -1422
rect 1094 -1426 1098 -1422
rect 1382 -1427 1386 -1423
rect -1249 -1434 -1245 -1430
rect -1209 -1434 -1205 -1430
rect -1189 -1434 -1185 -1430
rect -924 -1433 -920 -1429
rect -776 -1433 -772 -1429
rect -566 -1433 -562 -1429
rect -418 -1433 -414 -1429
rect -208 -1433 -204 -1429
rect -60 -1433 -56 -1429
rect 220 -1433 224 -1429
rect 368 -1433 372 -1429
rect 576 -1433 580 -1429
rect 724 -1433 728 -1429
rect 974 -1433 978 -1429
rect 1122 -1433 1126 -1429
rect 1332 -1434 1336 -1430
rect 1372 -1434 1376 -1430
rect 1392 -1434 1396 -1430
rect -1253 -1441 -1249 -1437
rect -1223 -1441 -1219 -1437
rect -1175 -1441 -1171 -1437
rect -902 -1440 -898 -1436
rect -794 -1440 -790 -1436
rect -760 -1440 -756 -1436
rect -544 -1440 -540 -1436
rect -436 -1440 -432 -1436
rect -402 -1440 -398 -1436
rect -186 -1440 -182 -1436
rect -78 -1440 -74 -1436
rect -44 -1440 -40 -1436
rect 242 -1440 246 -1436
rect 350 -1440 354 -1436
rect 384 -1440 388 -1436
rect 598 -1440 602 -1436
rect 706 -1440 710 -1436
rect 740 -1440 744 -1436
rect 996 -1440 1000 -1436
rect 1104 -1440 1108 -1436
rect 1138 -1440 1142 -1436
rect 1328 -1441 1332 -1437
rect 1358 -1441 1362 -1437
rect 1406 -1441 1410 -1437
rect -928 -1447 -924 -1443
rect -872 -1447 -868 -1443
rect -838 -1447 -834 -1443
rect -570 -1447 -566 -1443
rect -514 -1447 -510 -1443
rect -480 -1447 -476 -1443
rect -212 -1447 -208 -1443
rect -156 -1447 -152 -1443
rect -122 -1447 -118 -1443
rect 216 -1447 220 -1443
rect 272 -1447 276 -1443
rect 306 -1447 310 -1443
rect 572 -1447 576 -1443
rect 628 -1447 632 -1443
rect 662 -1447 666 -1443
rect 970 -1447 974 -1443
rect 1026 -1447 1030 -1443
rect 1060 -1447 1064 -1443
rect -1233 -1549 -1229 -1545
rect -1195 -1549 -1191 -1545
rect -1135 -1549 -1131 -1545
rect -1111 -1549 -1107 -1545
rect -908 -1549 -904 -1545
rect -870 -1549 -866 -1545
rect -810 -1549 -806 -1545
rect -786 -1549 -782 -1545
rect -550 -1549 -546 -1545
rect -512 -1549 -508 -1545
rect -452 -1549 -448 -1545
rect -428 -1549 -424 -1545
rect -192 -1549 -188 -1545
rect -154 -1549 -150 -1545
rect -94 -1549 -90 -1545
rect -70 -1549 -66 -1545
rect 236 -1549 240 -1545
rect 274 -1549 278 -1545
rect 334 -1549 338 -1545
rect 358 -1549 362 -1545
rect 592 -1549 596 -1545
rect 630 -1549 634 -1545
rect 690 -1549 694 -1545
rect 714 -1549 718 -1545
rect 990 -1549 994 -1545
rect 1028 -1549 1032 -1545
rect 1088 -1549 1092 -1545
rect 1112 -1549 1116 -1545
rect -1253 -1557 -1249 -1553
rect -1219 -1557 -1215 -1553
rect -1167 -1557 -1163 -1553
rect -1107 -1557 -1103 -1553
rect -1069 -1557 -1065 -1553
rect -928 -1557 -924 -1553
rect -894 -1557 -890 -1553
rect -842 -1557 -838 -1553
rect -782 -1557 -778 -1553
rect -744 -1557 -740 -1553
rect -570 -1557 -566 -1553
rect -536 -1557 -532 -1553
rect -484 -1557 -480 -1553
rect -424 -1557 -420 -1553
rect -386 -1557 -382 -1553
rect -212 -1557 -208 -1553
rect -178 -1557 -174 -1553
rect -126 -1557 -122 -1553
rect -66 -1557 -62 -1553
rect -28 -1557 -24 -1553
rect 216 -1557 220 -1553
rect 250 -1557 254 -1553
rect 302 -1557 306 -1553
rect 362 -1557 366 -1553
rect 400 -1557 404 -1553
rect 572 -1557 576 -1553
rect 606 -1557 610 -1553
rect 658 -1557 662 -1553
rect 718 -1557 722 -1553
rect 756 -1557 760 -1553
rect 970 -1557 974 -1553
rect 1004 -1557 1008 -1553
rect 1056 -1557 1060 -1553
rect 1116 -1557 1120 -1553
rect 1154 -1557 1158 -1553
rect -1209 -1564 -1205 -1560
rect -1177 -1564 -1173 -1560
rect -1125 -1564 -1121 -1560
rect -1093 -1564 -1089 -1560
rect -884 -1564 -880 -1560
rect -852 -1564 -848 -1560
rect -800 -1564 -796 -1560
rect -768 -1564 -764 -1560
rect -526 -1564 -522 -1560
rect -494 -1564 -490 -1560
rect -442 -1564 -438 -1560
rect -410 -1564 -406 -1560
rect -168 -1564 -164 -1560
rect -136 -1564 -132 -1560
rect -84 -1564 -80 -1560
rect -52 -1564 -48 -1560
rect 260 -1564 264 -1560
rect 292 -1564 296 -1560
rect 344 -1564 348 -1560
rect 376 -1564 380 -1560
rect 616 -1564 620 -1560
rect 648 -1564 652 -1560
rect 700 -1564 704 -1560
rect 732 -1564 736 -1560
rect 1014 -1564 1018 -1560
rect 1046 -1564 1050 -1560
rect 1098 -1564 1102 -1560
rect 1130 -1564 1134 -1560
rect -1249 -1571 -1245 -1567
rect -1135 -1571 -1131 -1567
rect -1083 -1571 -1079 -1567
rect -924 -1571 -920 -1567
rect -810 -1571 -806 -1567
rect -758 -1571 -754 -1567
rect -566 -1571 -562 -1567
rect -452 -1571 -448 -1567
rect -400 -1571 -396 -1567
rect -208 -1571 -204 -1567
rect -94 -1571 -90 -1567
rect -42 -1571 -38 -1567
rect 220 -1571 224 -1567
rect 334 -1571 338 -1567
rect 386 -1571 390 -1567
rect 576 -1571 580 -1567
rect 690 -1571 694 -1567
rect 742 -1571 746 -1567
rect 974 -1571 978 -1567
rect 1088 -1571 1092 -1567
rect 1140 -1571 1144 -1567
rect -1191 -1578 -1187 -1574
rect -1153 -1578 -1149 -1574
rect -866 -1578 -862 -1574
rect -828 -1578 -824 -1574
rect -508 -1578 -504 -1574
rect -470 -1578 -466 -1574
rect -150 -1578 -146 -1574
rect -112 -1578 -108 -1574
rect 278 -1578 282 -1574
rect 316 -1578 320 -1574
rect 634 -1578 638 -1574
rect 672 -1578 676 -1574
rect 1032 -1578 1036 -1574
rect 1070 -1578 1074 -1574
rect -1233 -1670 -1229 -1666
rect -1195 -1670 -1191 -1666
rect -1135 -1670 -1131 -1666
rect -1111 -1670 -1107 -1666
rect -908 -1670 -904 -1666
rect -870 -1670 -866 -1666
rect -810 -1670 -806 -1666
rect -786 -1670 -782 -1666
rect -550 -1670 -546 -1666
rect -512 -1670 -508 -1666
rect -452 -1670 -448 -1666
rect -428 -1670 -424 -1666
rect -192 -1670 -188 -1666
rect -154 -1670 -150 -1666
rect -94 -1670 -90 -1666
rect -70 -1670 -66 -1666
rect 236 -1670 240 -1666
rect 274 -1670 278 -1666
rect 334 -1670 338 -1666
rect 358 -1670 362 -1666
rect 592 -1670 596 -1666
rect 630 -1670 634 -1666
rect 690 -1670 694 -1666
rect 714 -1670 718 -1666
rect 990 -1670 994 -1666
rect 1028 -1670 1032 -1666
rect 1088 -1670 1092 -1666
rect 1112 -1670 1116 -1666
rect 1348 -1670 1352 -1666
rect 1386 -1670 1390 -1666
rect 1446 -1670 1450 -1666
rect 1470 -1670 1474 -1666
rect -1253 -1678 -1249 -1674
rect -1219 -1678 -1215 -1674
rect -1167 -1678 -1163 -1674
rect -1107 -1678 -1103 -1674
rect -1069 -1678 -1065 -1674
rect -928 -1678 -924 -1674
rect -894 -1678 -890 -1674
rect -842 -1678 -838 -1674
rect -782 -1678 -778 -1674
rect -744 -1678 -740 -1674
rect -570 -1678 -566 -1674
rect -536 -1678 -532 -1674
rect -484 -1678 -480 -1674
rect -424 -1678 -420 -1674
rect -386 -1678 -382 -1674
rect -212 -1678 -208 -1674
rect -178 -1678 -174 -1674
rect -126 -1678 -122 -1674
rect -66 -1678 -62 -1674
rect -28 -1678 -24 -1674
rect 216 -1678 220 -1674
rect 250 -1678 254 -1674
rect 302 -1678 306 -1674
rect 362 -1678 366 -1674
rect 400 -1678 404 -1674
rect 572 -1678 576 -1674
rect 606 -1678 610 -1674
rect 658 -1678 662 -1674
rect 718 -1678 722 -1674
rect 756 -1678 760 -1674
rect 970 -1678 974 -1674
rect 1004 -1678 1008 -1674
rect 1056 -1678 1060 -1674
rect 1116 -1678 1120 -1674
rect 1154 -1678 1158 -1674
rect 1328 -1678 1332 -1674
rect 1362 -1678 1366 -1674
rect 1414 -1678 1418 -1674
rect 1474 -1678 1478 -1674
rect 1512 -1678 1516 -1674
rect -1209 -1685 -1205 -1681
rect -1177 -1685 -1173 -1681
rect -1125 -1685 -1121 -1681
rect -1093 -1685 -1089 -1681
rect -884 -1685 -880 -1681
rect -852 -1685 -848 -1681
rect -800 -1685 -796 -1681
rect -768 -1685 -764 -1681
rect -526 -1685 -522 -1681
rect -494 -1685 -490 -1681
rect -442 -1685 -438 -1681
rect -410 -1685 -406 -1681
rect -168 -1685 -164 -1681
rect -136 -1685 -132 -1681
rect -84 -1685 -80 -1681
rect -52 -1685 -48 -1681
rect 260 -1685 264 -1681
rect 292 -1685 296 -1681
rect 344 -1685 348 -1681
rect 376 -1685 380 -1681
rect 616 -1685 620 -1681
rect 648 -1685 652 -1681
rect 700 -1685 704 -1681
rect 732 -1685 736 -1681
rect 1014 -1685 1018 -1681
rect 1046 -1685 1050 -1681
rect 1098 -1685 1102 -1681
rect 1130 -1685 1134 -1681
rect 1372 -1685 1376 -1681
rect 1404 -1685 1408 -1681
rect 1456 -1685 1460 -1681
rect 1488 -1685 1492 -1681
rect -1249 -1692 -1245 -1688
rect -1135 -1692 -1131 -1688
rect -1083 -1692 -1079 -1688
rect -924 -1692 -920 -1688
rect -810 -1692 -806 -1688
rect -758 -1692 -754 -1688
rect -566 -1692 -562 -1688
rect -452 -1692 -448 -1688
rect -400 -1692 -396 -1688
rect -208 -1692 -204 -1688
rect -94 -1692 -90 -1688
rect -42 -1692 -38 -1688
rect 220 -1692 224 -1688
rect 334 -1692 338 -1688
rect 386 -1692 390 -1688
rect 576 -1692 580 -1688
rect 690 -1692 694 -1688
rect 742 -1692 746 -1688
rect 974 -1692 978 -1688
rect 1088 -1692 1092 -1688
rect 1140 -1692 1144 -1688
rect 1332 -1692 1336 -1688
rect 1446 -1692 1450 -1688
rect 1498 -1692 1502 -1688
rect -1191 -1699 -1187 -1695
rect -1153 -1699 -1149 -1695
rect -866 -1699 -862 -1695
rect -828 -1699 -824 -1695
rect -508 -1699 -504 -1695
rect -470 -1699 -466 -1695
rect -150 -1699 -146 -1695
rect -112 -1699 -108 -1695
rect 278 -1699 282 -1695
rect 316 -1699 320 -1695
rect 634 -1699 638 -1695
rect 672 -1699 676 -1695
rect 1032 -1699 1036 -1695
rect 1070 -1699 1074 -1695
rect 1390 -1699 1394 -1695
rect 1428 -1699 1432 -1695
rect -1233 -1791 -1229 -1787
rect -1195 -1791 -1191 -1787
rect -1135 -1791 -1131 -1787
rect -1111 -1791 -1107 -1787
rect -1028 -1795 -1024 -1785
rect -908 -1791 -904 -1787
rect -870 -1791 -866 -1787
rect -810 -1791 -806 -1787
rect -786 -1791 -782 -1787
rect -550 -1791 -546 -1787
rect -512 -1791 -508 -1787
rect -452 -1791 -448 -1787
rect -428 -1791 -424 -1787
rect -331 -1795 -327 -1785
rect -192 -1791 -188 -1787
rect -154 -1791 -150 -1787
rect -94 -1791 -90 -1787
rect -70 -1791 -66 -1787
rect 236 -1791 240 -1787
rect 274 -1791 278 -1787
rect 334 -1791 338 -1787
rect 358 -1791 362 -1787
rect 465 -1795 469 -1785
rect 592 -1791 596 -1787
rect 630 -1791 634 -1787
rect 690 -1791 694 -1787
rect 714 -1791 718 -1787
rect 990 -1791 994 -1787
rect 1028 -1791 1032 -1787
rect 1088 -1791 1092 -1787
rect 1112 -1791 1116 -1787
rect 1204 -1795 1208 -1785
rect 1348 -1791 1352 -1787
rect 1386 -1791 1390 -1787
rect 1446 -1791 1450 -1787
rect 1470 -1791 1474 -1787
rect -1253 -1799 -1249 -1795
rect -1219 -1799 -1215 -1795
rect -1167 -1799 -1163 -1795
rect -1107 -1799 -1103 -1795
rect -1069 -1799 -1065 -1795
rect -928 -1799 -924 -1795
rect -894 -1799 -890 -1795
rect -842 -1799 -838 -1795
rect -782 -1799 -778 -1795
rect -744 -1799 -740 -1795
rect -570 -1799 -566 -1795
rect -536 -1799 -532 -1795
rect -484 -1799 -480 -1795
rect -424 -1799 -420 -1795
rect -386 -1799 -382 -1795
rect -212 -1799 -208 -1795
rect -178 -1799 -174 -1795
rect -126 -1799 -122 -1795
rect -66 -1799 -62 -1795
rect -28 -1799 -24 -1795
rect 216 -1799 220 -1795
rect 250 -1799 254 -1795
rect 302 -1799 306 -1795
rect 362 -1799 366 -1795
rect 400 -1799 404 -1795
rect 572 -1799 576 -1795
rect 606 -1799 610 -1795
rect 658 -1799 662 -1795
rect 718 -1799 722 -1795
rect 756 -1799 760 -1795
rect 970 -1799 974 -1795
rect 1004 -1799 1008 -1795
rect 1056 -1799 1060 -1795
rect 1116 -1799 1120 -1795
rect 1154 -1799 1158 -1795
rect 1328 -1799 1332 -1795
rect 1362 -1799 1366 -1795
rect 1414 -1799 1418 -1795
rect 1474 -1799 1478 -1795
rect 1512 -1799 1516 -1795
rect -1209 -1806 -1205 -1802
rect -1177 -1806 -1173 -1802
rect -1125 -1806 -1121 -1802
rect -1093 -1806 -1089 -1802
rect -884 -1806 -880 -1802
rect -852 -1806 -848 -1802
rect -800 -1806 -796 -1802
rect -768 -1806 -764 -1802
rect -526 -1806 -522 -1802
rect -494 -1806 -490 -1802
rect -442 -1806 -438 -1802
rect -410 -1806 -406 -1802
rect -168 -1806 -164 -1802
rect -136 -1806 -132 -1802
rect -84 -1806 -80 -1802
rect -52 -1806 -48 -1802
rect 260 -1806 264 -1802
rect 292 -1806 296 -1802
rect 344 -1806 348 -1802
rect 376 -1806 380 -1802
rect 616 -1806 620 -1802
rect 648 -1806 652 -1802
rect 700 -1806 704 -1802
rect 732 -1806 736 -1802
rect 1014 -1806 1018 -1802
rect 1046 -1806 1050 -1802
rect 1098 -1806 1102 -1802
rect 1130 -1806 1134 -1802
rect 1372 -1806 1376 -1802
rect 1404 -1806 1408 -1802
rect 1456 -1806 1460 -1802
rect 1488 -1806 1492 -1802
rect -1249 -1813 -1245 -1809
rect -1135 -1813 -1131 -1809
rect -1083 -1813 -1079 -1809
rect -924 -1813 -920 -1809
rect -810 -1813 -806 -1809
rect -758 -1813 -754 -1809
rect -566 -1813 -562 -1809
rect -452 -1813 -448 -1809
rect -400 -1813 -396 -1809
rect -208 -1813 -204 -1809
rect -94 -1813 -90 -1809
rect -42 -1813 -38 -1809
rect 220 -1813 224 -1809
rect 334 -1813 338 -1809
rect 386 -1813 390 -1809
rect 576 -1813 580 -1809
rect 690 -1813 694 -1809
rect 742 -1813 746 -1809
rect 974 -1813 978 -1809
rect 1088 -1813 1092 -1809
rect 1140 -1813 1144 -1809
rect 1332 -1813 1336 -1809
rect 1446 -1813 1450 -1809
rect 1498 -1813 1502 -1809
rect -1191 -1820 -1187 -1816
rect -1153 -1820 -1149 -1816
rect -866 -1820 -862 -1816
rect -828 -1820 -824 -1816
rect -508 -1820 -504 -1816
rect -470 -1820 -466 -1816
rect -150 -1820 -146 -1816
rect -112 -1820 -108 -1816
rect 278 -1820 282 -1816
rect 316 -1820 320 -1816
rect 634 -1820 638 -1816
rect 672 -1820 676 -1816
rect 1032 -1820 1036 -1816
rect 1070 -1820 1074 -1816
rect 1390 -1820 1394 -1816
rect 1428 -1820 1432 -1816
rect -1233 -1906 -1229 -1902
rect -1195 -1906 -1191 -1902
rect -1135 -1906 -1131 -1902
rect -1111 -1906 -1107 -1902
rect -1028 -1910 -1024 -1900
rect -672 -1910 -668 -1900
rect -331 -1910 -327 -1900
rect 465 -1910 469 -1900
rect 842 -1910 846 -1900
rect 1204 -1910 1208 -1900
rect -1253 -1914 -1249 -1910
rect -1219 -1914 -1215 -1910
rect -1167 -1914 -1163 -1910
rect -1107 -1914 -1103 -1910
rect -1069 -1914 -1065 -1910
rect -1209 -1921 -1205 -1917
rect -1177 -1921 -1173 -1917
rect -1125 -1921 -1121 -1917
rect -1093 -1921 -1089 -1917
rect -1249 -1928 -1245 -1924
rect -1135 -1928 -1131 -1924
rect -1083 -1928 -1079 -1924
rect -1191 -1935 -1187 -1931
rect -1153 -1935 -1149 -1931
rect -1338 -2002 -1334 -1998
rect -934 -2002 -930 -1998
rect -576 -2002 -572 -1998
rect -218 -2002 -214 -1998
rect 210 -2002 214 -1998
rect 566 -2002 570 -1998
rect 964 -2002 968 -1998
rect 1322 -2002 1326 -1998
rect -1327 -2010 -1323 -2006
rect -923 -2010 -919 -2006
rect -565 -2010 -561 -2006
rect -207 -2010 -203 -2006
rect 221 -2010 225 -2006
rect 577 -2010 581 -2006
rect 975 -2010 979 -2006
rect 1333 -2010 1337 -2006
rect -924 -2108 -920 -2104
rect -858 -2108 -854 -2104
rect -824 -2108 -820 -2104
rect -780 -2108 -776 -2104
rect -746 -2108 -742 -2104
rect -566 -2108 -562 -2104
rect -500 -2108 -496 -2104
rect -466 -2108 -462 -2104
rect -422 -2108 -418 -2104
rect -388 -2108 -384 -2104
rect -208 -2108 -204 -2104
rect -142 -2108 -138 -2104
rect -108 -2108 -104 -2104
rect -64 -2108 -60 -2104
rect -30 -2108 -26 -2104
rect 220 -2108 224 -2104
rect 286 -2108 290 -2104
rect 320 -2108 324 -2104
rect 364 -2108 368 -2104
rect 398 -2108 402 -2104
rect 576 -2108 580 -2104
rect 642 -2108 646 -2104
rect 676 -2108 680 -2104
rect 720 -2108 724 -2104
rect 754 -2108 758 -2104
rect 974 -2108 978 -2104
rect 1040 -2108 1044 -2104
rect 1074 -2108 1078 -2104
rect 1118 -2108 1122 -2104
rect 1152 -2108 1156 -2104
rect 1332 -2108 1336 -2104
rect 1398 -2108 1402 -2104
rect 1432 -2108 1436 -2104
rect 1476 -2108 1480 -2104
rect 1510 -2108 1514 -2104
rect -882 -2115 -878 -2111
rect -524 -2115 -520 -2111
rect -166 -2115 -162 -2111
rect 262 -2115 266 -2111
rect 618 -2115 622 -2111
rect 1016 -2115 1020 -2111
rect 1374 -2115 1378 -2111
rect -848 -2122 -844 -2118
rect -706 -2122 -702 -2118
rect -490 -2122 -486 -2118
rect -348 -2122 -344 -2118
rect -132 -2122 -128 -2118
rect 10 -2122 14 -2118
rect 296 -2122 300 -2118
rect 438 -2122 442 -2118
rect 652 -2122 656 -2118
rect 794 -2122 798 -2118
rect 1050 -2122 1054 -2118
rect 1192 -2122 1196 -2118
rect 1408 -2122 1412 -2118
rect 1550 -2122 1554 -2118
rect -928 -2129 -924 -2125
rect -898 -2129 -894 -2125
rect -780 -2129 -776 -2125
rect -570 -2129 -566 -2125
rect -540 -2129 -536 -2125
rect -422 -2129 -418 -2125
rect -212 -2129 -208 -2125
rect -182 -2129 -178 -2125
rect -64 -2129 -60 -2125
rect 216 -2129 220 -2125
rect 246 -2129 250 -2125
rect 364 -2129 368 -2125
rect 572 -2129 576 -2125
rect 602 -2129 606 -2125
rect 720 -2129 724 -2125
rect 970 -2129 974 -2125
rect 1000 -2129 1004 -2125
rect 1118 -2129 1122 -2125
rect 1328 -2129 1332 -2125
rect 1358 -2129 1362 -2125
rect 1476 -2129 1480 -2125
rect -1199 -2138 -1195 -2134
rect -902 -2137 -898 -2133
rect -804 -2137 -800 -2133
rect -544 -2137 -540 -2133
rect -446 -2137 -442 -2133
rect -186 -2137 -182 -2133
rect -88 -2137 -84 -2133
rect 242 -2137 246 -2133
rect 340 -2137 344 -2133
rect 598 -2137 602 -2133
rect 696 -2137 700 -2133
rect 996 -2137 1000 -2133
rect 1094 -2137 1098 -2133
rect 1354 -2137 1358 -2133
rect 1452 -2137 1456 -2133
rect -1249 -2145 -1245 -2141
rect -1209 -2145 -1205 -2141
rect -1189 -2145 -1185 -2141
rect -924 -2144 -920 -2140
rect -776 -2144 -772 -2140
rect -566 -2144 -562 -2140
rect -418 -2144 -414 -2140
rect -208 -2144 -204 -2140
rect -60 -2144 -56 -2140
rect 220 -2144 224 -2140
rect 368 -2144 372 -2140
rect 576 -2144 580 -2140
rect 724 -2144 728 -2140
rect 974 -2144 978 -2140
rect 1122 -2144 1126 -2140
rect 1332 -2144 1336 -2140
rect 1480 -2144 1484 -2140
rect -1253 -2152 -1249 -2148
rect -1223 -2152 -1219 -2148
rect -1175 -2152 -1171 -2148
rect -902 -2151 -898 -2147
rect -794 -2151 -790 -2147
rect -760 -2151 -756 -2147
rect -544 -2151 -540 -2147
rect -436 -2151 -432 -2147
rect -402 -2151 -398 -2147
rect -186 -2151 -182 -2147
rect -78 -2151 -74 -2147
rect -44 -2151 -40 -2147
rect 242 -2151 246 -2147
rect 350 -2151 354 -2147
rect 384 -2151 388 -2147
rect 598 -2151 602 -2147
rect 706 -2151 710 -2147
rect 740 -2151 744 -2147
rect 996 -2151 1000 -2147
rect 1104 -2151 1108 -2147
rect 1138 -2151 1142 -2147
rect 1354 -2151 1358 -2147
rect 1462 -2151 1466 -2147
rect 1496 -2151 1500 -2147
rect -928 -2158 -924 -2154
rect -872 -2158 -868 -2154
rect -838 -2158 -834 -2154
rect -570 -2158 -566 -2154
rect -514 -2158 -510 -2154
rect -480 -2158 -476 -2154
rect -212 -2158 -208 -2154
rect -156 -2158 -152 -2154
rect -122 -2158 -118 -2154
rect 216 -2158 220 -2154
rect 272 -2158 276 -2154
rect 306 -2158 310 -2154
rect 572 -2158 576 -2154
rect 628 -2158 632 -2154
rect 662 -2158 666 -2154
rect 970 -2158 974 -2154
rect 1026 -2158 1030 -2154
rect 1060 -2158 1064 -2154
rect 1328 -2158 1332 -2154
rect 1384 -2158 1388 -2154
rect 1418 -2158 1422 -2154
rect -1237 -2281 -1233 -2277
rect -1199 -2281 -1195 -2277
rect -1139 -2281 -1135 -2277
rect -1115 -2281 -1111 -2277
rect -908 -2281 -904 -2277
rect -870 -2281 -866 -2277
rect -810 -2281 -806 -2277
rect -786 -2281 -782 -2277
rect -550 -2281 -546 -2277
rect -512 -2281 -508 -2277
rect -452 -2281 -448 -2277
rect -428 -2281 -424 -2277
rect -192 -2281 -188 -2277
rect -154 -2281 -150 -2277
rect -94 -2281 -90 -2277
rect -70 -2281 -66 -2277
rect 236 -2281 240 -2277
rect 274 -2281 278 -2277
rect 334 -2281 338 -2277
rect 358 -2281 362 -2277
rect 592 -2281 596 -2277
rect 630 -2281 634 -2277
rect 690 -2281 694 -2277
rect 714 -2281 718 -2277
rect -1257 -2289 -1253 -2285
rect -1223 -2289 -1219 -2285
rect -1171 -2289 -1167 -2285
rect -1111 -2289 -1107 -2285
rect -1073 -2289 -1069 -2285
rect -928 -2289 -924 -2285
rect -894 -2289 -890 -2285
rect -842 -2289 -838 -2285
rect -782 -2289 -778 -2285
rect -744 -2289 -740 -2285
rect -570 -2289 -566 -2285
rect -536 -2289 -532 -2285
rect -484 -2289 -480 -2285
rect -424 -2289 -420 -2285
rect -386 -2289 -382 -2285
rect -212 -2289 -208 -2285
rect -178 -2289 -174 -2285
rect -126 -2289 -122 -2285
rect -66 -2289 -62 -2285
rect -28 -2289 -24 -2285
rect 216 -2289 220 -2285
rect 250 -2289 254 -2285
rect 302 -2289 306 -2285
rect 362 -2289 366 -2285
rect 400 -2289 404 -2285
rect 572 -2289 576 -2285
rect 606 -2289 610 -2285
rect 658 -2289 662 -2285
rect 718 -2289 722 -2285
rect 756 -2289 760 -2285
rect -1213 -2296 -1209 -2292
rect -1181 -2296 -1177 -2292
rect -1129 -2296 -1125 -2292
rect -1097 -2296 -1093 -2292
rect -884 -2296 -880 -2292
rect -852 -2296 -848 -2292
rect -800 -2296 -796 -2292
rect -768 -2296 -764 -2292
rect -526 -2296 -522 -2292
rect -494 -2296 -490 -2292
rect -442 -2296 -438 -2292
rect -410 -2296 -406 -2292
rect -168 -2296 -164 -2292
rect -136 -2296 -132 -2292
rect -84 -2296 -80 -2292
rect -52 -2296 -48 -2292
rect 260 -2296 264 -2292
rect 292 -2296 296 -2292
rect 344 -2296 348 -2292
rect 376 -2296 380 -2292
rect 616 -2296 620 -2292
rect 648 -2296 652 -2292
rect 700 -2296 704 -2292
rect 732 -2296 736 -2292
rect -1253 -2303 -1249 -2299
rect -1139 -2303 -1135 -2299
rect -1087 -2303 -1083 -2299
rect -924 -2303 -920 -2299
rect -810 -2303 -806 -2299
rect -758 -2303 -754 -2299
rect -566 -2303 -562 -2299
rect -452 -2303 -448 -2299
rect -400 -2303 -396 -2299
rect -208 -2303 -204 -2299
rect -94 -2303 -90 -2299
rect -42 -2303 -38 -2299
rect 220 -2303 224 -2299
rect 334 -2303 338 -2299
rect 386 -2303 390 -2299
rect 576 -2303 580 -2299
rect 690 -2303 694 -2299
rect 742 -2303 746 -2299
rect -1195 -2310 -1191 -2306
rect -1157 -2310 -1153 -2306
rect -866 -2310 -862 -2306
rect -828 -2310 -824 -2306
rect -508 -2310 -504 -2306
rect -470 -2310 -466 -2306
rect -150 -2310 -146 -2306
rect -112 -2310 -108 -2306
rect 278 -2310 282 -2306
rect 316 -2310 320 -2306
rect 634 -2310 638 -2306
rect 672 -2310 676 -2306
rect -1237 -2412 -1233 -2408
rect -1199 -2412 -1195 -2408
rect -1139 -2412 -1135 -2408
rect -1115 -2412 -1111 -2408
rect -908 -2412 -904 -2408
rect -870 -2412 -866 -2408
rect -810 -2412 -806 -2408
rect -786 -2412 -782 -2408
rect -550 -2412 -546 -2408
rect -512 -2412 -508 -2408
rect -452 -2412 -448 -2408
rect -428 -2412 -424 -2408
rect -192 -2412 -188 -2408
rect -154 -2412 -150 -2408
rect -94 -2412 -90 -2408
rect -70 -2412 -66 -2408
rect 236 -2412 240 -2408
rect 274 -2412 278 -2408
rect 334 -2412 338 -2408
rect 358 -2412 362 -2408
rect 592 -2412 596 -2408
rect 630 -2412 634 -2408
rect 690 -2412 694 -2408
rect 714 -2412 718 -2408
rect 990 -2412 994 -2408
rect 1028 -2412 1032 -2408
rect 1088 -2412 1092 -2408
rect 1112 -2412 1116 -2408
rect 1348 -2412 1352 -2408
rect 1386 -2412 1390 -2408
rect 1446 -2412 1450 -2408
rect 1470 -2412 1474 -2408
rect -1257 -2420 -1253 -2416
rect -1223 -2420 -1219 -2416
rect -1171 -2420 -1167 -2416
rect -1111 -2420 -1107 -2416
rect -1073 -2420 -1069 -2416
rect -928 -2420 -924 -2416
rect -894 -2420 -890 -2416
rect -842 -2420 -838 -2416
rect -782 -2420 -778 -2416
rect -744 -2420 -740 -2416
rect -570 -2420 -566 -2416
rect -536 -2420 -532 -2416
rect -484 -2420 -480 -2416
rect -424 -2420 -420 -2416
rect -386 -2420 -382 -2416
rect -212 -2420 -208 -2416
rect -178 -2420 -174 -2416
rect -126 -2420 -122 -2416
rect -66 -2420 -62 -2416
rect -28 -2420 -24 -2416
rect 216 -2420 220 -2416
rect 250 -2420 254 -2416
rect 302 -2420 306 -2416
rect 362 -2420 366 -2416
rect 400 -2420 404 -2416
rect 572 -2420 576 -2416
rect 606 -2420 610 -2416
rect 658 -2420 662 -2416
rect 718 -2420 722 -2416
rect 756 -2420 760 -2416
rect 970 -2420 974 -2416
rect 1004 -2420 1008 -2416
rect 1056 -2420 1060 -2416
rect 1116 -2420 1120 -2416
rect 1154 -2420 1158 -2416
rect 1328 -2420 1332 -2416
rect 1362 -2420 1366 -2416
rect 1414 -2420 1418 -2416
rect 1474 -2420 1478 -2416
rect 1512 -2420 1516 -2416
rect -1213 -2427 -1209 -2423
rect -1181 -2427 -1177 -2423
rect -1129 -2427 -1125 -2423
rect -1097 -2427 -1093 -2423
rect -884 -2427 -880 -2423
rect -852 -2427 -848 -2423
rect -800 -2427 -796 -2423
rect -768 -2427 -764 -2423
rect -526 -2427 -522 -2423
rect -494 -2427 -490 -2423
rect -442 -2427 -438 -2423
rect -410 -2427 -406 -2423
rect -168 -2427 -164 -2423
rect -136 -2427 -132 -2423
rect -84 -2427 -80 -2423
rect -52 -2427 -48 -2423
rect 260 -2427 264 -2423
rect 292 -2427 296 -2423
rect 344 -2427 348 -2423
rect 376 -2427 380 -2423
rect 616 -2427 620 -2423
rect 648 -2427 652 -2423
rect 700 -2427 704 -2423
rect 732 -2427 736 -2423
rect 1014 -2427 1018 -2423
rect 1046 -2427 1050 -2423
rect 1098 -2427 1102 -2423
rect 1130 -2427 1134 -2423
rect 1372 -2427 1376 -2423
rect 1404 -2427 1408 -2423
rect 1456 -2427 1460 -2423
rect 1488 -2427 1492 -2423
rect -1253 -2434 -1249 -2430
rect -1139 -2434 -1135 -2430
rect -1087 -2434 -1083 -2430
rect -924 -2434 -920 -2430
rect -810 -2434 -806 -2430
rect -758 -2434 -754 -2430
rect -566 -2434 -562 -2430
rect -452 -2434 -448 -2430
rect -400 -2434 -396 -2430
rect -208 -2434 -204 -2430
rect -94 -2434 -90 -2430
rect -42 -2434 -38 -2430
rect 220 -2434 224 -2430
rect 334 -2434 338 -2430
rect 386 -2434 390 -2430
rect 576 -2434 580 -2430
rect 690 -2434 694 -2430
rect 742 -2434 746 -2430
rect 974 -2434 978 -2430
rect 1088 -2434 1092 -2430
rect 1140 -2434 1144 -2430
rect 1332 -2434 1336 -2430
rect 1446 -2434 1450 -2430
rect 1498 -2434 1502 -2430
rect -1195 -2441 -1191 -2437
rect -1157 -2441 -1153 -2437
rect -866 -2441 -862 -2437
rect -828 -2441 -824 -2437
rect -508 -2441 -504 -2437
rect -470 -2441 -466 -2437
rect -150 -2441 -146 -2437
rect -112 -2441 -108 -2437
rect 278 -2441 282 -2437
rect 316 -2441 320 -2437
rect 634 -2441 638 -2437
rect 672 -2441 676 -2437
rect 1032 -2441 1036 -2437
rect 1070 -2441 1074 -2437
rect 1390 -2441 1394 -2437
rect 1428 -2441 1432 -2437
rect -1237 -2543 -1233 -2539
rect -1199 -2543 -1195 -2539
rect -1139 -2543 -1135 -2539
rect -1115 -2543 -1111 -2539
rect -908 -2543 -904 -2539
rect -870 -2543 -866 -2539
rect -810 -2543 -806 -2539
rect -786 -2543 -782 -2539
rect -550 -2543 -546 -2539
rect -512 -2543 -508 -2539
rect -452 -2543 -448 -2539
rect -428 -2543 -424 -2539
rect -192 -2543 -188 -2539
rect -154 -2543 -150 -2539
rect -94 -2543 -90 -2539
rect -70 -2543 -66 -2539
rect -1257 -2551 -1253 -2547
rect -1223 -2551 -1219 -2547
rect -1171 -2551 -1167 -2547
rect -1111 -2551 -1107 -2547
rect -1073 -2551 -1069 -2547
rect -928 -2551 -924 -2547
rect -894 -2551 -890 -2547
rect -842 -2551 -838 -2547
rect -782 -2551 -778 -2547
rect -744 -2551 -740 -2547
rect -570 -2551 -566 -2547
rect -536 -2551 -532 -2547
rect -484 -2551 -480 -2547
rect -424 -2551 -420 -2547
rect -386 -2551 -382 -2547
rect -212 -2551 -208 -2547
rect -178 -2551 -174 -2547
rect -126 -2551 -122 -2547
rect -66 -2551 -62 -2547
rect -28 -2551 -24 -2547
rect 91 -2551 95 -2537
rect 236 -2543 240 -2539
rect 274 -2543 278 -2539
rect 334 -2543 338 -2539
rect 358 -2543 362 -2539
rect 592 -2543 596 -2539
rect 630 -2543 634 -2539
rect 690 -2543 694 -2539
rect 714 -2543 718 -2539
rect 990 -2543 994 -2539
rect 1028 -2543 1032 -2539
rect 1088 -2543 1092 -2539
rect 1112 -2543 1116 -2539
rect 1348 -2543 1352 -2539
rect 1386 -2543 1390 -2539
rect 1446 -2543 1450 -2539
rect 1470 -2543 1474 -2539
rect 216 -2551 220 -2547
rect 250 -2551 254 -2547
rect 302 -2551 306 -2547
rect 362 -2551 366 -2547
rect 400 -2551 404 -2547
rect 572 -2551 576 -2547
rect 606 -2551 610 -2547
rect 658 -2551 662 -2547
rect 718 -2551 722 -2547
rect 756 -2551 760 -2547
rect 970 -2551 974 -2547
rect 1004 -2551 1008 -2547
rect 1056 -2551 1060 -2547
rect 1116 -2551 1120 -2547
rect 1154 -2551 1158 -2547
rect 1328 -2551 1332 -2547
rect 1362 -2551 1366 -2547
rect 1414 -2551 1418 -2547
rect 1474 -2551 1478 -2547
rect 1512 -2551 1516 -2547
rect -1213 -2558 -1209 -2554
rect -1181 -2558 -1177 -2554
rect -1129 -2558 -1125 -2554
rect -1097 -2558 -1093 -2554
rect -884 -2558 -880 -2554
rect -852 -2558 -848 -2554
rect -800 -2558 -796 -2554
rect -768 -2558 -764 -2554
rect -526 -2558 -522 -2554
rect -494 -2558 -490 -2554
rect -442 -2558 -438 -2554
rect -410 -2558 -406 -2554
rect -168 -2558 -164 -2554
rect -136 -2558 -132 -2554
rect -84 -2558 -80 -2554
rect -52 -2558 -48 -2554
rect 260 -2558 264 -2554
rect 292 -2558 296 -2554
rect 344 -2558 348 -2554
rect 376 -2558 380 -2554
rect 616 -2558 620 -2554
rect 648 -2558 652 -2554
rect 700 -2558 704 -2554
rect 732 -2558 736 -2554
rect 1014 -2558 1018 -2554
rect 1046 -2558 1050 -2554
rect 1098 -2558 1102 -2554
rect 1130 -2558 1134 -2554
rect 1372 -2558 1376 -2554
rect 1404 -2558 1408 -2554
rect 1456 -2558 1460 -2554
rect 1488 -2558 1492 -2554
rect -1253 -2565 -1249 -2561
rect -1139 -2565 -1135 -2561
rect -1087 -2565 -1083 -2561
rect -924 -2565 -920 -2561
rect -810 -2565 -806 -2561
rect -758 -2565 -754 -2561
rect -566 -2565 -562 -2561
rect -452 -2565 -448 -2561
rect -400 -2565 -396 -2561
rect -208 -2565 -204 -2561
rect -94 -2565 -90 -2561
rect -42 -2565 -38 -2561
rect 220 -2565 224 -2561
rect 334 -2565 338 -2561
rect 386 -2565 390 -2561
rect 576 -2565 580 -2561
rect 690 -2565 694 -2561
rect 742 -2565 746 -2561
rect 974 -2565 978 -2561
rect 1088 -2565 1092 -2561
rect 1140 -2565 1144 -2561
rect 1332 -2565 1336 -2561
rect 1446 -2565 1450 -2561
rect 1498 -2565 1502 -2561
rect -1195 -2572 -1191 -2568
rect -1157 -2572 -1153 -2568
rect -866 -2572 -862 -2568
rect -828 -2572 -824 -2568
rect -508 -2572 -504 -2568
rect -470 -2572 -466 -2568
rect -150 -2572 -146 -2568
rect -112 -2572 -108 -2568
rect 278 -2572 282 -2568
rect 316 -2572 320 -2568
rect 634 -2572 638 -2568
rect 672 -2572 676 -2568
rect 1032 -2572 1036 -2568
rect 1070 -2572 1074 -2568
rect 1390 -2572 1394 -2568
rect 1428 -2572 1432 -2568
rect -1237 -2655 -1233 -2651
rect -1199 -2655 -1195 -2651
rect -1139 -2655 -1135 -2651
rect -1115 -2655 -1111 -2651
rect -908 -2655 -904 -2651
rect -870 -2655 -866 -2651
rect -810 -2655 -806 -2651
rect -786 -2655 -782 -2651
rect -1257 -2663 -1253 -2659
rect -1223 -2663 -1219 -2659
rect -1171 -2663 -1167 -2659
rect -1111 -2663 -1107 -2659
rect -1073 -2663 -1069 -2659
rect -928 -2663 -924 -2659
rect -894 -2663 -890 -2659
rect -842 -2663 -838 -2659
rect -782 -2663 -778 -2659
rect -744 -2663 -740 -2659
rect -1213 -2670 -1209 -2666
rect -1181 -2670 -1177 -2666
rect -1129 -2670 -1125 -2666
rect -1097 -2670 -1093 -2666
rect -884 -2670 -880 -2666
rect -852 -2670 -848 -2666
rect -800 -2670 -796 -2666
rect -768 -2670 -764 -2666
rect -1253 -2677 -1249 -2673
rect -1139 -2677 -1135 -2673
rect -1087 -2677 -1083 -2673
rect -924 -2677 -920 -2673
rect -810 -2677 -806 -2673
rect -758 -2677 -754 -2673
rect -1195 -2684 -1191 -2680
rect -1157 -2684 -1153 -2680
rect -866 -2684 -862 -2680
rect -828 -2684 -824 -2680
rect -1338 -2752 -1334 -2748
rect -934 -2752 -930 -2748
rect -576 -2752 -572 -2748
rect -218 -2752 -214 -2748
rect 210 -2752 214 -2748
rect 566 -2752 570 -2748
rect 964 -2752 968 -2748
rect 1322 -2752 1326 -2748
rect -1327 -2760 -1323 -2756
rect -923 -2760 -919 -2756
rect -565 -2760 -561 -2756
rect -207 -2760 -203 -2756
rect 221 -2760 225 -2756
rect 577 -2760 581 -2756
rect 975 -2760 979 -2756
rect 1333 -2760 1337 -2756
rect -924 -2858 -920 -2854
rect -858 -2858 -854 -2854
rect -824 -2858 -820 -2854
rect -780 -2858 -776 -2854
rect -746 -2858 -742 -2854
rect -566 -2858 -562 -2854
rect -500 -2858 -496 -2854
rect -466 -2858 -462 -2854
rect -422 -2858 -418 -2854
rect -388 -2858 -384 -2854
rect -208 -2858 -204 -2854
rect -142 -2858 -138 -2854
rect -108 -2858 -104 -2854
rect -64 -2858 -60 -2854
rect -30 -2858 -26 -2854
rect 220 -2858 224 -2854
rect 286 -2858 290 -2854
rect 320 -2858 324 -2854
rect 364 -2858 368 -2854
rect 398 -2858 402 -2854
rect 576 -2858 580 -2854
rect 642 -2858 646 -2854
rect 676 -2858 680 -2854
rect 720 -2858 724 -2854
rect 754 -2858 758 -2854
rect 974 -2858 978 -2854
rect 1040 -2858 1044 -2854
rect 1074 -2858 1078 -2854
rect 1118 -2858 1122 -2854
rect 1152 -2858 1156 -2854
rect 1332 -2858 1336 -2854
rect 1398 -2858 1402 -2854
rect 1432 -2858 1436 -2854
rect 1476 -2858 1480 -2854
rect 1510 -2858 1514 -2854
rect -882 -2865 -878 -2861
rect -524 -2865 -520 -2861
rect -166 -2865 -162 -2861
rect 262 -2865 266 -2861
rect 618 -2865 622 -2861
rect 1016 -2865 1020 -2861
rect 1374 -2865 1378 -2861
rect -848 -2872 -844 -2868
rect -706 -2872 -702 -2868
rect -490 -2872 -486 -2868
rect -348 -2872 -344 -2868
rect -132 -2872 -128 -2868
rect 10 -2872 14 -2868
rect 296 -2872 300 -2868
rect 438 -2872 442 -2868
rect 652 -2872 656 -2868
rect 794 -2872 798 -2868
rect 1050 -2872 1054 -2868
rect 1192 -2872 1196 -2868
rect 1408 -2872 1412 -2868
rect 1550 -2872 1554 -2868
rect -928 -2879 -924 -2875
rect -898 -2879 -894 -2875
rect -780 -2879 -776 -2875
rect -570 -2879 -566 -2875
rect -540 -2879 -536 -2875
rect -422 -2879 -418 -2875
rect -212 -2879 -208 -2875
rect -182 -2879 -178 -2875
rect -64 -2879 -60 -2875
rect 216 -2879 220 -2875
rect 246 -2879 250 -2875
rect 364 -2879 368 -2875
rect 572 -2879 576 -2875
rect 602 -2879 606 -2875
rect 720 -2879 724 -2875
rect 970 -2879 974 -2875
rect 1000 -2879 1004 -2875
rect 1118 -2879 1122 -2875
rect 1328 -2879 1332 -2875
rect 1358 -2879 1362 -2875
rect 1476 -2879 1480 -2875
rect -1203 -2888 -1199 -2884
rect -902 -2887 -898 -2883
rect -804 -2887 -800 -2883
rect -544 -2887 -540 -2883
rect -446 -2887 -442 -2883
rect -186 -2887 -182 -2883
rect -88 -2887 -84 -2883
rect 242 -2887 246 -2883
rect 340 -2887 344 -2883
rect 598 -2887 602 -2883
rect 696 -2887 700 -2883
rect 996 -2887 1000 -2883
rect 1094 -2887 1098 -2883
rect 1354 -2887 1358 -2883
rect 1452 -2887 1456 -2883
rect -1253 -2895 -1249 -2891
rect -1213 -2895 -1209 -2891
rect -1193 -2895 -1189 -2891
rect -924 -2894 -920 -2890
rect -776 -2894 -772 -2890
rect -566 -2894 -562 -2890
rect -418 -2894 -414 -2890
rect -208 -2894 -204 -2890
rect -60 -2894 -56 -2890
rect 220 -2894 224 -2890
rect 368 -2894 372 -2890
rect 576 -2894 580 -2890
rect 724 -2894 728 -2890
rect 974 -2894 978 -2890
rect 1122 -2894 1126 -2890
rect 1332 -2894 1336 -2890
rect 1480 -2894 1484 -2890
rect -1257 -2902 -1253 -2898
rect -1227 -2902 -1223 -2898
rect -1179 -2902 -1175 -2898
rect -902 -2901 -898 -2897
rect -794 -2901 -790 -2897
rect -760 -2901 -756 -2897
rect -544 -2901 -540 -2897
rect -436 -2901 -432 -2897
rect -402 -2901 -398 -2897
rect -186 -2901 -182 -2897
rect -78 -2901 -74 -2897
rect -44 -2901 -40 -2897
rect 242 -2901 246 -2897
rect 350 -2901 354 -2897
rect 384 -2901 388 -2897
rect 598 -2901 602 -2897
rect 706 -2901 710 -2897
rect 740 -2901 744 -2897
rect 996 -2901 1000 -2897
rect 1104 -2901 1108 -2897
rect 1138 -2901 1142 -2897
rect 1354 -2901 1358 -2897
rect 1462 -2901 1466 -2897
rect 1496 -2901 1500 -2897
rect -928 -2908 -924 -2904
rect -872 -2908 -868 -2904
rect -838 -2908 -834 -2904
rect -570 -2908 -566 -2904
rect -514 -2908 -510 -2904
rect -480 -2908 -476 -2904
rect -212 -2908 -208 -2904
rect -156 -2908 -152 -2904
rect -122 -2908 -118 -2904
rect 216 -2908 220 -2904
rect 272 -2908 276 -2904
rect 306 -2908 310 -2904
rect 572 -2908 576 -2904
rect 628 -2908 632 -2904
rect 662 -2908 666 -2904
rect 970 -2908 974 -2904
rect 1026 -2908 1030 -2904
rect 1060 -2908 1064 -2904
rect 1328 -2908 1332 -2904
rect 1384 -2908 1388 -2904
rect 1418 -2908 1422 -2904
rect -1237 -3006 -1233 -3002
rect -1199 -3006 -1195 -3002
rect -1139 -3006 -1135 -3002
rect -1115 -3006 -1111 -3002
rect -1257 -3014 -1253 -3010
rect -1223 -3014 -1219 -3010
rect -1171 -3014 -1167 -3010
rect -1111 -3014 -1107 -3010
rect -1073 -3014 -1069 -3010
rect -1025 -3011 -1021 -3001
rect -908 -3006 -904 -3002
rect -870 -3006 -866 -3002
rect -810 -3006 -806 -3002
rect -786 -3006 -782 -3002
rect -671 -3010 -667 -3000
rect -550 -3006 -546 -3002
rect -512 -3006 -508 -3002
rect -452 -3006 -448 -3002
rect -428 -3006 -424 -3002
rect -928 -3014 -924 -3010
rect -894 -3014 -890 -3010
rect -842 -3014 -838 -3010
rect -782 -3014 -778 -3010
rect -744 -3014 -740 -3010
rect -570 -3014 -566 -3010
rect -536 -3014 -532 -3010
rect -484 -3014 -480 -3010
rect -424 -3014 -420 -3010
rect -386 -3014 -382 -3010
rect -328 -3012 -324 -3002
rect -192 -3006 -188 -3002
rect -154 -3006 -150 -3002
rect -94 -3006 -90 -3002
rect -70 -3006 -66 -3002
rect 236 -3006 240 -3002
rect 274 -3006 278 -3002
rect 334 -3006 338 -3002
rect 358 -3006 362 -3002
rect 473 -3010 477 -3000
rect 842 -3010 846 -3000
rect -212 -3014 -208 -3010
rect -178 -3014 -174 -3010
rect -126 -3014 -122 -3010
rect -66 -3014 -62 -3010
rect -28 -3014 -24 -3010
rect 216 -3014 220 -3010
rect 250 -3014 254 -3010
rect 302 -3014 306 -3010
rect 362 -3014 366 -3010
rect 400 -3014 404 -3010
rect 1200 -3011 1204 -3001
rect -1213 -3021 -1209 -3017
rect -1181 -3021 -1177 -3017
rect -1129 -3021 -1125 -3017
rect -1097 -3021 -1093 -3017
rect -884 -3021 -880 -3017
rect -852 -3021 -848 -3017
rect -800 -3021 -796 -3017
rect -768 -3021 -764 -3017
rect -526 -3021 -522 -3017
rect -494 -3021 -490 -3017
rect -442 -3021 -438 -3017
rect -410 -3021 -406 -3017
rect -168 -3021 -164 -3017
rect -136 -3021 -132 -3017
rect -84 -3021 -80 -3017
rect -52 -3021 -48 -3017
rect 260 -3021 264 -3017
rect 292 -3021 296 -3017
rect 344 -3021 348 -3017
rect 376 -3021 380 -3017
rect -1253 -3028 -1249 -3024
rect -1139 -3028 -1135 -3024
rect -1087 -3028 -1083 -3024
rect -924 -3028 -920 -3024
rect -810 -3028 -806 -3024
rect -758 -3028 -754 -3024
rect -566 -3028 -562 -3024
rect -452 -3028 -448 -3024
rect -400 -3028 -396 -3024
rect -208 -3028 -204 -3024
rect -94 -3028 -90 -3024
rect -42 -3028 -38 -3024
rect 220 -3028 224 -3024
rect 334 -3028 338 -3024
rect 386 -3028 390 -3024
rect -1195 -3035 -1191 -3031
rect -1157 -3035 -1153 -3031
rect -866 -3035 -862 -3031
rect -828 -3035 -824 -3031
rect -508 -3035 -504 -3031
rect -470 -3035 -466 -3031
rect -150 -3035 -146 -3031
rect -112 -3035 -108 -3031
rect 278 -3035 282 -3031
rect 316 -3035 320 -3031
rect -1237 -3122 -1233 -3118
rect -1199 -3122 -1195 -3118
rect -1139 -3122 -1135 -3118
rect -1115 -3122 -1111 -3118
rect -1025 -3126 -1021 -3116
rect -908 -3122 -904 -3118
rect -870 -3122 -866 -3118
rect -810 -3122 -806 -3118
rect -786 -3122 -782 -3118
rect -550 -3122 -546 -3118
rect -512 -3122 -508 -3118
rect -452 -3122 -448 -3118
rect -428 -3122 -424 -3118
rect -1257 -3130 -1253 -3126
rect -1223 -3130 -1219 -3126
rect -1171 -3130 -1167 -3126
rect -1111 -3130 -1107 -3126
rect -1073 -3130 -1069 -3126
rect -928 -3130 -924 -3126
rect -894 -3130 -890 -3126
rect -842 -3130 -838 -3126
rect -782 -3130 -778 -3126
rect -744 -3130 -740 -3126
rect -570 -3130 -566 -3126
rect -536 -3130 -532 -3126
rect -484 -3130 -480 -3126
rect -424 -3130 -420 -3126
rect -386 -3130 -382 -3126
rect -328 -3127 -324 -3117
rect -192 -3122 -188 -3118
rect -154 -3122 -150 -3118
rect -94 -3122 -90 -3118
rect -70 -3122 -66 -3118
rect 236 -3122 240 -3118
rect 274 -3122 278 -3118
rect 334 -3122 338 -3118
rect 358 -3122 362 -3118
rect 473 -3126 477 -3116
rect 592 -3122 596 -3118
rect 630 -3122 634 -3118
rect 690 -3122 694 -3118
rect 714 -3122 718 -3118
rect 990 -3122 994 -3118
rect 1028 -3122 1032 -3118
rect 1088 -3122 1092 -3118
rect 1112 -3122 1116 -3118
rect 1200 -3126 1204 -3116
rect 1348 -3122 1352 -3118
rect 1386 -3122 1390 -3118
rect 1446 -3122 1450 -3118
rect 1470 -3122 1474 -3118
rect -212 -3130 -208 -3126
rect -178 -3130 -174 -3126
rect -126 -3130 -122 -3126
rect -66 -3130 -62 -3126
rect -28 -3130 -24 -3126
rect 216 -3130 220 -3126
rect 250 -3130 254 -3126
rect 302 -3130 306 -3126
rect 362 -3130 366 -3126
rect 400 -3130 404 -3126
rect 572 -3130 576 -3126
rect 606 -3130 610 -3126
rect 658 -3130 662 -3126
rect 718 -3130 722 -3126
rect 756 -3130 760 -3126
rect 970 -3130 974 -3126
rect 1004 -3130 1008 -3126
rect 1056 -3130 1060 -3126
rect 1116 -3130 1120 -3126
rect 1154 -3130 1158 -3126
rect 1328 -3130 1332 -3126
rect 1362 -3130 1366 -3126
rect 1414 -3130 1418 -3126
rect 1474 -3130 1478 -3126
rect 1512 -3130 1516 -3126
rect -1213 -3137 -1209 -3133
rect -1181 -3137 -1177 -3133
rect -1129 -3137 -1125 -3133
rect -1097 -3137 -1093 -3133
rect -884 -3137 -880 -3133
rect -852 -3137 -848 -3133
rect -800 -3137 -796 -3133
rect -768 -3137 -764 -3133
rect -526 -3137 -522 -3133
rect -494 -3137 -490 -3133
rect -442 -3137 -438 -3133
rect -410 -3137 -406 -3133
rect -168 -3137 -164 -3133
rect -136 -3137 -132 -3133
rect -84 -3137 -80 -3133
rect -52 -3137 -48 -3133
rect 260 -3137 264 -3133
rect 292 -3137 296 -3133
rect 344 -3137 348 -3133
rect 376 -3137 380 -3133
rect 616 -3137 620 -3133
rect 648 -3137 652 -3133
rect 700 -3137 704 -3133
rect 732 -3137 736 -3133
rect 1014 -3137 1018 -3133
rect 1046 -3137 1050 -3133
rect 1098 -3137 1102 -3133
rect 1130 -3137 1134 -3133
rect 1372 -3137 1376 -3133
rect 1404 -3137 1408 -3133
rect 1456 -3137 1460 -3133
rect 1488 -3137 1492 -3133
rect -1253 -3144 -1249 -3140
rect -1139 -3144 -1135 -3140
rect -1087 -3144 -1083 -3140
rect -924 -3144 -920 -3140
rect -810 -3144 -806 -3140
rect -758 -3144 -754 -3140
rect -566 -3144 -562 -3140
rect -452 -3144 -448 -3140
rect -400 -3144 -396 -3140
rect -208 -3144 -204 -3140
rect -94 -3144 -90 -3140
rect -42 -3144 -38 -3140
rect 220 -3144 224 -3140
rect 334 -3144 338 -3140
rect 386 -3144 390 -3140
rect 576 -3144 580 -3140
rect 690 -3144 694 -3140
rect 742 -3144 746 -3140
rect 974 -3144 978 -3140
rect 1088 -3144 1092 -3140
rect 1140 -3144 1144 -3140
rect 1332 -3144 1336 -3140
rect 1446 -3144 1450 -3140
rect 1498 -3144 1502 -3140
rect -1195 -3151 -1191 -3147
rect -1157 -3151 -1153 -3147
rect -866 -3151 -862 -3147
rect -828 -3151 -824 -3147
rect -508 -3151 -504 -3147
rect -470 -3151 -466 -3147
rect -150 -3151 -146 -3147
rect -112 -3151 -108 -3147
rect 278 -3151 282 -3147
rect 316 -3151 320 -3147
rect 634 -3151 638 -3147
rect 672 -3151 676 -3147
rect 1032 -3151 1036 -3147
rect 1070 -3151 1074 -3147
rect 1390 -3151 1394 -3147
rect 1428 -3151 1432 -3147
rect -1237 -3243 -1233 -3239
rect -1199 -3243 -1195 -3239
rect -1139 -3243 -1135 -3239
rect -1115 -3243 -1111 -3239
rect -908 -3243 -904 -3239
rect -870 -3243 -866 -3239
rect -810 -3243 -806 -3239
rect -786 -3243 -782 -3239
rect -550 -3243 -546 -3239
rect -512 -3243 -508 -3239
rect -452 -3243 -448 -3239
rect -428 -3243 -424 -3239
rect -192 -3243 -188 -3239
rect -154 -3243 -150 -3239
rect -94 -3243 -90 -3239
rect -70 -3243 -66 -3239
rect 236 -3243 240 -3239
rect 274 -3243 278 -3239
rect 334 -3243 338 -3239
rect 358 -3243 362 -3239
rect 592 -3243 596 -3239
rect 630 -3243 634 -3239
rect 690 -3243 694 -3239
rect 714 -3243 718 -3239
rect 990 -3243 994 -3239
rect 1028 -3243 1032 -3239
rect 1088 -3243 1092 -3239
rect 1112 -3243 1116 -3239
rect 1348 -3243 1352 -3239
rect 1386 -3243 1390 -3239
rect 1446 -3243 1450 -3239
rect 1470 -3243 1474 -3239
rect -1257 -3251 -1253 -3247
rect -1223 -3251 -1219 -3247
rect -1171 -3251 -1167 -3247
rect -1111 -3251 -1107 -3247
rect -1073 -3251 -1069 -3247
rect -928 -3251 -924 -3247
rect -894 -3251 -890 -3247
rect -842 -3251 -838 -3247
rect -782 -3251 -778 -3247
rect -744 -3251 -740 -3247
rect -570 -3251 -566 -3247
rect -536 -3251 -532 -3247
rect -484 -3251 -480 -3247
rect -424 -3251 -420 -3247
rect -386 -3251 -382 -3247
rect -212 -3251 -208 -3247
rect -178 -3251 -174 -3247
rect -126 -3251 -122 -3247
rect -66 -3251 -62 -3247
rect -28 -3251 -24 -3247
rect 216 -3251 220 -3247
rect 250 -3251 254 -3247
rect 302 -3251 306 -3247
rect 362 -3251 366 -3247
rect 400 -3251 404 -3247
rect 572 -3251 576 -3247
rect 606 -3251 610 -3247
rect 658 -3251 662 -3247
rect 718 -3251 722 -3247
rect 756 -3251 760 -3247
rect 970 -3251 974 -3247
rect 1004 -3251 1008 -3247
rect 1056 -3251 1060 -3247
rect 1116 -3251 1120 -3247
rect 1154 -3251 1158 -3247
rect 1328 -3251 1332 -3247
rect 1362 -3251 1366 -3247
rect 1414 -3251 1418 -3247
rect 1474 -3251 1478 -3247
rect 1512 -3251 1516 -3247
rect -1213 -3258 -1209 -3254
rect -1181 -3258 -1177 -3254
rect -1129 -3258 -1125 -3254
rect -1097 -3258 -1093 -3254
rect -884 -3258 -880 -3254
rect -852 -3258 -848 -3254
rect -800 -3258 -796 -3254
rect -768 -3258 -764 -3254
rect -526 -3258 -522 -3254
rect -494 -3258 -490 -3254
rect -442 -3258 -438 -3254
rect -410 -3258 -406 -3254
rect -168 -3258 -164 -3254
rect -136 -3258 -132 -3254
rect -84 -3258 -80 -3254
rect -52 -3258 -48 -3254
rect 260 -3258 264 -3254
rect 292 -3258 296 -3254
rect 344 -3258 348 -3254
rect 376 -3258 380 -3254
rect 616 -3258 620 -3254
rect 648 -3258 652 -3254
rect 700 -3258 704 -3254
rect 732 -3258 736 -3254
rect 1014 -3258 1018 -3254
rect 1046 -3258 1050 -3254
rect 1098 -3258 1102 -3254
rect 1130 -3258 1134 -3254
rect 1372 -3258 1376 -3254
rect 1404 -3258 1408 -3254
rect 1456 -3258 1460 -3254
rect 1488 -3258 1492 -3254
rect -1253 -3265 -1249 -3261
rect -1139 -3265 -1135 -3261
rect -1087 -3265 -1083 -3261
rect -924 -3265 -920 -3261
rect -810 -3265 -806 -3261
rect -758 -3265 -754 -3261
rect -566 -3265 -562 -3261
rect -452 -3265 -448 -3261
rect -400 -3265 -396 -3261
rect -208 -3265 -204 -3261
rect -94 -3265 -90 -3261
rect -42 -3265 -38 -3261
rect 220 -3265 224 -3261
rect 334 -3265 338 -3261
rect 386 -3265 390 -3261
rect 576 -3265 580 -3261
rect 690 -3265 694 -3261
rect 742 -3265 746 -3261
rect 974 -3265 978 -3261
rect 1088 -3265 1092 -3261
rect 1140 -3265 1144 -3261
rect 1332 -3265 1336 -3261
rect 1446 -3265 1450 -3261
rect 1498 -3265 1502 -3261
rect -1195 -3272 -1191 -3268
rect -1157 -3272 -1153 -3268
rect -866 -3272 -862 -3268
rect -828 -3272 -824 -3268
rect -508 -3272 -504 -3268
rect -470 -3272 -466 -3268
rect -150 -3272 -146 -3268
rect -112 -3272 -108 -3268
rect 278 -3272 282 -3268
rect 316 -3272 320 -3268
rect 634 -3272 638 -3268
rect 672 -3272 676 -3268
rect 1032 -3272 1036 -3268
rect 1070 -3272 1074 -3268
rect 1390 -3272 1394 -3268
rect 1428 -3272 1432 -3268
rect -1237 -3357 -1233 -3353
rect -1199 -3357 -1195 -3353
rect -1139 -3357 -1135 -3353
rect -1115 -3357 -1111 -3353
rect -908 -3357 -904 -3353
rect -870 -3357 -866 -3353
rect -810 -3357 -806 -3353
rect -786 -3357 -782 -3353
rect -550 -3357 -546 -3353
rect -512 -3357 -508 -3353
rect -452 -3357 -448 -3353
rect -428 -3357 -424 -3353
rect -1257 -3365 -1253 -3361
rect -1223 -3365 -1219 -3361
rect -1171 -3365 -1167 -3361
rect -1111 -3365 -1107 -3361
rect -1073 -3365 -1069 -3361
rect -928 -3365 -924 -3361
rect -894 -3365 -890 -3361
rect -842 -3365 -838 -3361
rect -782 -3365 -778 -3361
rect -744 -3365 -740 -3361
rect -570 -3365 -566 -3361
rect -536 -3365 -532 -3361
rect -484 -3365 -480 -3361
rect -424 -3365 -420 -3361
rect -386 -3365 -382 -3361
rect -1213 -3372 -1209 -3368
rect -1181 -3372 -1177 -3368
rect -1129 -3372 -1125 -3368
rect -1097 -3372 -1093 -3368
rect -884 -3372 -880 -3368
rect -852 -3372 -848 -3368
rect -800 -3372 -796 -3368
rect -768 -3372 -764 -3368
rect -526 -3372 -522 -3368
rect -494 -3372 -490 -3368
rect -442 -3372 -438 -3368
rect -410 -3372 -406 -3368
rect -1253 -3379 -1249 -3375
rect -1139 -3379 -1135 -3375
rect -1087 -3379 -1083 -3375
rect -924 -3379 -920 -3375
rect -810 -3379 -806 -3375
rect -758 -3379 -754 -3375
rect -566 -3379 -562 -3375
rect -452 -3379 -448 -3375
rect -400 -3379 -396 -3375
rect -1195 -3386 -1191 -3382
rect -1157 -3386 -1153 -3382
rect -866 -3386 -862 -3382
rect -828 -3386 -824 -3382
rect -508 -3386 -504 -3382
rect -470 -3386 -466 -3382
rect -1338 -3458 -1334 -3454
rect -934 -3458 -930 -3454
rect -576 -3458 -572 -3454
rect -218 -3458 -214 -3454
rect 210 -3458 214 -3454
rect 566 -3458 570 -3454
rect 964 -3458 968 -3454
rect 1322 -3458 1326 -3454
rect -1327 -3466 -1323 -3462
rect -923 -3466 -919 -3462
rect -565 -3466 -561 -3462
rect -207 -3466 -203 -3462
rect 221 -3466 225 -3462
rect 577 -3466 581 -3462
rect 975 -3466 979 -3462
rect 1333 -3466 1337 -3462
rect -924 -3569 -920 -3565
rect -858 -3569 -854 -3565
rect -824 -3569 -820 -3565
rect -780 -3569 -776 -3565
rect -746 -3569 -742 -3565
rect -566 -3569 -562 -3565
rect -500 -3569 -496 -3565
rect -466 -3569 -462 -3565
rect -422 -3569 -418 -3565
rect -388 -3569 -384 -3565
rect -208 -3569 -204 -3565
rect -142 -3569 -138 -3565
rect -108 -3569 -104 -3565
rect -64 -3569 -60 -3565
rect -30 -3569 -26 -3565
rect 220 -3569 224 -3565
rect 286 -3569 290 -3565
rect 320 -3569 324 -3565
rect 364 -3569 368 -3565
rect 398 -3569 402 -3565
rect 576 -3569 580 -3565
rect 642 -3569 646 -3565
rect 676 -3569 680 -3565
rect 720 -3569 724 -3565
rect 754 -3569 758 -3565
rect 974 -3569 978 -3565
rect 1040 -3569 1044 -3565
rect 1074 -3569 1078 -3565
rect 1118 -3569 1122 -3565
rect 1152 -3569 1156 -3565
rect 1332 -3569 1336 -3565
rect 1398 -3569 1402 -3565
rect 1432 -3569 1436 -3565
rect 1476 -3569 1480 -3565
rect 1510 -3569 1514 -3565
rect -882 -3576 -878 -3572
rect -524 -3576 -520 -3572
rect -166 -3576 -162 -3572
rect 262 -3576 266 -3572
rect 618 -3576 622 -3572
rect 1016 -3576 1020 -3572
rect 1374 -3576 1378 -3572
rect -848 -3583 -844 -3579
rect -706 -3583 -702 -3579
rect -490 -3583 -486 -3579
rect -348 -3583 -344 -3579
rect -132 -3583 -128 -3579
rect 10 -3583 14 -3579
rect 296 -3583 300 -3579
rect 438 -3583 442 -3579
rect 652 -3583 656 -3579
rect 794 -3583 798 -3579
rect 1050 -3583 1054 -3579
rect 1192 -3583 1196 -3579
rect 1408 -3583 1412 -3579
rect 1550 -3583 1554 -3579
rect -928 -3590 -924 -3586
rect -898 -3590 -894 -3586
rect -780 -3590 -776 -3586
rect -570 -3590 -566 -3586
rect -540 -3590 -536 -3586
rect -422 -3590 -418 -3586
rect -212 -3590 -208 -3586
rect -182 -3590 -178 -3586
rect -64 -3590 -60 -3586
rect 216 -3590 220 -3586
rect 246 -3590 250 -3586
rect 364 -3590 368 -3586
rect 572 -3590 576 -3586
rect 602 -3590 606 -3586
rect 720 -3590 724 -3586
rect 970 -3590 974 -3586
rect 1000 -3590 1004 -3586
rect 1118 -3590 1122 -3586
rect 1328 -3590 1332 -3586
rect 1358 -3590 1362 -3586
rect 1476 -3590 1480 -3586
rect -1203 -3599 -1199 -3595
rect -902 -3598 -898 -3594
rect -804 -3598 -800 -3594
rect -544 -3598 -540 -3594
rect -446 -3598 -442 -3594
rect -186 -3598 -182 -3594
rect -88 -3598 -84 -3594
rect 242 -3598 246 -3594
rect 340 -3598 344 -3594
rect 598 -3598 602 -3594
rect 696 -3598 700 -3594
rect 996 -3598 1000 -3594
rect 1094 -3598 1098 -3594
rect 1354 -3598 1358 -3594
rect 1452 -3598 1456 -3594
rect -1253 -3606 -1249 -3602
rect -1213 -3606 -1209 -3602
rect -1193 -3606 -1189 -3602
rect -924 -3605 -920 -3601
rect -776 -3605 -772 -3601
rect -566 -3605 -562 -3601
rect -418 -3605 -414 -3601
rect -208 -3605 -204 -3601
rect -60 -3605 -56 -3601
rect 220 -3605 224 -3601
rect 368 -3605 372 -3601
rect 576 -3605 580 -3601
rect 724 -3605 728 -3601
rect 974 -3605 978 -3601
rect 1122 -3605 1126 -3601
rect 1332 -3605 1336 -3601
rect 1480 -3605 1484 -3601
rect -1257 -3613 -1253 -3609
rect -1227 -3613 -1223 -3609
rect -1179 -3613 -1175 -3609
rect -902 -3612 -898 -3608
rect -794 -3612 -790 -3608
rect -760 -3612 -756 -3608
rect -544 -3612 -540 -3608
rect -436 -3612 -432 -3608
rect -402 -3612 -398 -3608
rect -186 -3612 -182 -3608
rect -78 -3612 -74 -3608
rect -44 -3612 -40 -3608
rect 242 -3612 246 -3608
rect 350 -3612 354 -3608
rect 384 -3612 388 -3608
rect 598 -3612 602 -3608
rect 706 -3612 710 -3608
rect 740 -3612 744 -3608
rect 996 -3612 1000 -3608
rect 1104 -3612 1108 -3608
rect 1138 -3612 1142 -3608
rect 1354 -3612 1358 -3608
rect 1462 -3612 1466 -3608
rect 1496 -3612 1500 -3608
rect -928 -3619 -924 -3615
rect -872 -3619 -868 -3615
rect -838 -3619 -834 -3615
rect -570 -3619 -566 -3615
rect -514 -3619 -510 -3615
rect -480 -3619 -476 -3615
rect -212 -3619 -208 -3615
rect -156 -3619 -152 -3615
rect -122 -3619 -118 -3615
rect 216 -3619 220 -3615
rect 272 -3619 276 -3615
rect 306 -3619 310 -3615
rect 572 -3619 576 -3615
rect 628 -3619 632 -3615
rect 662 -3619 666 -3615
rect 970 -3619 974 -3615
rect 1026 -3619 1030 -3615
rect 1060 -3619 1064 -3615
rect 1328 -3619 1332 -3615
rect 1384 -3619 1388 -3615
rect 1418 -3619 1422 -3615
rect -1237 -3728 -1233 -3724
rect -1199 -3728 -1195 -3724
rect -1139 -3728 -1135 -3724
rect -1115 -3728 -1111 -3724
rect -908 -3728 -904 -3724
rect -870 -3728 -866 -3724
rect -810 -3728 -806 -3724
rect -786 -3728 -782 -3724
rect -550 -3728 -546 -3724
rect -512 -3728 -508 -3724
rect -452 -3728 -448 -3724
rect -428 -3728 -424 -3724
rect -192 -3728 -188 -3724
rect -154 -3728 -150 -3724
rect -94 -3728 -90 -3724
rect -70 -3728 -66 -3724
rect -1257 -3736 -1253 -3732
rect -1223 -3736 -1219 -3732
rect -1171 -3736 -1167 -3732
rect -1111 -3736 -1107 -3732
rect -1073 -3736 -1069 -3732
rect -928 -3736 -924 -3732
rect -894 -3736 -890 -3732
rect -842 -3736 -838 -3732
rect -782 -3736 -778 -3732
rect -744 -3736 -740 -3732
rect -570 -3736 -566 -3732
rect -536 -3736 -532 -3732
rect -484 -3736 -480 -3732
rect -424 -3736 -420 -3732
rect -386 -3736 -382 -3732
rect -212 -3736 -208 -3732
rect -178 -3736 -174 -3732
rect -126 -3736 -122 -3732
rect -66 -3736 -62 -3732
rect -28 -3736 -24 -3732
rect -1213 -3743 -1209 -3739
rect -1181 -3743 -1177 -3739
rect -1129 -3743 -1125 -3739
rect -1097 -3743 -1093 -3739
rect -884 -3743 -880 -3739
rect -852 -3743 -848 -3739
rect -800 -3743 -796 -3739
rect -768 -3743 -764 -3739
rect -526 -3743 -522 -3739
rect -494 -3743 -490 -3739
rect -442 -3743 -438 -3739
rect -410 -3743 -406 -3739
rect -168 -3743 -164 -3739
rect -136 -3743 -132 -3739
rect -84 -3743 -80 -3739
rect -52 -3743 -48 -3739
rect -1253 -3750 -1249 -3746
rect -1139 -3750 -1135 -3746
rect -1087 -3750 -1083 -3746
rect -924 -3750 -920 -3746
rect -810 -3750 -806 -3746
rect -758 -3750 -754 -3746
rect -566 -3750 -562 -3746
rect -452 -3750 -448 -3746
rect -400 -3750 -396 -3746
rect -208 -3750 -204 -3746
rect -94 -3750 -90 -3746
rect -42 -3750 -38 -3746
rect -1195 -3757 -1191 -3753
rect -1157 -3757 -1153 -3753
rect -866 -3757 -862 -3753
rect -828 -3757 -824 -3753
rect -508 -3757 -504 -3753
rect -470 -3757 -466 -3753
rect -150 -3757 -146 -3753
rect -112 -3757 -108 -3753
rect 69 -3852 73 -3836
rect -1237 -3959 -1233 -3955
rect -1199 -3959 -1195 -3955
rect -1139 -3959 -1135 -3955
rect -1115 -3959 -1111 -3955
rect -908 -3959 -904 -3955
rect -870 -3959 -866 -3955
rect -810 -3959 -806 -3955
rect -786 -3959 -782 -3955
rect -550 -3959 -546 -3955
rect -512 -3959 -508 -3955
rect -452 -3959 -448 -3955
rect -428 -3959 -424 -3955
rect -192 -3959 -188 -3955
rect -154 -3959 -150 -3955
rect -94 -3959 -90 -3955
rect -70 -3959 -66 -3955
rect 236 -3959 240 -3955
rect 274 -3959 278 -3955
rect 334 -3959 338 -3955
rect 358 -3959 362 -3955
rect 592 -3959 596 -3955
rect 630 -3959 634 -3955
rect 690 -3959 694 -3955
rect 714 -3959 718 -3955
rect 990 -3959 994 -3955
rect 1028 -3959 1032 -3955
rect 1088 -3959 1092 -3955
rect 1112 -3959 1116 -3955
rect 1348 -3959 1352 -3955
rect 1386 -3959 1390 -3955
rect 1446 -3959 1450 -3955
rect 1470 -3959 1474 -3955
rect -1257 -3967 -1253 -3963
rect -1223 -3967 -1219 -3963
rect -1171 -3967 -1167 -3963
rect -1111 -3967 -1107 -3963
rect -1073 -3967 -1069 -3963
rect -928 -3967 -924 -3963
rect -894 -3967 -890 -3963
rect -842 -3967 -838 -3963
rect -782 -3967 -778 -3963
rect -744 -3967 -740 -3963
rect -570 -3967 -566 -3963
rect -536 -3967 -532 -3963
rect -484 -3967 -480 -3963
rect -424 -3967 -420 -3963
rect -386 -3967 -382 -3963
rect -212 -3967 -208 -3963
rect -178 -3967 -174 -3963
rect -126 -3967 -122 -3963
rect -66 -3967 -62 -3963
rect -28 -3967 -24 -3963
rect 216 -3967 220 -3963
rect 250 -3967 254 -3963
rect 302 -3967 306 -3963
rect 362 -3967 366 -3963
rect 400 -3967 404 -3963
rect 572 -3967 576 -3963
rect 606 -3967 610 -3963
rect 658 -3967 662 -3963
rect 718 -3967 722 -3963
rect 756 -3967 760 -3963
rect 970 -3967 974 -3963
rect 1004 -3967 1008 -3963
rect 1056 -3967 1060 -3963
rect 1116 -3967 1120 -3963
rect 1154 -3967 1158 -3963
rect 1328 -3967 1332 -3963
rect 1362 -3967 1366 -3963
rect 1414 -3967 1418 -3963
rect 1474 -3967 1478 -3963
rect 1512 -3967 1516 -3963
rect -1213 -3974 -1209 -3970
rect -1181 -3974 -1177 -3970
rect -1129 -3974 -1125 -3970
rect -1097 -3974 -1093 -3970
rect -884 -3974 -880 -3970
rect -852 -3974 -848 -3970
rect -800 -3974 -796 -3970
rect -768 -3974 -764 -3970
rect -526 -3974 -522 -3970
rect -494 -3974 -490 -3970
rect -442 -3974 -438 -3970
rect -410 -3974 -406 -3970
rect -168 -3974 -164 -3970
rect -136 -3974 -132 -3970
rect -84 -3974 -80 -3970
rect -52 -3974 -48 -3970
rect 260 -3974 264 -3970
rect 292 -3974 296 -3970
rect 344 -3974 348 -3970
rect 376 -3974 380 -3970
rect 616 -3974 620 -3970
rect 648 -3974 652 -3970
rect 700 -3974 704 -3970
rect 732 -3974 736 -3970
rect 1014 -3974 1018 -3970
rect 1046 -3974 1050 -3970
rect 1098 -3974 1102 -3970
rect 1130 -3974 1134 -3970
rect 1372 -3974 1376 -3970
rect 1404 -3974 1408 -3970
rect 1456 -3974 1460 -3970
rect 1488 -3974 1492 -3970
rect -1253 -3981 -1249 -3977
rect -1139 -3981 -1135 -3977
rect -1087 -3981 -1083 -3977
rect -924 -3981 -920 -3977
rect -810 -3981 -806 -3977
rect -758 -3981 -754 -3977
rect -566 -3981 -562 -3977
rect -452 -3981 -448 -3977
rect -400 -3981 -396 -3977
rect -208 -3981 -204 -3977
rect -94 -3981 -90 -3977
rect -42 -3981 -38 -3977
rect 220 -3981 224 -3977
rect 334 -3981 338 -3977
rect 386 -3981 390 -3977
rect 576 -3981 580 -3977
rect 690 -3981 694 -3977
rect 742 -3981 746 -3977
rect 974 -3981 978 -3977
rect 1088 -3981 1092 -3977
rect 1140 -3981 1144 -3977
rect 1332 -3981 1336 -3977
rect 1446 -3981 1450 -3977
rect 1498 -3981 1502 -3977
rect -1195 -3988 -1191 -3984
rect -1157 -3988 -1153 -3984
rect -866 -3988 -862 -3984
rect -828 -3988 -824 -3984
rect -508 -3988 -504 -3984
rect -470 -3988 -466 -3984
rect -150 -3988 -146 -3984
rect -112 -3988 -108 -3984
rect 278 -3988 282 -3984
rect 316 -3988 320 -3984
rect 634 -3988 638 -3984
rect 672 -3988 676 -3984
rect 1032 -3988 1036 -3984
rect 1070 -3988 1074 -3984
rect 1390 -3988 1394 -3984
rect 1428 -3988 1432 -3984
rect -1237 -4084 -1233 -4080
rect -1199 -4084 -1195 -4080
rect -1139 -4084 -1135 -4080
rect -1115 -4084 -1111 -4080
rect -908 -4084 -904 -4080
rect -870 -4084 -866 -4080
rect -810 -4084 -806 -4080
rect -786 -4084 -782 -4080
rect -550 -4084 -546 -4080
rect -512 -4084 -508 -4080
rect -452 -4084 -448 -4080
rect -428 -4084 -424 -4080
rect -192 -4084 -188 -4080
rect -154 -4084 -150 -4080
rect -94 -4084 -90 -4080
rect -70 -4084 -66 -4080
rect 236 -4084 240 -4080
rect 274 -4084 278 -4080
rect 334 -4084 338 -4080
rect 358 -4084 362 -4080
rect 592 -4084 596 -4080
rect 630 -4084 634 -4080
rect 690 -4084 694 -4080
rect 714 -4084 718 -4080
rect 990 -4084 994 -4080
rect 1028 -4084 1032 -4080
rect 1088 -4084 1092 -4080
rect 1112 -4084 1116 -4080
rect 1348 -4084 1352 -4080
rect 1386 -4084 1390 -4080
rect 1446 -4084 1450 -4080
rect 1470 -4084 1474 -4080
rect -1257 -4092 -1253 -4088
rect -1223 -4092 -1219 -4088
rect -1171 -4092 -1167 -4088
rect -1111 -4092 -1107 -4088
rect -1073 -4092 -1069 -4088
rect -928 -4092 -924 -4088
rect -894 -4092 -890 -4088
rect -842 -4092 -838 -4088
rect -782 -4092 -778 -4088
rect -744 -4092 -740 -4088
rect -570 -4092 -566 -4088
rect -536 -4092 -532 -4088
rect -484 -4092 -480 -4088
rect -424 -4092 -420 -4088
rect -386 -4092 -382 -4088
rect -212 -4092 -208 -4088
rect -178 -4092 -174 -4088
rect -126 -4092 -122 -4088
rect -66 -4092 -62 -4088
rect -28 -4092 -24 -4088
rect 216 -4092 220 -4088
rect 250 -4092 254 -4088
rect 302 -4092 306 -4088
rect 362 -4092 366 -4088
rect 400 -4092 404 -4088
rect 572 -4092 576 -4088
rect 606 -4092 610 -4088
rect 658 -4092 662 -4088
rect 718 -4092 722 -4088
rect 756 -4092 760 -4088
rect 970 -4092 974 -4088
rect 1004 -4092 1008 -4088
rect 1056 -4092 1060 -4088
rect 1116 -4092 1120 -4088
rect 1154 -4092 1158 -4088
rect 1328 -4092 1332 -4088
rect 1362 -4092 1366 -4088
rect 1414 -4092 1418 -4088
rect 1474 -4092 1478 -4088
rect 1512 -4092 1516 -4088
rect -1213 -4099 -1209 -4095
rect -1181 -4099 -1177 -4095
rect -1129 -4099 -1125 -4095
rect -1097 -4099 -1093 -4095
rect -884 -4099 -880 -4095
rect -852 -4099 -848 -4095
rect -800 -4099 -796 -4095
rect -768 -4099 -764 -4095
rect -526 -4099 -522 -4095
rect -494 -4099 -490 -4095
rect -442 -4099 -438 -4095
rect -410 -4099 -406 -4095
rect -168 -4099 -164 -4095
rect -136 -4099 -132 -4095
rect -84 -4099 -80 -4095
rect -52 -4099 -48 -4095
rect 260 -4099 264 -4095
rect 292 -4099 296 -4095
rect 344 -4099 348 -4095
rect 376 -4099 380 -4095
rect 616 -4099 620 -4095
rect 648 -4099 652 -4095
rect 700 -4099 704 -4095
rect 732 -4099 736 -4095
rect 1014 -4099 1018 -4095
rect 1046 -4099 1050 -4095
rect 1098 -4099 1102 -4095
rect 1130 -4099 1134 -4095
rect 1372 -4099 1376 -4095
rect 1404 -4099 1408 -4095
rect 1456 -4099 1460 -4095
rect 1488 -4099 1492 -4095
rect -1253 -4106 -1249 -4102
rect -1139 -4106 -1135 -4102
rect -1087 -4106 -1083 -4102
rect -924 -4106 -920 -4102
rect -810 -4106 -806 -4102
rect -758 -4106 -754 -4102
rect -566 -4106 -562 -4102
rect -452 -4106 -448 -4102
rect -400 -4106 -396 -4102
rect -208 -4106 -204 -4102
rect -94 -4106 -90 -4102
rect -42 -4106 -38 -4102
rect 220 -4106 224 -4102
rect 334 -4106 338 -4102
rect 386 -4106 390 -4102
rect 576 -4106 580 -4102
rect 690 -4106 694 -4102
rect 742 -4106 746 -4102
rect 974 -4106 978 -4102
rect 1088 -4106 1092 -4102
rect 1140 -4106 1144 -4102
rect 1332 -4106 1336 -4102
rect 1446 -4106 1450 -4102
rect 1498 -4106 1502 -4102
rect -1195 -4113 -1191 -4109
rect -1157 -4113 -1153 -4109
rect -866 -4113 -862 -4109
rect -828 -4113 -824 -4109
rect -508 -4113 -504 -4109
rect -470 -4113 -466 -4109
rect -150 -4113 -146 -4109
rect -112 -4113 -108 -4109
rect 278 -4113 282 -4109
rect 316 -4113 320 -4109
rect 634 -4113 638 -4109
rect 672 -4113 676 -4109
rect 1032 -4113 1036 -4109
rect 1070 -4113 1074 -4109
rect 1390 -4113 1394 -4109
rect 1428 -4113 1432 -4109
rect -1237 -4208 -1233 -4204
rect -1199 -4208 -1195 -4204
rect -1139 -4208 -1135 -4204
rect -1115 -4208 -1111 -4204
rect -1028 -4208 -1024 -4198
rect -908 -4208 -904 -4204
rect -870 -4208 -866 -4204
rect -810 -4208 -806 -4204
rect -786 -4208 -782 -4204
rect -550 -4208 -546 -4204
rect -512 -4208 -508 -4204
rect -452 -4208 -448 -4204
rect -428 -4208 -424 -4204
rect -331 -4210 -327 -4200
rect -192 -4208 -188 -4204
rect -154 -4208 -150 -4204
rect -94 -4208 -90 -4204
rect -70 -4208 -66 -4204
rect 457 -4208 461 -4198
rect 1202 -4208 1206 -4198
rect -1257 -4216 -1253 -4212
rect -1223 -4216 -1219 -4212
rect -1171 -4216 -1167 -4212
rect -1111 -4216 -1107 -4212
rect -1073 -4216 -1069 -4212
rect -928 -4216 -924 -4212
rect -894 -4216 -890 -4212
rect -842 -4216 -838 -4212
rect -782 -4216 -778 -4212
rect -744 -4216 -740 -4212
rect -570 -4216 -566 -4212
rect -536 -4216 -532 -4212
rect -484 -4216 -480 -4212
rect -424 -4216 -420 -4212
rect -386 -4216 -382 -4212
rect -212 -4216 -208 -4212
rect -178 -4216 -174 -4212
rect -126 -4216 -122 -4212
rect -66 -4216 -62 -4212
rect -28 -4216 -24 -4212
rect -1213 -4223 -1209 -4219
rect -1181 -4223 -1177 -4219
rect -1129 -4223 -1125 -4219
rect -1097 -4223 -1093 -4219
rect -884 -4223 -880 -4219
rect -852 -4223 -848 -4219
rect -800 -4223 -796 -4219
rect -768 -4223 -764 -4219
rect -526 -4223 -522 -4219
rect -494 -4223 -490 -4219
rect -442 -4223 -438 -4219
rect -410 -4223 -406 -4219
rect -168 -4223 -164 -4219
rect -136 -4223 -132 -4219
rect -84 -4223 -80 -4219
rect -52 -4223 -48 -4219
rect -1253 -4230 -1249 -4226
rect -1139 -4230 -1135 -4226
rect -1087 -4230 -1083 -4226
rect -924 -4230 -920 -4226
rect -810 -4230 -806 -4226
rect -758 -4230 -754 -4226
rect -566 -4230 -562 -4226
rect -452 -4230 -448 -4226
rect -400 -4230 -396 -4226
rect -208 -4230 -204 -4226
rect -94 -4230 -90 -4226
rect -42 -4230 -38 -4226
rect -1195 -4237 -1191 -4233
rect -1157 -4237 -1153 -4233
rect -866 -4237 -862 -4233
rect -828 -4237 -824 -4233
rect -508 -4237 -504 -4233
rect -470 -4237 -466 -4233
rect -150 -4237 -146 -4233
rect -112 -4237 -108 -4233
rect -1338 -4303 -1334 -4299
rect -934 -4303 -930 -4299
rect -576 -4303 -572 -4299
rect -218 -4303 -214 -4299
rect 210 -4303 214 -4299
rect 566 -4303 570 -4299
rect 964 -4303 968 -4299
rect 1322 -4303 1326 -4299
rect -1327 -4311 -1323 -4307
rect -923 -4311 -919 -4307
rect -565 -4311 -561 -4307
rect -207 -4311 -203 -4307
rect 221 -4311 225 -4307
rect 577 -4311 581 -4307
rect 975 -4311 979 -4307
rect 1333 -4311 1337 -4307
rect -1028 -4324 -1024 -4314
rect -672 -4324 -668 -4314
rect -331 -4325 -327 -4315
rect 457 -4324 461 -4314
rect 861 -4324 865 -4314
rect 1202 -4324 1206 -4314
rect -924 -4409 -920 -4405
rect -858 -4409 -854 -4405
rect -824 -4409 -820 -4405
rect -780 -4409 -776 -4405
rect -746 -4409 -742 -4405
rect -566 -4409 -562 -4405
rect -500 -4409 -496 -4405
rect -466 -4409 -462 -4405
rect -422 -4409 -418 -4405
rect -388 -4409 -384 -4405
rect -208 -4409 -204 -4405
rect -142 -4409 -138 -4405
rect -108 -4409 -104 -4405
rect -64 -4409 -60 -4405
rect -30 -4409 -26 -4405
rect 220 -4409 224 -4405
rect 286 -4409 290 -4405
rect 320 -4409 324 -4405
rect 364 -4409 368 -4405
rect 398 -4409 402 -4405
rect 576 -4409 580 -4405
rect 642 -4409 646 -4405
rect 676 -4409 680 -4405
rect 720 -4409 724 -4405
rect 754 -4409 758 -4405
rect 974 -4409 978 -4405
rect 1040 -4409 1044 -4405
rect 1074 -4409 1078 -4405
rect 1118 -4409 1122 -4405
rect 1152 -4409 1156 -4405
rect 1332 -4409 1336 -4405
rect 1398 -4409 1402 -4405
rect 1432 -4409 1436 -4405
rect 1476 -4409 1480 -4405
rect 1510 -4409 1514 -4405
rect -882 -4416 -878 -4412
rect -524 -4416 -520 -4412
rect -166 -4416 -162 -4412
rect 262 -4416 266 -4412
rect 618 -4416 622 -4412
rect 1016 -4416 1020 -4412
rect 1374 -4416 1378 -4412
rect -848 -4423 -844 -4419
rect -706 -4423 -702 -4419
rect -490 -4423 -486 -4419
rect -348 -4423 -344 -4419
rect -132 -4423 -128 -4419
rect 10 -4423 14 -4419
rect 296 -4423 300 -4419
rect 438 -4423 442 -4419
rect 652 -4423 656 -4419
rect 794 -4423 798 -4419
rect 1050 -4423 1054 -4419
rect 1192 -4423 1196 -4419
rect 1408 -4423 1412 -4419
rect 1550 -4423 1554 -4419
rect -928 -4430 -924 -4426
rect -898 -4430 -894 -4426
rect -780 -4430 -776 -4426
rect -570 -4430 -566 -4426
rect -540 -4430 -536 -4426
rect -422 -4430 -418 -4426
rect -212 -4430 -208 -4426
rect -182 -4430 -178 -4426
rect -64 -4430 -60 -4426
rect 216 -4430 220 -4426
rect 246 -4430 250 -4426
rect 364 -4430 368 -4426
rect 572 -4430 576 -4426
rect 602 -4430 606 -4426
rect 720 -4430 724 -4426
rect 970 -4430 974 -4426
rect 1000 -4430 1004 -4426
rect 1118 -4430 1122 -4426
rect 1328 -4430 1332 -4426
rect 1358 -4430 1362 -4426
rect 1476 -4430 1480 -4426
rect -1203 -4439 -1199 -4435
rect -902 -4438 -898 -4434
rect -804 -4438 -800 -4434
rect -544 -4438 -540 -4434
rect -446 -4438 -442 -4434
rect -186 -4438 -182 -4434
rect -88 -4438 -84 -4434
rect 242 -4438 246 -4434
rect 340 -4438 344 -4434
rect 598 -4438 602 -4434
rect 696 -4438 700 -4434
rect 996 -4438 1000 -4434
rect 1094 -4438 1098 -4434
rect 1354 -4438 1358 -4434
rect 1452 -4438 1456 -4434
rect -1253 -4446 -1249 -4442
rect -1213 -4446 -1209 -4442
rect -1193 -4446 -1189 -4442
rect -924 -4445 -920 -4441
rect -776 -4445 -772 -4441
rect -566 -4445 -562 -4441
rect -418 -4445 -414 -4441
rect -208 -4445 -204 -4441
rect -60 -4445 -56 -4441
rect 220 -4445 224 -4441
rect 368 -4445 372 -4441
rect 576 -4445 580 -4441
rect 724 -4445 728 -4441
rect 974 -4445 978 -4441
rect 1122 -4445 1126 -4441
rect 1332 -4445 1336 -4441
rect 1480 -4445 1484 -4441
rect -1257 -4453 -1253 -4449
rect -1227 -4453 -1223 -4449
rect -1179 -4453 -1175 -4449
rect -902 -4452 -898 -4448
rect -794 -4452 -790 -4448
rect -760 -4452 -756 -4448
rect -544 -4452 -540 -4448
rect -436 -4452 -432 -4448
rect -402 -4452 -398 -4448
rect -186 -4452 -182 -4448
rect -78 -4452 -74 -4448
rect -44 -4452 -40 -4448
rect 242 -4452 246 -4448
rect 350 -4452 354 -4448
rect 384 -4452 388 -4448
rect 598 -4452 602 -4448
rect 706 -4452 710 -4448
rect 740 -4452 744 -4448
rect 996 -4452 1000 -4448
rect 1104 -4452 1108 -4448
rect 1138 -4452 1142 -4448
rect 1354 -4452 1358 -4448
rect 1462 -4452 1466 -4448
rect 1496 -4452 1500 -4448
rect -928 -4459 -924 -4455
rect -872 -4459 -868 -4455
rect -838 -4459 -834 -4455
rect -570 -4459 -566 -4455
rect -514 -4459 -510 -4455
rect -480 -4459 -476 -4455
rect -212 -4459 -208 -4455
rect -156 -4459 -152 -4455
rect -122 -4459 -118 -4455
rect 216 -4459 220 -4455
rect 272 -4459 276 -4455
rect 306 -4459 310 -4455
rect 572 -4459 576 -4455
rect 628 -4459 632 -4455
rect 662 -4459 666 -4455
rect 970 -4459 974 -4455
rect 1026 -4459 1030 -4455
rect 1060 -4459 1064 -4455
rect 1328 -4459 1332 -4455
rect 1384 -4459 1388 -4455
rect 1418 -4459 1422 -4455
rect -1237 -4561 -1233 -4557
rect -1199 -4561 -1195 -4557
rect -1139 -4561 -1135 -4557
rect -1115 -4561 -1111 -4557
rect -908 -4561 -904 -4557
rect -870 -4561 -866 -4557
rect -810 -4561 -806 -4557
rect -786 -4561 -782 -4557
rect -550 -4561 -546 -4557
rect -512 -4561 -508 -4557
rect -452 -4561 -448 -4557
rect -428 -4561 -424 -4557
rect -1257 -4569 -1253 -4565
rect -1223 -4569 -1219 -4565
rect -1171 -4569 -1167 -4565
rect -1111 -4569 -1107 -4565
rect -1073 -4569 -1069 -4565
rect -928 -4569 -924 -4565
rect -894 -4569 -890 -4565
rect -842 -4569 -838 -4565
rect -782 -4569 -778 -4565
rect -744 -4569 -740 -4565
rect -570 -4569 -566 -4565
rect -536 -4569 -532 -4565
rect -484 -4569 -480 -4565
rect -424 -4569 -420 -4565
rect -386 -4569 -382 -4565
rect -1213 -4576 -1209 -4572
rect -1181 -4576 -1177 -4572
rect -1129 -4576 -1125 -4572
rect -1097 -4576 -1093 -4572
rect -884 -4576 -880 -4572
rect -852 -4576 -848 -4572
rect -800 -4576 -796 -4572
rect -768 -4576 -764 -4572
rect -526 -4576 -522 -4572
rect -494 -4576 -490 -4572
rect -442 -4576 -438 -4572
rect -410 -4576 -406 -4572
rect -1253 -4583 -1249 -4579
rect -1139 -4583 -1135 -4579
rect -1087 -4583 -1083 -4579
rect -924 -4583 -920 -4579
rect -810 -4583 -806 -4579
rect -758 -4583 -754 -4579
rect -566 -4583 -562 -4579
rect -452 -4583 -448 -4579
rect -400 -4583 -396 -4579
rect -1195 -4590 -1191 -4586
rect -1157 -4590 -1153 -4586
rect -866 -4590 -862 -4586
rect -828 -4590 -824 -4586
rect -508 -4590 -504 -4586
rect -470 -4590 -466 -4586
rect -1237 -4682 -1233 -4678
rect -1199 -4682 -1195 -4678
rect -1139 -4682 -1135 -4678
rect -1115 -4682 -1111 -4678
rect -908 -4682 -904 -4678
rect -870 -4682 -866 -4678
rect -810 -4682 -806 -4678
rect -786 -4682 -782 -4678
rect -550 -4682 -546 -4678
rect -512 -4682 -508 -4678
rect -452 -4682 -448 -4678
rect -428 -4682 -424 -4678
rect -192 -4682 -188 -4678
rect -154 -4682 -150 -4678
rect -94 -4682 -90 -4678
rect -70 -4682 -66 -4678
rect 236 -4682 240 -4678
rect 274 -4682 278 -4678
rect 334 -4682 338 -4678
rect 358 -4682 362 -4678
rect 592 -4682 596 -4678
rect 630 -4682 634 -4678
rect 690 -4682 694 -4678
rect 714 -4682 718 -4678
rect 990 -4682 994 -4678
rect 1028 -4682 1032 -4678
rect 1088 -4682 1092 -4678
rect 1112 -4682 1116 -4678
rect 1348 -4682 1352 -4678
rect 1386 -4682 1390 -4678
rect 1446 -4682 1450 -4678
rect 1470 -4682 1474 -4678
rect -1257 -4690 -1253 -4686
rect -1223 -4690 -1219 -4686
rect -1171 -4690 -1167 -4686
rect -1111 -4690 -1107 -4686
rect -1073 -4690 -1069 -4686
rect -928 -4690 -924 -4686
rect -894 -4690 -890 -4686
rect -842 -4690 -838 -4686
rect -782 -4690 -778 -4686
rect -744 -4690 -740 -4686
rect -570 -4690 -566 -4686
rect -536 -4690 -532 -4686
rect -484 -4690 -480 -4686
rect -424 -4690 -420 -4686
rect -386 -4690 -382 -4686
rect -212 -4690 -208 -4686
rect -178 -4690 -174 -4686
rect -126 -4690 -122 -4686
rect -66 -4690 -62 -4686
rect -28 -4690 -24 -4686
rect 216 -4690 220 -4686
rect 250 -4690 254 -4686
rect 302 -4690 306 -4686
rect 362 -4690 366 -4686
rect 400 -4690 404 -4686
rect 572 -4690 576 -4686
rect 606 -4690 610 -4686
rect 658 -4690 662 -4686
rect 718 -4690 722 -4686
rect 756 -4690 760 -4686
rect 970 -4690 974 -4686
rect 1004 -4690 1008 -4686
rect 1056 -4690 1060 -4686
rect 1116 -4690 1120 -4686
rect 1154 -4690 1158 -4686
rect 1328 -4690 1332 -4686
rect 1362 -4690 1366 -4686
rect 1414 -4690 1418 -4686
rect 1474 -4690 1478 -4686
rect 1512 -4690 1516 -4686
rect -1213 -4697 -1209 -4693
rect -1181 -4697 -1177 -4693
rect -1129 -4697 -1125 -4693
rect -1097 -4697 -1093 -4693
rect -884 -4697 -880 -4693
rect -852 -4697 -848 -4693
rect -800 -4697 -796 -4693
rect -768 -4697 -764 -4693
rect -526 -4697 -522 -4693
rect -494 -4697 -490 -4693
rect -442 -4697 -438 -4693
rect -410 -4697 -406 -4693
rect -168 -4697 -164 -4693
rect -136 -4697 -132 -4693
rect -84 -4697 -80 -4693
rect -52 -4697 -48 -4693
rect 260 -4697 264 -4693
rect 292 -4697 296 -4693
rect 344 -4697 348 -4693
rect 376 -4697 380 -4693
rect 616 -4697 620 -4693
rect 648 -4697 652 -4693
rect 700 -4697 704 -4693
rect 732 -4697 736 -4693
rect 1014 -4697 1018 -4693
rect 1046 -4697 1050 -4693
rect 1098 -4697 1102 -4693
rect 1130 -4697 1134 -4693
rect 1372 -4697 1376 -4693
rect 1404 -4697 1408 -4693
rect 1456 -4697 1460 -4693
rect 1488 -4697 1492 -4693
rect -1253 -4704 -1249 -4700
rect -1139 -4704 -1135 -4700
rect -1087 -4704 -1083 -4700
rect -924 -4704 -920 -4700
rect -810 -4704 -806 -4700
rect -758 -4704 -754 -4700
rect -566 -4704 -562 -4700
rect -452 -4704 -448 -4700
rect -400 -4704 -396 -4700
rect -208 -4704 -204 -4700
rect -94 -4704 -90 -4700
rect -42 -4704 -38 -4700
rect 220 -4704 224 -4700
rect 334 -4704 338 -4700
rect 386 -4704 390 -4700
rect 576 -4704 580 -4700
rect 690 -4704 694 -4700
rect 742 -4704 746 -4700
rect 974 -4704 978 -4700
rect 1088 -4704 1092 -4700
rect 1140 -4704 1144 -4700
rect 1332 -4704 1336 -4700
rect 1446 -4704 1450 -4700
rect 1498 -4704 1502 -4700
rect -1195 -4711 -1191 -4707
rect -1157 -4711 -1153 -4707
rect -866 -4711 -862 -4707
rect -828 -4711 -824 -4707
rect -508 -4711 -504 -4707
rect -470 -4711 -466 -4707
rect -150 -4711 -146 -4707
rect -112 -4711 -108 -4707
rect 278 -4711 282 -4707
rect 316 -4711 320 -4707
rect 634 -4711 638 -4707
rect 672 -4711 676 -4707
rect 1032 -4711 1036 -4707
rect 1070 -4711 1074 -4707
rect 1390 -4711 1394 -4707
rect 1428 -4711 1432 -4707
rect -1237 -4803 -1233 -4799
rect -1199 -4803 -1195 -4799
rect -1139 -4803 -1135 -4799
rect -1115 -4803 -1111 -4799
rect -908 -4803 -904 -4799
rect -870 -4803 -866 -4799
rect -810 -4803 -806 -4799
rect -786 -4803 -782 -4799
rect -550 -4803 -546 -4799
rect -512 -4803 -508 -4799
rect -452 -4803 -448 -4799
rect -428 -4803 -424 -4799
rect -192 -4803 -188 -4799
rect -154 -4803 -150 -4799
rect -94 -4803 -90 -4799
rect -70 -4803 -66 -4799
rect -1257 -4811 -1253 -4807
rect -1223 -4811 -1219 -4807
rect -1171 -4811 -1167 -4807
rect -1111 -4811 -1107 -4807
rect -1073 -4811 -1069 -4807
rect -928 -4811 -924 -4807
rect -894 -4811 -890 -4807
rect -842 -4811 -838 -4807
rect -782 -4811 -778 -4807
rect -744 -4811 -740 -4807
rect -570 -4811 -566 -4807
rect -536 -4811 -532 -4807
rect -484 -4811 -480 -4807
rect -424 -4811 -420 -4807
rect -386 -4811 -382 -4807
rect -212 -4811 -208 -4807
rect -178 -4811 -174 -4807
rect -126 -4811 -122 -4807
rect -66 -4811 -62 -4807
rect -28 -4811 -24 -4807
rect 91 -4812 95 -4796
rect 236 -4803 240 -4799
rect 274 -4803 278 -4799
rect 334 -4803 338 -4799
rect 358 -4803 362 -4799
rect 592 -4803 596 -4799
rect 630 -4803 634 -4799
rect 690 -4803 694 -4799
rect 714 -4803 718 -4799
rect 990 -4803 994 -4799
rect 1028 -4803 1032 -4799
rect 1088 -4803 1092 -4799
rect 1112 -4803 1116 -4799
rect 1348 -4803 1352 -4799
rect 1386 -4803 1390 -4799
rect 1446 -4803 1450 -4799
rect 1470 -4803 1474 -4799
rect 216 -4811 220 -4807
rect 250 -4811 254 -4807
rect 302 -4811 306 -4807
rect 362 -4811 366 -4807
rect 400 -4811 404 -4807
rect 572 -4811 576 -4807
rect 606 -4811 610 -4807
rect 658 -4811 662 -4807
rect 718 -4811 722 -4807
rect 756 -4811 760 -4807
rect 970 -4811 974 -4807
rect 1004 -4811 1008 -4807
rect 1056 -4811 1060 -4807
rect 1116 -4811 1120 -4807
rect 1154 -4811 1158 -4807
rect 1328 -4811 1332 -4807
rect 1362 -4811 1366 -4807
rect 1414 -4811 1418 -4807
rect 1474 -4811 1478 -4807
rect 1512 -4811 1516 -4807
rect -1213 -4818 -1209 -4814
rect -1181 -4818 -1177 -4814
rect -1129 -4818 -1125 -4814
rect -1097 -4818 -1093 -4814
rect -884 -4818 -880 -4814
rect -852 -4818 -848 -4814
rect -800 -4818 -796 -4814
rect -768 -4818 -764 -4814
rect -526 -4818 -522 -4814
rect -494 -4818 -490 -4814
rect -442 -4818 -438 -4814
rect -410 -4818 -406 -4814
rect -168 -4818 -164 -4814
rect -136 -4818 -132 -4814
rect -84 -4818 -80 -4814
rect -52 -4818 -48 -4814
rect 260 -4818 264 -4814
rect 292 -4818 296 -4814
rect 344 -4818 348 -4814
rect 376 -4818 380 -4814
rect 616 -4818 620 -4814
rect 648 -4818 652 -4814
rect 700 -4818 704 -4814
rect 732 -4818 736 -4814
rect 1014 -4818 1018 -4814
rect 1046 -4818 1050 -4814
rect 1098 -4818 1102 -4814
rect 1130 -4818 1134 -4814
rect 1372 -4818 1376 -4814
rect 1404 -4818 1408 -4814
rect 1456 -4818 1460 -4814
rect 1488 -4818 1492 -4814
rect -1253 -4825 -1249 -4821
rect -1139 -4825 -1135 -4821
rect -1087 -4825 -1083 -4821
rect -924 -4825 -920 -4821
rect -810 -4825 -806 -4821
rect -758 -4825 -754 -4821
rect -566 -4825 -562 -4821
rect -452 -4825 -448 -4821
rect -400 -4825 -396 -4821
rect -208 -4825 -204 -4821
rect -94 -4825 -90 -4821
rect -42 -4825 -38 -4821
rect 220 -4825 224 -4821
rect 334 -4825 338 -4821
rect 386 -4825 390 -4821
rect 576 -4825 580 -4821
rect 690 -4825 694 -4821
rect 742 -4825 746 -4821
rect 974 -4825 978 -4821
rect 1088 -4825 1092 -4821
rect 1140 -4825 1144 -4821
rect 1332 -4825 1336 -4821
rect 1446 -4825 1450 -4821
rect 1498 -4825 1502 -4821
rect -1195 -4832 -1191 -4828
rect -1157 -4832 -1153 -4828
rect -866 -4832 -862 -4828
rect -828 -4832 -824 -4828
rect -508 -4832 -504 -4828
rect -470 -4832 -466 -4828
rect -150 -4832 -146 -4828
rect -112 -4832 -108 -4828
rect 278 -4832 282 -4828
rect 316 -4832 320 -4828
rect 634 -4832 638 -4828
rect 672 -4832 676 -4828
rect 1032 -4832 1036 -4828
rect 1070 -4832 1074 -4828
rect 1390 -4832 1394 -4828
rect 1428 -4832 1432 -4828
rect -1237 -4921 -1233 -4917
rect -1199 -4921 -1195 -4917
rect -1139 -4921 -1135 -4917
rect -1115 -4921 -1111 -4917
rect -908 -4921 -904 -4917
rect -870 -4921 -866 -4917
rect -810 -4921 -806 -4917
rect -786 -4921 -782 -4917
rect -550 -4921 -546 -4917
rect -512 -4921 -508 -4917
rect -452 -4921 -448 -4917
rect -428 -4921 -424 -4917
rect -192 -4921 -188 -4917
rect -154 -4921 -150 -4917
rect -94 -4921 -90 -4917
rect -70 -4921 -66 -4917
rect 236 -4921 240 -4917
rect 274 -4921 278 -4917
rect 334 -4921 338 -4917
rect 358 -4921 362 -4917
rect -1257 -4929 -1253 -4925
rect -1223 -4929 -1219 -4925
rect -1171 -4929 -1167 -4925
rect -1111 -4929 -1107 -4925
rect -1073 -4929 -1069 -4925
rect -928 -4929 -924 -4925
rect -894 -4929 -890 -4925
rect -842 -4929 -838 -4925
rect -782 -4929 -778 -4925
rect -744 -4929 -740 -4925
rect -570 -4929 -566 -4925
rect -536 -4929 -532 -4925
rect -484 -4929 -480 -4925
rect -424 -4929 -420 -4925
rect -386 -4929 -382 -4925
rect -212 -4929 -208 -4925
rect -178 -4929 -174 -4925
rect -126 -4929 -122 -4925
rect -66 -4929 -62 -4925
rect -28 -4929 -24 -4925
rect 216 -4929 220 -4925
rect 250 -4929 254 -4925
rect 302 -4929 306 -4925
rect 362 -4929 366 -4925
rect 400 -4929 404 -4925
rect -1213 -4936 -1209 -4932
rect -1181 -4936 -1177 -4932
rect -1129 -4936 -1125 -4932
rect -1097 -4936 -1093 -4932
rect -884 -4936 -880 -4932
rect -852 -4936 -848 -4932
rect -800 -4936 -796 -4932
rect -768 -4936 -764 -4932
rect -526 -4936 -522 -4932
rect -494 -4936 -490 -4932
rect -442 -4936 -438 -4932
rect -410 -4936 -406 -4932
rect -168 -4936 -164 -4932
rect -136 -4936 -132 -4932
rect -84 -4936 -80 -4932
rect -52 -4936 -48 -4932
rect 260 -4936 264 -4932
rect 292 -4936 296 -4932
rect 344 -4936 348 -4932
rect 376 -4936 380 -4932
rect -1253 -4943 -1249 -4939
rect -1139 -4943 -1135 -4939
rect -1087 -4943 -1083 -4939
rect -924 -4943 -920 -4939
rect -810 -4943 -806 -4939
rect -758 -4943 -754 -4939
rect -566 -4943 -562 -4939
rect -452 -4943 -448 -4939
rect -400 -4943 -396 -4939
rect -208 -4943 -204 -4939
rect -94 -4943 -90 -4939
rect -42 -4943 -38 -4939
rect 220 -4943 224 -4939
rect 334 -4943 338 -4939
rect 386 -4943 390 -4939
rect -1195 -4950 -1191 -4946
rect -1157 -4950 -1153 -4946
rect -866 -4950 -862 -4946
rect -828 -4950 -824 -4946
rect -508 -4950 -504 -4946
rect -470 -4950 -466 -4946
rect -150 -4950 -146 -4946
rect -112 -4950 -108 -4946
rect 278 -4950 282 -4946
rect 316 -4950 320 -4946
rect -1338 -5022 -1334 -5018
rect -934 -5022 -930 -5018
rect -576 -5022 -572 -5018
rect -218 -5022 -214 -5018
rect 210 -5022 214 -5018
rect 964 -5022 968 -5018
rect 1322 -5022 1326 -5018
rect -1327 -5030 -1323 -5026
rect -923 -5030 -919 -5026
rect -565 -5030 -561 -5026
rect -207 -5030 -203 -5026
rect 221 -5030 225 -5026
rect 577 -5030 581 -5026
rect 975 -5030 979 -5026
rect 1333 -5030 1337 -5026
rect -924 -5128 -920 -5124
rect -858 -5128 -854 -5124
rect -824 -5128 -820 -5124
rect -780 -5128 -776 -5124
rect -746 -5128 -742 -5124
rect -566 -5128 -562 -5124
rect -500 -5128 -496 -5124
rect -466 -5128 -462 -5124
rect -422 -5128 -418 -5124
rect -388 -5128 -384 -5124
rect -208 -5128 -204 -5124
rect -142 -5128 -138 -5124
rect -108 -5128 -104 -5124
rect -64 -5128 -60 -5124
rect -30 -5128 -26 -5124
rect 220 -5128 224 -5124
rect 286 -5128 290 -5124
rect 320 -5128 324 -5124
rect 364 -5128 368 -5124
rect 398 -5128 402 -5124
rect 576 -5128 580 -5124
rect 642 -5128 646 -5124
rect 676 -5128 680 -5124
rect 720 -5128 724 -5124
rect 754 -5128 758 -5124
rect 974 -5128 978 -5124
rect 1040 -5128 1044 -5124
rect 1074 -5128 1078 -5124
rect 1118 -5128 1122 -5124
rect 1152 -5128 1156 -5124
rect 1332 -5128 1336 -5124
rect 1398 -5128 1402 -5124
rect 1432 -5128 1436 -5124
rect 1476 -5128 1480 -5124
rect 1510 -5128 1514 -5124
rect -882 -5135 -878 -5131
rect -524 -5135 -520 -5131
rect -166 -5135 -162 -5131
rect 262 -5135 266 -5131
rect 618 -5135 622 -5131
rect 1016 -5135 1020 -5131
rect 1374 -5135 1378 -5131
rect -848 -5142 -844 -5138
rect -706 -5142 -702 -5138
rect -490 -5142 -486 -5138
rect -348 -5142 -344 -5138
rect -132 -5142 -128 -5138
rect 10 -5142 14 -5138
rect 296 -5142 300 -5138
rect 438 -5142 442 -5138
rect 652 -5142 656 -5138
rect 794 -5142 798 -5138
rect 1050 -5142 1054 -5138
rect 1192 -5142 1196 -5138
rect 1408 -5142 1412 -5138
rect 1550 -5142 1554 -5138
rect -928 -5149 -924 -5145
rect -898 -5149 -894 -5145
rect -780 -5149 -776 -5145
rect -570 -5149 -566 -5145
rect -540 -5149 -536 -5145
rect -422 -5149 -418 -5145
rect -212 -5149 -208 -5145
rect -182 -5149 -178 -5145
rect -64 -5149 -60 -5145
rect 216 -5149 220 -5145
rect 246 -5149 250 -5145
rect 364 -5149 368 -5145
rect 572 -5149 576 -5145
rect 602 -5149 606 -5145
rect 720 -5149 724 -5145
rect 970 -5149 974 -5145
rect 1000 -5149 1004 -5145
rect 1118 -5149 1122 -5145
rect 1328 -5149 1332 -5145
rect 1358 -5149 1362 -5145
rect 1476 -5149 1480 -5145
rect -1203 -5158 -1199 -5154
rect -902 -5157 -898 -5153
rect -804 -5157 -800 -5153
rect -544 -5157 -540 -5153
rect -446 -5157 -442 -5153
rect -186 -5157 -182 -5153
rect -88 -5157 -84 -5153
rect 242 -5157 246 -5153
rect 340 -5157 344 -5153
rect 598 -5157 602 -5153
rect 696 -5157 700 -5153
rect 996 -5157 1000 -5153
rect 1094 -5157 1098 -5153
rect 1354 -5157 1358 -5153
rect 1452 -5157 1456 -5153
rect -1253 -5165 -1249 -5161
rect -1213 -5165 -1209 -5161
rect -1193 -5165 -1189 -5161
rect -924 -5164 -920 -5160
rect -776 -5164 -772 -5160
rect -566 -5164 -562 -5160
rect -418 -5164 -414 -5160
rect -208 -5164 -204 -5160
rect -60 -5164 -56 -5160
rect 220 -5164 224 -5160
rect 368 -5164 372 -5160
rect 576 -5164 580 -5160
rect 724 -5164 728 -5160
rect 974 -5164 978 -5160
rect 1122 -5164 1126 -5160
rect 1332 -5164 1336 -5160
rect 1480 -5164 1484 -5160
rect -1257 -5172 -1253 -5168
rect -1227 -5172 -1223 -5168
rect -1179 -5172 -1175 -5168
rect -902 -5171 -898 -5167
rect -794 -5171 -790 -5167
rect -760 -5171 -756 -5167
rect -544 -5171 -540 -5167
rect -436 -5171 -432 -5167
rect -402 -5171 -398 -5167
rect -186 -5171 -182 -5167
rect -78 -5171 -74 -5167
rect -44 -5171 -40 -5167
rect 242 -5171 246 -5167
rect 350 -5171 354 -5167
rect 384 -5171 388 -5167
rect 598 -5171 602 -5167
rect 706 -5171 710 -5167
rect 740 -5171 744 -5167
rect 996 -5171 1000 -5167
rect 1104 -5171 1108 -5167
rect 1138 -5171 1142 -5167
rect 1354 -5171 1358 -5167
rect 1462 -5171 1466 -5167
rect 1496 -5171 1500 -5167
rect -928 -5178 -924 -5174
rect -872 -5178 -868 -5174
rect -838 -5178 -834 -5174
rect -570 -5178 -566 -5174
rect -514 -5178 -510 -5174
rect -480 -5178 -476 -5174
rect -212 -5178 -208 -5174
rect -156 -5178 -152 -5174
rect -122 -5178 -118 -5174
rect 216 -5178 220 -5174
rect 272 -5178 276 -5174
rect 306 -5178 310 -5174
rect 572 -5178 576 -5174
rect 628 -5178 632 -5174
rect 662 -5178 666 -5174
rect 970 -5178 974 -5174
rect 1026 -5178 1030 -5174
rect 1060 -5178 1064 -5174
rect 1328 -5178 1332 -5174
rect 1384 -5178 1388 -5174
rect 1418 -5178 1422 -5174
rect -1237 -5276 -1233 -5272
rect -1199 -5276 -1195 -5272
rect -1139 -5276 -1135 -5272
rect -1115 -5276 -1111 -5272
rect -908 -5276 -904 -5272
rect -870 -5276 -866 -5272
rect -810 -5276 -806 -5272
rect -786 -5276 -782 -5272
rect -1257 -5284 -1253 -5280
rect -1223 -5284 -1219 -5280
rect -1171 -5284 -1167 -5280
rect -1111 -5284 -1107 -5280
rect -1073 -5284 -1069 -5280
rect -928 -5284 -924 -5280
rect -894 -5284 -890 -5280
rect -842 -5284 -838 -5280
rect -782 -5284 -778 -5280
rect -744 -5284 -740 -5280
rect -1213 -5291 -1209 -5287
rect -1181 -5291 -1177 -5287
rect -1129 -5291 -1125 -5287
rect -1097 -5291 -1093 -5287
rect -884 -5291 -880 -5287
rect -852 -5291 -848 -5287
rect -800 -5291 -796 -5287
rect -768 -5291 -764 -5287
rect -1253 -5298 -1249 -5294
rect -1139 -5298 -1135 -5294
rect -1087 -5298 -1083 -5294
rect -924 -5298 -920 -5294
rect -810 -5298 -806 -5294
rect -758 -5298 -754 -5294
rect -1195 -5305 -1191 -5301
rect -1157 -5305 -1153 -5301
rect -866 -5305 -862 -5301
rect -828 -5305 -824 -5301
rect -1237 -5397 -1233 -5393
rect -1199 -5397 -1195 -5393
rect -1139 -5397 -1135 -5393
rect -1115 -5397 -1111 -5393
rect -1025 -5397 -1021 -5387
rect -908 -5397 -904 -5393
rect -870 -5397 -866 -5393
rect -810 -5397 -806 -5393
rect -786 -5397 -782 -5393
rect -1257 -5405 -1253 -5401
rect -1223 -5405 -1219 -5401
rect -1171 -5405 -1167 -5401
rect -1111 -5405 -1107 -5401
rect -1073 -5405 -1069 -5401
rect -928 -5405 -924 -5401
rect -894 -5405 -890 -5401
rect -842 -5405 -838 -5401
rect -782 -5405 -778 -5401
rect -744 -5405 -740 -5401
rect -672 -5402 -668 -5392
rect -550 -5397 -546 -5393
rect -512 -5397 -508 -5393
rect -452 -5397 -448 -5393
rect -428 -5397 -424 -5393
rect -570 -5405 -566 -5401
rect -536 -5405 -532 -5401
rect -484 -5405 -480 -5401
rect -424 -5405 -420 -5401
rect -386 -5405 -382 -5401
rect -326 -5403 -322 -5393
rect -192 -5397 -188 -5393
rect -154 -5397 -150 -5393
rect -94 -5397 -90 -5393
rect -70 -5397 -66 -5393
rect 236 -5397 240 -5393
rect 274 -5397 278 -5393
rect 334 -5397 338 -5393
rect 358 -5397 362 -5393
rect 467 -5397 471 -5387
rect 592 -5397 596 -5393
rect 630 -5397 634 -5393
rect 690 -5397 694 -5393
rect 714 -5397 718 -5393
rect -212 -5405 -208 -5401
rect -178 -5405 -174 -5401
rect -126 -5405 -122 -5401
rect -66 -5405 -62 -5401
rect -28 -5405 -24 -5401
rect 216 -5405 220 -5401
rect 250 -5405 254 -5401
rect 302 -5405 306 -5401
rect 362 -5405 366 -5401
rect 400 -5405 404 -5401
rect 572 -5405 576 -5401
rect 606 -5405 610 -5401
rect 658 -5405 662 -5401
rect 718 -5405 722 -5401
rect 756 -5405 760 -5401
rect 868 -5402 872 -5392
rect 990 -5397 994 -5393
rect 1028 -5397 1032 -5393
rect 1088 -5397 1092 -5393
rect 1112 -5397 1116 -5393
rect 970 -5405 974 -5401
rect 1004 -5405 1008 -5401
rect 1056 -5405 1060 -5401
rect 1116 -5405 1120 -5401
rect 1154 -5405 1158 -5401
rect 1211 -5406 1215 -5396
rect 1348 -5397 1352 -5393
rect 1386 -5397 1390 -5393
rect 1446 -5397 1450 -5393
rect 1470 -5397 1474 -5393
rect 1328 -5405 1332 -5401
rect 1362 -5405 1366 -5401
rect 1414 -5405 1418 -5401
rect 1474 -5405 1478 -5401
rect 1512 -5405 1516 -5401
rect -1213 -5412 -1209 -5408
rect -1181 -5412 -1177 -5408
rect -1129 -5412 -1125 -5408
rect -1097 -5412 -1093 -5408
rect -884 -5412 -880 -5408
rect -852 -5412 -848 -5408
rect -800 -5412 -796 -5408
rect -768 -5412 -764 -5408
rect -526 -5412 -522 -5408
rect -494 -5412 -490 -5408
rect -442 -5412 -438 -5408
rect -410 -5412 -406 -5408
rect -168 -5412 -164 -5408
rect -136 -5412 -132 -5408
rect -84 -5412 -80 -5408
rect -52 -5412 -48 -5408
rect 260 -5412 264 -5408
rect 292 -5412 296 -5408
rect 344 -5412 348 -5408
rect 376 -5412 380 -5408
rect 616 -5412 620 -5408
rect 648 -5412 652 -5408
rect 700 -5412 704 -5408
rect 732 -5412 736 -5408
rect 1014 -5412 1018 -5408
rect 1046 -5412 1050 -5408
rect 1098 -5412 1102 -5408
rect 1130 -5412 1134 -5408
rect 1372 -5412 1376 -5408
rect 1404 -5412 1408 -5408
rect 1456 -5412 1460 -5408
rect 1488 -5412 1492 -5408
rect -1253 -5419 -1249 -5415
rect -1139 -5419 -1135 -5415
rect -1087 -5419 -1083 -5415
rect -924 -5419 -920 -5415
rect -810 -5419 -806 -5415
rect -758 -5419 -754 -5415
rect -566 -5419 -562 -5415
rect -452 -5419 -448 -5415
rect -400 -5419 -396 -5415
rect -208 -5419 -204 -5415
rect -94 -5419 -90 -5415
rect -42 -5419 -38 -5415
rect 220 -5419 224 -5415
rect 334 -5419 338 -5415
rect 386 -5419 390 -5415
rect 576 -5419 580 -5415
rect 690 -5419 694 -5415
rect 742 -5419 746 -5415
rect 974 -5419 978 -5415
rect 1088 -5419 1092 -5415
rect 1140 -5419 1144 -5415
rect 1332 -5419 1336 -5415
rect 1446 -5419 1450 -5415
rect 1498 -5419 1502 -5415
rect -1195 -5426 -1191 -5422
rect -1157 -5426 -1153 -5422
rect -866 -5426 -862 -5422
rect -828 -5426 -824 -5422
rect -508 -5426 -504 -5422
rect -470 -5426 -466 -5422
rect -150 -5426 -146 -5422
rect -112 -5426 -108 -5422
rect 278 -5426 282 -5422
rect 316 -5426 320 -5422
rect 634 -5426 638 -5422
rect 672 -5426 676 -5422
rect 1032 -5426 1036 -5422
rect 1070 -5426 1074 -5422
rect 1390 -5426 1394 -5422
rect 1428 -5426 1432 -5422
rect -1237 -5517 -1233 -5513
rect -1199 -5517 -1195 -5513
rect -1139 -5517 -1135 -5513
rect -1115 -5517 -1111 -5513
rect -1257 -5525 -1253 -5521
rect -1223 -5525 -1219 -5521
rect -1171 -5525 -1167 -5521
rect -1111 -5525 -1107 -5521
rect -1073 -5525 -1069 -5521
rect -1025 -5522 -1021 -5512
rect -908 -5517 -904 -5513
rect -870 -5517 -866 -5513
rect -810 -5517 -806 -5513
rect -786 -5517 -782 -5513
rect -550 -5517 -546 -5513
rect -512 -5517 -508 -5513
rect -452 -5517 -448 -5513
rect -428 -5517 -424 -5513
rect -326 -5518 -322 -5508
rect -192 -5517 -188 -5513
rect -154 -5517 -150 -5513
rect -94 -5517 -90 -5513
rect -70 -5517 -66 -5513
rect 236 -5517 240 -5513
rect 274 -5517 278 -5513
rect 334 -5517 338 -5513
rect 358 -5517 362 -5513
rect -928 -5525 -924 -5521
rect -894 -5525 -890 -5521
rect -842 -5525 -838 -5521
rect -782 -5525 -778 -5521
rect -744 -5525 -740 -5521
rect -570 -5525 -566 -5521
rect -536 -5525 -532 -5521
rect -484 -5525 -480 -5521
rect -424 -5525 -420 -5521
rect -386 -5525 -382 -5521
rect -212 -5525 -208 -5521
rect -178 -5525 -174 -5521
rect -126 -5525 -122 -5521
rect -66 -5525 -62 -5521
rect -28 -5525 -24 -5521
rect 216 -5525 220 -5521
rect 250 -5525 254 -5521
rect 302 -5525 306 -5521
rect 362 -5525 366 -5521
rect 400 -5525 404 -5521
rect 467 -5522 471 -5512
rect 592 -5517 596 -5513
rect 630 -5517 634 -5513
rect 690 -5517 694 -5513
rect 714 -5517 718 -5513
rect 990 -5517 994 -5513
rect 1028 -5517 1032 -5513
rect 1088 -5517 1092 -5513
rect 1112 -5517 1116 -5513
rect 572 -5525 576 -5521
rect 606 -5525 610 -5521
rect 658 -5525 662 -5521
rect 718 -5525 722 -5521
rect 756 -5525 760 -5521
rect 970 -5525 974 -5521
rect 1004 -5525 1008 -5521
rect 1056 -5525 1060 -5521
rect 1116 -5525 1120 -5521
rect 1154 -5525 1158 -5521
rect 1211 -5522 1215 -5512
rect 1348 -5517 1352 -5513
rect 1386 -5517 1390 -5513
rect 1446 -5517 1450 -5513
rect 1470 -5517 1474 -5513
rect 1328 -5525 1332 -5521
rect 1362 -5525 1366 -5521
rect 1414 -5525 1418 -5521
rect 1474 -5525 1478 -5521
rect 1512 -5525 1516 -5521
rect -1213 -5532 -1209 -5528
rect -1181 -5532 -1177 -5528
rect -1129 -5532 -1125 -5528
rect -1097 -5532 -1093 -5528
rect -884 -5532 -880 -5528
rect -852 -5532 -848 -5528
rect -800 -5532 -796 -5528
rect -768 -5532 -764 -5528
rect -526 -5532 -522 -5528
rect -494 -5532 -490 -5528
rect -442 -5532 -438 -5528
rect -410 -5532 -406 -5528
rect -168 -5532 -164 -5528
rect -136 -5532 -132 -5528
rect -84 -5532 -80 -5528
rect -52 -5532 -48 -5528
rect 260 -5532 264 -5528
rect 292 -5532 296 -5528
rect 344 -5532 348 -5528
rect 376 -5532 380 -5528
rect 616 -5532 620 -5528
rect 648 -5532 652 -5528
rect 700 -5532 704 -5528
rect 732 -5532 736 -5528
rect 1014 -5532 1018 -5528
rect 1046 -5532 1050 -5528
rect 1098 -5532 1102 -5528
rect 1130 -5532 1134 -5528
rect 1372 -5532 1376 -5528
rect 1404 -5532 1408 -5528
rect 1456 -5532 1460 -5528
rect 1488 -5532 1492 -5528
rect -1253 -5539 -1249 -5535
rect -1139 -5539 -1135 -5535
rect -1087 -5539 -1083 -5535
rect -924 -5539 -920 -5535
rect -810 -5539 -806 -5535
rect -758 -5539 -754 -5535
rect -566 -5539 -562 -5535
rect -452 -5539 -448 -5535
rect -400 -5539 -396 -5535
rect -208 -5539 -204 -5535
rect -94 -5539 -90 -5535
rect -42 -5539 -38 -5535
rect 220 -5539 224 -5535
rect 334 -5539 338 -5535
rect 386 -5539 390 -5535
rect 576 -5539 580 -5535
rect 690 -5539 694 -5535
rect 742 -5539 746 -5535
rect 974 -5539 978 -5535
rect 1088 -5539 1092 -5535
rect 1140 -5539 1144 -5535
rect 1332 -5539 1336 -5535
rect 1446 -5539 1450 -5535
rect 1498 -5539 1502 -5535
rect -1195 -5546 -1191 -5542
rect -1157 -5546 -1153 -5542
rect -866 -5546 -862 -5542
rect -828 -5546 -824 -5542
rect -508 -5546 -504 -5542
rect -470 -5546 -466 -5542
rect -150 -5546 -146 -5542
rect -112 -5546 -108 -5542
rect 278 -5546 282 -5542
rect 316 -5546 320 -5542
rect 634 -5546 638 -5542
rect 672 -5546 676 -5542
rect 1032 -5546 1036 -5542
rect 1070 -5546 1074 -5542
rect 1390 -5546 1394 -5542
rect 1428 -5546 1432 -5542
rect -1237 -5634 -1233 -5630
rect -1199 -5634 -1195 -5630
rect -1139 -5634 -1135 -5630
rect -1115 -5634 -1111 -5630
rect -908 -5634 -904 -5630
rect -870 -5634 -866 -5630
rect -810 -5634 -806 -5630
rect -786 -5634 -782 -5630
rect -550 -5634 -546 -5630
rect -512 -5634 -508 -5630
rect -452 -5634 -448 -5630
rect -428 -5634 -424 -5630
rect -192 -5634 -188 -5630
rect -154 -5634 -150 -5630
rect -94 -5634 -90 -5630
rect -70 -5634 -66 -5630
rect 236 -5634 240 -5630
rect 274 -5634 278 -5630
rect 334 -5634 338 -5630
rect 358 -5634 362 -5630
rect 592 -5634 596 -5630
rect 630 -5634 634 -5630
rect 690 -5634 694 -5630
rect 714 -5634 718 -5630
rect -1257 -5642 -1253 -5638
rect -1223 -5642 -1219 -5638
rect -1171 -5642 -1167 -5638
rect -1111 -5642 -1107 -5638
rect -1073 -5642 -1069 -5638
rect -928 -5642 -924 -5638
rect -894 -5642 -890 -5638
rect -842 -5642 -838 -5638
rect -782 -5642 -778 -5638
rect -744 -5642 -740 -5638
rect -570 -5642 -566 -5638
rect -536 -5642 -532 -5638
rect -484 -5642 -480 -5638
rect -424 -5642 -420 -5638
rect -386 -5642 -382 -5638
rect -212 -5642 -208 -5638
rect -178 -5642 -174 -5638
rect -126 -5642 -122 -5638
rect -66 -5642 -62 -5638
rect -28 -5642 -24 -5638
rect 216 -5642 220 -5638
rect 250 -5642 254 -5638
rect 302 -5642 306 -5638
rect 362 -5642 366 -5638
rect 400 -5642 404 -5638
rect 572 -5642 576 -5638
rect 606 -5642 610 -5638
rect 658 -5642 662 -5638
rect 718 -5642 722 -5638
rect 756 -5642 760 -5638
rect -1213 -5649 -1209 -5645
rect -1181 -5649 -1177 -5645
rect -1129 -5649 -1125 -5645
rect -1097 -5649 -1093 -5645
rect -884 -5649 -880 -5645
rect -852 -5649 -848 -5645
rect -800 -5649 -796 -5645
rect -768 -5649 -764 -5645
rect -526 -5649 -522 -5645
rect -494 -5649 -490 -5645
rect -442 -5649 -438 -5645
rect -410 -5649 -406 -5645
rect -168 -5649 -164 -5645
rect -136 -5649 -132 -5645
rect -84 -5649 -80 -5645
rect -52 -5649 -48 -5645
rect 260 -5649 264 -5645
rect 292 -5649 296 -5645
rect 344 -5649 348 -5645
rect 376 -5649 380 -5645
rect 616 -5649 620 -5645
rect 648 -5649 652 -5645
rect 700 -5649 704 -5645
rect 732 -5649 736 -5645
rect -1253 -5656 -1249 -5652
rect -1139 -5656 -1135 -5652
rect -1087 -5656 -1083 -5652
rect -924 -5656 -920 -5652
rect -810 -5656 -806 -5652
rect -758 -5656 -754 -5652
rect -566 -5656 -562 -5652
rect -452 -5656 -448 -5652
rect -400 -5656 -396 -5652
rect -208 -5656 -204 -5652
rect -94 -5656 -90 -5652
rect -42 -5656 -38 -5652
rect 220 -5656 224 -5652
rect 334 -5656 338 -5652
rect 386 -5656 390 -5652
rect 576 -5656 580 -5652
rect 690 -5656 694 -5652
rect 742 -5656 746 -5652
rect -1195 -5663 -1191 -5659
rect -1157 -5663 -1153 -5659
rect -866 -5663 -862 -5659
rect -828 -5663 -824 -5659
rect -508 -5663 -504 -5659
rect -470 -5663 -466 -5659
rect -150 -5663 -146 -5659
rect -112 -5663 -108 -5659
rect 278 -5663 282 -5659
rect 316 -5663 320 -5659
rect 634 -5663 638 -5659
rect 672 -5663 676 -5659
rect -1338 -5735 -1334 -5731
rect -934 -5735 -930 -5731
rect -576 -5735 -572 -5731
rect -218 -5735 -214 -5731
rect 210 -5735 214 -5731
rect 566 -5735 570 -5731
rect 964 -5735 968 -5731
rect 1322 -5735 1326 -5731
rect -1327 -5743 -1323 -5739
rect -923 -5743 -919 -5739
rect -565 -5743 -561 -5739
rect -207 -5743 -203 -5739
rect 221 -5743 225 -5739
rect 577 -5743 581 -5739
rect 975 -5743 979 -5739
rect 1333 -5743 1337 -5739
rect -924 -5841 -920 -5837
rect -858 -5841 -854 -5837
rect -824 -5841 -820 -5837
rect -780 -5841 -776 -5837
rect -746 -5841 -742 -5837
rect -566 -5841 -562 -5837
rect -500 -5841 -496 -5837
rect -466 -5841 -462 -5837
rect -422 -5841 -418 -5837
rect -388 -5841 -384 -5837
rect -208 -5841 -204 -5837
rect -142 -5841 -138 -5837
rect -108 -5841 -104 -5837
rect -64 -5841 -60 -5837
rect -30 -5841 -26 -5837
rect 220 -5841 224 -5837
rect 286 -5841 290 -5837
rect 320 -5841 324 -5837
rect 364 -5841 368 -5837
rect 398 -5841 402 -5837
rect 576 -5841 580 -5837
rect 642 -5841 646 -5837
rect 676 -5841 680 -5837
rect 720 -5841 724 -5837
rect 754 -5841 758 -5837
rect 974 -5841 978 -5837
rect 1040 -5841 1044 -5837
rect 1074 -5841 1078 -5837
rect 1118 -5841 1122 -5837
rect 1152 -5841 1156 -5837
rect 1332 -5841 1336 -5837
rect 1398 -5841 1402 -5837
rect 1432 -5841 1436 -5837
rect 1476 -5841 1480 -5837
rect 1510 -5841 1514 -5837
rect -882 -5848 -878 -5844
rect -524 -5848 -520 -5844
rect -166 -5848 -162 -5844
rect 262 -5848 266 -5844
rect 618 -5848 622 -5844
rect 1016 -5848 1020 -5844
rect 1374 -5848 1378 -5844
rect -848 -5855 -844 -5851
rect -706 -5855 -702 -5851
rect -490 -5855 -486 -5851
rect -348 -5855 -344 -5851
rect -132 -5855 -128 -5851
rect 10 -5855 14 -5851
rect 296 -5855 300 -5851
rect 438 -5855 442 -5851
rect 652 -5855 656 -5851
rect 794 -5855 798 -5851
rect 1050 -5855 1054 -5851
rect 1192 -5855 1196 -5851
rect 1408 -5855 1412 -5851
rect 1550 -5855 1554 -5851
rect -928 -5862 -924 -5858
rect -898 -5862 -894 -5858
rect -780 -5862 -776 -5858
rect -570 -5862 -566 -5858
rect -540 -5862 -536 -5858
rect -422 -5862 -418 -5858
rect -212 -5862 -208 -5858
rect -182 -5862 -178 -5858
rect -64 -5862 -60 -5858
rect 216 -5862 220 -5858
rect 246 -5862 250 -5858
rect 364 -5862 368 -5858
rect 572 -5862 576 -5858
rect 602 -5862 606 -5858
rect 720 -5862 724 -5858
rect 970 -5862 974 -5858
rect 1000 -5862 1004 -5858
rect 1118 -5862 1122 -5858
rect 1328 -5862 1332 -5858
rect 1358 -5862 1362 -5858
rect 1476 -5862 1480 -5858
rect -1203 -5871 -1199 -5867
rect -902 -5870 -898 -5866
rect -804 -5870 -800 -5866
rect -544 -5870 -540 -5866
rect -446 -5870 -442 -5866
rect -186 -5870 -182 -5866
rect -88 -5870 -84 -5866
rect 242 -5870 246 -5866
rect 340 -5870 344 -5866
rect 598 -5870 602 -5866
rect 696 -5870 700 -5866
rect 996 -5870 1000 -5866
rect 1094 -5870 1098 -5866
rect 1354 -5870 1358 -5866
rect 1452 -5870 1456 -5866
rect -1253 -5878 -1249 -5874
rect -1213 -5878 -1209 -5874
rect -1193 -5878 -1189 -5874
rect -924 -5877 -920 -5873
rect -776 -5877 -772 -5873
rect -566 -5877 -562 -5873
rect -418 -5877 -414 -5873
rect -208 -5877 -204 -5873
rect -60 -5877 -56 -5873
rect 220 -5877 224 -5873
rect 368 -5877 372 -5873
rect 576 -5877 580 -5873
rect 724 -5877 728 -5873
rect 974 -5877 978 -5873
rect 1122 -5877 1126 -5873
rect 1332 -5877 1336 -5873
rect 1480 -5877 1484 -5873
rect -1257 -5885 -1253 -5881
rect -1227 -5885 -1223 -5881
rect -1179 -5885 -1175 -5881
rect -902 -5884 -898 -5880
rect -794 -5884 -790 -5880
rect -760 -5884 -756 -5880
rect -544 -5884 -540 -5880
rect -436 -5884 -432 -5880
rect -402 -5884 -398 -5880
rect -186 -5884 -182 -5880
rect -78 -5884 -74 -5880
rect -44 -5884 -40 -5880
rect 242 -5884 246 -5880
rect 350 -5884 354 -5880
rect 384 -5884 388 -5880
rect 598 -5884 602 -5880
rect 706 -5884 710 -5880
rect 740 -5884 744 -5880
rect 996 -5884 1000 -5880
rect 1104 -5884 1108 -5880
rect 1138 -5884 1142 -5880
rect 1354 -5884 1358 -5880
rect 1462 -5884 1466 -5880
rect 1496 -5884 1500 -5880
rect -928 -5891 -924 -5887
rect -872 -5891 -868 -5887
rect -838 -5891 -834 -5887
rect -570 -5891 -566 -5887
rect -514 -5891 -510 -5887
rect -480 -5891 -476 -5887
rect -212 -5891 -208 -5887
rect -156 -5891 -152 -5887
rect -122 -5891 -118 -5887
rect 216 -5891 220 -5887
rect 272 -5891 276 -5887
rect 306 -5891 310 -5887
rect 572 -5891 576 -5887
rect 628 -5891 632 -5887
rect 662 -5891 666 -5887
rect 970 -5891 974 -5887
rect 1026 -5891 1030 -5887
rect 1060 -5891 1064 -5887
rect 1328 -5891 1332 -5887
rect 1384 -5891 1388 -5887
rect 1418 -5891 1422 -5887
rect -1237 -5993 -1233 -5989
rect -1199 -5993 -1195 -5989
rect -1139 -5993 -1135 -5989
rect -1115 -5993 -1111 -5989
rect -908 -5993 -904 -5989
rect -870 -5993 -866 -5989
rect -810 -5993 -806 -5989
rect -786 -5993 -782 -5989
rect -550 -5993 -546 -5989
rect -512 -5993 -508 -5989
rect -452 -5993 -448 -5989
rect -428 -5993 -424 -5989
rect -192 -5993 -188 -5989
rect -154 -5993 -150 -5989
rect -94 -5993 -90 -5989
rect -70 -5993 -66 -5989
rect 236 -5993 240 -5989
rect 274 -5993 278 -5989
rect 334 -5993 338 -5989
rect 358 -5993 362 -5989
rect 592 -5993 596 -5989
rect 630 -5993 634 -5989
rect 690 -5993 694 -5989
rect 714 -5993 718 -5989
rect 990 -5993 994 -5989
rect 1028 -5993 1032 -5989
rect 1088 -5993 1092 -5989
rect 1112 -5993 1116 -5989
rect 1348 -5993 1352 -5989
rect 1386 -5993 1390 -5989
rect 1446 -5993 1450 -5989
rect 1470 -5993 1474 -5989
rect -1257 -6001 -1253 -5997
rect -1223 -6001 -1219 -5997
rect -1171 -6001 -1167 -5997
rect -1111 -6001 -1107 -5997
rect -1073 -6001 -1069 -5997
rect -928 -6001 -924 -5997
rect -894 -6001 -890 -5997
rect -842 -6001 -838 -5997
rect -782 -6001 -778 -5997
rect -744 -6001 -740 -5997
rect -570 -6001 -566 -5997
rect -536 -6001 -532 -5997
rect -484 -6001 -480 -5997
rect -424 -6001 -420 -5997
rect -386 -6001 -382 -5997
rect -212 -6001 -208 -5997
rect -178 -6001 -174 -5997
rect -126 -6001 -122 -5997
rect -66 -6001 -62 -5997
rect -28 -6001 -24 -5997
rect 216 -6001 220 -5997
rect 250 -6001 254 -5997
rect 302 -6001 306 -5997
rect 362 -6001 366 -5997
rect 400 -6001 404 -5997
rect 572 -6001 576 -5997
rect 606 -6001 610 -5997
rect 658 -6001 662 -5997
rect 718 -6001 722 -5997
rect 756 -6001 760 -5997
rect 970 -6001 974 -5997
rect 1004 -6001 1008 -5997
rect 1056 -6001 1060 -5997
rect 1116 -6001 1120 -5997
rect 1154 -6001 1158 -5997
rect 1328 -6001 1332 -5997
rect 1362 -6001 1366 -5997
rect 1414 -6001 1418 -5997
rect 1474 -6001 1478 -5997
rect 1512 -6001 1516 -5997
rect -1213 -6008 -1209 -6004
rect -1181 -6008 -1177 -6004
rect -1129 -6008 -1125 -6004
rect -1097 -6008 -1093 -6004
rect -884 -6008 -880 -6004
rect -852 -6008 -848 -6004
rect -800 -6008 -796 -6004
rect -768 -6008 -764 -6004
rect -526 -6008 -522 -6004
rect -494 -6008 -490 -6004
rect -442 -6008 -438 -6004
rect -410 -6008 -406 -6004
rect -168 -6008 -164 -6004
rect -136 -6008 -132 -6004
rect -84 -6008 -80 -6004
rect -52 -6008 -48 -6004
rect 260 -6008 264 -6004
rect 292 -6008 296 -6004
rect 344 -6008 348 -6004
rect 376 -6008 380 -6004
rect 616 -6008 620 -6004
rect 648 -6008 652 -6004
rect 700 -6008 704 -6004
rect 732 -6008 736 -6004
rect 1014 -6008 1018 -6004
rect 1046 -6008 1050 -6004
rect 1098 -6008 1102 -6004
rect 1130 -6008 1134 -6004
rect 1372 -6008 1376 -6004
rect 1404 -6008 1408 -6004
rect 1456 -6008 1460 -6004
rect 1488 -6008 1492 -6004
rect -1253 -6015 -1249 -6011
rect -1139 -6015 -1135 -6011
rect -1087 -6015 -1083 -6011
rect -924 -6015 -920 -6011
rect -810 -6015 -806 -6011
rect -758 -6015 -754 -6011
rect -566 -6015 -562 -6011
rect -452 -6015 -448 -6011
rect -400 -6015 -396 -6011
rect -208 -6015 -204 -6011
rect -94 -6015 -90 -6011
rect -42 -6015 -38 -6011
rect 220 -6015 224 -6011
rect 334 -6015 338 -6011
rect 386 -6015 390 -6011
rect 576 -6015 580 -6011
rect 690 -6015 694 -6011
rect 742 -6015 746 -6011
rect 974 -6015 978 -6011
rect 1088 -6015 1092 -6011
rect 1140 -6015 1144 -6011
rect 1332 -6015 1336 -6011
rect 1446 -6015 1450 -6011
rect 1498 -6015 1502 -6011
rect -1195 -6022 -1191 -6018
rect -1157 -6022 -1153 -6018
rect -866 -6022 -862 -6018
rect -828 -6022 -824 -6018
rect -508 -6022 -504 -6018
rect -470 -6022 -466 -6018
rect -150 -6022 -146 -6018
rect -112 -6022 -108 -6018
rect 278 -6022 282 -6018
rect 316 -6022 320 -6018
rect 634 -6022 638 -6018
rect 672 -6022 676 -6018
rect 1032 -6022 1036 -6018
rect 1070 -6022 1074 -6018
rect 1390 -6022 1394 -6018
rect 1428 -6022 1432 -6018
rect 1348 -6111 1352 -6107
rect 1386 -6111 1390 -6107
rect 1446 -6111 1450 -6107
rect 1470 -6111 1474 -6107
rect 1328 -6119 1332 -6115
rect 1362 -6119 1366 -6115
rect 1414 -6119 1418 -6115
rect 1474 -6119 1478 -6115
rect 1512 -6119 1516 -6115
rect 1372 -6126 1376 -6122
rect 1404 -6126 1408 -6122
rect 1456 -6126 1460 -6122
rect 1488 -6126 1492 -6122
rect 1332 -6133 1336 -6129
rect 1446 -6133 1450 -6129
rect 1498 -6133 1502 -6129
rect 1390 -6140 1394 -6136
rect 1428 -6140 1432 -6136
<< labels >>
rlabel metal1 -942 -998 -938 -998 5 X1
rlabel metal1 -583 -999 -579 -999 5 X2
rlabel metal2 -19 -3728 -19 -3724 1 Z4
rlabel metal1 -225 -998 -221 -998 5 X3
rlabel metal2 409 -3006 409 -3002 1 Z3
rlabel metal1 203 -998 207 -998 5 X4
rlabel metal2 765 -2281 765 -2277 1 Z2
rlabel metal1 559 -998 563 -998 5 X5
rlabel metal2 765 -5993 765 -5989 1 Z12
rlabel metal2 409 -5993 409 -5989 1 Z11
rlabel metal2 -19 -5993 -19 -5989 1 Z10
rlabel metal2 -377 -4561 -377 -4557 1 Z5
rlabel metal2 -377 -5993 -377 -5989 1 Z9
rlabel metal2 -735 -5276 -735 -5272 1 Z6
rlabel metal2 -735 -5993 -735 -5989 1 Z8
rlabel metal2 1163 -5993 1163 -5989 1 Z13
rlabel metal2 1521 -5993 1521 -5989 1 Z14
rlabel metal2 1521 -6111 1521 -6107 1 Z15
rlabel metal1 1315 -998 1319 -998 5 X7
rlabel metal2 1665 -3461 1665 -3461 1 GND!
rlabel metal1 957 -998 961 -998 5 X6
rlabel metal2 1163 -1196 1163 -1192 1 Z0
rlabel metal2 1163 -1549 1163 -1545 1 Z1
rlabel metal2 -1064 -5993 -1064 -5989 1 Z7
rlabel metal2 -1421 -4216 -1421 -4212 1 Y5
rlabel metal2 -1421 -4929 -1421 -4925 1 Y6
rlabel metal2 -1421 -5642 -1421 -5638 1 Y7
rlabel metal2 -1421 -3365 -1421 -3361 1 Y4
rlabel metal2 -1421 -2663 -1421 -2659 1 Y3
rlabel metal2 -1421 -1914 -1421 -1910 1 Y2
rlabel metal2 -1421 -1304 -1421 -1300 1 Y1
rlabel metal2 -1421 -1074 -1421 -1070 1 Y0
rlabel metal2 -1464 -3462 -1464 -3462 1 VDD!
rlabel metal1 -1349 -998 -1345 -998 5 X0
rlabel metal1 -1629 -3851 -1629 -3837 3 CLK
<< end >>
