magic
tech scmos
timestamp 1612988437
<< ntransistor >>
rect 47 3 49 7
rect 55 3 57 7
rect 75 3 77 7
<< ptransistor >>
rect 47 24 49 33
rect 55 24 57 33
rect 75 24 77 33
<< ndiffusion >>
rect 46 3 47 7
rect 49 3 55 7
rect 57 3 58 7
rect 74 3 75 7
rect 77 3 78 7
<< pdiffusion >>
rect 46 24 47 33
rect 49 24 50 33
rect 54 24 55 33
rect 57 24 58 33
rect 74 24 75 33
rect 77 24 78 33
<< ndcontact >>
rect 42 3 46 7
rect 58 3 62 7
rect 70 3 74 7
rect 78 3 82 7
<< pdcontact >>
rect 42 24 46 33
rect 50 24 54 33
rect 58 24 62 33
rect 70 24 74 33
rect 78 24 82 33
<< psubstratepcontact >>
rect 42 -5 46 -1
rect 70 -5 74 -1
<< nsubstratencontact >>
rect 42 37 46 41
rect 58 37 62 41
rect 70 37 74 41
<< polysilicon >>
rect 47 33 49 35
rect 55 33 57 35
rect 75 33 77 35
rect 47 7 49 24
rect 55 14 57 24
rect 75 16 77 24
rect 74 12 77 16
rect 55 7 57 10
rect 75 7 77 12
rect 47 1 49 3
rect 55 1 57 3
rect 75 1 77 3
<< polycontact >>
rect 43 17 47 21
rect 53 10 57 14
rect 70 12 74 16
<< metal1 >>
rect 38 37 42 41
rect 46 37 58 41
rect 62 37 70 41
rect 74 37 86 41
rect 42 33 46 37
rect 58 33 62 37
rect 70 33 74 37
rect 50 21 54 24
rect 42 17 43 21
rect 50 17 66 21
rect 62 16 66 17
rect 78 16 82 24
rect 42 10 53 14
rect 62 12 70 16
rect 78 12 86 16
rect 62 3 66 12
rect 78 7 82 12
rect 42 -1 46 3
rect 70 -1 74 3
rect 38 -5 42 -1
rect 46 -5 70 -1
rect 74 -5 86 -1
<< labels >>
rlabel metal1 42 17 42 21 3 a
rlabel metal1 42 10 42 14 3 b
rlabel metal1 86 12 86 16 7 out
rlabel metal1 61 -3 61 -3 1 GND!
rlabel metal1 66 39 66 39 5 VDD!
<< end >>
