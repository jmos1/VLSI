magic
tech scmos
timestamp 1615651426
<< ntransistor >>
rect -100 -18 -98 -14
rect -84 -18 -82 -14
rect -68 -18 -66 -14
rect -60 -18 -58 -14
rect -41 -18 -39 -14
rect -33 -18 -31 -14
rect -14 -18 -12 -14
rect -6 -18 -4 -14
rect 13 -18 15 -14
rect 21 -18 23 -14
rect 40 -18 42 -14
rect 48 -18 50 -14
rect 67 -18 69 -14
rect 75 -18 77 -14
rect 94 -18 96 -14
rect 102 -18 104 -14
rect 121 -18 123 -14
rect 129 -18 131 -14
<< ptransistor >>
rect -100 38 -98 47
rect -84 38 -82 47
rect -68 38 -66 47
rect -60 38 -58 47
rect -41 38 -39 47
rect -33 38 -31 47
rect -14 38 -12 47
rect -6 38 -4 47
rect 13 38 15 47
rect 21 38 23 47
rect 40 38 42 47
rect 48 38 50 47
rect 67 38 69 47
rect 75 38 77 47
rect 94 38 96 47
rect 102 38 104 47
rect 121 38 123 47
rect 129 38 131 47
<< ndiffusion >>
rect -101 -18 -100 -14
rect -98 -18 -97 -14
rect -85 -18 -84 -14
rect -82 -18 -81 -14
rect -69 -18 -68 -14
rect -66 -18 -60 -14
rect -58 -18 -57 -14
rect -42 -18 -41 -14
rect -39 -18 -33 -14
rect -31 -18 -30 -14
rect -15 -18 -14 -14
rect -12 -18 -6 -14
rect -4 -18 -3 -14
rect 12 -18 13 -14
rect 15 -18 21 -14
rect 23 -18 24 -14
rect 39 -18 40 -14
rect 42 -18 48 -14
rect 50 -18 51 -14
rect 66 -18 67 -14
rect 69 -18 75 -14
rect 77 -18 78 -14
rect 93 -18 94 -14
rect 96 -18 102 -14
rect 104 -18 105 -14
rect 120 -18 121 -14
rect 123 -18 129 -14
rect 131 -18 132 -14
<< pdiffusion >>
rect -101 38 -100 47
rect -98 38 -97 47
rect -85 38 -84 47
rect -82 38 -81 47
rect -69 38 -68 47
rect -66 38 -65 47
rect -61 38 -60 47
rect -58 38 -51 47
rect -47 38 -41 47
rect -39 38 -38 47
rect -34 38 -33 47
rect -31 38 -24 47
rect -20 38 -14 47
rect -12 38 -11 47
rect -7 38 -6 47
rect -4 38 3 47
rect 7 38 13 47
rect 15 38 16 47
rect 20 38 21 47
rect 23 38 31 47
rect 35 38 40 47
rect 42 38 43 47
rect 47 38 48 47
rect 50 38 58 47
rect 62 38 67 47
rect 69 38 70 47
rect 74 38 75 47
rect 77 38 84 47
rect 88 38 94 47
rect 96 38 97 47
rect 101 38 102 47
rect 104 38 111 47
rect 115 38 121 47
rect 123 38 124 47
rect 128 38 129 47
rect 131 38 132 47
<< ndcontact >>
rect -105 -18 -101 -14
rect -97 -18 -93 -14
rect -89 -18 -85 -14
rect -81 -18 -77 -14
rect -73 -18 -69 -14
rect -57 -18 -53 -14
rect -46 -18 -42 -14
rect -30 -18 -26 -14
rect -19 -18 -15 -14
rect -3 -18 1 -14
rect 8 -18 12 -14
rect 24 -18 28 -14
rect 35 -18 39 -14
rect 51 -18 55 -14
rect 62 -18 66 -14
rect 78 -18 82 -14
rect 89 -18 93 -14
rect 105 -18 109 -14
rect 116 -18 120 -14
rect 132 -18 136 -14
<< pdcontact >>
rect -105 38 -101 47
rect -97 38 -93 47
rect -89 38 -85 47
rect -81 38 -77 47
rect -73 38 -69 47
rect -65 38 -61 47
rect -51 38 -47 47
rect -38 38 -34 47
rect -24 38 -20 47
rect -11 38 -7 47
rect 3 38 7 47
rect 16 38 20 47
rect 31 38 35 47
rect 43 38 47 47
rect 58 38 62 47
rect 70 38 74 47
rect 84 38 88 47
rect 97 38 101 47
rect 111 38 115 47
rect 124 38 128 47
rect 132 38 136 47
<< psubstratepcontact >>
rect -105 -26 -101 -22
rect -89 -26 -85 -22
rect -73 -26 -69 -22
rect -46 -26 -42 -22
rect -19 -26 -15 -22
rect 8 -26 12 -22
rect 35 -26 39 -22
rect 62 -26 66 -22
rect 89 -26 93 -22
rect 116 -26 120 -22
<< nsubstratencontact >>
rect -105 51 -101 55
rect -89 51 -85 55
rect -73 51 -69 55
rect -51 51 -47 55
rect -24 51 -20 55
rect 3 51 7 55
rect 31 51 35 55
rect 58 51 62 55
rect 84 51 88 55
rect 111 51 115 55
rect 132 51 136 55
<< polysilicon >>
rect -100 47 -98 49
rect -84 47 -82 49
rect -68 47 -66 49
rect -60 47 -58 49
rect -41 47 -39 49
rect -33 47 -31 49
rect -14 47 -12 49
rect -6 47 -4 49
rect 13 47 15 49
rect 21 47 23 49
rect 40 47 42 49
rect 48 47 50 49
rect 67 47 69 49
rect 75 47 77 49
rect 94 47 96 49
rect 102 47 104 49
rect 121 47 123 49
rect 129 47 131 49
rect -100 11 -98 38
rect -84 18 -82 38
rect -85 14 -82 18
rect -101 7 -98 11
rect -100 -14 -98 7
rect -84 -14 -82 14
rect -68 -14 -66 38
rect -60 11 -58 38
rect -60 -14 -58 7
rect -41 -14 -39 38
rect -33 11 -31 38
rect -33 -14 -31 7
rect -14 -14 -12 38
rect -6 11 -4 38
rect -6 -14 -4 7
rect 13 -14 15 38
rect 21 11 23 38
rect 21 -14 23 7
rect 40 -14 42 38
rect 48 11 50 38
rect 48 -14 50 7
rect 67 -14 69 38
rect 75 11 77 38
rect 75 -14 77 7
rect 94 -14 96 38
rect 102 11 104 38
rect 102 -14 104 7
rect 121 -14 123 38
rect 129 11 131 38
rect 129 -14 131 7
rect -100 -20 -98 -18
rect -84 -20 -82 -18
rect -68 -20 -66 -18
rect -60 -20 -58 -18
rect -41 -20 -39 -18
rect -33 -20 -31 -18
rect -14 -20 -12 -18
rect -6 -20 -4 -18
rect 13 -20 15 -18
rect 21 -20 23 -18
rect 40 -20 42 -18
rect 48 -20 50 -18
rect 67 -20 69 -18
rect 75 -20 77 -18
rect 94 -20 96 -18
rect 102 -20 104 -18
rect 121 -20 123 -18
rect 129 -20 131 -18
<< polycontact >>
rect 19 7 23 11
rect 127 7 131 11
<< metal1 >>
rect -109 51 -105 55
rect -101 51 -89 55
rect -85 51 -73 55
rect -69 51 -51 55
rect -47 51 -24 55
rect -20 51 3 55
rect 7 51 31 55
rect 35 51 58 55
rect 62 51 84 55
rect 88 51 111 55
rect 115 51 132 55
rect 136 51 140 55
rect -105 47 -101 51
rect -89 47 -85 51
rect -73 47 -69 51
rect -51 47 -47 51
rect -24 47 -20 51
rect 3 47 7 51
rect 31 47 35 51
rect 58 47 62 51
rect 84 47 88 51
rect 111 47 115 51
rect 132 47 136 51
rect -97 11 -93 38
rect -81 25 -77 38
rect -65 25 -61 38
rect -38 25 -34 38
rect -11 25 -7 38
rect 16 25 20 38
rect 43 25 47 38
rect 70 25 74 38
rect 97 25 101 38
rect -81 21 -73 25
rect -65 21 -46 25
rect -38 21 -19 25
rect -11 21 8 25
rect 16 21 35 25
rect 43 21 62 25
rect 70 21 89 25
rect 97 21 116 25
rect -97 7 -89 11
rect -97 -14 -93 7
rect -81 -14 -77 21
rect -65 18 -61 21
rect -38 18 -34 21
rect -11 18 -7 21
rect 16 18 20 21
rect 43 18 47 21
rect 70 18 74 21
rect 97 18 101 21
rect 124 18 128 38
rect -65 14 -49 18
rect -38 14 -22 18
rect -11 14 5 18
rect 16 14 32 18
rect 43 14 59 18
rect 70 14 86 18
rect 97 14 113 18
rect 124 14 140 18
rect -53 -18 -49 14
rect -26 -18 -22 14
rect 1 11 5 14
rect 28 11 32 14
rect 1 7 19 11
rect 1 -18 5 7
rect 28 -18 32 7
rect 55 -18 59 14
rect 82 -18 86 14
rect 109 11 113 14
rect 136 11 140 14
rect 109 7 127 11
rect 109 -18 113 7
rect 136 -18 140 7
rect -105 -22 -101 -18
rect -89 -22 -85 -18
rect -73 -22 -69 -18
rect -46 -22 -42 -18
rect -19 -22 -15 -18
rect 8 -22 12 -18
rect 35 -22 39 -18
rect 62 -22 66 -18
rect 89 -22 93 -18
rect 116 -22 120 -18
rect -109 -26 -105 -22
rect -101 -26 -89 -22
rect -85 -26 -73 -22
rect -69 -26 -46 -22
rect -42 -26 -19 -22
rect -15 -26 8 -22
rect 12 -26 35 -22
rect 39 -26 62 -22
rect 66 -26 89 -22
rect 93 -26 116 -22
rect 120 -26 140 -22
<< m2contact >>
rect -73 21 -69 25
rect -46 21 -42 25
rect -19 21 -15 25
rect 8 21 12 25
rect 35 21 39 25
rect 62 21 66 25
rect 89 21 93 25
rect 116 21 120 25
rect -89 7 -85 11
rect 28 7 32 11
rect 136 7 140 11
<< pm12contact >>
rect -89 14 -85 18
rect -105 7 -101 11
rect -72 14 -68 18
rect -45 14 -41 18
rect -18 14 -14 18
rect 9 14 13 18
rect 36 14 40 18
rect 63 14 67 18
rect 90 14 94 18
rect 117 14 121 18
rect -62 7 -58 11
rect -35 7 -31 11
rect -8 7 -4 11
rect 46 7 50 11
rect 73 7 77 11
rect 100 7 104 11
<< metal2 >>
rect -69 21 -61 25
rect -42 21 -34 25
rect -15 21 -7 25
rect 12 21 20 25
rect 39 21 47 25
rect 66 21 74 25
rect 93 21 101 25
rect 120 21 128 25
rect -65 18 -61 21
rect -38 18 -34 21
rect -11 18 -7 21
rect 16 18 20 21
rect 43 18 47 21
rect 70 18 74 21
rect 97 18 101 21
rect 124 18 128 21
rect -109 14 -89 18
rect -85 14 -72 18
rect -65 14 -45 18
rect -38 14 -18 18
rect -11 14 9 18
rect 16 14 36 18
rect 43 14 63 18
rect 70 14 90 18
rect 97 14 117 18
rect 124 14 140 18
rect -109 7 -105 11
rect -101 7 -93 11
rect -85 7 -62 11
rect -58 7 -35 11
rect -4 7 28 11
rect 36 7 46 11
rect 50 7 73 11
rect 104 7 136 11
rect -97 4 -93 7
rect 36 4 40 7
rect -97 0 40 4
<< labels >>
rlabel metal2 -109 7 -109 11 1 CLK
rlabel metal2 -109 14 -109 18 1 D
rlabel metal1 -9 -24 -9 -24 1 GND!
rlabel metal1 -9 53 -9 53 5 VDD!
rlabel metal2 140 14 140 18 1 Q
rlabel m2contact 140 7 140 11 1 QN
<< end >>
