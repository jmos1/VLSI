magic
tech scmos
timestamp 1613058019
<< ntransistor >>
rect -101 -13 -99 -9
rect -80 -13 -78 -9
rect -59 -13 -57 -9
rect -51 -13 -49 -9
rect -43 -13 -41 -9
rect -35 -13 -33 -9
rect -19 -13 -17 -9
rect -11 -13 -9 -9
rect 8 -13 10 -9
rect 38 -13 40 -9
rect 59 -13 61 -9
rect 80 -13 82 -9
rect 88 -13 90 -9
rect 96 -13 98 -9
rect 104 -13 106 -9
rect 120 -13 122 -9
rect 128 -13 130 -9
rect 147 -13 149 -9
rect 177 -17 179 -13
rect 185 -17 187 -13
rect 204 -17 206 -13
<< ptransistor >>
rect -101 28 -99 37
rect -80 28 -78 37
rect -59 28 -57 37
rect -51 28 -49 37
rect -43 28 -41 37
rect -35 28 -33 37
rect -19 28 -17 37
rect -11 28 -9 37
rect 8 28 10 37
rect 38 28 40 37
rect 59 28 61 37
rect 80 28 82 37
rect 88 28 90 37
rect 96 28 98 37
rect 104 28 106 37
rect 120 28 122 37
rect 128 28 130 37
rect 147 28 149 37
rect 177 28 179 37
rect 185 28 187 37
rect 204 28 206 37
<< ndiffusion >>
rect -102 -13 -101 -9
rect -99 -13 -98 -9
rect -81 -13 -80 -9
rect -78 -13 -77 -9
rect -60 -13 -59 -9
rect -57 -13 -51 -9
rect -49 -13 -48 -9
rect -44 -13 -43 -9
rect -41 -13 -35 -9
rect -33 -13 -32 -9
rect -20 -13 -19 -9
rect -17 -13 -11 -9
rect -9 -13 -8 -9
rect 7 -13 8 -9
rect 10 -13 11 -9
rect 37 -13 38 -9
rect 40 -13 41 -9
rect 58 -13 59 -9
rect 61 -13 62 -9
rect 79 -13 80 -9
rect 82 -13 88 -9
rect 90 -13 91 -9
rect 95 -13 96 -9
rect 98 -13 104 -9
rect 106 -13 107 -9
rect 119 -13 120 -9
rect 122 -13 128 -9
rect 130 -13 131 -9
rect 146 -13 147 -9
rect 149 -13 150 -9
rect 176 -17 177 -13
rect 179 -17 180 -13
rect 184 -17 185 -13
rect 187 -17 188 -13
rect 203 -17 204 -13
rect 206 -17 207 -13
<< pdiffusion >>
rect -102 28 -101 37
rect -99 28 -98 37
rect -81 28 -80 37
rect -78 28 -77 37
rect -60 28 -59 37
rect -57 28 -51 37
rect -49 28 -48 37
rect -44 28 -43 37
rect -41 28 -35 37
rect -33 28 -32 37
rect -20 28 -19 37
rect -17 28 -16 37
rect -12 28 -11 37
rect -9 28 -8 37
rect 7 28 8 37
rect 10 28 11 37
rect 37 28 38 37
rect 40 28 41 37
rect 58 28 59 37
rect 61 28 62 37
rect 79 28 80 37
rect 82 28 88 37
rect 90 28 91 37
rect 95 28 96 37
rect 98 28 104 37
rect 106 28 107 37
rect 119 28 120 37
rect 122 28 123 37
rect 127 28 128 37
rect 130 28 131 37
rect 146 28 147 37
rect 149 28 150 37
rect 176 28 177 37
rect 179 28 185 37
rect 187 28 188 37
rect 203 28 204 37
rect 206 28 207 37
<< ndcontact >>
rect -106 -13 -102 -9
rect -98 -13 -94 -9
rect -85 -13 -81 -9
rect -77 -13 -73 -9
rect -64 -13 -60 -9
rect -32 -13 -28 -9
rect -24 -13 -20 -9
rect -8 -13 -4 -9
rect 3 -13 7 -9
rect 11 -13 15 -9
rect 33 -13 37 -9
rect 41 -13 45 -9
rect 54 -13 58 -9
rect 62 -13 66 -9
rect 75 -13 79 -9
rect 107 -13 111 -9
rect 115 -13 119 -9
rect 131 -13 135 -9
rect 142 -13 146 -9
rect 150 -13 154 -9
rect 172 -17 176 -13
rect 180 -17 184 -13
rect 188 -17 192 -13
rect 199 -17 203 -13
rect 207 -17 211 -13
<< pdcontact >>
rect -106 28 -102 37
rect -98 28 -94 37
rect -85 28 -81 37
rect -77 28 -73 37
rect -64 28 -60 37
rect -32 28 -28 37
rect -24 28 -20 37
rect -16 28 -12 37
rect -8 28 -4 37
rect 3 28 7 37
rect 11 28 15 37
rect 33 28 37 37
rect 41 28 45 37
rect 54 28 58 37
rect 62 28 66 37
rect 75 28 79 37
rect 107 28 111 37
rect 115 28 119 37
rect 123 28 127 37
rect 131 28 135 37
rect 142 28 146 37
rect 150 28 154 37
rect 172 28 176 37
rect 188 28 192 37
rect 199 28 203 37
rect 207 28 211 37
<< psubstratepcontact >>
rect -106 -25 -102 -21
rect -85 -25 -81 -21
rect -64 -25 -60 -21
rect -32 -25 -28 -21
rect -24 -25 -20 -21
rect 3 -25 7 -21
rect 33 -25 37 -21
rect 54 -25 58 -21
rect 75 -25 79 -21
rect 107 -25 111 -21
rect 115 -25 119 -21
rect 142 -25 146 -21
rect 172 -25 176 -21
rect 188 -25 192 -21
rect 199 -25 203 -21
<< nsubstratencontact >>
rect -106 50 -102 54
rect -85 50 -81 54
rect -64 50 -60 54
rect -32 50 -28 54
rect -24 50 -20 54
rect -8 50 -4 54
rect 3 50 7 54
rect 33 50 37 54
rect 54 50 58 54
rect 75 50 79 54
rect 107 50 111 54
rect 115 50 119 54
rect 131 50 135 54
rect 142 50 146 54
rect 172 50 176 54
rect 199 50 203 54
<< polysilicon >>
rect -101 47 -33 49
rect -101 37 -99 47
rect -80 42 -49 44
rect -80 37 -78 42
rect -59 37 -57 39
rect -51 37 -49 42
rect -43 37 -41 39
rect -35 37 -33 47
rect 38 47 106 49
rect -19 37 -17 39
rect -11 37 -9 39
rect 8 37 10 39
rect 38 37 40 47
rect 59 42 90 44
rect 59 37 61 42
rect 80 37 82 39
rect 88 37 90 42
rect 96 37 98 39
rect 104 37 106 47
rect 120 37 122 39
rect 128 37 130 39
rect 147 37 149 39
rect 177 37 179 39
rect 185 37 187 39
rect 204 37 206 39
rect -101 20 -99 28
rect -80 20 -78 28
rect -59 25 -57 28
rect -51 26 -49 28
rect -102 16 -99 20
rect -81 16 -78 20
rect -101 -9 -99 16
rect -80 -9 -78 16
rect -59 15 -57 21
rect -43 20 -41 28
rect -35 25 -33 28
rect -35 23 -25 25
rect -43 18 -33 20
rect -59 13 -41 15
rect -59 -9 -57 -7
rect -51 -9 -49 -7
rect -43 -9 -41 13
rect -35 -9 -33 14
rect -101 -15 -99 -13
rect -80 -16 -78 -13
rect -59 -16 -57 -13
rect -80 -18 -57 -16
rect -51 -18 -49 -13
rect -43 -15 -41 -13
rect -35 -15 -33 -13
rect -27 -18 -25 23
rect -19 11 -17 28
rect -19 -9 -17 7
rect -11 4 -9 28
rect 8 25 10 28
rect 7 21 10 25
rect -11 -9 -9 0
rect 8 -9 10 21
rect 38 20 40 28
rect 59 20 61 28
rect 80 25 82 28
rect 88 26 90 28
rect 37 16 40 20
rect 58 16 61 20
rect 38 -9 40 16
rect 59 -9 61 16
rect 80 15 82 21
rect 96 20 98 28
rect 104 25 106 28
rect 104 23 114 25
rect 96 18 106 20
rect 80 13 98 15
rect 80 -9 82 -7
rect 88 -9 90 -7
rect 96 -9 98 13
rect 104 -9 106 14
rect -19 -15 -17 -13
rect -11 -15 -9 -13
rect 8 -15 10 -13
rect 38 -15 40 -13
rect 59 -16 61 -13
rect 80 -16 82 -13
rect 59 -18 82 -16
rect 88 -18 90 -13
rect 96 -15 98 -13
rect 104 -15 106 -13
rect 112 -18 114 23
rect 120 11 122 28
rect 120 -9 122 7
rect 128 4 130 28
rect 147 25 149 28
rect 146 21 149 25
rect 128 -9 130 0
rect 147 -9 149 21
rect 177 20 179 28
rect 177 -13 179 16
rect 185 13 187 28
rect 204 15 206 28
rect 203 11 206 15
rect 185 -13 187 9
rect 204 -13 206 11
rect 120 -15 122 -13
rect 128 -15 130 -13
rect 147 -15 149 -13
rect -51 -20 -25 -18
rect 88 -20 114 -18
rect 177 -19 179 -17
rect 185 -19 187 -17
rect 204 -19 206 -17
<< polycontact >>
rect -85 16 -81 20
rect -37 14 -33 18
rect 3 21 7 25
rect 54 16 58 20
rect 102 14 106 18
rect 142 21 146 25
rect 183 9 187 13
rect 199 11 203 15
<< metal1 >>
rect -110 50 -106 54
rect -102 50 -85 54
rect -81 50 -64 54
rect -60 50 -32 54
rect -28 50 -24 54
rect -20 50 -8 54
rect -4 50 3 54
rect 7 50 33 54
rect 37 50 54 54
rect 58 50 75 54
rect 79 50 107 54
rect 111 50 115 54
rect 119 50 131 54
rect 135 50 142 54
rect 146 50 172 54
rect 176 50 199 54
rect 203 50 215 54
rect -106 37 -102 50
rect -85 37 -81 50
rect -64 37 -60 50
rect -32 37 -28 50
rect -24 37 -20 50
rect -8 37 -4 50
rect 3 37 7 50
rect 33 37 37 50
rect 54 37 58 50
rect 75 37 79 50
rect 107 37 111 50
rect 115 37 119 50
rect 131 37 135 50
rect 142 37 146 50
rect 172 37 176 50
rect 199 37 203 50
rect -98 -9 -94 28
rect -85 4 -81 16
rect -77 18 -73 28
rect -16 25 -12 28
rect -16 21 3 25
rect -77 14 -37 18
rect -77 -9 -73 14
rect -106 -21 -102 -13
rect -85 -21 -81 -13
rect -64 -21 -60 -13
rect -32 -21 -28 -13
rect -4 -13 0 21
rect 11 -9 15 28
rect 41 -9 45 28
rect 54 4 58 16
rect 62 18 66 28
rect 123 25 127 28
rect 123 21 142 25
rect 62 14 102 18
rect 62 -9 66 14
rect -24 -21 -20 -13
rect 3 -21 7 -13
rect 33 -21 37 -13
rect 54 -21 58 -13
rect 75 -21 79 -13
rect 107 -21 111 -13
rect 135 -13 139 21
rect 150 13 154 28
rect 192 15 196 37
rect 207 15 211 28
rect 150 9 183 13
rect 192 11 199 15
rect 207 11 215 15
rect 150 -9 154 9
rect 192 6 196 11
rect 180 2 196 6
rect 180 -13 184 2
rect 207 -13 211 11
rect 115 -21 119 -13
rect 142 -21 146 -13
rect 172 -21 176 -17
rect 188 -21 192 -17
rect 199 -21 203 -17
rect -110 -25 -106 -21
rect -102 -25 -85 -21
rect -81 -25 -64 -21
rect -60 -25 -32 -21
rect -28 -25 -24 -21
rect -20 -25 3 -21
rect 7 -25 33 -21
rect 37 -25 54 -21
rect 58 -25 75 -21
rect 79 -25 107 -21
rect 111 -25 115 -21
rect 119 -25 142 -21
rect 146 -25 172 -21
rect 176 -25 188 -21
rect 192 -25 199 -21
rect 203 -25 215 -21
<< m2contact >>
rect -94 21 -90 25
rect -85 0 -81 4
rect 45 21 49 25
rect 54 0 58 4
<< pm12contact >>
rect -106 16 -102 20
rect -61 21 -57 25
rect -21 7 -17 11
rect -13 0 -9 4
rect 15 20 19 24
rect 33 16 37 20
rect 78 21 82 25
rect 118 7 122 11
rect 126 0 130 4
rect 175 16 179 20
<< pdm12contact >>
rect -48 28 -44 37
rect 91 28 95 37
<< ndm12contact >>
rect -48 -13 -44 -9
rect 91 -13 95 -9
<< metal2 >>
rect 19 41 159 45
rect -48 25 -44 28
rect -90 21 -61 25
rect -48 21 0 25
rect -106 11 -102 16
rect -4 11 0 21
rect 19 20 23 41
rect 91 25 95 28
rect 49 21 78 25
rect 91 21 139 25
rect 33 11 37 16
rect -110 7 -21 11
rect -4 7 118 11
rect -110 0 -85 4
rect -81 0 -13 4
rect -4 -3 0 7
rect 135 6 139 21
rect 155 20 159 41
rect 155 16 175 20
rect -48 -7 0 -3
rect 19 0 54 4
rect 58 0 126 4
rect 135 2 215 6
rect -48 -9 -44 -7
rect 19 -16 23 0
rect 135 -3 139 2
rect 91 -7 139 -3
rect 91 -9 95 -7
rect -110 -20 23 -16
<< labels >>
rlabel metal2 -110 0 -110 4 3 b
rlabel metal2 -110 7 -110 11 3 a
rlabel metal2 215 2 215 6 7 sum
rlabel metal2 -110 -20 -110 -16 3 cin
rlabel metal1 67 53 67 53 5 VDD!
rlabel metal1 68 -24 68 -24 1 GND!
rlabel metal1 215 11 215 15 7 cout
<< end >>
